module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n201 , n202 , n203 , n204 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n273 , n274 , n275 , n276 , n277 ;
  assign n65 = x59 ^ x27 ;
  assign n69 = x25 & x57 ;
  assign n67 = x27 & ~x59 ;
  assign n66 = x58 ^ x57 ;
  assign n68 = n67 ^ n66 ;
  assign n70 = n69 ^ n68 ;
  assign n73 = x59 ^ x26 ;
  assign n71 = x59 ^ x58 ;
  assign n72 = n71 ^ n67 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~n70 & ~n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = ~n65 & n76 ;
  assign n78 = n77 ^ x27 ;
  assign n79 = x28 & ~x60 ;
  assign n80 = n79 ^ x29 ;
  assign n81 = ~x31 & x63 ;
  assign n82 = ~n79 & n81 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = ~x61 & ~n83 ;
  assign n85 = n80 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = x30 & ~x62 ;
  assign n88 = ~n86 & n87 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = n78 & ~n89 ;
  assign n138 = n69 ^ x25 ;
  assign n139 = ~n67 & ~n138 ;
  assign n140 = x26 & ~x58 ;
  assign n141 = n139 & n140 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = ~x24 & n142 ;
  assign n91 = x51 ^ x19 ;
  assign n94 = x16 & ~x48 ;
  assign n93 = x48 ^ x16 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = n95 ^ x50 ;
  assign n92 = x50 ^ x17 ;
  assign n97 = n96 ^ n92 ;
  assign n98 = x50 ^ x49 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = ~n97 & n99 ;
  assign n101 = n100 ^ n96 ;
  assign n103 = x51 ^ x18 ;
  assign n102 = x51 ^ x50 ;
  assign n104 = n103 ^ n102 ;
  assign n105 = ~n101 & ~n104 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = ~n91 & n106 ;
  assign n108 = n107 ^ x19 ;
  assign n109 = x20 & ~x52 ;
  assign n110 = x21 & ~x53 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = n111 ^ n109 ;
  assign n113 = x22 & ~x54 ;
  assign n114 = ~n112 & n113 ;
  assign n115 = n114 ^ n112 ;
  assign n116 = x23 & ~x55 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = ~n108 & ~n118 ;
  assign n120 = x55 ^ x23 ;
  assign n122 = x52 ^ x20 ;
  assign n123 = n122 ^ n109 ;
  assign n124 = n123 ^ x54 ;
  assign n121 = x54 ^ x21 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = x54 ^ x53 ;
  assign n127 = n126 ^ n124 ;
  assign n128 = ~n125 & n127 ;
  assign n129 = n128 ^ n124 ;
  assign n131 = x55 ^ x22 ;
  assign n130 = x55 ^ x54 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = ~n129 & ~n132 ;
  assign n134 = n133 ^ n131 ;
  assign n135 = ~n120 & n134 ;
  assign n136 = n135 ^ x23 ;
  assign n137 = ~n119 & n136 ;
  assign n144 = n143 ^ n137 ;
  assign n145 = x56 & n142 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = ~n144 & n146 ;
  assign n148 = n147 ^ n143 ;
  assign n149 = n90 & ~n148 ;
  assign n150 = n149 ^ n89 ;
  assign n151 = x63 ^ x31 ;
  assign n155 = x62 ^ x61 ;
  assign n152 = x60 ^ x28 ;
  assign n153 = n152 ^ n79 ;
  assign n154 = n153 ^ x62 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = x62 ^ x29 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n156 & ~n158 ;
  assign n160 = n159 ^ n154 ;
  assign n162 = x63 ^ x30 ;
  assign n161 = x63 ^ x62 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = ~n160 & ~n163 ;
  assign n165 = n164 ^ n162 ;
  assign n166 = ~n151 & ~n165 ;
  assign n167 = n166 ^ x31 ;
  assign n168 = x47 ^ x15 ;
  assign n170 = x14 & ~x46 ;
  assign n169 = x46 ^ x14 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = n171 ^ x47 ;
  assign n173 = ~n168 & ~n172 ;
  assign n174 = n173 ^ x15 ;
  assign n175 = x45 ^ x13 ;
  assign n177 = x12 & ~x44 ;
  assign n176 = x44 ^ x12 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n178 ^ x45 ;
  assign n180 = ~n175 & ~n179 ;
  assign n181 = n180 ^ x13 ;
  assign n182 = ~n175 & ~n177 ;
  assign n183 = ~n168 & ~n170 ;
  assign n184 = x42 ^ x10 ;
  assign n185 = x43 ^ x11 ;
  assign n186 = ~n184 & ~n185 ;
  assign n188 = ~x9 & x41 ;
  assign n187 = x41 ^ x9 ;
  assign n189 = n188 ^ n187 ;
  assign n192 = ~x8 & ~n189 ;
  assign n193 = n186 & n192 ;
  assign n190 = x40 & ~n189 ;
  assign n191 = n186 & n190 ;
  assign n194 = n193 ^ n191 ;
  assign n229 = n191 ^ x39 ;
  assign n195 = x38 ^ x6 ;
  assign n196 = x5 & x37 ;
  assign n197 = n196 ^ x5 ;
  assign n198 = x36 ^ x4 ;
  assign n201 = x34 ^ x2 ;
  assign n203 = x34 ^ x1 ;
  assign n202 = x34 ^ x33 ;
  assign n204 = n203 ^ n202 ;
  assign n206 = x0 & ~x32 ;
  assign n207 = n206 ^ x1 ;
  assign n208 = ~n204 & n207 ;
  assign n209 = n208 ^ n203 ;
  assign n210 = ~n201 & n209 ;
  assign n199 = x35 ^ x2 ;
  assign n211 = n210 ^ n199 ;
  assign n213 = x36 ^ x3 ;
  assign n212 = x36 ^ x35 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n211 & ~n214 ;
  assign n216 = n215 ^ n213 ;
  assign n217 = ~n198 & n216 ;
  assign n218 = n217 ^ x4 ;
  assign n219 = ~n197 & ~n218 ;
  assign n220 = ~n195 & n219 ;
  assign n221 = x7 & ~x39 ;
  assign n222 = n221 ^ n195 ;
  assign n223 = n196 ^ x37 ;
  assign n224 = n223 ^ x6 ;
  assign n225 = ~n222 & ~n224 ;
  assign n226 = n225 ^ x6 ;
  assign n227 = ~n220 & n226 ;
  assign n228 = n227 ^ n191 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n191 ^ x7 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = ~n230 & ~n232 ;
  assign n234 = n233 ^ n229 ;
  assign n235 = n194 & ~n234 ;
  assign n236 = n235 ^ n193 ;
  assign n240 = n188 ^ x43 ;
  assign n237 = x43 ^ x42 ;
  assign n241 = n240 ^ n237 ;
  assign n242 = ~n184 & n241 ;
  assign n243 = n242 ^ n237 ;
  assign n244 = ~n185 & n243 ;
  assign n245 = n244 ^ x43 ;
  assign n246 = ~n236 & ~n245 ;
  assign n247 = n183 & ~n246 ;
  assign n248 = n182 & n247 ;
  assign n249 = n248 ^ n183 ;
  assign n250 = n181 & n249 ;
  assign n251 = n250 ^ n183 ;
  assign n252 = n174 & ~n251 ;
  assign n253 = ~n94 & ~n252 ;
  assign n254 = ~n118 & n253 ;
  assign n255 = ~n89 & n254 ;
  assign n256 = ~n167 & n255 ;
  assign n257 = x17 & ~x49 ;
  assign n258 = n256 & n257 ;
  assign n259 = n258 ^ n256 ;
  assign n260 = x18 & ~x50 ;
  assign n261 = n259 & n260 ;
  assign n262 = n261 ^ n259 ;
  assign n263 = x19 & ~x51 ;
  assign n264 = n262 & n263 ;
  assign n265 = n264 ^ n262 ;
  assign n273 = ~n145 & n265 ;
  assign n274 = ~n143 & n273 ;
  assign n275 = n274 ^ n143 ;
  assign n266 = n265 ^ n167 ;
  assign n267 = n266 ^ n143 ;
  assign n276 = n275 ^ n267 ;
  assign n277 = n150 & ~n276 ;
  assign y0 = ~n277 ;
endmodule
