module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n348 , n349 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n600 , n601 , n602 , n603 , n604 , n605 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3242 , n3243 , n3244 , n3245 , n3246 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3724 , n3725 , n3726 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4416 , n4417 , n4418 , n4419 , n4420 , n4423 , n4424 , n4425 , n4426 , n4427 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4536 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4610 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4896 , n4897 , n4898 , n4899 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5696 , n5697 , n5698 , n5699 , n5700 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5875 , n5876 , n5877 , n5878 , n5879 , n5881 , n5882 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5946 , n5947 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6087 , n6088 , n6089 , n6091 , n6092 , n6093 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6350 , n6351 , n6352 , n6353 , n6354 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6446 , n6447 , n6448 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6652 , n6653 , n6655 , n6656 , n6657 , n6658 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6679 , n6680 , n6681 , n6683 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6849 , n6850 , n6851 , n6852 , n6853 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6947 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7090 , n7091 , n7092 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7140 , n7141 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7224 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7611 , n7612 , n7613 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7640 , n7641 , n7642 , n7643 , n7644 , n7647 , n7648 , n7649 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7982 , n7983 , n7984 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8074 , n8075 , n8076 , n8077 , n8078 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8420 , n8421 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8469 , n8470 , n8471 , n8472 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8508 , n8509 , n8510 , n8511 , n8512 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8550 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8574 , n8575 , n8576 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8601 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8622 , n8623 , n8624 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8654 , n8655 , n8656 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8684 , n8685 , n8686 , n8689 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8796 , n8797 , n8798 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8829 , n8830 , n8831 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8909 , n8910 , n8911 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8943 , n8944 , n8945 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8995 , n8996 , n8997 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9293 , n9295 , n9297 , n9298 , n9301 , n9302 , n9303 , n9304 , n9308 , n9310 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9337 , n9365 , n9366 , n9367 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9577 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9821 , n9823 , n9825 , n9826 , n9829 , n9830 , n9831 , n9832 , n9836 , n9838 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9865 , n9893 , n9894 , n9895 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10364 , n10365 , n10366 , n10367 , n10369 , n10370 , n10375 , n10408 , n10411 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10421 , n10422 , n10424 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10712 , n10713 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10743 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10778 , n10779 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10799 , n10800 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10817 , n10818 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10877 , n10878 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10895 , n10896 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10930 , n10931 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10976 , n10977 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11008 , n11009 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11026 , n11027 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11058 , n11059 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11077 , n11078 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11113 , n11114 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11130 , n11131 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11196 , n11197 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11229 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11991 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12065 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12600 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12674 , n12675 , n12676 , n12677 , n12678 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12854 , n12855 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12945 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12961 , n12962 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14376 , n14377 , n14378 , n14379 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14921 , n14922 , n14923 , n14924 , n14925 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15442 , n15443 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16391 , n16392 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17495 , n17496 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17541 , n17542 , n17548 , n17549 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17568 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17626 , n17629 , n17630 , n17631 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17694 , n17698 , n17699 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17719 , n17725 , n17726 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17951 , n17956 , n17957 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19414 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19861 , n19862 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19898 , n19899 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19931 , n19932 , n19933 , n19934 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19975 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20726 , n20727 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21318 , n21319 , n21320 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22640 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22878 , n22879 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23066 , n23067 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23086 , n23087 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23102 , n23103 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23120 , n23121 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23136 , n23137 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23173 , n23174 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23191 , n23192 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23208 , n23209 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23226 , n23227 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23303 , n23304 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23456 , n23458 , n23459 , n23460 , n23461 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23952 , n23953 , n23956 , n23957 , n23958 , n23959 , n23960 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24476 , n24478 , n24479 , n24480 , n24482 , n24483 , n24490 , n24491 , n24492 , n24493 , n24494 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24510 , n24513 , n24515 , n24516 , n24517 , n24521 , n24522 , n24523 , n24524 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24543 , n24544 , n24545 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24555 , n24556 , n24557 , n24558 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24573 , n24577 , n24578 , n24584 , n24585 , n24586 , n24587 , n24590 , n24593 , n24594 , n24595 , n24597 , n24598 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24622 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25121 , n25122 , n25123 , n25124 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26874 , n26875 , n26876 , n26877 , n26878 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27690 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28319 , n28320 , n28321 , n28322 , n28323 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28500 , n28501 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28966 , n28967 , n28968 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29179 , n29180 , n29181 , n29182 , n29183 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29525 , n29526 , n29527 , n29528 , n29529 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29660 , n29661 , n29662 , n29663 , n29664 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 ;
  assign n10850 = ~x0 & x1 ;
  assign n825 = x26 & x27 ;
  assign n829 = x28 & n825 ;
  assign n826 = n825 ^ x28 ;
  assign n650 = x27 ^ x26 ;
  assign n654 = ~x28 & n650 ;
  assign n827 = n826 ^ n654 ;
  assign n24688 = n829 ^ n827 ;
  assign n33 = ~x29 & ~x30 ;
  assign n44 = x27 & x28 ;
  assign n45 = n33 & n44 ;
  assign n262 = x26 & n45 ;
  assign n24694 = n24688 ^ n262 ;
  assign n36 = x25 & ~x26 ;
  assign n37 = n36 ^ x25 ;
  assign n38 = n37 ^ x26 ;
  assign n77 = n38 ^ x25 ;
  assign n39 = ~x23 & ~x24 ;
  assign n73 = ~x25 & n39 ;
  assign n53 = x24 & x25 ;
  assign n52 = x25 ^ x24 ;
  assign n54 = n53 ^ n52 ;
  assign n74 = n73 ^ n54 ;
  assign n72 = ~x23 & ~x25 ;
  assign n75 = n74 ^ n72 ;
  assign n40 = n39 ^ x24 ;
  assign n41 = n40 ^ x23 ;
  assign n42 = n38 & n41 ;
  assign n76 = n75 ^ n42 ;
  assign n78 = n77 ^ n76 ;
  assign n69 = ~x26 & n39 ;
  assign n64 = x24 ^ x23 ;
  assign n65 = x26 & ~n64 ;
  assign n66 = n65 ^ x26 ;
  assign n67 = n66 ^ n64 ;
  assign n68 = n67 ^ x26 ;
  assign n70 = n69 ^ n68 ;
  assign n60 = ~x24 & ~x26 ;
  assign n61 = n60 ^ x26 ;
  assign n57 = x26 & n54 ;
  assign n58 = n57 ^ x26 ;
  assign n55 = n54 ^ x26 ;
  assign n56 = n55 ^ n36 ;
  assign n59 = n58 ^ n56 ;
  assign n62 = n61 ^ n59 ;
  assign n71 = n70 ^ n62 ;
  assign n79 = n78 ^ n71 ;
  assign n80 = n79 ^ n62 ;
  assign n34 = n33 ^ x29 ;
  assign n35 = n34 ^ x30 ;
  assign n95 = n35 ^ x29 ;
  assign n248 = n44 & ~n95 ;
  assign n703 = ~n80 & n248 ;
  assign n81 = x23 & n36 ;
  assign n533 = n81 & n248 ;
  assign n1148 = n703 ^ n533 ;
  assign n50 = n44 ^ x27 ;
  assign n51 = n33 & n50 ;
  assign n47 = ~x28 & n33 ;
  assign n254 = n51 ^ n47 ;
  assign n428 = n81 & n254 ;
  assign n1050 = x24 & n428 ;
  assign n429 = n1050 ^ n428 ;
  assign n46 = n45 ^ n33 ;
  assign n48 = n47 ^ n46 ;
  assign n138 = n74 ^ x24 ;
  assign n139 = n138 ^ n39 ;
  assign n82 = n81 ^ n80 ;
  assign n140 = n139 ^ n82 ;
  assign n186 = n48 & ~n140 ;
  assign n720 = n429 ^ n186 ;
  assign n722 = n1148 ^ n720 ;
  assign n89 = ~n35 & n44 ;
  assign n126 = n53 ^ x26 ;
  assign n127 = n126 ^ n62 ;
  assign n111 = n75 ^ x25 ;
  assign n112 = n111 ^ n41 ;
  assign n113 = n112 ^ x26 ;
  assign n114 = n113 ^ n80 ;
  assign n128 = n127 ^ n114 ;
  assign n212 = n89 & ~n128 ;
  assign n12859 = ~n73 & ~n114 ;
  assign n12858 = n114 ^ n73 ;
  assign n12860 = n12859 ^ n12858 ;
  assign n86 = ~n12860 ^ n58 ;
  assign n90 = n86 & n89 ;
  assign n716 = n212 ^ n90 ;
  assign n98 = n69 ^ n39 ;
  assign n105 = ~n12860 ^ n98 ;
  assign n94 = n44 ^ x28 ;
  assign n341 = ~n35 & n94 ;
  assign n426 = n105 & n341 ;
  assign n425 = ~n128 & n341 ;
  assign n427 = n426 ^ n425 ;
  assign n141 = n89 & ~n140 ;
  assign n715 = n427 ^ n141 ;
  assign n717 = n716 ^ n715 ;
  assign n269 = n254 & ~n12860 ;
  assign n718 = n717 ^ n269 ;
  assign n612 = n79 & n248 ;
  assign n241 = n50 & ~n95 ;
  assign n242 = ~n128 & n241 ;
  assign n712 = n612 ^ n242 ;
  assign n169 = n69 ^ n60 ;
  assign n170 = n169 ^ n82 ;
  assign n416 = ~n170 & n241 ;
  assign n96 = n94 & ~n95 ;
  assign n115 = n114 ^ x26 ;
  assign n291 = n96 & n115 ;
  assign n710 = n416 ^ n291 ;
  assign n406 = n48 & n169 ;
  assign n396 = n48 & ~n82 ;
  assign n407 = n406 ^ n396 ;
  assign n405 = n51 & ~n128 ;
  assign n408 = n407 ^ n405 ;
  assign n711 = n710 ^ n408 ;
  assign n713 = n712 ^ n711 ;
  assign n107 = n57 ^ n37 ;
  assign n43 = n42 ^ n38 ;
  assign n108 = n107 ^ n43 ;
  assign n171 = ~n34 & n44 ;
  assign n321 = n108 & n171 ;
  assign n245 = n78 & n171 ;
  assign n322 = n321 ^ n245 ;
  assign n63 = n62 ^ n36 ;
  assign n83 = n82 ^ n63 ;
  assign n130 = n83 & n96 ;
  assign n708 = n322 ^ n130 ;
  assign n292 = n83 & n248 ;
  assign n205 = n96 & n111 ;
  assign n204 = n43 & n96 ;
  assign n206 = n205 ^ n204 ;
  assign n705 = n292 ^ n206 ;
  assign n129 = n96 & ~n128 ;
  assign n704 = n703 ^ n129 ;
  assign n706 = n705 ^ n704 ;
  assign n702 = n108 & n241 ;
  assign n707 = n706 ^ n702 ;
  assign n709 = n708 ^ n707 ;
  assign n714 = n713 ^ n709 ;
  assign n719 = n718 ^ n714 ;
  assign n723 = n722 ^ n719 ;
  assign n661 = n79 & n241 ;
  assign n660 = n43 & n241 ;
  assign n662 = n661 ^ n660 ;
  assign n259 = n83 & n171 ;
  assign n258 = n115 & n241 ;
  assign n260 = n259 ^ n258 ;
  assign n12690 = n662 ^ n260 ;
  assign n309 = n58 & n171 ;
  assign n12691 = n12690 ^ n309 ;
  assign n281 = ~n62 & n171 ;
  assign n12692 = n12691 ^ n281 ;
  assign n438 = n48 & ~n70 ;
  assign n228 = n48 & n107 ;
  assign n3925 = n438 ^ n228 ;
  assign n409 = n51 & n115 ;
  assign n3926 = n3925 ^ n409 ;
  assign n3927 = n3926 ^ n48 ;
  assign n3928 = ~x23 & ~n77 ;
  assign n3929 = n45 & n3928 ;
  assign n239 = n51 & ~n140 ;
  assign n216 = n48 & ~n128 ;
  assign n2627 = n239 ^ n216 ;
  assign n3930 = n3929 ^ n2627 ;
  assign n3931 = ~n3927 & ~n3930 ;
  assign n12693 = n12692 ^ n3931 ;
  assign n394 = n48 & n78 ;
  assign n176 = n45 & ~n170 ;
  assign n5012 = n394 ^ n176 ;
  assign n308 = ~n82 & n171 ;
  assign n5010 = n308 ^ n228 ;
  assign n122 = n96 & n108 ;
  assign n5011 = n5010 ^ n122 ;
  assign n5013 = n5012 ^ n5011 ;
  assign n433 = n79 & n254 ;
  assign n400 = n83 & n241 ;
  assign n1513 = n433 ^ n400 ;
  assign n1029 = n241 & ~n12860 ;
  assign n244 = n96 & ~n170 ;
  assign n1030 = n1029 ^ n244 ;
  assign n5008 = n1513 ^ n1030 ;
  assign n298 = n86 & n254 ;
  assign n84 = n83 ^ n69 ;
  assign n268 = n84 & n96 ;
  assign n5006 = n298 ^ n268 ;
  assign n549 = x26 & n248 ;
  assign n626 = ~n73 & n549 ;
  assign n627 = n626 ^ n549 ;
  assign n203 = n79 & n96 ;
  assign n1876 = n627 ^ n203 ;
  assign n5007 = n5006 ^ n1876 ;
  assign n5009 = n5008 ^ n5007 ;
  assign n5014 = n5013 ^ n5009 ;
  assign n12694 = n12693 ^ n5014 ;
  assign n12695 = ~n723 & n12694 ;
  assign n456 = n105 & n241 ;
  assign n455 = ~n140 & n241 ;
  assign n457 = n456 ^ n455 ;
  assign n133 = n39 ^ x23 ;
  assign n134 = n133 ^ n59 ;
  assign n135 = n134 ^ n78 ;
  assign n136 = n135 ^ n133 ;
  assign n279 = n96 & n136 ;
  assign n458 = n457 ^ n279 ;
  assign n402 = n59 & n241 ;
  assign n459 = n458 ^ n402 ;
  assign n431 = n81 & n241 ;
  assign n99 = n96 & n98 ;
  assign n453 = n431 ^ n99 ;
  assign n450 = n86 & n241 ;
  assign n293 = n69 & n248 ;
  assign n294 = n293 ^ n248 ;
  assign n295 = n294 ^ n292 ;
  assign n296 = n295 ^ n248 ;
  assign n451 = n450 ^ n296 ;
  assign n191 = x23 & n96 ;
  assign n452 = n451 ^ n191 ;
  assign n454 = n453 ^ n452 ;
  assign n460 = n459 ^ n454 ;
  assign n117 = n43 & n89 ;
  assign n116 = n89 & n115 ;
  assign n118 = n117 ^ n116 ;
  assign n109 = n89 & n108 ;
  assign n106 = n89 & n105 ;
  assign n110 = n109 ^ n106 ;
  assign n119 = n118 ^ n110 ;
  assign n12697 = n460 ^ n119 ;
  assign n1355 = x25 & n438 ;
  assign n252 = n136 & n248 ;
  assign n250 = ~n170 & n248 ;
  assign n249 = n78 & n248 ;
  assign n251 = n250 ^ n249 ;
  assign n253 = n252 ^ n251 ;
  assign n12631 = n1355 ^ n253 ;
  assign n351 = n79 & n89 ;
  assign n352 = n1050 ^ n351 ;
  assign n335 = x26 & ~n72 ;
  assign n345 = n89 & n135 ;
  assign n348 = n335 & n345 ;
  assign n337 = ~x27 & ~n35 ;
  assign n336 = n89 ^ n35 ;
  assign n338 = n337 ^ n336 ;
  assign n342 = n341 ^ n338 ;
  assign n343 = n37 & ~n342 ;
  assign n339 = ~n37 & ~n338 ;
  assign n340 = n339 ^ n338 ;
  assign n344 = n343 ^ n340 ;
  assign n346 = n345 ^ n344 ;
  assign n349 = n348 ^ n346 ;
  assign n353 = n352 ^ n349 ;
  assign n12632 = n12631 ^ n353 ;
  assign n358 = n341 ^ n337 ;
  assign n385 = x26 & n358 ;
  assign n386 = n385 ^ n339 ;
  assign n384 = ~n77 & n254 ;
  assign n387 = n386 ^ n384 ;
  assign n380 = n78 & n358 ;
  assign n379 = ~n170 & n358 ;
  assign n381 = n380 ^ n379 ;
  assign n378 = n83 & n254 ;
  assign n382 = n381 ^ n378 ;
  assign n376 = n136 & n358 ;
  assign n375 = ~n80 & n358 ;
  assign n377 = n376 ^ n375 ;
  assign n383 = n382 ^ n377 ;
  assign n388 = n387 ^ n383 ;
  assign n372 = n343 ^ n341 ;
  assign n370 = n84 & n358 ;
  assign n369 = n79 & n358 ;
  assign n371 = n370 ^ n369 ;
  assign n373 = n372 ^ n371 ;
  assign n364 = n105 & n171 ;
  assign n363 = ~n82 & n358 ;
  assign n365 = n364 ^ n363 ;
  assign n362 = n115 & n171 ;
  assign n366 = n365 ^ n362 ;
  assign n360 = ~n128 & n171 ;
  assign n359 = n83 & n358 ;
  assign n361 = n360 ^ n359 ;
  assign n367 = n366 ^ n361 ;
  assign n356 = ~n140 & n171 ;
  assign n355 = n43 & n171 ;
  assign n357 = n356 ^ n355 ;
  assign n368 = n367 ^ n357 ;
  assign n374 = n373 ^ n368 ;
  assign n389 = n388 ^ n374 ;
  assign n12696 = n12632 ^ n389 ;
  assign n12698 = n12697 ^ n12696 ;
  assign n12699 = n12695 & n12698 ;
  assign n499 = n45 & n136 ;
  assign n1789 = n499 ^ n249 ;
  assign n123 = ~n34 & n94 ;
  assign n954 = n43 & n123 ;
  assign n263 = n53 & n262 ;
  assign n261 = n45 & n115 ;
  assign n264 = n263 ^ n261 ;
  assign n1788 = n954 ^ n264 ;
  assign n1790 = n1789 ^ n1788 ;
  assign n102 = n94 ^ x27 ;
  assign n448 = ~n34 & ~n102 ;
  assign n1116 = n448 & ~n12860 ;
  assign n1785 = n1116 ^ n627 ;
  assign n728 = n123 & ~n128 ;
  assign n1205 = n728 ^ n702 ;
  assign n1786 = n1785 ^ n1205 ;
  assign n981 = n86 & n358 ;
  assign n1783 = n981 ^ n375 ;
  assign n210 = n45 & n84 ;
  assign n183 = n78 & n123 ;
  assign n1674 = n210 ^ n183 ;
  assign n1784 = n1783 ^ n1674 ;
  assign n1787 = n1786 ^ n1784 ;
  assign n1791 = n1790 ^ n1787 ;
  assign n103 = ~n95 & ~n102 ;
  assign n506 = n103 & ~n140 ;
  assign n505 = n51 & n84 ;
  assign n507 = n506 ^ n505 ;
  assign n1780 = n507 ^ n244 ;
  assign n745 = n51 & n136 ;
  assign n1781 = n1780 ^ n745 ;
  assign n1775 = ~x23 & n37 ;
  assign n1776 = n448 & n1775 ;
  assign n782 = n79 & n123 ;
  assign n635 = ~n140 & n358 ;
  assign n1774 = n782 ^ n635 ;
  assign n1777 = n1776 ^ n1774 ;
  assign n392 = n48 & n83 ;
  assign n153 = ~n80 & n123 ;
  assign n1772 = n392 ^ n153 ;
  assign n270 = n269 ^ n268 ;
  assign n1773 = n1772 ^ n270 ;
  assign n1778 = n1777 ^ n1773 ;
  assign n87 = n51 & n86 ;
  assign n1233 = n1050 ^ n87 ;
  assign n226 = n83 & n123 ;
  assign n1231 = n226 ^ n110 ;
  assign n1232 = n1231 ^ n456 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1779 = n1778 ^ n1234 ;
  assign n1782 = n1781 ^ n1779 ;
  assign n1792 = n1791 ^ n1782 ;
  assign n848 = n115 & n448 ;
  assign n275 = ~n34 & n50 ;
  assign n483 = n84 & n275 ;
  assign n1224 = n848 ^ n483 ;
  assign n772 = n115 & n123 ;
  assign n255 = n84 & n254 ;
  assign n1153 = n772 ^ n255 ;
  assign n1225 = n1224 ^ n1153 ;
  assign n897 = n45 & n108 ;
  assign n197 = n136 & n171 ;
  assign n1222 = n897 ^ n197 ;
  assign n1223 = n1222 ^ n716 ;
  assign n1226 = n1225 ^ n1223 ;
  assign n1219 = n89 & ~n12860 ;
  assign n1058 = n108 & n123 ;
  assign n1218 = n1058 ^ n292 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n497 = n83 & ~n338 ;
  assign n219 = n86 & n103 ;
  assign n1215 = n497 ^ n219 ;
  assign n778 = ~n41 & ~n338 ;
  assign n779 = n36 & n778 ;
  assign n1216 = n1215 ^ n779 ;
  assign n302 = n69 & n103 ;
  assign n196 = n83 & n103 ;
  assign n303 = n302 ^ n196 ;
  assign n1217 = n1216 ^ n303 ;
  assign n1221 = n1220 ^ n1217 ;
  assign n1227 = n1226 ^ n1221 ;
  assign n1793 = n1792 ^ n1227 ;
  assign n5225 = n394 ^ n351 ;
  assign n391 = n48 & n79 ;
  assign n5224 = n433 ^ n391 ;
  assign n5226 = n5225 ^ n5224 ;
  assign n579 = n43 & n358 ;
  assign n200 = n96 & ~n140 ;
  assign n2899 = n579 ^ n200 ;
  assign n5227 = n5226 ^ n2899 ;
  assign n2987 = n660 ^ n369 ;
  assign n2988 = n2987 ^ n455 ;
  assign n217 = n123 & n136 ;
  assign n4344 = n2988 ^ n217 ;
  assign n12567 = n5227 ^ n4344 ;
  assign n793 = n108 & n448 ;
  assign n521 = n78 & ~n338 ;
  assign n5101 = n793 ^ n521 ;
  assign n12565 = n5101 ^ n176 ;
  assign n597 = ~n170 & ~n338 ;
  assign n12563 = n597 ^ n291 ;
  assign n1494 = n123 & ~n140 ;
  assign n2315 = n1494 ^ n252 ;
  assign n1014 = n79 & n448 ;
  assign n230 = n48 & n115 ;
  assign n2313 = n1014 ^ n230 ;
  assign n161 = n105 & n123 ;
  assign n2314 = n2313 ^ n161 ;
  assign n2316 = n2315 ^ n2314 ;
  assign n12564 = n12563 ^ n2316 ;
  assign n12566 = n12565 ^ n12564 ;
  assign n12568 = n12567 ^ n12566 ;
  assign n762 = ~n338 & ~n12860 ;
  assign n180 = n51 & n108 ;
  assign n4185 = n762 ^ n180 ;
  assign n541 = ~n128 & n358 ;
  assign n495 = n103 & ~n112 ;
  assign n181 = ~n80 & n103 ;
  assign n496 = n495 ^ n181 ;
  assign n2509 = n541 ^ n496 ;
  assign n12559 = n4185 ^ n2509 ;
  assign n542 = n84 & ~n338 ;
  assign n417 = n48 & n136 ;
  assign n5218 = n542 ^ n417 ;
  assign n774 = n108 & ~n338 ;
  assign n742 = n123 & ~n12860 ;
  assign n3603 = n774 ^ n742 ;
  assign n12558 = n5218 ^ n3603 ;
  assign n12560 = n12559 ^ n12558 ;
  assign n272 = ~n170 & n254 ;
  assign n922 = n279 ^ n272 ;
  assign n12555 = n922 ^ n250 ;
  assign n221 = n103 & n105 ;
  assign n12556 = n12555 ^ n221 ;
  assign n726 = n86 & ~n338 ;
  assign n624 = n136 & ~n338 ;
  assign n2592 = n726 ^ n624 ;
  assign n237 = n43 & n51 ;
  assign n12554 = n2592 ^ n237 ;
  assign n12557 = n12556 ^ n12554 ;
  assign n12561 = n12560 ^ n12557 ;
  assign n1982 = n261 ^ n129 ;
  assign n172 = ~n170 & n171 ;
  assign n12551 = n1982 ^ n172 ;
  assign n490 = n115 & n254 ;
  assign n1798 = n490 ^ n186 ;
  assign n6374 = n1798 ^ n118 ;
  assign n12552 = n12551 ^ n6374 ;
  assign n1074 = n45 & ~n140 ;
  assign n414 = n84 & n241 ;
  assign n2035 = n1074 ^ n414 ;
  assign n194 = n84 & n171 ;
  assign n3855 = n2035 ^ n194 ;
  assign n838 = ~n80 & n448 ;
  assign n836 = ~n140 & n448 ;
  assign n124 = n86 & n123 ;
  assign n837 = n836 ^ n124 ;
  assign n839 = n838 ^ n837 ;
  assign n12550 = n3855 ^ n839 ;
  assign n12553 = n12552 ^ n12550 ;
  assign n12562 = n12561 ^ n12553 ;
  assign n12569 = n12568 ^ n12562 ;
  assign n1273 = n298 ^ n216 ;
  assign n1128 = ~n62 & n89 ;
  assign n1129 = n1128 ^ n351 ;
  assign n489 = n51 & ~n170 ;
  assign n1272 = n1129 ^ n489 ;
  assign n1274 = n1273 ^ n1272 ;
  assign n799 = n79 & ~n338 ;
  assign n547 = n358 & ~n12860 ;
  assign n1269 = n799 ^ n547 ;
  assign n760 = n86 & n448 ;
  assign n1270 = n1269 ^ n760 ;
  assign n819 = ~n82 & n123 ;
  assign n614 = n105 & n358 ;
  assign n1266 = n819 ^ n614 ;
  assign n1267 = n1266 ^ n242 ;
  assign n678 = n43 & ~n338 ;
  assign n1268 = n1267 ^ n678 ;
  assign n1271 = n1270 ^ n1268 ;
  assign n1275 = n1274 ^ n1271 ;
  assign n785 = n43 & n45 ;
  assign n1276 = n1275 ^ n785 ;
  assign n12570 = n12569 ^ n1276 ;
  assign n697 = n45 & n105 ;
  assign n222 = n103 & n108 ;
  assign n12547 = n697 ^ n222 ;
  assign n236 = n51 & n105 ;
  assign n12548 = n12547 ^ n236 ;
  assign n285 = n136 & n275 ;
  assign n284 = ~n170 & n275 ;
  assign n286 = n285 ^ n284 ;
  assign n3279 = n703 ^ n286 ;
  assign n557 = ~n112 & n358 ;
  assign n558 = n557 ^ n375 ;
  assign n190 = n43 & n103 ;
  assign n1024 = n558 ^ n190 ;
  assign n12544 = n3279 ^ n1024 ;
  assign n565 = n108 & n358 ;
  assign n225 = n51 & ~n12860 ;
  assign n5595 = n565 ^ n225 ;
  assign n737 = n43 & n448 ;
  assign n3117 = n737 ^ n141 ;
  assign n12542 = n5595 ^ n3117 ;
  assign n814 = ~n82 & ~n338 ;
  assign n12539 = n814 ^ n296 ;
  assign n12540 = n12539 ^ n258 ;
  assign n12541 = n12540 ^ n396 ;
  assign n12543 = n12542 ^ n12541 ;
  assign n12545 = n12544 ^ n12543 ;
  assign n413 = n103 & ~n128 ;
  assign n1149 = n1148 ^ n413 ;
  assign n4273 = n1149 ^ n612 ;
  assign n526 = ~n82 & n448 ;
  assign n4274 = n4273 ^ n526 ;
  assign n12546 = n12545 ^ n4274 ;
  assign n12549 = n12548 ^ n12546 ;
  assign n12571 = n12570 ^ n12549 ;
  assign n12572 = ~n1793 & ~n12571 ;
  assign n12686 = n12572 ^ x29 ;
  assign n238 = n237 ^ n236 ;
  assign n12633 = n12632 ^ n238 ;
  assign n276 = n76 & n275 ;
  assign n277 = n276 ^ n123 ;
  assign n12638 = n496 ^ n277 ;
  assign n12634 = ~n12860 ^ n36 ;
  assign n12635 = n248 & n12634 ;
  assign n510 = n55 & n254 ;
  assign n12636 = n12635 ^ n510 ;
  assign n12637 = n12636 ^ n506 ;
  assign n12639 = n12638 ^ n12637 ;
  assign n682 = n51 & n83 ;
  assign n265 = n103 & ~n170 ;
  assign n1961 = n682 ^ n265 ;
  assign n12640 = n1961 ^ n427 ;
  assign n297 = n296 ^ n291 ;
  assign n299 = n298 ^ n297 ;
  assign n12641 = n12640 ^ n299 ;
  assign n12642 = n12641 ^ n372 ;
  assign n12643 = ~n12639 & ~n12642 ;
  assign n12644 = n12633 & n12643 ;
  assign n478 = n51 & ~n82 ;
  assign n1605 = n478 ^ n413 ;
  assign n6422 = n1605 ^ n499 ;
  assign n871 = n51 & n78 ;
  assign n5257 = n871 ^ n414 ;
  assign n12645 = n6422 ^ n5257 ;
  assign n1085 = x23 & n228 ;
  assign n229 = n1085 ^ n228 ;
  assign n231 = n230 ^ n229 ;
  assign n227 = n226 ^ n225 ;
  assign n232 = n231 ^ n227 ;
  assign n223 = n222 ^ n221 ;
  assign n218 = n217 ^ n216 ;
  assign n220 = n219 ^ n218 ;
  assign n224 = n223 ^ n220 ;
  assign n233 = n232 ^ n224 ;
  assign n97 = n96 & ~n12860 ;
  assign n211 = n210 ^ n97 ;
  assign n213 = n212 ^ n211 ;
  assign n214 = n213 ^ n204 ;
  assign n207 = n206 ^ n203 ;
  assign n201 = n51 & n79 ;
  assign n202 = n201 ^ n200 ;
  assign n208 = n207 ^ n202 ;
  assign n198 = n197 ^ n196 ;
  assign n192 = ~n62 & n191 ;
  assign n193 = n192 ^ n190 ;
  assign n195 = n194 ^ n193 ;
  assign n199 = n198 ^ n195 ;
  assign n209 = n208 ^ n199 ;
  assign n215 = n214 ^ n209 ;
  assign n234 = n233 ^ n215 ;
  assign n155 = n48 & n84 ;
  assign n154 = n48 & n73 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n156 ^ n153 ;
  assign n151 = n51 & ~n80 ;
  assign n149 = n48 & n105 ;
  assign n148 = n103 & ~n12860 ;
  assign n150 = n149 ^ n148 ;
  assign n152 = n151 ^ n150 ;
  assign n158 = n157 ^ n152 ;
  assign n144 = ~n82 & n96 ;
  assign n143 = n86 & n96 ;
  assign n145 = n144 ^ n143 ;
  assign n137 = n103 & n136 ;
  assign n142 = n141 ^ n137 ;
  assign n146 = n145 ^ n142 ;
  assign n131 = n130 ^ n129 ;
  assign n125 = n124 ^ n122 ;
  assign n132 = n131 ^ n125 ;
  assign n147 = n146 ^ n132 ;
  assign n159 = n158 ^ n147 ;
  assign n104 = n78 & n103 ;
  assign n120 = n119 ^ n104 ;
  assign n100 = n99 ^ n97 ;
  assign n88 = n48 & n86 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = n1085 ^ n92 ;
  assign n101 = n100 ^ n93 ;
  assign n121 = n120 ^ n101 ;
  assign n160 = n159 ^ n121 ;
  assign n182 = n181 ^ n180 ;
  assign n184 = n183 ^ n182 ;
  assign n178 = ~n82 & n103 ;
  assign n175 = n79 & n103 ;
  assign n177 = n176 ^ n175 ;
  assign n179 = n178 ^ n177 ;
  assign n185 = n184 ^ n179 ;
  assign n187 = n186 ^ n185 ;
  assign n162 = n60 ^ x24 ;
  assign n163 = ~n12860 ^ n162 ;
  assign n164 = n163 ^ x26 ;
  assign n165 = n139 ^ n53 ;
  assign n166 = n123 & ~n165 ;
  assign n167 = n164 & n166 ;
  assign n168 = n167 ^ n123 ;
  assign n173 = n172 ^ n168 ;
  assign n174 = n173 ^ n161 ;
  assign n188 = n187 ^ n174 ;
  assign n189 = ~n160 & ~n188 ;
  assign n235 = n234 ^ n189 ;
  assign n12646 = n12645 ^ n235 ;
  assign n12647 = n12644 & n12646 ;
  assign n12687 = n12647 ^ n12572 ;
  assign n12688 = n12686 & ~n12687 ;
  assign n12689 = n12688 ^ x29 ;
  assign n12700 = n12699 ^ n12689 ;
  assign n3520 = x30 ^ x29 ;
  assign n326 = n285 ^ n183 ;
  assign n280 = n79 & n171 ;
  assign n282 = n281 ^ n280 ;
  assign n325 = n282 ^ n217 ;
  assign n327 = n326 ^ n325 ;
  assign n328 = ~n277 & ~n327 ;
  assign n323 = n322 ^ n197 ;
  assign n310 = n309 ^ n280 ;
  assign n311 = n310 ^ n308 ;
  assign n320 = n311 ^ n259 ;
  assign n324 = n323 ^ n320 ;
  assign n329 = n328 ^ n324 ;
  assign n330 = n284 ^ n194 ;
  assign n331 = n330 ^ n124 ;
  assign n332 = n331 ^ n226 ;
  assign n333 = n332 ^ n173 ;
  assign n334 = n329 & ~n333 ;
  assign n354 = n353 ^ n334 ;
  assign n390 = n389 ^ n354 ;
  assign n440 = n62 ^ n42 ;
  assign n441 = n51 & ~n440 ;
  assign n442 = n1355 ^ n441 ;
  assign n435 = n127 ^ n79 ;
  assign n436 = n241 & ~n435 ;
  assign n430 = n429 ^ n427 ;
  assign n432 = n431 ^ n430 ;
  assign n434 = n433 ^ n432 ;
  assign n437 = n436 ^ n434 ;
  assign n443 = n442 ^ n437 ;
  assign n397 = n396 ^ n222 ;
  assign n393 = n392 ^ n391 ;
  assign n395 = n394 ^ n393 ;
  assign n398 = n397 ^ n395 ;
  assign n399 = n263 ^ n103 ;
  assign n418 = n417 ^ n416 ;
  assign n401 = n78 & n241 ;
  assign n419 = n418 ^ n401 ;
  assign n415 = n414 ^ n413 ;
  assign n420 = n419 ^ n415 ;
  assign n410 = n409 ^ n155 ;
  assign n411 = n410 ^ n408 ;
  assign n403 = n402 ^ n401 ;
  assign n404 = n403 ^ n400 ;
  assign n412 = n411 ^ n404 ;
  assign n421 = n420 ^ n412 ;
  assign n422 = ~n399 & ~n421 ;
  assign n423 = ~n398 & n422 ;
  assign n240 = n239 ^ n238 ;
  assign n424 = n423 ^ n240 ;
  assign n444 = n443 ^ n424 ;
  assign n445 = ~n390 & n444 ;
  assign n313 = ~n140 & n254 ;
  assign n312 = n311 ^ n261 ;
  assign n314 = n313 ^ n312 ;
  assign n304 = n47 & n105 ;
  assign n305 = n304 ^ n236 ;
  assign n306 = n305 ^ n303 ;
  assign n300 = n107 & n254 ;
  assign n301 = n300 ^ n299 ;
  assign n307 = n306 ^ n301 ;
  assign n315 = n314 ^ n307 ;
  assign n283 = n282 ^ n279 ;
  assign n287 = n286 ^ n283 ;
  assign n273 = ~n128 & n254 ;
  assign n274 = n273 ^ n272 ;
  assign n278 = n277 ^ n274 ;
  assign n288 = n287 ^ n278 ;
  assign n266 = n265 ^ n264 ;
  assign n267 = n266 ^ n260 ;
  assign n271 = n270 ^ n267 ;
  assign n289 = n288 ^ n271 ;
  assign n256 = n255 ^ n253 ;
  assign n246 = n245 ^ n244 ;
  assign n243 = n242 ^ n240 ;
  assign n247 = n246 ^ n243 ;
  assign n257 = n256 ^ n247 ;
  assign n290 = n289 ^ n257 ;
  assign n316 = n315 ^ n290 ;
  assign n317 = n235 & ~n316 ;
  assign n525 = n169 & n448 ;
  assign n527 = n526 ^ n525 ;
  assign n528 = n527 ^ n130 ;
  assign n529 = n528 ^ n207 ;
  assign n520 = n45 & n79 ;
  assign n522 = n521 ^ n520 ;
  assign n523 = n522 ^ n97 ;
  assign n518 = n45 & ~n82 ;
  assign n519 = n518 ^ n144 ;
  assign n524 = n523 ^ n519 ;
  assign n530 = n529 ^ n524 ;
  assign n531 = n530 ^ n421 ;
  assign n513 = n45 & n83 ;
  assign n512 = n45 & n78 ;
  assign n514 = n513 ^ n512 ;
  assign n508 = ~n57 & n254 ;
  assign n509 = n508 ^ n384 ;
  assign n511 = n510 ^ n509 ;
  assign n515 = n514 ^ n511 ;
  assign n516 = n515 ^ n507 ;
  assign n500 = n45 & ~n80 ;
  assign n501 = n500 ^ n499 ;
  assign n502 = n501 ^ n192 ;
  assign n498 = n497 ^ n496 ;
  assign n503 = n502 ^ n498 ;
  assign n491 = n490 ^ n378 ;
  assign n492 = n491 ^ n489 ;
  assign n493 = n492 ^ n321 ;
  assign n494 = n493 ^ n286 ;
  assign n504 = n503 ^ n494 ;
  assign n517 = n516 ^ n504 ;
  assign n532 = n531 ^ n517 ;
  assign n642 = n123 & ~n170 ;
  assign n641 = n115 & n275 ;
  assign n643 = n642 ^ n641 ;
  assign n644 = n643 ^ n149 ;
  assign n645 = n644 ^ n302 ;
  assign n636 = ~n128 & n275 ;
  assign n637 = n636 ^ n355 ;
  assign n638 = n637 ^ n379 ;
  assign n639 = n638 ^ n635 ;
  assign n632 = n380 ^ n363 ;
  assign n633 = n632 ^ n156 ;
  assign n628 = n627 ^ n292 ;
  assign n625 = n43 & n275 ;
  assign n629 = n628 ^ n625 ;
  assign n630 = n629 ^ n624 ;
  assign n622 = n105 & n248 ;
  assign n621 = ~n128 & n248 ;
  assign n623 = n622 ^ n621 ;
  assign n631 = n630 ^ n623 ;
  assign n634 = n633 ^ n631 ;
  assign n640 = n639 ^ n634 ;
  assign n646 = n645 ^ n640 ;
  assign n613 = n79 & n275 ;
  assign n615 = n614 ^ n613 ;
  assign n616 = n615 ^ n212 ;
  assign n617 = n616 ^ n268 ;
  assign n618 = n617 ^ n279 ;
  assign n619 = n618 ^ n612 ;
  assign n667 = x23 & n300 ;
  assign n607 = n667 ^ n300 ;
  assign n608 = n607 ^ n137 ;
  assign n609 = n608 ^ n244 ;
  assign n610 = n609 ^ n110 ;
  assign n602 = n275 & ~n12860 ;
  assign n603 = n602 ^ n261 ;
  assign n604 = n603 ^ n201 ;
  assign n600 = n981 ^ n356 ;
  assign n601 = n600 ^ n597 ;
  assign n605 = n604 ^ n601 ;
  assign n611 = n610 ^ n605 ;
  assign n620 = n619 ^ n611 ;
  assign n647 = n646 ^ n620 ;
  assign n592 = ~n140 & n248 ;
  assign n593 = n592 ^ n151 ;
  assign n590 = n217 ^ n117 ;
  assign n589 = n105 & n275 ;
  assign n591 = n590 ^ n589 ;
  assign n594 = n593 ^ n591 ;
  assign n584 = n115 & n248 ;
  assign n583 = n108 & n275 ;
  assign n585 = n584 ^ n583 ;
  assign n586 = n585 ^ n104 ;
  assign n587 = n586 ^ n377 ;
  assign n580 = n579 ^ n116 ;
  assign n578 = n359 ^ n225 ;
  assign n581 = n580 ^ n578 ;
  assign n577 = n108 & n248 ;
  assign n582 = n581 ^ n577 ;
  assign n588 = n587 ^ n582 ;
  assign n595 = n594 ^ n588 ;
  assign n571 = n78 & n275 ;
  assign n572 = n571 ^ n360 ;
  assign n570 = ~n140 & n275 ;
  assign n573 = n572 ^ n570 ;
  assign n567 = n83 & n275 ;
  assign n568 = n567 ^ n141 ;
  assign n566 = n565 ^ n298 ;
  assign n569 = n568 ^ n566 ;
  assign n574 = n573 ^ n569 ;
  assign n560 = n84 & n448 ;
  assign n559 = n84 & n123 ;
  assign n561 = n560 ^ n559 ;
  assign n562 = n561 ^ n364 ;
  assign n563 = n562 ^ n558 ;
  assign n554 = n370 ^ n269 ;
  assign n555 = n554 ^ n362 ;
  assign n556 = n555 ^ n258 ;
  assign n564 = n563 ^ n556 ;
  assign n575 = n574 ^ n564 ;
  assign n550 = n111 & n549 ;
  assign n551 = n550 ^ n228 ;
  assign n548 = n547 ^ n266 ;
  assign n552 = n551 ^ n548 ;
  assign n543 = n542 ^ n369 ;
  assign n544 = n543 ^ n541 ;
  assign n540 = n86 & n275 ;
  assign n545 = n544 ^ n540 ;
  assign n841 = ~n74 & n549 ;
  assign n537 = n841 ^ n242 ;
  assign n535 = n81 & n275 ;
  assign n538 = n537 ^ n535 ;
  assign n534 = n533 ^ n92 ;
  assign n539 = n538 ^ n534 ;
  assign n546 = n545 ^ n539 ;
  assign n553 = n552 ^ n546 ;
  assign n576 = n575 ^ n553 ;
  assign n596 = n595 ^ n576 ;
  assign n648 = n647 ^ n596 ;
  assign n649 = ~n532 & ~n648 ;
  assign n2948 = n394 ^ n178 ;
  assign n3418 = n2948 ^ n577 ;
  assign n3415 = n495 ^ n204 ;
  assign n739 = n45 & n86 ;
  assign n3416 = n3415 ^ n739 ;
  assign n912 = n200 ^ n186 ;
  assign n3417 = n3416 ^ n912 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n1249 = ~n82 & n341 ;
  assign n467 = x26 ^ x25 ;
  assign n1098 = n467 & n778 ;
  assign n1097 = n778 ^ n521 ;
  assign n1099 = n1098 ^ n1097 ;
  assign n1250 = n1249 ^ n1099 ;
  assign n3412 = n1273 ^ n1250 ;
  assign n2745 = n122 ^ n106 ;
  assign n3413 = n3412 ^ n2745 ;
  assign n3408 = n819 ^ n244 ;
  assign n3409 = n3408 ^ n226 ;
  assign n1093 = ~n170 & n341 ;
  assign n3410 = n3409 ^ n1093 ;
  assign n1122 = n83 & n341 ;
  assign n673 = n45 & ~n12860 ;
  assign n1359 = n1122 ^ n673 ;
  assign n3406 = n1359 ^ n183 ;
  assign n1130 = n78 & n254 ;
  assign n3407 = n3406 ^ n1130 ;
  assign n3411 = n3410 ^ n3407 ;
  assign n3414 = n3413 ^ n3411 ;
  assign n3420 = n3419 ^ n3414 ;
  assign n3401 = n897 ^ n415 ;
  assign n3402 = n3401 ^ n268 ;
  assign n3403 = n3402 ^ n667 ;
  assign n3398 = n286 ^ n212 ;
  assign n797 = ~n133 & n384 ;
  assign n3399 = n3398 ^ n797 ;
  assign n3397 = n745 ^ n537 ;
  assign n3400 = n3399 ^ n3397 ;
  assign n3404 = n3403 ^ n3400 ;
  assign n1088 = n84 & n341 ;
  assign n3321 = n1088 ^ n258 ;
  assign n867 = n78 & n341 ;
  assign n1311 = n867 ^ n180 ;
  assign n3394 = n3321 ^ n1311 ;
  assign n2888 = n279 ^ n100 ;
  assign n1480 = n175 ^ n141 ;
  assign n3393 = n2888 ^ n1480 ;
  assign n3395 = n3394 ^ n3393 ;
  assign n952 = n136 & n341 ;
  assign n3390 = n952 ^ n392 ;
  assign n3391 = n3390 ^ n118 ;
  assign n1236 = n871 ^ n321 ;
  assign n1188 = n305 ^ n237 ;
  assign n3389 = n1236 ^ n1188 ;
  assign n3392 = n3391 ^ n3389 ;
  assign n3396 = n3395 ^ n3392 ;
  assign n3405 = n3404 ^ n3396 ;
  assign n3421 = n3420 ^ n3405 ;
  assign n804 = n136 & n448 ;
  assign n1658 = n804 ^ n499 ;
  assign n1659 = n1658 ^ n201 ;
  assign n1176 = n838 ^ n567 ;
  assign n1602 = n1176 ^ n954 ;
  assign n3469 = n1659 ^ n1602 ;
  assign n880 = ~n62 & n275 ;
  assign n881 = n880 ^ n613 ;
  assign n1728 = n881 ^ n513 ;
  assign n1015 = n1014 ^ n762 ;
  assign n3466 = n1728 ^ n1015 ;
  assign n3464 = n774 ^ n370 ;
  assign n3465 = n3464 ^ n1785 ;
  assign n3467 = n3466 ^ n3465 ;
  assign n3468 = n3467 ^ n367 ;
  assign n3470 = n3469 ^ n3468 ;
  assign n1069 = n814 ^ n109 ;
  assign n3459 = n1069 ^ n431 ;
  assign n3460 = n3459 ^ n410 ;
  assign n3458 = n726 ^ n266 ;
  assign n3461 = n3460 ^ n3458 ;
  assign n3456 = n1148 ^ n303 ;
  assign n743 = n571 ^ n153 ;
  assign n3455 = n743 ^ n91 ;
  assign n3457 = n3456 ^ n3455 ;
  assign n3462 = n3461 ^ n3457 ;
  assign n1181 = n433 ^ n379 ;
  assign n3453 = n1181 ^ n613 ;
  assign n882 = n881 ^ n535 ;
  assign n1495 = n1494 ^ n882 ;
  assign n3451 = n1495 ^ n1029 ;
  assign n773 = n105 & ~n338 ;
  assign n3448 = n773 ^ n161 ;
  assign n3449 = n3448 ^ n429 ;
  assign n3450 = n3449 ^ n490 ;
  assign n3452 = n3451 ^ n3450 ;
  assign n3454 = n3453 ^ n3452 ;
  assign n3463 = n3462 ^ n3454 ;
  assign n3471 = n3470 ^ n3463 ;
  assign n3444 = n678 ^ n612 ;
  assign n1756 = n661 ^ n405 ;
  assign n3445 = n3444 ^ n1756 ;
  assign n3442 = n782 ^ n512 ;
  assign n932 = ~n128 & ~n338 ;
  assign n3440 = n932 ^ n540 ;
  assign n3441 = n3440 ^ n269 ;
  assign n3443 = n3442 ^ n3441 ;
  assign n3446 = n3445 ^ n3443 ;
  assign n677 = n83 & n448 ;
  assign n1759 = n677 ^ n151 ;
  assign n3436 = n1759 ^ n602 ;
  assign n3437 = n3436 ^ n507 ;
  assign n3433 = n292 ^ n148 ;
  assign n3432 = n1058 ^ n143 ;
  assign n3434 = n3433 ^ n3432 ;
  assign n3431 = n450 ^ n380 ;
  assign n3435 = n3434 ^ n3431 ;
  assign n3438 = n3437 ^ n3435 ;
  assign n3428 = n742 ^ n357 ;
  assign n945 = ~n140 & ~n338 ;
  assign n1150 = n945 ^ n156 ;
  assign n3427 = n1150 ^ n261 ;
  assign n3429 = n3428 ^ n3427 ;
  assign n1060 = n779 ^ n526 ;
  assign n3425 = n1060 ^ n255 ;
  assign n725 = n78 & n448 ;
  assign n3423 = n725 ^ n376 ;
  assign n1802 = n799 ^ n124 ;
  assign n3422 = n1802 ^ n703 ;
  assign n3424 = n3423 ^ n3422 ;
  assign n3426 = n3425 ^ n3424 ;
  assign n3430 = n3429 ^ n3426 ;
  assign n3439 = n3438 ^ n3430 ;
  assign n3447 = n3446 ^ n3439 ;
  assign n3472 = n3471 ^ n3447 ;
  assign n3473 = ~n3421 & ~n3472 ;
  assign n899 = n725 ^ n401 ;
  assign n898 = n897 ^ n117 ;
  assign n900 = n899 ^ n898 ;
  assign n901 = n900 ^ n196 ;
  assign n893 = n89 & ~n170 ;
  assign n894 = n893 ^ n192 ;
  assign n895 = n894 ^ n782 ;
  assign n896 = n895 ^ n391 ;
  assign n902 = n901 ^ n896 ;
  assign n890 = n565 ^ n394 ;
  assign n764 = ~n80 & n241 ;
  assign n888 = n1050 ^ n764 ;
  assign n889 = n888 ^ n745 ;
  assign n891 = n890 ^ n889 ;
  assign n885 = n351 ^ n183 ;
  assign n886 = n885 ^ n426 ;
  assign n883 = n882 ^ n785 ;
  assign n878 = n500 ^ n176 ;
  assign n877 = n760 ^ n642 ;
  assign n879 = n878 ^ n877 ;
  assign n884 = n883 ^ n879 ;
  assign n887 = n886 ^ n884 ;
  assign n892 = n891 ^ n887 ;
  assign n903 = n902 ^ n892 ;
  assign n872 = n871 ^ n230 ;
  assign n873 = n872 ^ n250 ;
  assign n868 = n867 ^ n226 ;
  assign n869 = n868 ^ n321 ;
  assign n865 = n298 ^ n239 ;
  assign n866 = n865 ^ n203 ;
  assign n870 = n869 ^ n866 ;
  assign n874 = n873 ^ n870 ;
  assign n863 = n804 ^ n181 ;
  assign n862 = n774 ^ n641 ;
  assign n864 = n863 ^ n862 ;
  assign n875 = n874 ^ n864 ;
  assign n856 = ~n82 & n89 ;
  assign n857 = n856 ^ n489 ;
  assign n858 = n857 ^ n175 ;
  assign n853 = n206 ^ n122 ;
  assign n854 = n853 ^ n541 ;
  assign n765 = n764 ^ n431 ;
  assign n855 = n854 ^ n765 ;
  assign n859 = n858 ^ n855 ;
  assign n850 = n737 ^ n282 ;
  assign n849 = n848 ^ n261 ;
  assign n851 = n850 ^ n849 ;
  assign n845 = n84 & n89 ;
  assign n846 = n845 ^ n264 ;
  assign n844 = n799 ^ n728 ;
  assign n847 = n846 ^ n844 ;
  assign n852 = n851 ^ n847 ;
  assign n860 = n859 ^ n852 ;
  assign n842 = n841 ^ n456 ;
  assign n835 = n624 ^ n579 ;
  assign n840 = n839 ^ n835 ;
  assign n843 = n842 ^ n840 ;
  assign n861 = n860 ^ n843 ;
  assign n876 = n875 ^ n861 ;
  assign n904 = n903 ^ n876 ;
  assign n818 = n375 ^ n356 ;
  assign n964 = n818 ^ n242 ;
  assign n961 = n550 ^ n513 ;
  assign n962 = n961 ^ n526 ;
  assign n959 = n589 ^ n455 ;
  assign n960 = n959 ^ n400 ;
  assign n963 = n962 ^ n960 ;
  assign n965 = n964 ^ n963 ;
  assign n955 = n954 ^ n417 ;
  assign n953 = n952 ^ n259 ;
  assign n956 = n955 ^ n953 ;
  assign n950 = n814 ^ n571 ;
  assign n949 = n661 ^ n129 ;
  assign n951 = n950 ^ n949 ;
  assign n957 = n956 ^ n951 ;
  assign n946 = n945 ^ n90 ;
  assign n947 = n946 ^ n623 ;
  assign n747 = ~n80 & n341 ;
  assign n748 = n747 ^ n116 ;
  assign n948 = n947 ^ n748 ;
  assign n958 = n957 ^ n948 ;
  assign n966 = n965 ^ n958 ;
  assign n940 = n378 ^ n273 ;
  assign n941 = n940 ^ n178 ;
  assign n810 = n79 & n341 ;
  assign n937 = n810 ^ n380 ;
  assign n938 = n937 ^ n405 ;
  assign n939 = n938 ^ n403 ;
  assign n942 = n941 ^ n939 ;
  assign n935 = n520 ^ n280 ;
  assign n672 = n43 & n341 ;
  assign n933 = n932 ^ n672 ;
  assign n931 = n371 ^ n172 ;
  assign n934 = n933 ^ n931 ;
  assign n936 = n935 ^ n934 ;
  assign n943 = n942 ^ n936 ;
  assign n927 = n1085 ^ n597 ;
  assign n926 = n612 ^ n148 ;
  assign n928 = n927 ^ n926 ;
  assign n923 = n922 ^ n244 ;
  assign n924 = n923 ^ n409 ;
  assign n920 = n284 ^ n255 ;
  assign n918 = n83 & n89 ;
  assign n919 = n918 ^ n726 ;
  assign n921 = n920 ^ n919 ;
  assign n925 = n924 ^ n921 ;
  assign n929 = n928 ^ n925 ;
  assign n914 = ~n41 & ~n344 ;
  assign n915 = n914 ^ n667 ;
  assign n911 = n249 ^ n109 ;
  assign n913 = n912 ^ n911 ;
  assign n916 = n915 ^ n913 ;
  assign n909 = n583 ^ n293 ;
  assign n906 = n560 ^ n161 ;
  assign n907 = n906 ^ n88 ;
  assign n905 = n602 ^ n359 ;
  assign n908 = n907 ^ n905 ;
  assign n910 = n909 ^ n908 ;
  assign n917 = n916 ^ n910 ;
  assign n930 = n929 ^ n917 ;
  assign n944 = n943 ^ n930 ;
  assign n967 = n966 ^ n944 ;
  assign n968 = ~n904 & ~n967 ;
  assign n698 = n697 ^ n360 ;
  assign n699 = n698 ^ n231 ;
  assign n693 = n284 ^ n144 ;
  assign n694 = n693 ^ n625 ;
  assign n695 = n694 ^ n210 ;
  assign n690 = n369 ^ n264 ;
  assign n691 = n690 ^ n236 ;
  assign n689 = ~n140 & n341 ;
  assign n692 = n691 ^ n689 ;
  assign n696 = n695 ^ n692 ;
  assign n700 = n699 ^ n696 ;
  assign n683 = n682 ^ n490 ;
  assign n684 = n683 ^ n183 ;
  assign n685 = n684 ^ n570 ;
  assign n681 = n622 ^ n197 ;
  assign n686 = n685 ^ n681 ;
  assign n679 = n678 ^ n677 ;
  assign n675 = n518 ^ n109 ;
  assign n674 = n673 ^ n672 ;
  assign n676 = n675 ^ n674 ;
  assign n680 = n679 ^ n676 ;
  assign n687 = n686 ^ n680 ;
  assign n668 = n667 ^ n285 ;
  assign n669 = n668 ^ n222 ;
  assign n666 = n589 ^ n565 ;
  assign n670 = n669 ^ n666 ;
  assign n663 = n547 ^ n396 ;
  assign n664 = n663 ^ n662 ;
  assign n658 = n614 ^ n355 ;
  assign n659 = n658 ^ n499 ;
  assign n665 = n664 ^ n659 ;
  assign n671 = n670 ^ n665 ;
  assign n688 = n687 ^ n671 ;
  assign n701 = n700 ^ n688 ;
  assign n724 = n723 ^ n701 ;
  assign n820 = n819 ^ n818 ;
  assign n815 = n814 ^ n204 ;
  assign n816 = n815 ^ n258 ;
  assign n811 = n810 ^ n506 ;
  assign n812 = n811 ^ n117 ;
  assign n809 = n105 & n448 ;
  assign n813 = n812 ^ n809 ;
  assign n817 = n816 ^ n813 ;
  assign n821 = n820 ^ n817 ;
  assign n805 = n804 ^ n313 ;
  assign n806 = n805 ^ n137 ;
  assign n803 = n156 ^ n143 ;
  assign n807 = n806 ^ n803 ;
  assign n798 = n797 ^ n394 ;
  assign n800 = n799 ^ n798 ;
  assign n796 = n362 ^ n201 ;
  assign n801 = n800 ^ n796 ;
  assign n794 = n793 ^ n122 ;
  assign n790 = n341 & ~n12860 ;
  assign n791 = n790 ^ n635 ;
  assign n792 = n791 ^ n227 ;
  assign n795 = n794 ^ n792 ;
  assign n802 = n801 ^ n795 ;
  assign n808 = n807 ^ n802 ;
  assign n822 = n821 ^ n808 ;
  assign n786 = n785 ^ n403 ;
  assign n787 = n981 ^ n786 ;
  assign n783 = n782 ^ n106 ;
  assign n780 = n779 ^ n550 ;
  assign n775 = n774 ^ n773 ;
  assign n776 = n775 ^ n772 ;
  assign n777 = n776 ^ n579 ;
  assign n781 = n780 ^ n777 ;
  assign n784 = n783 ^ n781 ;
  assign n788 = n787 ^ n784 ;
  assign n768 = n86 & n341 ;
  assign n769 = n768 ^ n512 ;
  assign n761 = n760 ^ n583 ;
  assign n763 = n762 ^ n761 ;
  assign n766 = n765 ^ n763 ;
  assign n759 = n567 ^ n413 ;
  assign n767 = n766 ^ n759 ;
  assign n770 = n769 ^ n767 ;
  assign n753 = n592 ^ n261 ;
  assign n754 = n753 ^ n172 ;
  assign n755 = n754 ^ n178 ;
  assign n751 = n194 ^ n104 ;
  assign n752 = n751 ^ n219 ;
  assign n756 = n755 ^ n752 ;
  assign n749 = n748 ^ n180 ;
  assign n744 = n743 ^ n742 ;
  assign n746 = n745 ^ n744 ;
  assign n750 = n749 ^ n746 ;
  assign n757 = n756 ^ n750 ;
  assign n736 = n636 ^ n364 ;
  assign n738 = n737 ^ n736 ;
  assign n740 = n739 ^ n738 ;
  assign n732 = n108 & n341 ;
  assign n733 = n732 ^ n607 ;
  assign n731 = n296 ^ n268 ;
  assign n734 = n733 ^ n731 ;
  assign n729 = n728 ^ n175 ;
  assign n727 = n726 ^ n725 ;
  assign n730 = n729 ^ n727 ;
  assign n735 = n734 ^ n730 ;
  assign n741 = n740 ^ n735 ;
  assign n758 = n757 ^ n741 ;
  assign n771 = n770 ^ n758 ;
  assign n789 = n788 ^ n771 ;
  assign n823 = n822 ^ n789 ;
  assign n824 = ~n724 & ~n823 ;
  assign n969 = n968 ^ n824 ;
  assign n1044 = n321 ^ n272 ;
  assign n1043 = n932 ^ n799 ;
  assign n1045 = n1044 ^ n1043 ;
  assign n1041 = n836 ^ n584 ;
  assign n1042 = n1041 ^ n682 ;
  assign n1046 = n1045 ^ n1042 ;
  assign n1038 = n881 ^ n499 ;
  assign n1039 = n1038 ^ n180 ;
  assign n1036 = n845 ^ n151 ;
  assign n1037 = n1036 ^ n129 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n1047 = n1046 ^ n1040 ;
  assign n1032 = n613 ^ n269 ;
  assign n1033 = n1032 ^ n506 ;
  assign n1028 = n303 ^ n225 ;
  assign n1031 = n1030 ^ n1028 ;
  assign n1034 = n1033 ^ n1031 ;
  assign n1023 = n401 ^ n117 ;
  assign n1025 = n1024 ^ n1023 ;
  assign n1021 = n183 ^ n141 ;
  assign n1020 = n518 ^ n489 ;
  assign n1022 = n1021 ^ n1020 ;
  assign n1026 = n1025 ^ n1022 ;
  assign n1017 = n370 ^ n242 ;
  assign n1018 = n1017 ^ n621 ;
  assign n1012 = n810 ^ n673 ;
  assign n1013 = n1012 ^ n143 ;
  assign n1016 = n1015 ^ n1013 ;
  assign n1019 = n1018 ^ n1016 ;
  assign n1027 = n1026 ^ n1019 ;
  assign n1035 = n1034 ^ n1027 ;
  assign n1048 = n1047 ^ n1035 ;
  assign n1008 = n409 ^ n378 ;
  assign n1007 = n804 ^ n768 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1004 = n541 ^ n355 ;
  assign n1005 = n1004 ^ n790 ;
  assign n1001 = n89 & n136 ;
  assign n1002 = n1001 ^ n456 ;
  assign n999 = n264 ^ n238 ;
  assign n1000 = n999 ^ n106 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n1006 = n1005 ^ n1003 ;
  assign n1010 = n1009 ^ n1006 ;
  assign n994 = n625 ^ n313 ;
  assign n995 = n994 ^ n291 ;
  assign n996 = n995 ^ n732 ;
  assign n990 = n559 ^ n258 ;
  assign n991 = n990 ^ n478 ;
  assign n992 = n1148 ^ n991 ;
  assign n993 = n992 ^ n239 ;
  assign n997 = n996 ^ n993 ;
  assign n987 = n785 ^ n667 ;
  assign n983 = n772 ^ n376 ;
  assign n984 = n983 ^ n130 ;
  assign n985 = n984 ^ n819 ;
  assign n982 = n981 ^ n203 ;
  assign n986 = n985 ^ n982 ;
  assign n988 = n987 ^ n986 ;
  assign n978 = n550 ^ n308 ;
  assign n976 = n745 ^ n137 ;
  assign n977 = n976 ^ n405 ;
  assign n979 = n978 ^ n977 ;
  assign n973 = n728 ^ n369 ;
  assign n971 = n78 & n89 ;
  assign n972 = n971 ^ n364 ;
  assign n974 = n973 ^ n972 ;
  assign n970 = n914 ^ n285 ;
  assign n975 = n974 ^ n970 ;
  assign n980 = n979 ^ n975 ;
  assign n989 = n988 ^ n980 ;
  assign n998 = n997 ^ n989 ;
  assign n1011 = n1010 ^ n998 ;
  assign n1049 = n1048 ^ n1011 ;
  assign n1104 = n226 ^ n178 ;
  assign n1105 = n1104 ^ n330 ;
  assign n1106 = n1105 ^ n628 ;
  assign n1100 = n1099 ^ n583 ;
  assign n1101 = n1100 ^ n229 ;
  assign n1102 = n1101 ^ n893 ;
  assign n1094 = n1093 ^ n87 ;
  assign n1095 = n1094 ^ n429 ;
  assign n1096 = n1095 ^ n305 ;
  assign n1103 = n1102 ^ n1096 ;
  assign n1107 = n1106 ^ n1103 ;
  assign n1086 = n1085 ^ n747 ;
  assign n1087 = n1086 ^ n201 ;
  assign n1089 = n1088 ^ n1087 ;
  assign n1090 = n1089 ^ n873 ;
  assign n1081 = n765 ^ n206 ;
  assign n1082 = n1081 ^ n641 ;
  assign n1078 = n416 ^ n216 ;
  assign n1079 = n1078 ^ n219 ;
  assign n1080 = n1079 ^ n520 ;
  assign n1083 = n1082 ^ n1080 ;
  assign n1076 = n393 ^ n379 ;
  assign n1075 = n1074 ^ n946 ;
  assign n1077 = n1076 ^ n1075 ;
  assign n1084 = n1083 ^ n1077 ;
  assign n1091 = n1090 ^ n1084 ;
  assign n1070 = n1069 ^ n702 ;
  assign n1068 = n495 ^ n212 ;
  assign n1071 = n1070 ^ n1068 ;
  assign n1066 = n882 ^ n542 ;
  assign n1064 = n760 ^ n259 ;
  assign n1065 = n1064 ^ n793 ;
  assign n1067 = n1066 ^ n1065 ;
  assign n1072 = n1071 ^ n1067 ;
  assign n1059 = n1058 ^ n252 ;
  assign n1061 = n1060 ^ n1059 ;
  assign n1062 = n1061 ^ n663 ;
  assign n1054 = ~n128 & n448 ;
  assign n1055 = n1054 ^ n375 ;
  assign n1056 = n1055 ^ n797 ;
  assign n1051 = n1050 ^ n124 ;
  assign n1052 = n1051 ^ n100 ;
  assign n1053 = n1052 ^ n764 ;
  assign n1057 = n1056 ^ n1053 ;
  assign n1063 = n1062 ^ n1057 ;
  assign n1073 = n1072 ^ n1063 ;
  assign n1092 = n1091 ^ n1073 ;
  assign n1108 = n1107 ^ n1092 ;
  assign n1109 = ~n1049 & ~n1108 ;
  assign n1110 = n1109 ^ n824 ;
  assign n1111 = ~n969 & n1110 ;
  assign n1112 = n743 ^ n701 ;
  assign n1159 = n809 ^ n760 ;
  assign n1160 = n1159 ^ n952 ;
  assign n1157 = n219 ^ n90 ;
  assign n1158 = n1157 ^ n1014 ;
  assign n1161 = n1160 ^ n1158 ;
  assign n1152 = n845 ^ n627 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1151 = n1150 ^ n1149 ;
  assign n1155 = n1154 ^ n1151 ;
  assign n1144 = n48 & ~n77 ;
  assign n1145 = x23 & n1144 ;
  assign n1142 = n954 ^ n725 ;
  assign n1143 = n1142 ^ n217 ;
  assign n1146 = n1145 ^ n1143 ;
  assign n1140 = n221 ^ n190 ;
  assign n1141 = n1140 ^ n370 ;
  assign n1147 = n1146 ^ n1141 ;
  assign n1156 = n1155 ^ n1147 ;
  assign n1162 = n1161 ^ n1156 ;
  assign n1136 = n888 ^ n129 ;
  assign n1135 = n506 ^ n363 ;
  assign n1137 = n1136 ^ n1135 ;
  assign n1131 = n1130 ^ n1129 ;
  assign n1132 = n1131 ^ n178 ;
  assign n1133 = n1132 ^ n521 ;
  assign n1134 = n1133 ^ n918 ;
  assign n1138 = n1137 ^ n1134 ;
  assign n1125 = n882 ^ n810 ;
  assign n1123 = n1122 ^ n206 ;
  assign n1121 = n409 ^ n196 ;
  assign n1124 = n1123 ^ n1121 ;
  assign n1126 = n1125 ^ n1124 ;
  assign n1118 = n483 ^ n308 ;
  assign n1117 = n1116 ^ n292 ;
  assign n1119 = n1118 ^ n1117 ;
  assign n1113 = n914 ^ n143 ;
  assign n1114 = n1113 ^ n242 ;
  assign n1115 = n1114 ^ n116 ;
  assign n1120 = n1119 ^ n1115 ;
  assign n1127 = n1126 ^ n1120 ;
  assign n1139 = n1138 ^ n1127 ;
  assign n1163 = n1162 ^ n1139 ;
  assign n1208 = n1054 ^ n520 ;
  assign n1206 = n814 ^ n414 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1209 = n1208 ^ n1207 ;
  assign n1202 = n836 ^ n613 ;
  assign n1201 = n1099 ^ n250 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1199 = n455 ^ n265 ;
  assign n1197 = n171 & ~n12860 ;
  assign n1198 = n1197 ^ n1001 ;
  assign n1200 = n1199 ^ n1198 ;
  assign n1204 = n1203 ^ n1200 ;
  assign n1210 = n1209 ^ n1204 ;
  assign n1194 = n737 ^ n592 ;
  assign n1195 = n1194 ^ n790 ;
  assign n1190 = n897 ^ n541 ;
  assign n1191 = n1190 ^ n280 ;
  assign n1192 = n1191 ^ n621 ;
  assign n1189 = n1188 ^ n558 ;
  assign n1193 = n1192 ^ n1189 ;
  assign n1196 = n1195 ^ n1193 ;
  assign n1211 = n1210 ^ n1196 ;
  assign n1184 = n793 ^ n272 ;
  assign n1185 = n1184 ^ n303 ;
  assign n1182 = n1181 ^ n478 ;
  assign n1180 = n841 ^ n100 ;
  assign n1183 = n1182 ^ n1180 ;
  assign n1186 = n1185 ^ n1183 ;
  assign n1177 = n1176 ^ n192 ;
  assign n1178 = n1177 ^ n1060 ;
  assign n1172 = n597 ^ n496 ;
  assign n1171 = n416 ^ n88 ;
  assign n1173 = n1172 ^ n1171 ;
  assign n1169 = n726 ^ n642 ;
  assign n1170 = n1169 ^ n857 ;
  assign n1174 = n1173 ^ n1170 ;
  assign n1166 = n1085 ^ n380 ;
  assign n1167 = n1166 ^ n268 ;
  assign n1164 = n783 ^ n176 ;
  assign n1165 = n1164 ^ n848 ;
  assign n1168 = n1167 ^ n1165 ;
  assign n1175 = n1174 ^ n1168 ;
  assign n1179 = n1178 ^ n1175 ;
  assign n1187 = n1186 ^ n1179 ;
  assign n1212 = n1211 ^ n1187 ;
  assign n1213 = ~n1163 & ~n1212 ;
  assign n1214 = ~n1112 & n1213 ;
  assign n1467 = n660 ^ n577 ;
  assign n1465 = n612 ^ n180 ;
  assign n1466 = n1465 ^ n499 ;
  assign n1468 = n1467 ^ n1466 ;
  assign n1461 = n521 ^ n183 ;
  assign n1462 = n1461 ^ n583 ;
  assign n1463 = n1462 ^ n982 ;
  assign n1457 = n505 ^ n129 ;
  assign n1458 = n1457 ^ n1058 ;
  assign n1459 = n1458 ^ n87 ;
  assign n1456 = n567 ^ n513 ;
  assign n1460 = n1459 ^ n1456 ;
  assign n1464 = n1463 ^ n1460 ;
  assign n1469 = n1468 ^ n1464 ;
  assign n1453 = n1219 ^ n397 ;
  assign n1450 = n678 ^ n607 ;
  assign n1451 = n1450 ^ n983 ;
  assign n1452 = n1451 ^ n820 ;
  assign n1454 = n1453 ^ n1452 ;
  assign n1447 = n940 ^ n489 ;
  assign n1444 = n526 ^ n414 ;
  assign n1445 = n1444 ^ n450 ;
  assign n1446 = n1445 ^ n597 ;
  assign n1448 = n1447 ^ n1446 ;
  assign n1441 = n613 ^ n186 ;
  assign n1440 = n1045 ^ n292 ;
  assign n1442 = n1441 ^ n1440 ;
  assign n1437 = n790 ^ n500 ;
  assign n1438 = n1437 ^ n431 ;
  assign n1435 = n622 ^ n130 ;
  assign n1428 = n303 ^ n252 ;
  assign n1436 = n1435 ^ n1428 ;
  assign n1439 = n1438 ^ n1436 ;
  assign n1443 = n1442 ^ n1439 ;
  assign n1449 = n1448 ^ n1443 ;
  assign n1455 = n1454 ^ n1449 ;
  assign n1470 = n1469 ^ n1455 ;
  assign n1534 = n1099 ^ n416 ;
  assign n1535 = n1534 ^ n937 ;
  assign n1533 = n919 ^ n572 ;
  assign n1536 = n1535 ^ n1533 ;
  assign n1531 = n945 ^ n624 ;
  assign n1527 = n511 ^ n269 ;
  assign n1528 = n1527 ^ n1024 ;
  assign n1529 = n1528 ^ n291 ;
  assign n1530 = n1529 ^ n261 ;
  assign n1532 = n1531 ^ n1530 ;
  assign n1537 = n1536 ^ n1532 ;
  assign n1523 = n773 ^ n768 ;
  assign n1524 = n1523 ^ n283 ;
  assign n1521 = n176 ^ n91 ;
  assign n1522 = n1521 ^ n145 ;
  assign n1525 = n1524 ^ n1522 ;
  assign n1518 = n853 ^ n547 ;
  assign n1516 = n725 ^ n259 ;
  assign n1517 = n1516 ^ n242 ;
  assign n1519 = n1518 ^ n1517 ;
  assign n1512 = n747 ^ n627 ;
  assign n1514 = n1513 ^ n1512 ;
  assign n1510 = n219 ^ n151 ;
  assign n1509 = n540 ^ n305 ;
  assign n1511 = n1510 ^ n1509 ;
  assign n1515 = n1514 ^ n1511 ;
  assign n1520 = n1519 ^ n1515 ;
  assign n1526 = n1525 ^ n1520 ;
  assign n1538 = n1537 ^ n1526 ;
  assign n1504 = n592 ^ n391 ;
  assign n1505 = n1504 ^ n236 ;
  assign n1506 = n1505 ^ n570 ;
  assign n1502 = n779 ^ n280 ;
  assign n1500 = n425 ^ n225 ;
  assign n1501 = n1500 ^ n201 ;
  assign n1503 = n1502 ^ n1501 ;
  assign n1507 = n1506 ^ n1503 ;
  assign n1492 = n762 ^ n196 ;
  assign n1493 = n1492 ^ n498 ;
  assign n1496 = n1495 ^ n1493 ;
  assign n1490 = n971 ^ n543 ;
  assign n1489 = n379 ^ n157 ;
  assign n1491 = n1490 ^ n1489 ;
  assign n1497 = n1496 ^ n1491 ;
  assign n1487 = n914 ^ n172 ;
  assign n1488 = n1487 ^ n774 ;
  assign n1498 = n1497 ^ n1488 ;
  assign n1482 = n682 ^ n97 ;
  assign n1483 = n1482 ^ n561 ;
  assign n1481 = n1480 ^ n1273 ;
  assign n1484 = n1483 ^ n1481 ;
  assign n1485 = n1484 ^ n977 ;
  assign n1476 = n584 ^ n250 ;
  assign n1477 = n1476 ^ n814 ;
  assign n1478 = n1477 ^ n520 ;
  assign n1472 = n490 ^ n106 ;
  assign n1473 = n1472 ^ n1088 ;
  assign n1474 = n1473 ^ n192 ;
  assign n1471 = n677 ^ n149 ;
  assign n1475 = n1474 ^ n1471 ;
  assign n1479 = n1478 ^ n1475 ;
  assign n1486 = n1485 ^ n1479 ;
  assign n1499 = n1498 ^ n1486 ;
  assign n1508 = n1507 ^ n1499 ;
  assign n1539 = n1538 ^ n1508 ;
  assign n1540 = ~n1470 & ~n1539 ;
  assign n1375 = n662 ^ n116 ;
  assign n1372 = n1197 ^ n409 ;
  assign n1373 = n1372 ^ n1129 ;
  assign n1371 = n970 ^ n623 ;
  assign n1374 = n1373 ^ n1371 ;
  assign n1376 = n1375 ^ n1374 ;
  assign n1377 = n1376 ^ n1084 ;
  assign n1366 = n1001 ^ n954 ;
  assign n1367 = n1366 ^ n506 ;
  assign n1368 = n1367 ^ n149 ;
  assign n1363 = n518 ^ n369 ;
  assign n1364 = n1363 ^ n456 ;
  assign n1365 = n1364 ^ n579 ;
  assign n1369 = n1368 ^ n1365 ;
  assign n1358 = n1116 ^ n356 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1356 = n1355 ^ n186 ;
  assign n1357 = n1356 ^ n803 ;
  assign n1361 = n1360 ^ n1357 ;
  assign n1353 = n1021 ^ n197 ;
  assign n1352 = n1032 ^ n769 ;
  assign n1354 = n1353 ^ n1352 ;
  assign n1362 = n1361 ^ n1354 ;
  assign n1370 = n1369 ^ n1362 ;
  assign n1378 = n1377 ^ n1370 ;
  assign n1429 = n1428 ^ n584 ;
  assign n1425 = n932 ^ n624 ;
  assign n1426 = n1425 ^ n499 ;
  assign n1423 = n279 ^ n182 ;
  assign n1422 = n838 ^ n362 ;
  assign n1424 = n1423 ^ n1422 ;
  assign n1427 = n1426 ^ n1424 ;
  assign n1430 = n1429 ^ n1427 ;
  assign n1418 = n583 ^ n249 ;
  assign n1419 = n1418 ^ n1014 ;
  assign n1414 = n1249 ^ n401 ;
  assign n1415 = n1414 ^ n1058 ;
  assign n1416 = n1415 ^ n597 ;
  assign n1417 = n1416 ^ n273 ;
  assign n1420 = n1419 ^ n1417 ;
  assign n1339 = n221 ^ n217 ;
  assign n1411 = n1339 ^ n375 ;
  assign n1412 = n1411 ^ n229 ;
  assign n1408 = ~n74 & n254 ;
  assign n1409 = n1408 ^ n745 ;
  assign n1405 = n739 ^ n200 ;
  assign n1406 = n1405 ^ n308 ;
  assign n1407 = n1406 ^ n607 ;
  assign n1410 = n1409 ^ n1407 ;
  assign n1413 = n1412 ^ n1410 ;
  assign n1421 = n1420 ^ n1413 ;
  assign n1431 = n1430 ^ n1421 ;
  assign n1399 = n280 ^ n151 ;
  assign n1400 = n1399 ^ n1088 ;
  assign n1401 = n1400 ^ n565 ;
  assign n1396 = n542 ^ n172 ;
  assign n1397 = n1396 ^ n558 ;
  assign n1394 = n918 ^ n355 ;
  assign n1395 = n1394 ^ n905 ;
  assign n1398 = n1397 ^ n1395 ;
  assign n1402 = n1401 ^ n1398 ;
  assign n1318 = n689 ^ n291 ;
  assign n1392 = n1318 ^ n961 ;
  assign n1389 = n527 ^ n426 ;
  assign n1388 = n201 ^ n117 ;
  assign n1390 = n1389 ^ n1388 ;
  assign n1387 = n284 ^ n124 ;
  assign n1391 = n1390 ^ n1387 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n1403 = n1402 ^ n1393 ;
  assign n1383 = n1099 ^ n264 ;
  assign n1384 = n1383 ^ n413 ;
  assign n1381 = n725 ^ n677 ;
  assign n1379 = n589 ^ n258 ;
  assign n1380 = n1379 ^ n122 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1385 = n1384 ^ n1382 ;
  assign n1386 = n1385 ^ n882 ;
  assign n1404 = n1403 ^ n1386 ;
  assign n1432 = n1431 ^ n1404 ;
  assign n1433 = ~n1378 & ~n1432 ;
  assign n1260 = n893 ^ n266 ;
  assign n1261 = n1260 ^ n672 ;
  assign n1259 = n697 ^ n405 ;
  assign n1262 = n1261 ^ n1259 ;
  assign n1257 = n1206 ^ n364 ;
  assign n1254 = n1088 ^ n673 ;
  assign n1255 = n1254 ^ n577 ;
  assign n1256 = n1255 ^ n355 ;
  assign n1258 = n1257 ^ n1256 ;
  assign n1263 = n1262 ^ n1258 ;
  assign n1251 = n1250 ^ n1148 ;
  assign n1247 = n526 ^ n210 ;
  assign n1248 = n1247 ^ n131 ;
  assign n1252 = n1251 ^ n1248 ;
  assign n1244 = n269 ^ n178 ;
  assign n1243 = n280 ^ n222 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1241 = n279 ^ n149 ;
  assign n1240 = n726 ^ n378 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1246 = n1245 ^ n1242 ;
  assign n1253 = n1252 ^ n1246 ;
  assign n1264 = n1263 ^ n1253 ;
  assign n1235 = n1142 ^ n521 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1238 = n1237 ^ n1234 ;
  assign n1229 = n268 ^ n141 ;
  assign n1228 = n702 ^ n683 ;
  assign n1230 = n1229 ^ n1228 ;
  assign n1239 = n1238 ^ n1230 ;
  assign n1265 = n1264 ^ n1239 ;
  assign n1277 = n1276 ^ n1265 ;
  assign n1343 = n1135 ^ n186 ;
  assign n1344 = n1343 ^ n622 ;
  assign n1345 = n1344 ^ n668 ;
  assign n1340 = n1339 ^ n570 ;
  assign n1341 = n1340 ^ n804 ;
  assign n1342 = n1341 ^ n225 ;
  assign n1346 = n1345 ^ n1342 ;
  assign n1336 = n1029 ^ n117 ;
  assign n1335 = n379 ^ n175 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1331 = n559 ^ n124 ;
  assign n1332 = n1331 ^ n1014 ;
  assign n1330 = n558 ^ n194 ;
  assign n1333 = n1332 ^ n1330 ;
  assign n1334 = n1333 ^ n451 ;
  assign n1338 = n1337 ^ n1334 ;
  assign n1347 = n1346 ^ n1338 ;
  assign n1326 = n391 ^ n252 ;
  assign n1325 = n762 ^ n369 ;
  assign n1327 = n1326 ^ n1325 ;
  assign n1324 = n994 ^ n775 ;
  assign n1328 = n1327 ^ n1324 ;
  assign n1321 = n765 ^ n362 ;
  assign n1322 = n1321 ^ n192 ;
  assign n1319 = n1318 ^ n413 ;
  assign n1317 = n305 ^ n144 ;
  assign n1320 = n1319 ^ n1317 ;
  assign n1323 = n1322 ^ n1320 ;
  assign n1329 = n1328 ^ n1323 ;
  assign n1348 = n1347 ^ n1329 ;
  assign n1312 = n1311 ^ n527 ;
  assign n1308 = n565 ^ n376 ;
  assign n1309 = n1308 ^ n584 ;
  assign n1310 = n1309 ^ n520 ;
  assign n1313 = n1312 ^ n1310 ;
  assign n1305 = n764 ^ n200 ;
  assign n1306 = n1305 ^ n360 ;
  assign n1303 = n793 ^ n589 ;
  assign n1304 = n1303 ^ n1001 ;
  assign n1307 = n1306 ^ n1304 ;
  assign n1314 = n1313 ^ n1307 ;
  assign n1301 = n602 ^ n181 ;
  assign n1302 = n1301 ^ n258 ;
  assign n1315 = n1314 ^ n1302 ;
  assign n1297 = n768 ^ n425 ;
  assign n1298 = n1297 ^ n560 ;
  assign n1294 = n567 ^ n261 ;
  assign n1293 = n841 ^ n122 ;
  assign n1295 = n1294 ^ n1293 ;
  assign n1290 = n607 ^ n478 ;
  assign n1291 = n1290 ^ n201 ;
  assign n1292 = n1291 ^ n156 ;
  assign n1296 = n1295 ^ n1292 ;
  assign n1299 = n1298 ^ n1296 ;
  assign n1286 = n613 ^ n500 ;
  assign n1287 = n1286 ^ n881 ;
  assign n1283 = n790 ^ n259 ;
  assign n1284 = n1283 ^ n282 ;
  assign n1282 = n540 ^ n116 ;
  assign n1285 = n1284 ^ n1282 ;
  assign n1288 = n1287 ^ n1285 ;
  assign n1280 = n356 ^ n237 ;
  assign n1278 = n370 ^ n351 ;
  assign n1279 = n1278 ^ n99 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n1289 = n1288 ^ n1281 ;
  assign n1300 = n1299 ^ n1289 ;
  assign n1316 = n1315 ^ n1300 ;
  assign n1349 = n1348 ^ n1316 ;
  assign n1350 = ~n1277 & ~n1349 ;
  assign n1351 = ~n1227 & n1350 ;
  assign n1434 = n1433 ^ n1351 ;
  assign n1541 = n1540 ^ n1433 ;
  assign n1564 = n489 ^ n363 ;
  assign n1565 = n1564 ^ n1122 ;
  assign n1566 = n1565 ^ n210 ;
  assign n1561 = n764 ^ n239 ;
  assign n1562 = n1561 ^ n682 ;
  assign n1560 = n672 ^ n91 ;
  assign n1563 = n1562 ^ n1560 ;
  assign n1567 = n1566 ^ n1563 ;
  assign n1555 = n1355 ^ n203 ;
  assign n1556 = n1555 ^ n221 ;
  assign n1553 = n1206 ^ n118 ;
  assign n1554 = n1553 ^ n500 ;
  assign n1557 = n1556 ^ n1554 ;
  assign n1558 = n1557 ^ n1517 ;
  assign n1549 = n1014 ^ n527 ;
  assign n1550 = n1549 ^ n1172 ;
  assign n1548 = n1205 ^ n983 ;
  assign n1551 = n1550 ^ n1548 ;
  assign n1545 = n565 ^ n226 ;
  assign n1546 = n1545 ^ n690 ;
  assign n1543 = n512 ^ n391 ;
  assign n1542 = n351 ^ n124 ;
  assign n1544 = n1543 ^ n1542 ;
  assign n1547 = n1546 ^ n1544 ;
  assign n1552 = n1551 ^ n1547 ;
  assign n1559 = n1558 ^ n1552 ;
  assign n1568 = n1567 ^ n1559 ;
  assign n1624 = n897 ^ n613 ;
  assign n1625 = n1624 ^ n153 ;
  assign n1626 = n1625 ^ n1494 ;
  assign n1621 = n952 ^ n429 ;
  assign n1622 = n1621 ^ n635 ;
  assign n1623 = n1622 ^ n918 ;
  assign n1627 = n1626 ^ n1623 ;
  assign n1618 = n628 ^ n400 ;
  assign n1617 = n1335 ^ n313 ;
  assign n1619 = n1618 ^ n1617 ;
  assign n1614 = n642 ^ n148 ;
  assign n1615 = n1614 ^ n697 ;
  assign n1616 = n1615 ^ n773 ;
  assign n1620 = n1619 ^ n1616 ;
  assign n1628 = n1627 ^ n1620 ;
  assign n1610 = n976 ^ n677 ;
  assign n1608 = n560 ^ n268 ;
  assign n1609 = n1608 ^ n330 ;
  assign n1611 = n1610 ^ n1609 ;
  assign n1606 = n1605 ^ n1318 ;
  assign n1607 = n1606 ^ n238 ;
  assign n1612 = n1611 ^ n1607 ;
  assign n1600 = n747 ^ n641 ;
  assign n1601 = n1600 ^ n230 ;
  assign n1603 = n1602 ^ n1601 ;
  assign n1597 = n577 ^ n149 ;
  assign n1598 = n1597 ^ n87 ;
  assign n1599 = n1598 ^ n396 ;
  assign n1604 = n1603 ^ n1599 ;
  assign n1613 = n1612 ^ n1604 ;
  assign n1629 = n1628 ^ n1613 ;
  assign n1592 = n935 ^ n583 ;
  assign n1593 = n1592 ^ n156 ;
  assign n1590 = n1219 ^ n774 ;
  assign n1591 = n1590 ^ n110 ;
  assign n1594 = n1593 ^ n1591 ;
  assign n1588 = n1085 ^ n355 ;
  assign n1586 = n589 ^ n497 ;
  assign n1587 = n1586 ^ n300 ;
  assign n1589 = n1588 ^ n1587 ;
  assign n1595 = n1594 ^ n1589 ;
  assign n1582 = n1058 ^ n244 ;
  assign n1581 = n258 ^ n97 ;
  assign n1583 = n1582 ^ n1581 ;
  assign n1578 = ~n64 & n1144 ;
  assign n1577 = n542 ^ n200 ;
  assign n1579 = n1578 ^ n1577 ;
  assign n1576 = n981 ^ n245 ;
  assign n1580 = n1579 ^ n1576 ;
  assign n1584 = n1583 ^ n1580 ;
  assign n1574 = n1199 ^ n1039 ;
  assign n1571 = n1054 ^ n197 ;
  assign n1569 = n790 ^ n141 ;
  assign n1570 = n1569 ^ n250 ;
  assign n1572 = n1571 ^ n1570 ;
  assign n1573 = n1572 ^ n217 ;
  assign n1575 = n1574 ^ n1573 ;
  assign n1585 = n1584 ^ n1575 ;
  assign n1596 = n1595 ^ n1585 ;
  assign n1630 = n1629 ^ n1596 ;
  assign n1631 = ~n1568 & ~n1630 ;
  assign n1632 = n1631 ^ n1434 ;
  assign n1633 = n1632 ^ n1541 ;
  assign n1677 = n836 ^ n689 ;
  assign n1678 = n1677 ^ n438 ;
  assign n1675 = n932 ^ n570 ;
  assign n1676 = n1675 ^ n1674 ;
  assign n1679 = n1678 ^ n1676 ;
  assign n1671 = n971 ^ n483 ;
  assign n1672 = n1671 ^ n867 ;
  assign n1668 = n369 ^ n265 ;
  assign n1669 = n1668 ^ n550 ;
  assign n1670 = n1669 ^ n673 ;
  assign n1673 = n1672 ^ n1670 ;
  assign n1680 = n1679 ^ n1673 ;
  assign n1666 = n882 ^ n280 ;
  assign n1667 = n1666 ^ n296 ;
  assign n1681 = n1680 ^ n1667 ;
  assign n1660 = n1659 ^ n226 ;
  assign n1661 = n1660 ^ n1129 ;
  assign n1657 = n760 ^ n222 ;
  assign n1662 = n1661 ^ n1657 ;
  assign n1654 = n838 ^ n258 ;
  assign n1655 = n1654 ^ n1435 ;
  assign n1652 = n542 ^ n100 ;
  assign n1653 = n1652 ^ n1208 ;
  assign n1656 = n1655 ^ n1653 ;
  assign n1663 = n1662 ^ n1656 ;
  assign n1649 = n203 ^ n155 ;
  assign n1650 = n1649 ^ n667 ;
  assign n1648 = n1195 ^ n940 ;
  assign n1651 = n1650 ^ n1648 ;
  assign n1664 = n1663 ^ n1651 ;
  assign n1644 = n703 ^ n196 ;
  assign n1645 = n1644 ^ n518 ;
  assign n1641 = n782 ^ n773 ;
  assign n1642 = n1641 ^ n641 ;
  assign n1640 = n893 ^ n308 ;
  assign n1643 = n1642 ^ n1640 ;
  assign n1646 = n1645 ^ n1643 ;
  assign n1636 = n952 ^ n547 ;
  assign n1637 = n1636 ^ n507 ;
  assign n1638 = n1637 ^ n1450 ;
  assign n1634 = n728 ^ n416 ;
  assign n1635 = n1634 ^ n617 ;
  assign n1639 = n1638 ^ n1635 ;
  assign n1647 = n1646 ^ n1639 ;
  assign n1665 = n1664 ^ n1647 ;
  assign n1682 = n1681 ^ n1665 ;
  assign n1698 = n1487 ^ n712 ;
  assign n1697 = n1605 ^ n1372 ;
  assign n1699 = n1698 ^ n1697 ;
  assign n1700 = n1699 ^ n1237 ;
  assign n1694 = n1512 ^ n216 ;
  assign n1695 = n1694 ^ n1140 ;
  assign n1696 = n1695 ^ n1333 ;
  assign n1701 = n1700 ^ n1696 ;
  assign n1690 = n809 ^ n426 ;
  assign n1689 = n1527 ^ n635 ;
  assign n1691 = n1690 ^ n1689 ;
  assign n1687 = n1058 ^ n976 ;
  assign n1683 = n175 ^ n87 ;
  assign n1684 = n1683 ^ n351 ;
  assign n1685 = n1684 ^ n1088 ;
  assign n1686 = n1685 ^ n148 ;
  assign n1688 = n1687 ^ n1686 ;
  assign n1692 = n1691 ^ n1688 ;
  assign n1693 = n1692 ^ n588 ;
  assign n1702 = n1701 ^ n1693 ;
  assign n1703 = ~n1682 & ~n1702 ;
  assign n1704 = n1703 ^ n1351 ;
  assign n1705 = n1704 ^ n1631 ;
  assign n1706 = n1705 ^ n1541 ;
  assign n1708 = n1703 ^ n1434 ;
  assign n1709 = ~n1706 & ~n1708 ;
  assign n1710 = ~n1633 & n1709 ;
  assign n1711 = n1710 ^ n1704 ;
  assign n1712 = n1711 ^ n1434 ;
  assign n1713 = n1541 & n1712 ;
  assign n1714 = n1434 & n1713 ;
  assign n1715 = n1714 ^ n1433 ;
  assign n1828 = n403 ^ n279 ;
  assign n1829 = n1828 ^ n954 ;
  assign n1826 = n1494 ^ n732 ;
  assign n1827 = n1826 ^ n1029 ;
  assign n1830 = n1829 ^ n1827 ;
  assign n1822 = n321 ^ n190 ;
  assign n1823 = n1822 ^ n330 ;
  assign n1824 = n1823 ^ n972 ;
  assign n1819 = n636 ^ n500 ;
  assign n1820 = n1819 ^ n392 ;
  assign n1818 = n981 ^ n296 ;
  assign n1821 = n1820 ^ n1818 ;
  assign n1825 = n1824 ^ n1821 ;
  assign n1831 = n1830 ^ n1825 ;
  assign n1813 = n407 ^ n249 ;
  assign n1814 = n1813 ^ n1222 ;
  assign n1815 = n1814 ^ n1549 ;
  assign n1809 = n871 ^ n660 ;
  assign n1810 = n1809 ^ n497 ;
  assign n1808 = n541 ^ n237 ;
  assign n1811 = n1810 ^ n1808 ;
  assign n1806 = n1085 ^ n143 ;
  assign n1807 = n1806 ^ n499 ;
  assign n1812 = n1811 ^ n1807 ;
  assign n1816 = n1815 ^ n1812 ;
  assign n1803 = n1802 ^ n425 ;
  assign n1804 = n1803 ^ n1780 ;
  assign n1799 = n1798 ^ n848 ;
  assign n1800 = n1799 ^ n496 ;
  assign n1796 = n1683 ^ n785 ;
  assign n1797 = n1796 ^ n1050 ;
  assign n1801 = n1800 ^ n1797 ;
  assign n1805 = n1804 ^ n1801 ;
  assign n1817 = n1816 ^ n1805 ;
  assign n1832 = n1831 ^ n1817 ;
  assign n1745 = n747 ^ n285 ;
  assign n1746 = n1745 ^ n560 ;
  assign n1743 = n642 ^ n141 ;
  assign n1742 = n370 ^ n181 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1747 = n1746 ^ n1744 ;
  assign n1739 = n597 ^ n518 ;
  assign n1740 = n1739 ^ n537 ;
  assign n1737 = n583 ^ n149 ;
  assign n1736 = n739 ^ n379 ;
  assign n1738 = n1737 ^ n1736 ;
  assign n1741 = n1740 ^ n1738 ;
  assign n1748 = n1747 ^ n1741 ;
  assign n1732 = n819 ^ n612 ;
  assign n1733 = n1732 ^ n1339 ;
  assign n1731 = n204 ^ n148 ;
  assign n1734 = n1733 ^ n1731 ;
  assign n1729 = n1728 ^ n230 ;
  assign n1725 = n359 ^ n97 ;
  assign n1726 = n1725 ^ n380 ;
  assign n1727 = n1726 ^ n521 ;
  assign n1730 = n1729 ^ n1727 ;
  assign n1735 = n1734 ^ n1730 ;
  assign n1749 = n1748 ^ n1735 ;
  assign n1750 = n1749 ^ n1651 ;
  assign n1833 = n1832 ^ n1750 ;
  assign n1863 = n1513 ^ n1202 ;
  assign n1864 = n1863 ^ n397 ;
  assign n1861 = n764 ^ n176 ;
  assign n1859 = n1093 ^ n976 ;
  assign n1860 = n1859 ^ n571 ;
  assign n1862 = n1861 ^ n1860 ;
  assign n1865 = n1864 ^ n1862 ;
  assign n1856 = n1396 ^ n375 ;
  assign n1855 = n245 ^ n236 ;
  assign n1857 = n1856 ^ n1855 ;
  assign n1853 = n1290 ^ n570 ;
  assign n1852 = n797 ^ n450 ;
  assign n1854 = n1853 ^ n1852 ;
  assign n1858 = n1857 ^ n1854 ;
  assign n1866 = n1865 ^ n1858 ;
  assign n1849 = n706 ^ n303 ;
  assign n1847 = n1219 ^ n369 ;
  assign n1848 = n1847 ^ n1355 ;
  assign n1850 = n1849 ^ n1848 ;
  assign n1844 = n945 ^ n259 ;
  assign n1842 = n782 ^ n614 ;
  assign n1843 = n1842 ^ n565 ;
  assign n1845 = n1844 ^ n1843 ;
  assign n1839 = n455 ^ n161 ;
  assign n1840 = n1839 ^ n210 ;
  assign n1837 = n702 ^ n697 ;
  assign n1838 = n1837 ^ n602 ;
  assign n1841 = n1840 ^ n1838 ;
  assign n1846 = n1845 ^ n1841 ;
  assign n1851 = n1850 ^ n1846 ;
  assign n1867 = n1866 ^ n1851 ;
  assign n1836 = n1408 ^ n726 ;
  assign n1868 = n1867 ^ n1836 ;
  assign n1835 = n838 ^ n483 ;
  assign n1869 = n1868 ^ n1835 ;
  assign n1834 = n584 ^ n268 ;
  assign n1870 = n1869 ^ n1834 ;
  assign n1871 = ~n1833 & ~n1870 ;
  assign n1722 = n899 ^ n764 ;
  assign n1721 = n1249 ^ n621 ;
  assign n1723 = n1722 ^ n1721 ;
  assign n1718 = n607 ^ n282 ;
  assign n1719 = n1718 ^ n88 ;
  assign n1716 = n672 ^ n236 ;
  assign n1717 = n1716 ^ n100 ;
  assign n1720 = n1719 ^ n1717 ;
  assign n1724 = n1723 ^ n1720 ;
  assign n1751 = n1750 ^ n1724 ;
  assign n1767 = n914 ^ n137 ;
  assign n1765 = n624 ^ n417 ;
  assign n1766 = n1765 ^ n239 ;
  assign n1768 = n1767 ^ n1766 ;
  assign n1763 = n1644 ^ n206 ;
  assign n1764 = n1763 ^ n1001 ;
  assign n1769 = n1768 ^ n1764 ;
  assign n1758 = n1074 ^ n265 ;
  assign n1760 = n1759 ^ n1758 ;
  assign n1757 = n1756 ^ n1272 ;
  assign n1761 = n1760 ^ n1757 ;
  assign n1754 = n613 ^ n409 ;
  assign n1752 = n1394 ^ n1355 ;
  assign n1753 = n1752 ^ n542 ;
  assign n1755 = n1754 ^ n1753 ;
  assign n1762 = n1761 ^ n1755 ;
  assign n1770 = n1769 ^ n1762 ;
  assign n1771 = n1770 ^ n1329 ;
  assign n1794 = n1793 ^ n1771 ;
  assign n1795 = ~n1751 & ~n1794 ;
  assign n1872 = n1871 ^ n1795 ;
  assign n1873 = n1795 ^ n1631 ;
  assign n1943 = n779 ^ n512 ;
  assign n1944 = n1943 ^ n426 ;
  assign n1945 = n1944 ^ n971 ;
  assign n1941 = n1008 ^ n841 ;
  assign n1942 = n1941 ^ n742 ;
  assign n1946 = n1945 ^ n1942 ;
  assign n1937 = n1122 ^ n201 ;
  assign n1938 = n1937 ^ n268 ;
  assign n1936 = n1739 ^ n292 ;
  assign n1939 = n1938 ^ n1936 ;
  assign n1933 = n678 ^ n149 ;
  assign n1934 = n1933 ^ n785 ;
  assign n1931 = n762 ^ n450 ;
  assign n1932 = n1931 ^ n308 ;
  assign n1935 = n1934 ^ n1932 ;
  assign n1940 = n1939 ^ n1935 ;
  assign n1947 = n1946 ^ n1940 ;
  assign n1927 = n745 ^ n282 ;
  assign n1928 = n1927 ^ n612 ;
  assign n1925 = n765 ^ n401 ;
  assign n1926 = n1925 ^ n396 ;
  assign n1929 = n1928 ^ n1926 ;
  assign n1921 = n661 ^ n144 ;
  assign n1920 = n882 ^ n702 ;
  assign n1922 = n1921 ^ n1920 ;
  assign n1919 = n1545 ^ n950 ;
  assign n1923 = n1922 ^ n1919 ;
  assign n1916 = n751 ^ n541 ;
  assign n1917 = n1916 ^ n641 ;
  assign n1914 = n1254 ^ n838 ;
  assign n1915 = n1914 ^ n379 ;
  assign n1918 = n1917 ^ n1915 ;
  assign n1924 = n1923 ^ n1918 ;
  assign n1930 = n1929 ^ n1924 ;
  assign n1948 = n1947 ^ n1930 ;
  assign n1908 = n764 ^ n359 ;
  assign n1906 = n1494 ^ n1054 ;
  assign n1907 = n1906 ^ n400 ;
  assign n1909 = n1908 ^ n1907 ;
  assign n1903 = n507 ^ n483 ;
  assign n1904 = n1903 ^ n186 ;
  assign n1905 = n1904 ^ n542 ;
  assign n1910 = n1909 ^ n1905 ;
  assign n1899 = n689 ^ n607 ;
  assign n1898 = n881 ^ n559 ;
  assign n1900 = n1899 ^ n1898 ;
  assign n1896 = n809 ^ n363 ;
  assign n1897 = n1896 ^ n1461 ;
  assign n1901 = n1900 ^ n1897 ;
  assign n1902 = n1901 ^ n1281 ;
  assign n1911 = n1910 ^ n1902 ;
  assign n1893 = n623 ^ n513 ;
  assign n1894 = n1893 ^ n225 ;
  assign n1889 = n1129 ^ n589 ;
  assign n1888 = n726 ^ n376 ;
  assign n1890 = n1889 ^ n1888 ;
  assign n1891 = n1890 ^ n497 ;
  assign n1892 = n1891 ^ n192 ;
  assign n1895 = n1894 ^ n1892 ;
  assign n1912 = n1911 ^ n1895 ;
  assign n1883 = n1085 ^ n197 ;
  assign n1884 = n1883 ^ n1074 ;
  assign n1882 = n550 ^ n269 ;
  assign n1885 = n1884 ^ n1882 ;
  assign n1880 = n1249 ^ n490 ;
  assign n1879 = n221 ^ n156 ;
  assign n1881 = n1880 ^ n1879 ;
  assign n1886 = n1885 ^ n1881 ;
  assign n1875 = n259 ^ n117 ;
  assign n1877 = n1876 ^ n1875 ;
  assign n1874 = n1157 ^ n932 ;
  assign n1878 = n1877 ^ n1874 ;
  assign n1887 = n1886 ^ n1878 ;
  assign n1913 = n1912 ^ n1887 ;
  assign n1949 = n1948 ^ n1913 ;
  assign n1989 = n250 ^ n210 ;
  assign n1990 = n1989 ^ n428 ;
  assign n1987 = n478 ^ n425 ;
  assign n1986 = n1130 ^ n296 ;
  assign n1988 = n1987 ^ n1986 ;
  assign n1991 = n1990 ^ n1988 ;
  assign n1984 = n1302 ^ n222 ;
  assign n1980 = n1041 ^ n298 ;
  assign n1981 = n1980 ^ n279 ;
  assign n1983 = n1982 ^ n1981 ;
  assign n1985 = n1984 ^ n1983 ;
  assign n1992 = n1991 ^ n1985 ;
  assign n1976 = n797 ^ n413 ;
  assign n1974 = n935 ^ n239 ;
  assign n1975 = n1974 ^ n229 ;
  assign n1977 = n1976 ^ n1975 ;
  assign n1970 = n952 ^ n732 ;
  assign n1971 = n1970 ^ n355 ;
  assign n1969 = n853 ^ n172 ;
  assign n1972 = n1971 ^ n1969 ;
  assign n1967 = n819 ^ n176 ;
  assign n1968 = n1967 ^ n583 ;
  assign n1973 = n1972 ^ n1968 ;
  assign n1978 = n1977 ^ n1973 ;
  assign n1963 = n1819 ^ n1184 ;
  assign n1964 = n1963 ^ n1059 ;
  assign n1960 = n783 ^ n739 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1965 = n1964 ^ n1962 ;
  assign n1956 = n1197 ^ n309 ;
  assign n1957 = n1956 ^ n1116 ;
  assign n1955 = n1195 ^ n856 ;
  assign n1958 = n1957 ^ n1955 ;
  assign n1952 = n768 ^ n635 ;
  assign n1953 = n1952 ^ n155 ;
  assign n1950 = n1802 ^ n137 ;
  assign n1951 = n1950 ^ n570 ;
  assign n1954 = n1953 ^ n1951 ;
  assign n1959 = n1958 ^ n1954 ;
  assign n1966 = n1965 ^ n1959 ;
  assign n1979 = n1978 ^ n1966 ;
  assign n1993 = n1992 ^ n1979 ;
  assign n1994 = ~n1949 & ~n1993 ;
  assign n2024 = n426 ^ n88 ;
  assign n2025 = n2024 ^ n265 ;
  assign n2022 = n1847 ^ n918 ;
  assign n2023 = n2022 ^ n512 ;
  assign n2026 = n2025 ^ n2023 ;
  assign n2018 = n577 ^ n296 ;
  assign n2019 = n2018 ^ n236 ;
  assign n2016 = n642 ^ n456 ;
  assign n2017 = n2016 ^ n425 ;
  assign n2020 = n2019 ^ n2017 ;
  assign n2014 = n1259 ^ n624 ;
  assign n2015 = n2014 ^ n592 ;
  assign n2021 = n2020 ^ n2015 ;
  assign n2027 = n2026 ^ n2021 ;
  assign n2010 = n1739 ^ n393 ;
  assign n2009 = n1906 ^ n1247 ;
  assign n2011 = n2010 ^ n2009 ;
  assign n2005 = n1093 ^ n292 ;
  assign n2006 = n2005 ^ n602 ;
  assign n2007 = n2006 ^ n641 ;
  assign n2002 = n376 ^ n194 ;
  assign n2003 = n2002 ^ n178 ;
  assign n2004 = n2003 ^ n375 ;
  assign n2008 = n2007 ^ n2004 ;
  assign n2012 = n2011 ^ n2008 ;
  assign n1998 = n1001 ^ n245 ;
  assign n1999 = n1998 ^ n971 ;
  assign n1997 = n589 ^ n99 ;
  assign n2000 = n1999 ^ n1997 ;
  assign n2001 = n2000 ^ n1685 ;
  assign n2013 = n2012 ^ n2001 ;
  assign n2028 = n2027 ^ n2013 ;
  assign n2029 = n2028 ^ n940 ;
  assign n2092 = n1731 ^ n661 ;
  assign n2090 = n933 ^ n527 ;
  assign n2091 = n2090 ^ n1340 ;
  assign n2093 = n2092 ^ n2091 ;
  assign n2085 = n774 ^ n636 ;
  assign n2086 = n2085 ^ n558 ;
  assign n2082 = n380 ^ n258 ;
  assign n2083 = n2082 ^ n279 ;
  assign n2084 = n2083 ^ n410 ;
  assign n2087 = n2086 ^ n2084 ;
  assign n2080 = n321 ^ n156 ;
  assign n2077 = n881 ^ n313 ;
  assign n2076 = n308 ^ n255 ;
  assign n2078 = n2077 ^ n2076 ;
  assign n2079 = n2078 ^ n737 ;
  assign n2081 = n2080 ^ n2079 ;
  assign n2088 = n2087 ^ n2081 ;
  assign n2072 = n742 ^ n400 ;
  assign n2073 = n2072 ^ n1135 ;
  assign n2074 = n2073 ^ n899 ;
  assign n2069 = n1116 ^ n130 ;
  assign n2070 = n2069 ^ n1355 ;
  assign n2067 = n809 ^ n478 ;
  assign n2068 = n2067 ^ n1197 ;
  assign n2071 = n2070 ^ n2068 ;
  assign n2075 = n2074 ^ n2071 ;
  assign n2089 = n2088 ^ n2075 ;
  assign n2094 = n2093 ^ n2089 ;
  assign n2062 = n1321 ^ n848 ;
  assign n2060 = n893 ^ n550 ;
  assign n2059 = n945 ^ n116 ;
  assign n2061 = n2060 ^ n2059 ;
  assign n2063 = n2062 ^ n2061 ;
  assign n2056 = n428 ^ n141 ;
  assign n2057 = n2056 ^ n200 ;
  assign n2054 = n673 ^ n364 ;
  assign n2055 = n2054 ^ n303 ;
  assign n2058 = n2057 ^ n2055 ;
  assign n2064 = n2063 ^ n2058 ;
  assign n2051 = n1636 ^ n726 ;
  assign n2050 = n1472 ^ n416 ;
  assign n2052 = n2051 ^ n2050 ;
  assign n2048 = n635 ^ n228 ;
  assign n2045 = n1029 ^ n237 ;
  assign n2046 = n2045 ^ n747 ;
  assign n2047 = n2046 ^ n153 ;
  assign n2049 = n2048 ^ n2047 ;
  assign n2053 = n2052 ^ n2049 ;
  assign n2065 = n2064 ^ n2053 ;
  assign n2042 = n521 ^ n225 ;
  assign n2041 = n739 ^ n413 ;
  assign n2043 = n2042 ^ n2041 ;
  assign n2037 = n497 ^ n407 ;
  assign n2038 = n2037 ^ n1875 ;
  assign n2036 = n2035 ^ n846 ;
  assign n2039 = n2038 ^ n2036 ;
  assign n2032 = n1059 ^ n144 ;
  assign n2033 = n2032 ^ n677 ;
  assign n2030 = n566 ^ n212 ;
  assign n2031 = n2030 ^ n559 ;
  assign n2034 = n2033 ^ n2031 ;
  assign n2040 = n2039 ^ n2034 ;
  assign n2044 = n2043 ^ n2040 ;
  assign n2066 = n2065 ^ n2044 ;
  assign n2095 = n2094 ^ n2066 ;
  assign n2096 = ~n2029 & ~n2095 ;
  assign n2151 = n945 ^ n396 ;
  assign n2150 = n409 ^ n229 ;
  assign n2152 = n2151 ^ n2150 ;
  assign n2148 = n635 ^ n100 ;
  assign n2147 = n1576 ^ n190 ;
  assign n2149 = n2148 ^ n2147 ;
  assign n2153 = n2152 ^ n2149 ;
  assign n2141 = n893 ^ n222 ;
  assign n2142 = n2141 ^ n244 ;
  assign n2143 = n2142 ^ n765 ;
  assign n2138 = n407 ^ n149 ;
  assign n2139 = n2138 ^ n793 ;
  assign n2140 = n2139 ^ n1199 ;
  assign n2144 = n2143 ^ n2140 ;
  assign n2145 = n2144 ^ n2071 ;
  assign n2135 = n971 ^ n401 ;
  assign n2133 = n841 ^ n810 ;
  assign n2132 = n773 ^ n87 ;
  assign n2134 = n2133 ^ n2132 ;
  assign n2136 = n2135 ^ n2134 ;
  assign n2129 = n364 ^ n249 ;
  assign n2130 = n2129 ^ n227 ;
  assign n2126 = n1989 ^ n641 ;
  assign n2127 = n2126 ^ n867 ;
  assign n2124 = n1219 ^ n1129 ;
  assign n2123 = n614 ^ n137 ;
  assign n2125 = n2124 ^ n2123 ;
  assign n2128 = n2127 ^ n2125 ;
  assign n2131 = n2130 ^ n2128 ;
  assign n2137 = n2136 ^ n2131 ;
  assign n2146 = n2145 ^ n2137 ;
  assign n2154 = n2153 ^ n2146 ;
  assign n2119 = n425 ^ n175 ;
  assign n2117 = n678 ^ n236 ;
  assign n2118 = n2117 ^ n392 ;
  assign n2120 = n2119 ^ n2118 ;
  assign n2114 = n702 ^ n558 ;
  assign n2111 = n565 ^ n433 ;
  assign n2112 = n2111 ^ n495 ;
  assign n2113 = n2112 ^ n1269 ;
  assign n2115 = n2114 ^ n2113 ;
  assign n2109 = n1834 ^ n751 ;
  assign n2108 = n1828 ^ n623 ;
  assign n2110 = n2109 ^ n2108 ;
  assign n2116 = n2115 ^ n2110 ;
  assign n2121 = n2120 ^ n2116 ;
  assign n2104 = n1457 ^ n151 ;
  assign n2101 = n1732 ^ n291 ;
  assign n2102 = n2101 ^ n871 ;
  assign n2103 = n2102 ^ n88 ;
  assign n2105 = n2104 ^ n2103 ;
  assign n2099 = n2016 ^ n1122 ;
  assign n2097 = n1015 ^ n116 ;
  assign n2098 = n2097 ^ n252 ;
  assign n2100 = n2099 ^ n2098 ;
  assign n2106 = n2105 ^ n2100 ;
  assign n2107 = n2106 ^ n1887 ;
  assign n2122 = n2121 ^ n2107 ;
  assign n2155 = n2154 ^ n2122 ;
  assign n2179 = n1058 ^ n272 ;
  assign n2180 = n2179 ^ n745 ;
  assign n2181 = n2180 ^ n400 ;
  assign n2177 = n321 ^ n303 ;
  assign n2178 = n2177 ^ n914 ;
  assign n2182 = n2181 ^ n2178 ;
  assign n2173 = n1363 ^ n351 ;
  assign n2174 = n2173 ^ n804 ;
  assign n2171 = n772 ^ n764 ;
  assign n2172 = n2171 ^ n513 ;
  assign n2175 = n2174 ^ n2172 ;
  assign n2169 = n416 ^ n380 ;
  assign n2167 = n742 ^ n737 ;
  assign n2168 = n2167 ^ n2018 ;
  assign n2170 = n2169 ^ n2168 ;
  assign n2176 = n2175 ^ n2170 ;
  assign n2183 = n2182 ^ n2176 ;
  assign n2164 = n1177 ^ n239 ;
  assign n2161 = n559 ^ n176 ;
  assign n2162 = n2161 ^ n378 ;
  assign n2163 = n2162 ^ n662 ;
  assign n2165 = n2164 ^ n2163 ;
  assign n2157 = n857 ^ n217 ;
  assign n2158 = n2157 ^ n798 ;
  assign n2156 = n1625 ^ n145 ;
  assign n2159 = n2158 ^ n2156 ;
  assign n2160 = n2159 ^ n1386 ;
  assign n2166 = n2165 ^ n2160 ;
  assign n2184 = n2183 ^ n2166 ;
  assign n2185 = ~n2155 & ~n2184 ;
  assign n2222 = n987 ^ n284 ;
  assign n2223 = n2222 ^ n603 ;
  assign n2220 = n1023 ^ n176 ;
  assign n2221 = n2220 ^ n658 ;
  assign n2224 = n2223 ^ n2221 ;
  assign n2218 = n1255 ^ n251 ;
  assign n2215 = n856 ^ n660 ;
  assign n2216 = n2215 ^ n1135 ;
  assign n2213 = n613 ^ n512 ;
  assign n2214 = n2213 ^ n2016 ;
  assign n2217 = n2216 ^ n2214 ;
  assign n2219 = n2218 ^ n2217 ;
  assign n2225 = n2224 ^ n2219 ;
  assign n2226 = n2225 ^ n1253 ;
  assign n2208 = n483 ^ n229 ;
  assign n2209 = n2208 ^ n558 ;
  assign n2206 = n1122 ^ n1058 ;
  assign n2205 = n1085 ^ n1029 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2210 = n2209 ^ n2207 ;
  assign n2203 = n848 ^ n513 ;
  assign n2200 = n1129 ^ n742 ;
  assign n2201 = n2200 ^ n426 ;
  assign n2202 = n2201 ^ n265 ;
  assign n2204 = n2203 ^ n2202 ;
  assign n2211 = n2210 ^ n2204 ;
  assign n2196 = n1970 ^ n794 ;
  assign n2195 = n409 ^ n403 ;
  assign n2197 = n2196 ^ n2195 ;
  assign n2198 = n2197 ^ n1980 ;
  assign n2191 = n489 ^ n285 ;
  assign n2192 = n2191 ^ n1450 ;
  assign n2190 = n1001 ^ n212 ;
  assign n2193 = n2192 ^ n2190 ;
  assign n2187 = n973 ^ n116 ;
  assign n2188 = n2187 ^ n745 ;
  assign n2186 = n1157 ^ n303 ;
  assign n2189 = n2188 ^ n2186 ;
  assign n2194 = n2193 ^ n2189 ;
  assign n2199 = n2198 ^ n2194 ;
  assign n2212 = n2211 ^ n2199 ;
  assign n2227 = n2226 ^ n2212 ;
  assign n2262 = n244 ^ n201 ;
  assign n2263 = n2262 ^ n359 ;
  assign n2264 = n2263 ^ n914 ;
  assign n2261 = n1956 ^ n505 ;
  assign n2265 = n2264 ^ n2261 ;
  assign n2259 = n527 ^ n252 ;
  assign n2258 = n1117 ^ n239 ;
  assign n2260 = n2259 ^ n2258 ;
  assign n2266 = n2265 ^ n2260 ;
  assign n2254 = n2169 ^ n417 ;
  assign n2253 = n413 ^ n124 ;
  assign n2255 = n2254 ^ n2253 ;
  assign n2251 = n1759 ^ n1658 ;
  assign n2249 = n451 ^ n273 ;
  assign n2250 = n2249 ^ n1195 ;
  assign n2252 = n2251 ^ n2250 ;
  assign n2256 = n2255 ^ n2252 ;
  assign n2245 = n1172 ^ n197 ;
  assign n2243 = n392 ^ n245 ;
  assign n2244 = n2243 ^ n225 ;
  assign n2246 = n2245 ^ n2244 ;
  assign n2240 = n567 ^ n542 ;
  assign n2241 = n2240 ^ n237 ;
  assign n2242 = n2241 ^ n918 ;
  assign n2247 = n2246 ^ n2242 ;
  assign n2236 = n1130 ^ n932 ;
  assign n2237 = n2236 ^ n990 ;
  assign n2234 = n1074 ^ n153 ;
  assign n2233 = n1219 ^ n175 ;
  assign n2235 = n2234 ^ n2233 ;
  assign n2238 = n2237 ^ n2235 ;
  assign n2231 = n912 ^ n192 ;
  assign n2228 = n809 ^ n144 ;
  assign n2229 = n2228 ^ n782 ;
  assign n2230 = n2229 ^ n845 ;
  assign n2232 = n2231 ^ n2230 ;
  assign n2239 = n2238 ^ n2232 ;
  assign n2248 = n2247 ^ n2239 ;
  assign n2257 = n2256 ^ n2248 ;
  assign n2267 = n2266 ^ n2257 ;
  assign n2268 = ~n2227 & ~n2267 ;
  assign n2310 = n506 ^ n425 ;
  assign n2311 = n2310 ^ n568 ;
  assign n2308 = n1001 ^ n945 ;
  assign n2307 = n726 ^ n148 ;
  assign n2309 = n2308 ^ n2307 ;
  assign n2312 = n2311 ^ n2309 ;
  assign n2317 = n2316 ^ n2312 ;
  assign n2303 = n520 ^ n359 ;
  assign n2301 = n732 ^ n689 ;
  assign n2302 = n2301 ^ n1206 ;
  assign n2304 = n2303 ^ n2302 ;
  assign n2305 = n2304 ^ n185 ;
  assign n2298 = n298 ^ n197 ;
  assign n2299 = n2298 ^ n284 ;
  assign n2296 = n1668 ^ n583 ;
  assign n2295 = n2046 ^ n308 ;
  assign n2297 = n2296 ^ n2295 ;
  assign n2300 = n2299 ^ n2297 ;
  assign n2306 = n2305 ^ n2300 ;
  assign n2318 = n2317 ^ n2306 ;
  assign n2291 = n790 ^ n200 ;
  assign n2289 = n2129 ^ n499 ;
  assign n2290 = n2289 ^ n313 ;
  assign n2292 = n2291 ^ n2290 ;
  assign n2286 = n1644 ^ n1054 ;
  assign n2285 = n1785 ^ n849 ;
  assign n2287 = n2286 ^ n2285 ;
  assign n2282 = n673 ^ n264 ;
  assign n2283 = n2282 ^ n1215 ;
  assign n2284 = n2283 ^ n2213 ;
  assign n2288 = n2287 ^ n2284 ;
  assign n2293 = n2292 ^ n2288 ;
  assign n2278 = n819 ^ n725 ;
  assign n2277 = n1893 ^ n737 ;
  assign n2279 = n2278 ^ n2277 ;
  assign n2276 = n542 ^ n405 ;
  assign n2280 = n2279 ^ n2276 ;
  assign n2274 = n1085 ^ n661 ;
  assign n2272 = n590 ^ n273 ;
  assign n2269 = n760 ^ n156 ;
  assign n2270 = n2269 ^ n279 ;
  assign n2271 = n2270 ^ n1956 ;
  assign n2273 = n2272 ^ n2271 ;
  assign n2275 = n2274 ^ n2273 ;
  assign n2281 = n2280 ^ n2275 ;
  assign n2294 = n2293 ^ n2281 ;
  assign n2319 = n2318 ^ n2294 ;
  assign n2360 = n1798 ^ n679 ;
  assign n2361 = n2360 ^ n2141 ;
  assign n2358 = n500 ^ n269 ;
  assign n2355 = n641 ^ n109 ;
  assign n2356 = n2355 ^ n565 ;
  assign n2354 = n526 ^ n305 ;
  assign n2357 = n2356 ^ n2354 ;
  assign n2359 = n2358 ^ n2357 ;
  assign n2362 = n2361 ^ n2359 ;
  assign n2348 = n845 ^ n321 ;
  assign n2349 = n2348 ^ n1355 ;
  assign n2347 = n1649 ^ n1504 ;
  assign n2350 = n2349 ^ n2347 ;
  assign n2351 = n2350 ^ n2181 ;
  assign n2345 = n871 ^ n413 ;
  assign n2343 = n559 ^ n87 ;
  assign n2341 = n1330 ^ n612 ;
  assign n2342 = n2341 ^ n153 ;
  assign n2344 = n2343 ^ n2342 ;
  assign n2346 = n2345 ^ n2344 ;
  assign n2352 = n2351 ^ n2346 ;
  assign n2336 = n625 ^ n255 ;
  assign n2334 = n577 ^ n282 ;
  assign n2335 = n2334 ^ n705 ;
  assign n2337 = n2336 ^ n2335 ;
  assign n2332 = n570 ^ n216 ;
  assign n2330 = n971 ^ n360 ;
  assign n2331 = n2330 ^ n1074 ;
  assign n2333 = n2332 ^ n2331 ;
  assign n2338 = n2337 ^ n2333 ;
  assign n2327 = n1099 ^ n212 ;
  assign n2325 = n954 ^ n379 ;
  assign n2326 = n2325 ^ n614 ;
  assign n2328 = n2327 ^ n2326 ;
  assign n2320 = n407 ^ n250 ;
  assign n2321 = n2320 ^ n130 ;
  assign n2322 = n2321 ^ n856 ;
  assign n2323 = n2322 ^ n1148 ;
  assign n2324 = n2323 ^ n1130 ;
  assign n2329 = n2328 ^ n2324 ;
  assign n2339 = n2338 ^ n2329 ;
  assign n2340 = n2339 ^ n788 ;
  assign n2353 = n2352 ^ n2340 ;
  assign n2363 = n2362 ^ n2353 ;
  assign n2364 = ~n2319 & ~n2363 ;
  assign n2392 = n753 ^ n661 ;
  assign n2390 = n987 ^ n881 ;
  assign n2389 = n1088 ^ n194 ;
  assign n2391 = n2390 ^ n2389 ;
  assign n2393 = n2392 ^ n2391 ;
  assign n2386 = n862 ^ n425 ;
  assign n2387 = n2386 ^ n237 ;
  assign n2384 = n1358 ^ n223 ;
  assign n2385 = n2384 ^ n283 ;
  assign n2388 = n2387 ^ n2385 ;
  assign n2394 = n2393 ^ n2388 ;
  assign n2379 = n400 ^ n151 ;
  assign n2380 = n2379 ^ n2320 ;
  assign n2377 = n500 ^ n212 ;
  assign n2378 = n2377 ^ n1021 ;
  assign n2381 = n2380 ^ n2378 ;
  assign n2374 = n1093 ^ n137 ;
  assign n2375 = n2374 ^ n814 ;
  assign n2371 = n779 ^ n129 ;
  assign n2372 = n2371 ^ n292 ;
  assign n2373 = n2372 ^ n732 ;
  assign n2376 = n2375 ^ n2373 ;
  assign n2382 = n2381 ^ n2376 ;
  assign n2368 = n554 ^ n375 ;
  assign n2369 = n2368 ^ n760 ;
  assign n2365 = n589 ^ n429 ;
  assign n2366 = n2365 ^ n392 ;
  assign n2367 = n2366 ^ n1494 ;
  assign n2370 = n2369 ^ n2367 ;
  assign n2383 = n2382 ^ n2370 ;
  assign n2395 = n2394 ^ n2383 ;
  assign n2396 = n2395 ^ n1388 ;
  assign n2442 = n391 ^ n236 ;
  assign n2443 = n2442 ^ n478 ;
  assign n2444 = n2443 ^ n683 ;
  assign n2440 = n945 ^ n920 ;
  assign n2441 = n2440 ^ n1521 ;
  assign n2445 = n2444 ^ n2441 ;
  assign n2436 = n893 ^ n882 ;
  assign n2435 = n505 ^ n426 ;
  assign n2437 = n2436 ^ n2435 ;
  assign n2433 = n954 ^ n376 ;
  assign n2432 = n622 ^ n104 ;
  assign n2434 = n2433 ^ n2432 ;
  assign n2438 = n2437 ^ n2434 ;
  assign n2430 = n1148 ^ n952 ;
  assign n2429 = n1523 ^ n558 ;
  assign n2431 = n2430 ^ n2429 ;
  assign n2439 = n2438 ^ n2431 ;
  assign n2446 = n2445 ^ n2439 ;
  assign n2447 = n2446 ^ n1584 ;
  assign n2423 = n351 ^ n249 ;
  assign n2424 = n2423 ^ n1487 ;
  assign n2425 = n2424 ^ n854 ;
  assign n2426 = n2425 ^ n942 ;
  assign n2419 = n672 ^ n303 ;
  assign n2420 = n2419 ^ n726 ;
  assign n2417 = n703 ^ n602 ;
  assign n2418 = n2417 ^ n819 ;
  assign n2421 = n2420 ^ n2418 ;
  assign n2414 = n1224 ^ n521 ;
  assign n2413 = n1608 ^ n495 ;
  assign n2415 = n2414 ^ n2413 ;
  assign n2411 = n1176 ^ n265 ;
  assign n2408 = n856 ^ n677 ;
  assign n2409 = n2408 ^ n130 ;
  assign n2410 = n2409 ^ n1197 ;
  assign n2412 = n2411 ^ n2410 ;
  assign n2416 = n2415 ^ n2412 ;
  assign n2422 = n2421 ^ n2416 ;
  assign n2427 = n2426 ^ n2422 ;
  assign n2405 = n1765 ^ n230 ;
  assign n2404 = n1683 ^ n364 ;
  assign n2406 = n2405 ^ n2404 ;
  assign n2401 = n799 ^ n747 ;
  assign n2397 = n570 ^ n456 ;
  assign n2398 = n2397 ^ n790 ;
  assign n2399 = n2398 ^ n409 ;
  assign n2400 = n2399 ^ n512 ;
  assign n2402 = n2401 ^ n2400 ;
  assign n2403 = n2402 ^ n638 ;
  assign n2407 = n2406 ^ n2403 ;
  assign n2428 = n2427 ^ n2407 ;
  assign n2448 = n2447 ^ n2428 ;
  assign n2449 = ~n2396 & ~n2448 ;
  assign n2450 = n1948 ^ n1596 ;
  assign n2481 = n496 ^ n456 ;
  assign n2482 = n2481 ^ n1387 ;
  assign n2483 = n2482 ^ n2141 ;
  assign n2478 = n1130 ^ n737 ;
  assign n2476 = n973 ^ n375 ;
  assign n2477 = n2476 ^ n636 ;
  assign n2479 = n2478 ^ n2477 ;
  assign n2474 = n614 ^ n143 ;
  assign n2473 = n1148 ^ n540 ;
  assign n2475 = n2474 ^ n2473 ;
  assign n2480 = n2479 ^ n2475 ;
  assign n2484 = n2483 ^ n2480 ;
  assign n2469 = n567 ^ n362 ;
  assign n2466 = n954 ^ n433 ;
  assign n2467 = n2466 ^ n2215 ;
  assign n2465 = n579 ^ n547 ;
  assign n2468 = n2467 ^ n2465 ;
  assign n2470 = n2469 ^ n2468 ;
  assign n2471 = n2470 ^ n1769 ;
  assign n2462 = n212 ^ n190 ;
  assign n2459 = n867 ^ n635 ;
  assign n2458 = n848 ^ n305 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2461 = n2460 ^ n272 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2455 = n1967 ^ n526 ;
  assign n2456 = n2455 ^ n1029 ;
  assign n2453 = n1093 ^ n172 ;
  assign n2451 = n697 ^ n273 ;
  assign n2452 = n2451 ^ n1050 ;
  assign n2454 = n2453 ^ n2452 ;
  assign n2457 = n2456 ^ n2454 ;
  assign n2464 = n2463 ^ n2457 ;
  assign n2472 = n2471 ^ n2464 ;
  assign n2485 = n2484 ^ n2472 ;
  assign n2486 = ~n2450 & ~n2485 ;
  assign n2521 = n2379 ^ n1456 ;
  assign n2520 = n2196 ^ n991 ;
  assign n2522 = n2521 ^ n2520 ;
  assign n2516 = n624 ^ n370 ;
  assign n2517 = n2516 ^ n1219 ;
  assign n2518 = n2517 ^ n401 ;
  assign n2515 = n178 ^ n91 ;
  assign n2519 = n2518 ^ n2515 ;
  assign n2523 = n2522 ^ n2519 ;
  assign n2511 = n1088 ^ n841 ;
  assign n2510 = n2509 ^ n273 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2507 = n1640 ^ n391 ;
  assign n2506 = n1054 ^ n983 ;
  assign n2508 = n2507 ^ n2506 ;
  assign n2513 = n2512 ^ n2508 ;
  assign n2503 = n871 ^ n804 ;
  assign n2502 = n1116 ^ n106 ;
  assign n2504 = n2503 ^ n2502 ;
  assign n2500 = n867 ^ n407 ;
  assign n2499 = n1839 ^ n268 ;
  assign n2501 = n2500 ^ n2499 ;
  assign n2505 = n2504 ^ n2501 ;
  assign n2514 = n2513 ^ n2505 ;
  assign n2524 = n2523 ^ n2514 ;
  assign n2495 = n971 ^ n219 ;
  assign n2496 = n2495 ^ n1783 ;
  assign n2497 = n2496 ^ n1683 ;
  assign n2492 = n450 ^ n297 ;
  assign n2493 = n2492 ^ n819 ;
  assign n2490 = n1099 ^ n124 ;
  assign n2487 = n540 ^ n117 ;
  assign n2488 = n2487 ^ n521 ;
  assign n2489 = n2488 ^ n506 ;
  assign n2491 = n2490 ^ n2489 ;
  assign n2494 = n2493 ^ n2491 ;
  assign n2498 = n2497 ^ n2494 ;
  assign n2525 = n2524 ^ n2498 ;
  assign n2551 = n740 ^ n272 ;
  assign n2546 = n511 ^ n379 ;
  assign n2544 = n363 ^ n244 ;
  assign n2545 = n2544 ^ n403 ;
  assign n2547 = n2546 ^ n2545 ;
  assign n2541 = n1774 ^ n1129 ;
  assign n2542 = n2541 ^ n394 ;
  assign n2543 = n2542 ^ n313 ;
  assign n2548 = n2547 ^ n2543 ;
  assign n2539 = n1555 ^ n621 ;
  assign n2536 = n897 ^ n417 ;
  assign n2537 = n2536 ^ n627 ;
  assign n2538 = n2537 ^ n1597 ;
  assign n2540 = n2539 ^ n2538 ;
  assign n2549 = n2548 ^ n2540 ;
  assign n2533 = n1634 ^ n602 ;
  assign n2534 = n2533 ^ n2099 ;
  assign n2530 = n2177 ^ n196 ;
  assign n2531 = n2530 ^ n768 ;
  assign n2526 = n1592 ^ n255 ;
  assign n2527 = n2526 ^ n932 ;
  assign n2528 = n2527 ^ n192 ;
  assign n2529 = n2528 ^ n1085 ;
  assign n2532 = n2531 ^ n2529 ;
  assign n2535 = n2534 ^ n2532 ;
  assign n2550 = n2549 ^ n2535 ;
  assign n2552 = n2551 ^ n2550 ;
  assign n2553 = n2552 ^ n701 ;
  assign n2554 = ~n2525 & ~n2553 ;
  assign n2555 = n2256 ^ n765 ;
  assign n2556 = n2555 ^ n2225 ;
  assign n2605 = n872 ^ n203 ;
  assign n2603 = n2356 ^ n186 ;
  assign n2604 = n2603 ^ n621 ;
  assign n2606 = n2605 ^ n2604 ;
  assign n2599 = n1104 ^ n608 ;
  assign n2598 = n2171 ^ n751 ;
  assign n2600 = n2599 ^ n2598 ;
  assign n2596 = n2348 ^ n959 ;
  assign n2597 = n2596 ^ n2435 ;
  assign n2601 = n2600 ^ n2597 ;
  assign n2593 = n2592 ^ n571 ;
  assign n2594 = n2593 ^ n682 ;
  assign n2595 = n2594 ^ n2333 ;
  assign n2602 = n2601 ^ n2595 ;
  assign n2607 = n2606 ^ n2602 ;
  assign n2589 = n1509 ^ n519 ;
  assign n2586 = n1355 ^ n625 ;
  assign n2584 = n636 ^ n204 ;
  assign n2583 = n478 ^ n100 ;
  assign n2585 = n2584 ^ n2583 ;
  assign n2587 = n2586 ^ n2585 ;
  assign n2580 = n1826 ^ n496 ;
  assign n2581 = n2580 ^ n175 ;
  assign n2578 = n1472 ^ n703 ;
  assign n2579 = n2578 ^ n222 ;
  assign n2582 = n2581 ^ n2579 ;
  assign n2588 = n2587 ^ n2582 ;
  assign n2590 = n2589 ^ n2588 ;
  assign n2574 = n793 ^ n584 ;
  assign n2575 = n2574 ^ n918 ;
  assign n2571 = n513 ^ n266 ;
  assign n2572 = n2571 ^ n672 ;
  assign n2569 = n768 ^ n559 ;
  assign n2570 = n2569 ^ n2371 ;
  assign n2573 = n2572 ^ n2570 ;
  assign n2576 = n2575 ^ n2573 ;
  assign n2565 = n1549 ^ n255 ;
  assign n2566 = n2565 ^ n1125 ;
  assign n2567 = n2566 ^ n801 ;
  assign n2562 = n897 ^ n378 ;
  assign n2560 = n697 ^ n245 ;
  assign n2561 = n2560 ^ n206 ;
  assign n2563 = n2562 ^ n2561 ;
  assign n2558 = n1636 ^ n1064 ;
  assign n2557 = n1828 ^ n1783 ;
  assign n2559 = n2558 ^ n2557 ;
  assign n2564 = n2563 ^ n2559 ;
  assign n2568 = n2567 ^ n2564 ;
  assign n2577 = n2576 ^ n2568 ;
  assign n2591 = n2590 ^ n2577 ;
  assign n2608 = n2607 ^ n2591 ;
  assign n2609 = ~n2556 & ~n2608 ;
  assign n2641 = n2467 ^ n689 ;
  assign n2642 = n2641 ^ n658 ;
  assign n2638 = n537 ^ n110 ;
  assign n2639 = n2638 ^ n1222 ;
  assign n2640 = n2639 ^ n1424 ;
  assign n2643 = n2642 ^ n2640 ;
  assign n2634 = n1967 ^ n1450 ;
  assign n2632 = n291 ^ n117 ;
  assign n2633 = n2632 ^ n2348 ;
  assign n2635 = n2634 ^ n2633 ;
  assign n2636 = n2635 ^ n1230 ;
  assign n2628 = n2627 ^ n937 ;
  assign n2629 = n2628 ^ n201 ;
  assign n2630 = n2629 ^ n1159 ;
  assign n2625 = n1007 ^ n799 ;
  assign n2626 = n2625 ^ n520 ;
  assign n2631 = n2630 ^ n2626 ;
  assign n2637 = n2636 ^ n2631 ;
  assign n2644 = n2643 ^ n2637 ;
  assign n2621 = n981 ^ n183 ;
  assign n2622 = n2621 ^ n1123 ;
  assign n2623 = n2622 ^ n1929 ;
  assign n2618 = n400 ^ n361 ;
  assign n2616 = n667 ^ n90 ;
  assign n2614 = n1731 ^ n161 ;
  assign n2615 = n2614 ^ n303 ;
  assign n2617 = n2616 ^ n2615 ;
  assign n2619 = n2618 ^ n2617 ;
  assign n2611 = n1956 ^ n881 ;
  assign n2610 = n742 ^ n363 ;
  assign n2612 = n2611 ^ n2610 ;
  assign n2613 = n2612 ^ n2463 ;
  assign n2620 = n2619 ^ n2613 ;
  assign n2624 = n2623 ^ n2620 ;
  assign n2645 = n2644 ^ n2624 ;
  assign n2646 = ~n2029 & ~n2645 ;
  assign n2654 = n1050 ^ n558 ;
  assign n2655 = n2654 ^ n1086 ;
  assign n2656 = n2655 ^ n1020 ;
  assign n2651 = n881 ^ n703 ;
  assign n2652 = n2651 ^ n305 ;
  assign n2649 = n579 ^ n292 ;
  assign n2647 = n809 ^ n521 ;
  assign n2648 = n2647 ^ n678 ;
  assign n2650 = n2649 ^ n2648 ;
  assign n2653 = n2652 ^ n2650 ;
  assign n2657 = n2656 ^ n2653 ;
  assign n2658 = n2657 ^ n1857 ;
  assign n2683 = n778 ^ n514 ;
  assign n2681 = n743 ^ n405 ;
  assign n2682 = n2681 ^ n1054 ;
  assign n2684 = n2683 ^ n2682 ;
  assign n2679 = n954 ^ n804 ;
  assign n2677 = n356 ^ n151 ;
  assign n2678 = n2677 ^ n762 ;
  assign n2680 = n2679 ^ n2678 ;
  assign n2685 = n2684 ^ n2680 ;
  assign n2674 = n844 ^ n378 ;
  assign n2673 = n2541 ^ n149 ;
  assign n2675 = n2674 ^ n2673 ;
  assign n2670 = n570 ^ n376 ;
  assign n2671 = n2670 ^ n364 ;
  assign n2672 = n2671 ^ n1145 ;
  assign n2676 = n2675 ^ n2672 ;
  assign n2686 = n2685 ^ n2676 ;
  assign n2667 = n945 ^ n933 ;
  assign n2668 = n2667 ^ n886 ;
  assign n2663 = n819 ^ n230 ;
  assign n2662 = n636 ^ n106 ;
  assign n2664 = n2663 ^ n2662 ;
  assign n2660 = n952 ^ n602 ;
  assign n2659 = n597 ^ n298 ;
  assign n2661 = n2660 ^ n2659 ;
  assign n2665 = n2664 ^ n2661 ;
  assign n2666 = n2665 ^ n1292 ;
  assign n2669 = n2668 ^ n2666 ;
  assign n2687 = n2686 ^ n2669 ;
  assign n2688 = ~n2658 & ~n2687 ;
  assign n2734 = n127 ^ n58 ;
  assign n2731 = n108 ^ n98 ;
  assign n2732 = n2731 ^ x23 ;
  assign n2733 = n2732 ^ n73 ;
  assign n2735 = n2734 ^ n2733 ;
  assign n2736 = n103 & ~n2735 ;
  assign n2726 = n682 ^ n560 ;
  assign n2724 = n785 ^ n429 ;
  assign n2723 = n1088 ^ n871 ;
  assign n2725 = n2724 ^ n2723 ;
  assign n2727 = n2726 ^ n2725 ;
  assign n2720 = n838 ^ n547 ;
  assign n2721 = n2720 ^ n1001 ;
  assign n2722 = n2721 ^ n585 ;
  assign n2728 = n2727 ^ n2722 ;
  assign n2717 = n2161 ^ n361 ;
  assign n2718 = n2717 ^ n862 ;
  assign n2713 = n732 ^ n499 ;
  assign n2714 = n2713 ^ n370 ;
  assign n2715 = n2714 ^ n161 ;
  assign n2711 = n632 ^ n197 ;
  assign n2708 = n642 ^ n210 ;
  assign n2709 = n2708 ^ n396 ;
  assign n2710 = n2709 ^ n848 ;
  assign n2712 = n2711 ^ n2710 ;
  assign n2716 = n2715 ^ n2712 ;
  assign n2719 = n2718 ^ n2716 ;
  assign n2729 = n2728 ^ n2719 ;
  assign n463 = x26 ^ x24 ;
  assign n466 = n463 ^ n65 ;
  assign n468 = n467 ^ x23 ;
  assign n469 = n468 ^ n65 ;
  assign n470 = n466 & ~n469 ;
  assign n471 = n470 ^ n65 ;
  assign n472 = n96 & ~n471 ;
  assign n461 = n81 ^ n62 ;
  assign n462 = n461 ^ n73 ;
  assign n464 = n463 ^ n462 ;
  assign n465 = n241 & n464 ;
  assign n473 = n472 ^ n465 ;
  assign n2703 = n1148 ^ n473 ;
  assign n2702 = n836 ^ n222 ;
  assign n2704 = n2703 ^ n2702 ;
  assign n2701 = n1381 ^ n1064 ;
  assign n2705 = n2704 ^ n2701 ;
  assign n2699 = n2377 ^ n577 ;
  assign n2697 = n1387 ^ n541 ;
  assign n2698 = n2697 ^ n773 ;
  assign n2700 = n2699 ^ n2698 ;
  assign n2706 = n2705 ^ n2700 ;
  assign n2693 = n1074 ^ n225 ;
  assign n2694 = n2693 ^ n772 ;
  assign n2690 = n868 ^ n414 ;
  assign n2691 = n2690 ^ n263 ;
  assign n2689 = n527 ^ n90 ;
  assign n2692 = n2691 ^ n2689 ;
  assign n2695 = n2694 ^ n2692 ;
  assign n2696 = n2695 ^ n1977 ;
  assign n2707 = n2706 ^ n2696 ;
  assign n2730 = n2729 ^ n2707 ;
  assign n2737 = n2736 ^ n2730 ;
  assign n2738 = n2688 & ~n2737 ;
  assign n2774 = n945 ^ n579 ;
  assign n2775 = n2774 ^ n148 ;
  assign n2776 = n2775 ^ n720 ;
  assign n2771 = n1956 ^ n1355 ;
  assign n2772 = n2771 ^ n130 ;
  assign n2773 = n2772 ^ n513 ;
  assign n2777 = n2776 ^ n2773 ;
  assign n2768 = n636 ^ n417 ;
  assign n2769 = n2768 ^ n742 ;
  assign n2764 = n739 ^ n405 ;
  assign n2765 = n2764 ^ n689 ;
  assign n2766 = n2765 ^ n180 ;
  assign n2767 = n2766 ^ n1190 ;
  assign n2770 = n2769 ^ n2767 ;
  assign n2778 = n2777 ^ n2770 ;
  assign n2760 = n592 ^ n396 ;
  assign n2759 = n2320 ^ n1982 ;
  assign n2761 = n2760 ^ n2759 ;
  assign n2755 = n370 ^ n198 ;
  assign n2756 = n2755 ^ n88 ;
  assign n2753 = n321 ^ n104 ;
  assign n2754 = n2753 ^ n726 ;
  assign n2757 = n2756 ^ n2754 ;
  assign n2752 = n1317 ^ n270 ;
  assign n2758 = n2757 ^ n2752 ;
  assign n2762 = n2761 ^ n2758 ;
  assign n2748 = n1054 ^ n893 ;
  assign n2749 = n2748 ^ n1767 ;
  assign n2750 = n2749 ^ n1903 ;
  assign n2744 = n282 ^ n219 ;
  assign n2746 = n2745 ^ n2744 ;
  assign n2741 = n845 ^ n703 ;
  assign n2742 = n2741 ^ n391 ;
  assign n2739 = n2720 ^ n313 ;
  assign n2740 = n2739 ^ n667 ;
  assign n2743 = n2742 ^ n2740 ;
  assign n2747 = n2746 ^ n2743 ;
  assign n2751 = n2750 ^ n2747 ;
  assign n2763 = n2762 ^ n2751 ;
  assign n2779 = n2778 ^ n2763 ;
  assign n2830 = n797 ^ n522 ;
  assign n2831 = n2830 ^ n765 ;
  assign n2829 = n1001 ^ n392 ;
  assign n2832 = n2831 ^ n2829 ;
  assign n2827 = n1746 ^ n403 ;
  assign n2824 = n799 ^ n194 ;
  assign n2825 = n2824 ^ n1997 ;
  assign n2826 = n2825 ^ n1098 ;
  assign n2828 = n2827 ^ n2826 ;
  assign n2833 = n2832 ^ n2828 ;
  assign n2820 = n675 ^ n527 ;
  assign n2821 = n2820 ^ n1068 ;
  assign n2818 = n862 ^ n768 ;
  assign n2819 = n2818 ^ n2102 ;
  assign n2822 = n2821 ^ n2819 ;
  assign n2814 = n1148 ^ n559 ;
  assign n2815 = n2814 ^ n202 ;
  assign n2816 = n2815 ^ n1588 ;
  assign n2812 = n1197 ^ n360 ;
  assign n2809 = n737 ^ n143 ;
  assign n2810 = n2809 ^ n226 ;
  assign n2811 = n2810 ^ n856 ;
  assign n2813 = n2812 ^ n2811 ;
  assign n2817 = n2816 ^ n2813 ;
  assign n2823 = n2822 ^ n2817 ;
  assign n2834 = n2833 ^ n2823 ;
  assign n2805 = n1014 ^ n614 ;
  assign n2806 = n2805 ^ n1205 ;
  assign n2801 = n809 ^ n284 ;
  assign n2800 = n2659 ^ n1219 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2799 = n380 ^ n264 ;
  assign n2803 = n2802 ^ n2799 ;
  assign n2797 = ~x29 & n50 ;
  assign n2798 = n83 & n2797 ;
  assign n2804 = n2803 ^ n2798 ;
  assign n2807 = n2806 ^ n2804 ;
  assign n2794 = n1683 ^ n204 ;
  assign n2791 = n1074 ^ n362 ;
  assign n2792 = n2791 ^ n292 ;
  assign n2788 = n455 ^ n236 ;
  assign n2789 = n2788 ^ n409 ;
  assign n2790 = n2789 ^ n356 ;
  assign n2793 = n2792 ^ n2790 ;
  assign n2795 = n2794 ^ n2793 ;
  assign n2785 = n918 ^ n280 ;
  assign n2786 = n2785 ^ n585 ;
  assign n2782 = n1122 ^ n90 ;
  assign n2783 = n2782 ^ n401 ;
  assign n2780 = n982 ^ n782 ;
  assign n2781 = n2780 ^ n622 ;
  assign n2784 = n2783 ^ n2781 ;
  assign n2787 = n2786 ^ n2784 ;
  assign n2796 = n2795 ^ n2787 ;
  assign n2808 = n2807 ^ n2796 ;
  assign n2835 = n2834 ^ n2808 ;
  assign n2836 = ~n2779 & ~n2835 ;
  assign n2877 = n1967 ^ n1099 ;
  assign n2878 = n2877 ^ n1578 ;
  assign n2874 = n557 ^ n252 ;
  assign n2875 = n2874 ^ n793 ;
  assign n2872 = n1093 ^ n280 ;
  assign n2873 = n2872 ^ n728 ;
  assign n2876 = n2875 ^ n2873 ;
  assign n2879 = n2878 ^ n2876 ;
  assign n2869 = n2768 ^ n359 ;
  assign n2870 = n2869 ^ n518 ;
  assign n2868 = n765 ^ n456 ;
  assign n2871 = n2870 ^ n2868 ;
  assign n2880 = n2879 ^ n2871 ;
  assign n2864 = n667 ^ n506 ;
  assign n2865 = n2864 ^ n1746 ;
  assign n2863 = n1130 ^ n658 ;
  assign n2866 = n2865 ^ n2863 ;
  assign n2860 = n1927 ^ n1355 ;
  assign n2861 = n2860 ^ n673 ;
  assign n2858 = n898 ^ n351 ;
  assign n2856 = n547 ^ n303 ;
  assign n2857 = n2856 ^ n255 ;
  assign n2859 = n2858 ^ n2857 ;
  assign n2862 = n2861 ^ n2859 ;
  assign n2867 = n2866 ^ n2862 ;
  assign n2881 = n2880 ^ n2867 ;
  assign n2852 = n1543 ^ n455 ;
  assign n2853 = n2852 ^ n683 ;
  assign n2849 = n726 ^ n450 ;
  assign n2850 = n2849 ^ n500 ;
  assign n2848 = n662 ^ n216 ;
  assign n2851 = n2850 ^ n2848 ;
  assign n2854 = n2853 ^ n2851 ;
  assign n2845 = n809 ^ n425 ;
  assign n2846 = n2845 ^ n1237 ;
  assign n2843 = n779 ^ n720 ;
  assign n2840 = n272 ^ n222 ;
  assign n2839 = n764 ^ n762 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2837 = n291 ^ n249 ;
  assign n2838 = n2837 ^ n837 ;
  assign n2842 = n2841 ^ n2838 ;
  assign n2844 = n2843 ^ n2842 ;
  assign n2847 = n2846 ^ n2844 ;
  assign n2855 = n2854 ^ n2847 ;
  assign n2882 = n2881 ^ n2855 ;
  assign n2920 = n1683 ^ n1389 ;
  assign n2918 = n768 ^ n244 ;
  assign n2916 = n1182 ^ n296 ;
  assign n2917 = n2916 ^ n867 ;
  assign n2919 = n2918 ^ n2917 ;
  assign n2921 = n2920 ^ n2919 ;
  assign n2912 = n1054 ^ n400 ;
  assign n2913 = n2912 ^ n1772 ;
  assign n2910 = n772 ^ n370 ;
  assign n2911 = n2910 ^ n1149 ;
  assign n2914 = n2913 ^ n2911 ;
  assign n2907 = n239 ^ n161 ;
  assign n2908 = n2907 ^ n1129 ;
  assign n2909 = n2908 ^ n142 ;
  assign n2915 = n2914 ^ n2909 ;
  assign n2922 = n2921 ^ n2915 ;
  assign n2901 = n520 ^ n401 ;
  assign n2902 = n2901 ^ n109 ;
  assign n2903 = n2902 ^ n144 ;
  assign n2900 = n2899 ^ n799 ;
  assign n2904 = n2903 ^ n2900 ;
  assign n2905 = n2904 ^ n505 ;
  assign n2894 = n1194 ^ n804 ;
  assign n2895 = n2894 ^ n1176 ;
  assign n2896 = n2895 ^ n605 ;
  assign n2890 = n236 ^ n180 ;
  assign n2891 = n2890 ^ n266 ;
  assign n2889 = n2888 ^ n2670 ;
  assign n2892 = n2891 ^ n2889 ;
  assign n2886 = n2509 ^ n814 ;
  assign n2883 = n1956 ^ n230 ;
  assign n2884 = n2883 ^ n405 ;
  assign n2885 = n2884 ^ n313 ;
  assign n2887 = n2886 ^ n2885 ;
  assign n2893 = n2892 ^ n2887 ;
  assign n2897 = n2896 ^ n2893 ;
  assign n2898 = n2897 ^ n1127 ;
  assign n2906 = n2905 ^ n2898 ;
  assign n2923 = n2922 ^ n2906 ;
  assign n2924 = ~n2882 & ~n2923 ;
  assign n2952 = n1085 ^ n914 ;
  assign n2951 = n1099 ^ n845 ;
  assign n2953 = n2952 ^ n2951 ;
  assign n2949 = n2948 ^ n455 ;
  assign n2946 = n1381 ^ n429 ;
  assign n2947 = n2946 ^ n414 ;
  assign n2950 = n2949 ^ n2947 ;
  assign n2954 = n2953 ^ n2950 ;
  assign n2942 = n550 ^ n137 ;
  assign n2943 = n2942 ^ n2723 ;
  assign n2940 = n1555 ^ n359 ;
  assign n2941 = n2940 ^ n2451 ;
  assign n2944 = n2943 ^ n2941 ;
  assign n2937 = n810 ^ n541 ;
  assign n2938 = n2937 ^ n2667 ;
  assign n2935 = n1494 ^ n364 ;
  assign n2936 = n2935 ^ n2072 ;
  assign n2939 = n2938 ^ n2936 ;
  assign n2945 = n2944 ^ n2939 ;
  assign n2955 = n2954 ^ n2945 ;
  assign n2932 = n579 ^ n172 ;
  assign n2931 = n2760 ^ n129 ;
  assign n2933 = n2932 ^ n2931 ;
  assign n2928 = n2024 ^ n836 ;
  assign n2929 = n2928 ^ n2627 ;
  assign n2925 = n658 ^ n155 ;
  assign n2926 = n2925 ^ n856 ;
  assign n2927 = n2926 ^ n1399 ;
  assign n2930 = n2929 ^ n2927 ;
  assign n2934 = n2933 ^ n2930 ;
  assign n2956 = n2955 ^ n2934 ;
  assign n2957 = n2956 ^ n1316 ;
  assign n2958 = ~n1793 & ~n2957 ;
  assign n2979 = n2397 ^ n1783 ;
  assign n2975 = n1808 ^ n1085 ;
  assign n2974 = n1140 ^ n392 ;
  assign n2976 = n2975 ^ n2974 ;
  assign n2972 = n762 ^ n404 ;
  assign n2969 = n856 ^ n621 ;
  assign n2970 = n2969 ^ n572 ;
  assign n2968 = n1785 ^ n211 ;
  assign n2971 = n2970 ^ n2968 ;
  assign n2973 = n2972 ^ n2971 ;
  assign n2977 = n2976 ^ n2973 ;
  assign n2963 = n1093 ^ n1014 ;
  assign n2964 = n2963 ^ n527 ;
  assign n2962 = n417 ^ n260 ;
  assign n2965 = n2964 ^ n2962 ;
  assign n2960 = n773 ^ n178 ;
  assign n2959 = n2078 ^ n148 ;
  assign n2961 = n2960 ^ n2959 ;
  assign n2966 = n2965 ^ n2961 ;
  assign n2967 = n2966 ^ n2804 ;
  assign n2978 = n2977 ^ n2967 ;
  assign n2980 = n2979 ^ n2978 ;
  assign n3021 = n897 ^ n261 ;
  assign n3020 = n760 ^ n268 ;
  assign n3022 = n3021 ^ n3020 ;
  assign n3019 = n2928 ^ n2674 ;
  assign n3023 = n3022 ^ n3019 ;
  assign n3016 = n1780 ^ n1746 ;
  assign n3014 = n1756 ^ n250 ;
  assign n3011 = n607 ^ n291 ;
  assign n3012 = n3011 ^ n117 ;
  assign n3013 = n3012 ^ n413 ;
  assign n3015 = n3014 ^ n3013 ;
  assign n3017 = n3016 ^ n3015 ;
  assign n3006 = n78 ^ n69 ;
  assign n3007 = n3006 ^ n58 ;
  assign n3008 = n341 & n3007 ;
  assign n3009 = n3008 ^ n1099 ;
  assign n3010 = n3009 ^ n2810 ;
  assign n3018 = n3017 ^ n3010 ;
  assign n3024 = n3023 ^ n3018 ;
  assign n3002 = n1074 ^ n703 ;
  assign n3003 = n3002 ^ n245 ;
  assign n3001 = n2883 ^ n841 ;
  assign n3004 = n3003 ^ n3001 ;
  assign n2998 = n689 ^ n425 ;
  assign n2997 = n212 ^ n104 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n2995 = n2610 ^ n513 ;
  assign n2994 = n1652 ^ n149 ;
  assign n2996 = n2995 ^ n2994 ;
  assign n3000 = n2999 ^ n2996 ;
  assign n3005 = n3004 ^ n3000 ;
  assign n3025 = n3024 ^ n3005 ;
  assign n2990 = n2575 ^ n1070 ;
  assign n2989 = n2988 ^ n220 ;
  assign n2991 = n2990 ^ n2989 ;
  assign n2984 = n2890 ^ n1649 ;
  assign n2985 = n2984 ^ n2303 ;
  assign n2982 = n589 ^ n249 ;
  assign n2981 = n2249 ^ n1826 ;
  assign n2983 = n2982 ^ n2981 ;
  assign n2986 = n2985 ^ n2983 ;
  assign n2992 = n2991 ^ n2986 ;
  assign n2993 = n2992 ^ n2064 ;
  assign n3026 = n3025 ^ n2993 ;
  assign n3027 = ~n2980 & ~n3026 ;
  assign n3059 = n554 ^ n414 ;
  assign n3057 = n2771 ^ n122 ;
  assign n3058 = n3057 ^ n571 ;
  assign n3060 = n3059 ^ n3058 ;
  assign n3055 = n1658 ^ n178 ;
  assign n598 = n86 & n337 ;
  assign n3053 = n899 ^ n598 ;
  assign n3052 = n2538 ^ n305 ;
  assign n3054 = n3053 ^ n3052 ;
  assign n3056 = n3055 ^ n3054 ;
  assign n3061 = n3060 ^ n3056 ;
  assign n3046 = n797 ^ n261 ;
  assign n3047 = n3046 ^ n518 ;
  assign n3048 = n3047 ^ n882 ;
  assign n3045 = n2228 ^ n513 ;
  assign n3049 = n3048 ^ n3045 ;
  assign n3041 = n186 ^ n172 ;
  assign n3042 = n3041 ^ n745 ;
  assign n3043 = n3042 ^ n689 ;
  assign n4228 = n667 ^ n602 ;
  assign n3039 = n4228 ^ n1330 ;
  assign n3040 = n3039 ^ n205 ;
  assign n3044 = n3043 ^ n3040 ;
  assign n3050 = n3049 ^ n3044 ;
  assign n3034 = n953 ^ n932 ;
  assign n3035 = n3034 ^ n2435 ;
  assign n3031 = n625 ^ n533 ;
  assign n3030 = n360 ^ n258 ;
  assign n3032 = n3031 ^ n3030 ;
  assign n3028 = n739 ^ n363 ;
  assign n3029 = n3028 ^ n291 ;
  assign n3033 = n3032 ^ n3029 ;
  assign n3036 = n3035 ^ n3033 ;
  assign n3037 = n3036 ^ n777 ;
  assign n3051 = n3050 ^ n3037 ;
  assign n3062 = n3061 ^ n3051 ;
  assign n3093 = n819 ^ n356 ;
  assign n3094 = n3093 ^ n624 ;
  assign n3091 = n1177 ^ n1037 ;
  assign n3092 = n3091 ^ n641 ;
  assign n3095 = n3094 ^ n3092 ;
  assign n3088 = n1549 ^ n397 ;
  assign n3086 = n196 ^ n148 ;
  assign n3087 = n3086 ^ n266 ;
  assign n3089 = n3088 ^ n3087 ;
  assign n3084 = n1504 ^ n622 ;
  assign n3082 = n2907 ^ n282 ;
  assign n3083 = n3082 ^ n211 ;
  assign n3085 = n3084 ^ n3083 ;
  assign n3090 = n3089 ^ n3085 ;
  assign n3096 = n3095 ^ n3090 ;
  assign n3078 = n1001 ^ n175 ;
  assign n3079 = n3078 ^ n880 ;
  assign n3076 = n2179 ^ n490 ;
  assign n3075 = n764 ^ n124 ;
  assign n3077 = n3076 ^ n3075 ;
  assign n3080 = n3079 ^ n3077 ;
  assign n3072 = n1129 ^ n540 ;
  assign n3070 = n1197 ^ n394 ;
  assign n3071 = n3070 ^ n156 ;
  assign n3073 = n3072 ^ n3071 ;
  assign n3066 = n1029 ^ n785 ;
  assign n3067 = n3066 ^ n280 ;
  assign n3068 = n3067 ^ n183 ;
  assign n3063 = n559 ^ n90 ;
  assign n3064 = n3063 ^ n137 ;
  assign n3065 = n3064 ^ n483 ;
  assign n3069 = n3068 ^ n3065 ;
  assign n3074 = n3073 ^ n3069 ;
  assign n3081 = n3080 ^ n3074 ;
  assign n3097 = n3096 ^ n3081 ;
  assign n3098 = n3097 ^ n2993 ;
  assign n3099 = ~n3062 & ~n3098 ;
  assign n3100 = ~n3027 & ~n3099 ;
  assign n3101 = n2958 & ~n3100 ;
  assign n3102 = ~n2924 & ~n3101 ;
  assign n3129 = n1408 ^ n122 ;
  assign n3130 = n3129 ^ n250 ;
  assign n3127 = n1029 ^ n313 ;
  assign n3128 = n3127 ^ n782 ;
  assign n3131 = n3130 ^ n3128 ;
  assign n3132 = n3131 ^ n406 ;
  assign n3125 = n47 & ~n12860 ;
  assign n3121 = n433 ^ n183 ;
  assign n3122 = n3121 ^ n550 ;
  assign n3119 = n1249 ^ n867 ;
  assign n3120 = n3119 ^ n499 ;
  assign n3123 = n3122 ^ n3120 ;
  assign n3115 = n677 ^ n197 ;
  assign n3116 = n3115 ^ n292 ;
  assign n3118 = n3117 ^ n3116 ;
  assign n3124 = n3123 ^ n3118 ;
  assign n3126 = n3125 ^ n3124 ;
  assign n3133 = n3132 ^ n3126 ;
  assign n3111 = n258 ^ n242 ;
  assign n3112 = n3111 ^ n857 ;
  assign n3110 = n2132 ^ n863 ;
  assign n3113 = n3112 ^ n3110 ;
  assign n3107 = n790 ^ n401 ;
  assign n3106 = n1488 ^ n932 ;
  assign n3108 = n3107 ^ n3106 ;
  assign n3103 = n1050 ^ n450 ;
  assign n3104 = n3103 ^ n393 ;
  assign n3105 = n3104 ^ n928 ;
  assign n3109 = n3108 ^ n3105 ;
  assign n3114 = n3113 ^ n3109 ;
  assign n3134 = n3133 ^ n3114 ;
  assign n3135 = n3134 ^ n2881 ;
  assign n3149 = n2607 ^ n577 ;
  assign n3144 = n661 ^ n217 ;
  assign n3145 = n3144 ^ n2451 ;
  assign n3146 = n3145 ^ n2069 ;
  assign n3141 = n514 ^ n376 ;
  assign n3142 = n3141 ^ n540 ;
  assign n3139 = n365 ^ n284 ;
  assign n3140 = n3139 ^ n416 ;
  assign n3143 = n3142 ^ n3140 ;
  assign n3147 = n3146 ^ n3143 ;
  assign n3136 = n779 ^ n214 ;
  assign n3137 = n3136 ^ n797 ;
  assign n3138 = n3137 ^ n1161 ;
  assign n3148 = n3147 ^ n3138 ;
  assign n3150 = n3149 ^ n3148 ;
  assign n3151 = ~n3135 & ~n3150 ;
  assign n3152 = ~n3102 & n3151 ;
  assign n3153 = ~n2836 & ~n3152 ;
  assign n3154 = n2738 & ~n3153 ;
  assign n3155 = ~n2646 & ~n3154 ;
  assign n3187 = n1667 ^ n638 ;
  assign n3188 = n3187 ^ n2972 ;
  assign n3182 = n1970 ^ n836 ;
  assign n3183 = n3182 ^ n175 ;
  assign n3181 = n1982 ^ n526 ;
  assign n3184 = n3183 ^ n3181 ;
  assign n3185 = n3184 ^ n560 ;
  assign n3186 = n3185 ^ n1099 ;
  assign n3189 = n3188 ^ n3186 ;
  assign n3177 = n675 ^ n375 ;
  assign n3176 = n1308 ^ n361 ;
  assign n3178 = n3177 ^ n3176 ;
  assign n3174 = n1521 ^ n1074 ;
  assign n3175 = n3174 ^ n1728 ;
  assign n3179 = n3178 ^ n3175 ;
  assign n3180 = n3179 ^ n3126 ;
  assign n3190 = n3189 ^ n3180 ;
  assign n3171 = n773 ^ n282 ;
  assign n3172 = n3171 ^ n2236 ;
  assign n3167 = n624 ^ n305 ;
  assign n3165 = n3111 ^ n298 ;
  assign n3166 = n3165 ^ n1494 ;
  assign n3168 = n3167 ^ n3166 ;
  assign n3169 = n3168 ^ n1962 ;
  assign n3161 = n1135 ^ n116 ;
  assign n3162 = n3161 ^ n394 ;
  assign n3159 = n614 ^ n285 ;
  assign n3160 = n3159 ^ n249 ;
  assign n3163 = n3162 ^ n3160 ;
  assign n3156 = n1576 ^ n206 ;
  assign n3157 = n3156 ^ n1159 ;
  assign n3158 = n3157 ^ n1435 ;
  assign n3164 = n3163 ^ n3158 ;
  assign n3170 = n3169 ^ n3164 ;
  assign n3173 = n3172 ^ n3170 ;
  assign n3191 = n3190 ^ n3173 ;
  assign n3223 = n4228 ^ n2814 ;
  assign n3219 = n747 ^ n216 ;
  assign n3220 = n3219 ^ n264 ;
  assign n3217 = n2654 ^ n1116 ;
  assign n3218 = n3217 ^ n236 ;
  assign n3221 = n3220 ^ n3218 ;
  assign n3215 = n635 ^ n291 ;
  assign n3213 = n1732 ^ n772 ;
  assign n3212 = n589 ^ n255 ;
  assign n3214 = n3213 ^ n3212 ;
  assign n3216 = n3215 ^ n3214 ;
  assign n3222 = n3221 ^ n3216 ;
  assign n3224 = n3223 ^ n3222 ;
  assign n3225 = n3224 ^ n2374 ;
  assign n3207 = n810 ^ n229 ;
  assign n3206 = n583 ^ n362 ;
  assign n3208 = n3207 ^ n3206 ;
  assign n3204 = n641 ^ n237 ;
  assign n3203 = n1197 ^ n571 ;
  assign n3205 = n3204 ^ n3203 ;
  assign n3209 = n3208 ^ n3205 ;
  assign n3201 = n2774 ^ n1577 ;
  assign n3202 = n3201 ^ n2022 ;
  assign n3210 = n3209 ^ n3202 ;
  assign n3199 = n2614 ^ n2207 ;
  assign n3197 = n1007 ^ n872 ;
  assign n3194 = n814 ^ n678 ;
  assign n3195 = n3194 ^ n259 ;
  assign n3192 = n856 ^ n672 ;
  assign n3193 = n3192 ^ n2451 ;
  assign n3196 = n3195 ^ n3193 ;
  assign n3198 = n3197 ^ n3196 ;
  assign n3200 = n3199 ^ n3198 ;
  assign n3211 = n3210 ^ n3200 ;
  assign n3226 = n3225 ^ n3211 ;
  assign n3227 = ~n3191 & ~n3226 ;
  assign n3228 = ~n3155 & n3227 ;
  assign n3229 = ~n2609 & ~n3228 ;
  assign n3230 = n2554 & ~n3229 ;
  assign n3231 = ~n2486 & ~n3230 ;
  assign n3232 = n2449 & ~n3231 ;
  assign n3233 = ~n2364 & ~n3232 ;
  assign n3234 = n2268 & ~n3233 ;
  assign n3235 = ~n2185 & ~n3234 ;
  assign n3236 = n2096 & ~n3235 ;
  assign n3237 = ~n1994 & ~n3236 ;
  assign n3238 = n3237 ^ n1795 ;
  assign n1995 = n1994 ^ n1795 ;
  assign n3239 = n3238 ^ n1995 ;
  assign n3242 = ~n1871 & ~n3239 ;
  assign n3243 = n3242 ^ n1995 ;
  assign n3244 = ~n1873 & n3243 ;
  assign n3349 = n3154 ^ n3153 ;
  assign n3277 = n3119 ^ n760 ;
  assign n3276 = n1731 ^ n810 ;
  assign n3278 = n3277 ^ n3276 ;
  assign n3280 = n3279 ^ n3278 ;
  assign n3273 = n893 ^ n455 ;
  assign n3274 = n3273 ^ n558 ;
  assign n3271 = n1282 ^ n505 ;
  assign n3272 = n3271 ^ n725 ;
  assign n3275 = n3274 ^ n3272 ;
  assign n3281 = n3280 ^ n3275 ;
  assign n3267 = n1396 ^ n400 ;
  assign n3268 = n3267 ^ n3128 ;
  assign n3265 = n2901 ^ n203 ;
  assign n3263 = n1036 ^ n283 ;
  assign n3264 = n3263 ^ n579 ;
  assign n3266 = n3265 ^ n3264 ;
  assign n3269 = n3268 ^ n3266 ;
  assign n3259 = n363 ^ n124 ;
  assign n3260 = n3259 ^ n762 ;
  assign n3261 = n3260 ^ n1471 ;
  assign n3256 = n1512 ^ n87 ;
  assign n3253 = n613 ^ n483 ;
  assign n3254 = n3253 ^ n309 ;
  assign n3255 = n3254 ^ n745 ;
  assign n3257 = n3256 ^ n3255 ;
  assign n3251 = n379 ^ n298 ;
  assign n3250 = n2442 ^ n1986 ;
  assign n3252 = n3251 ^ n3250 ;
  assign n3258 = n3257 ^ n3252 ;
  assign n3262 = n3261 ^ n3258 ;
  assign n3270 = n3269 ^ n3262 ;
  assign n3282 = n3281 ^ n3270 ;
  assign n3332 = n3194 ^ n2693 ;
  assign n3331 = n496 ^ n255 ;
  assign n3333 = n3332 ^ n3331 ;
  assign n3328 = n418 ^ n361 ;
  assign n3326 = n407 ^ n176 ;
  assign n3327 = n3326 ^ n264 ;
  assign n3329 = n3328 ^ n3327 ;
  assign n3323 = n732 ^ n183 ;
  assign n3324 = n3323 ^ n818 ;
  assign n3322 = n3321 ^ n853 ;
  assign n3325 = n3324 ^ n3322 ;
  assign n3330 = n3329 ^ n3325 ;
  assign n3334 = n3333 ^ n3330 ;
  assign n3318 = n1121 ^ n104 ;
  assign n3316 = n2358 ^ n793 ;
  assign n3317 = n3316 ^ n1322 ;
  assign n3319 = n3318 ^ n3317 ;
  assign n3313 = n2837 ^ n1588 ;
  assign n3312 = n2228 ^ n1339 ;
  assign n3314 = n3313 ^ n3312 ;
  assign n3310 = n547 ^ n190 ;
  assign n3307 = n2016 ^ n394 ;
  assign n3308 = n3307 ^ n259 ;
  assign n3309 = n3308 ^ n161 ;
  assign n3311 = n3310 ^ n3309 ;
  assign n3315 = n3314 ^ n3311 ;
  assign n3320 = n3319 ^ n3315 ;
  assign n3335 = n3334 ^ n3320 ;
  assign n3303 = n983 ^ n201 ;
  assign n3302 = n2662 ^ n1906 ;
  assign n3304 = n3303 ^ n3302 ;
  assign n3301 = n2848 ^ n1560 ;
  assign n3305 = n3304 ^ n3301 ;
  assign n3298 = n2785 ^ n785 ;
  assign n3296 = n2233 ^ n961 ;
  assign n3297 = n3296 ^ n305 ;
  assign n3299 = n3298 ^ n3297 ;
  assign n3292 = n521 ^ n178 ;
  assign n3291 = n405 ^ n181 ;
  assign n3293 = n3292 ^ n3291 ;
  assign n3289 = n585 ^ n97 ;
  assign n3290 = n3289 ^ n673 ;
  assign n3294 = n3293 ^ n3290 ;
  assign n3286 = n351 ^ n200 ;
  assign n3285 = n497 ^ n245 ;
  assign n3287 = n3286 ^ n3285 ;
  assign n3283 = n726 ^ n226 ;
  assign n3284 = n3283 ^ n129 ;
  assign n3288 = n3287 ^ n3284 ;
  assign n3295 = n3294 ^ n3288 ;
  assign n3300 = n3299 ^ n3295 ;
  assign n3306 = n3305 ^ n3300 ;
  assign n3336 = n3335 ^ n3306 ;
  assign n3337 = ~n3282 & ~n3336 ;
  assign n3338 = n3027 & n3337 ;
  assign n3339 = n3338 ^ n3337 ;
  assign n3340 = n3339 ^ n3027 ;
  assign n3341 = n3099 & n3340 ;
  assign n3342 = ~n2958 & ~n3341 ;
  assign n3343 = n2924 & ~n3342 ;
  assign n3344 = ~n3152 & ~n3343 ;
  assign n3345 = n3344 ^ n3151 ;
  assign n3346 = n2836 & n3345 ;
  assign n3347 = n3346 ^ n3152 ;
  assign n3348 = ~n2738 & ~n3347 ;
  assign n3350 = n3349 ^ n3348 ;
  assign n3351 = n2646 & n3350 ;
  assign n3352 = ~n3227 & ~n3351 ;
  assign n3353 = n2609 & ~n3352 ;
  assign n3354 = ~n2554 & ~n3353 ;
  assign n3355 = n2486 & ~n3354 ;
  assign n3356 = ~n2449 & ~n3355 ;
  assign n3357 = n2364 & ~n3356 ;
  assign n3358 = ~n2268 & ~n3357 ;
  assign n3359 = n2185 & ~n3358 ;
  assign n3360 = ~n2096 & ~n3359 ;
  assign n3363 = n3244 & n3360 ;
  assign n3364 = ~n1631 & n3363 ;
  assign n3365 = n3364 ^ n1631 ;
  assign n3245 = n3244 ^ n1873 ;
  assign n3246 = n3245 ^ n1631 ;
  assign n3366 = n3365 ^ n3246 ;
  assign n3367 = n1872 & ~n3366 ;
  assign n3368 = n3367 ^ n1871 ;
  assign n3369 = ~n1715 & n3368 ;
  assign n3372 = n1433 & n1703 ;
  assign n3370 = n1351 & n1631 ;
  assign n3371 = n1540 & n3370 ;
  assign n3373 = n3372 ^ n3371 ;
  assign n3374 = n3369 & n3373 ;
  assign n3375 = n3374 ^ n1715 ;
  assign n3377 = ~n1540 & ~n3375 ;
  assign n3380 = n1214 & ~n3377 ;
  assign n3376 = n3375 ^ n1540 ;
  assign n3378 = n3377 ^ n3376 ;
  assign n3379 = ~n1214 & n3378 ;
  assign n3381 = n3380 ^ n3379 ;
  assign n3382 = n3380 ^ n1109 ;
  assign n3383 = n3382 ^ n3380 ;
  assign n3384 = n3381 & ~n3383 ;
  assign n3385 = n3384 ^ n3380 ;
  assign n3386 = n1111 & ~n3385 ;
  assign n3387 = n3386 ^ n1109 ;
  assign n3388 = n3387 ^ n824 ;
  assign n3474 = n3473 ^ n824 ;
  assign n3475 = ~n3388 & n3474 ;
  assign n3491 = n3473 & ~n3475 ;
  assign n3492 = n3491 ^ n3475 ;
  assign n3493 = n649 & n3492 ;
  assign n3494 = ~n317 & ~n3493 ;
  assign n3495 = n445 & ~n3494 ;
  assign n480 = ~x26 & n51 ;
  assign n481 = ~n165 & n480 ;
  assign n482 = n481 ^ n254 ;
  assign n484 = n483 ^ n482 ;
  assign n474 = n473 ^ n399 ;
  assign n475 = n474 ^ n414 ;
  assign n476 = ~n460 & ~n475 ;
  assign n449 = n448 ^ n295 ;
  assign n477 = n476 ^ n449 ;
  assign n479 = n478 ^ n477 ;
  assign n485 = n484 ^ n479 ;
  assign n3496 = ~n649 & ~n3491 ;
  assign n3497 = n317 & ~n3496 ;
  assign n3498 = ~n445 & ~n3497 ;
  assign n3920 = n485 & ~n3498 ;
  assign n3921 = ~n3495 & ~n3920 ;
  assign n3922 = n3921 ^ n3920 ;
  assign n3923 = n3922 ^ n485 ;
  assign n3924 = n3923 ^ n3920 ;
  assign n3941 = n478 ^ n441 ;
  assign n3933 = n111 ^ n36 ;
  assign n3934 = n3933 ^ n2731 ;
  assign n3935 = n45 & n3934 ;
  assign n3936 = n3935 ^ n3326 ;
  assign n3937 = n3936 ^ n238 ;
  assign n3932 = n3925 ^ n2764 ;
  assign n3938 = n3937 ^ n3932 ;
  assign n3939 = n3931 & ~n3938 ;
  assign n3940 = n3939 ^ n1074 ;
  assign n3942 = n3941 ^ n3940 ;
  assign n3943 = n3942 ^ n482 ;
  assign n4514 = n3924 & n3943 ;
  assign n4515 = n4514 ^ n3920 ;
  assign n12683 = n3520 & n4515 ;
  assign n12684 = n12683 ^ n3943 ;
  assign n12685 = x31 & ~n12684 ;
  assign n12744 = n12689 ^ n12685 ;
  assign n12745 = ~n12700 & n12744 ;
  assign n12746 = n12745 ^ n12699 ;
  assign n12701 = n12700 ^ n12685 ;
  assign n830 = n829 ^ x29 ;
  assign n828 = x29 & n827 ;
  assign n831 = n830 ^ n828 ;
  assign n12584 = n831 & ~n3943 ;
  assign n3720 = n35 ^ x31 ;
  assign n3721 = ~n3520 & n3720 ;
  assign n3513 = ~x31 & n33 ;
  assign n3514 = n3513 ^ x31 ;
  assign n3722 = n3721 ^ n3514 ;
  assign n24214 = x31 & ~n3722 ;
  assign n3724 = n24214 ^ n35 ;
  assign n3732 = n3724 ^ n33 ;
  assign n3733 = n3732 ^ n3513 ;
  assign n12580 = ~n445 & ~n3733 ;
  assign n12579 = ~n317 & n24214 ;
  assign n12581 = n12580 ^ n12579 ;
  assign n3499 = n3498 ^ n3495 ;
  assign n12576 = x31 & ~n3499 ;
  assign n12577 = n12576 ^ n485 ;
  assign n12578 = n3520 & ~n12577 ;
  assign n12582 = n12581 ^ n12578 ;
  assign n12583 = n12582 ^ x29 ;
  assign n12585 = n12584 ^ n12583 ;
  assign n12055 = n728 ^ n682 ;
  assign n12053 = n636 ^ n100 ;
  assign n6208 = n1116 ^ n971 ;
  assign n6209 = n6208 ^ n1122 ;
  assign n12054 = n12053 ^ n6209 ;
  assign n12056 = n12055 ^ n12054 ;
  assign n5572 = n541 ^ n197 ;
  assign n5573 = n5572 ^ n244 ;
  assign n5570 = n2190 ^ n359 ;
  assign n5571 = n5570 ^ n726 ;
  assign n5574 = n5573 ^ n5571 ;
  assign n5575 = n5574 ^ n3307 ;
  assign n12057 = n12056 ^ n5575 ;
  assign n5048 = n856 ^ n141 ;
  assign n12049 = n5048 ^ n1184 ;
  assign n12048 = n1898 ^ n791 ;
  assign n12050 = n12049 ^ n12048 ;
  assign n12046 = n742 ^ n678 ;
  assign n3631 = n2035 ^ n190 ;
  assign n12045 = n3631 ^ n237 ;
  assign n12047 = n12046 ^ n12045 ;
  assign n12051 = n12050 ^ n12047 ;
  assign n12052 = n12051 ^ n864 ;
  assign n12058 = n12057 ^ n12052 ;
  assign n12040 = n764 ^ n612 ;
  assign n12039 = n623 ^ n221 ;
  assign n12041 = n12040 ^ n12039 ;
  assign n12037 = n4228 ^ n751 ;
  assign n12035 = n697 ^ n407 ;
  assign n12036 = n12035 ^ n658 ;
  assign n12038 = n12037 ^ n12036 ;
  assign n12042 = n12041 ^ n12038 ;
  assign n4242 = n848 ^ n192 ;
  assign n12032 = n4242 ^ n230 ;
  assign n4244 = n918 ^ n496 ;
  assign n5567 = n4244 ^ n1772 ;
  assign n12033 = n12032 ^ n5567 ;
  assign n12030 = n2178 ^ n673 ;
  assign n12029 = n3103 ^ n737 ;
  assign n12031 = n12030 ^ n12029 ;
  assign n12034 = n12033 ^ n12031 ;
  assign n12043 = n12042 ^ n12034 ;
  assign n4804 = n380 ^ n250 ;
  assign n12025 = n4804 ^ n518 ;
  assign n12024 = n983 ^ n499 ;
  assign n12026 = n12025 ^ n12024 ;
  assign n12022 = n1621 ^ n196 ;
  assign n12021 = n753 ^ n252 ;
  assign n12023 = n12022 ^ n12021 ;
  assign n12027 = n12026 ^ n12023 ;
  assign n4017 = n2764 ^ n88 ;
  assign n4018 = n4017 ^ n273 ;
  assign n4019 = n4018 ^ n779 ;
  assign n12028 = n12027 ^ n4019 ;
  assign n12044 = n12043 ^ n12028 ;
  assign n12059 = n12058 ^ n12044 ;
  assign n12060 = ~n3282 & ~n12059 ;
  assign n12061 = n12060 ^ x26 ;
  assign n11830 = n401 ^ n360 ;
  assign n11831 = n11830 ^ n375 ;
  assign n11832 = n11831 ^ n3323 ;
  assign n11828 = n881 ^ n149 ;
  assign n11829 = n11828 ^ n144 ;
  assign n11833 = n11832 ^ n11829 ;
  assign n11825 = n1135 ^ n894 ;
  assign n11823 = n737 ^ n216 ;
  assign n11824 = n11823 ^ n1394 ;
  assign n11826 = n11825 ^ n11824 ;
  assign n11821 = n3086 ^ n2745 ;
  assign n11820 = n2451 ^ n418 ;
  assign n11822 = n11821 ^ n11820 ;
  assign n11827 = n11826 ^ n11822 ;
  assign n11834 = n11833 ^ n11827 ;
  assign n11816 = n1159 ^ n743 ;
  assign n11817 = n11816 ^ n3001 ;
  assign n4785 = n882 ^ n521 ;
  assign n5565 = n4785 ^ n660 ;
  assign n11818 = n11817 ^ n5565 ;
  assign n5605 = n785 ^ n376 ;
  assign n5606 = n5605 ^ n2276 ;
  assign n5607 = n5606 ^ n2262 ;
  assign n5602 = n1437 ^ n356 ;
  assign n5603 = n5602 ^ n520 ;
  assign n5600 = n1219 ^ n1094 ;
  assign n5601 = n5600 ^ n682 ;
  assign n5604 = n5603 ^ n5601 ;
  assign n5608 = n5607 ^ n5604 ;
  assign n11819 = n11818 ^ n5608 ;
  assign n11835 = n11834 ^ n11819 ;
  assign n5369 = n625 ^ n429 ;
  assign n5370 = n5369 ^ n1243 ;
  assign n5371 = n5370 ^ n1835 ;
  assign n5367 = n3192 ^ n635 ;
  assign n5364 = n772 ^ n190 ;
  assign n5365 = n5364 ^ n180 ;
  assign n5366 = n5365 ^ n413 ;
  assign n5368 = n5367 ^ n5366 ;
  assign n5372 = n5371 ^ n5368 ;
  assign n3563 = n624 ^ n204 ;
  assign n5359 = n3563 ^ n178 ;
  assign n5360 = n5359 ^ n1600 ;
  assign n3851 = n391 ^ n285 ;
  assign n5358 = n3851 ^ n1206 ;
  assign n5361 = n5360 ^ n5358 ;
  assign n5354 = n570 ^ n499 ;
  assign n5355 = n5354 ^ n527 ;
  assign n5356 = n5355 ^ n1906 ;
  assign n5352 = n1051 ^ n370 ;
  assign n5353 = n5352 ^ n677 ;
  assign n5357 = n5356 ^ n5353 ;
  assign n5362 = n5361 ^ n5357 ;
  assign n5350 = n3431 ^ n1366 ;
  assign n5349 = n2473 ^ n155 ;
  assign n5351 = n5350 ^ n5349 ;
  assign n5363 = n5362 ^ n5351 ;
  assign n5373 = n5372 ^ n5363 ;
  assign n11836 = n11835 ^ n5373 ;
  assign n11837 = ~n2122 & ~n11836 ;
  assign n12342 = n12060 ^ n11837 ;
  assign n12343 = n12061 & ~n12342 ;
  assign n12344 = n12343 ^ x26 ;
  assign n4192 = n2584 ^ n1206 ;
  assign n4188 = n570 ^ n362 ;
  assign n4189 = n4188 ^ n122 ;
  assign n4190 = n4189 ^ n954 ;
  assign n4191 = n4190 ^ n1487 ;
  assign n4193 = n4192 ^ n4191 ;
  assign n3596 = n672 ^ n313 ;
  assign n4186 = n4185 ^ n3596 ;
  assign n4183 = n728 ^ n703 ;
  assign n4184 = n4183 ^ n1297 ;
  assign n4187 = n4186 ^ n4184 ;
  assign n4194 = n4193 ^ n4187 ;
  assign n4181 = n1605 ^ n1029 ;
  assign n4180 = n3168 ^ n2826 ;
  assign n4182 = n4181 ^ n4180 ;
  assign n4195 = n4194 ^ n4182 ;
  assign n4196 = n4195 ^ n2719 ;
  assign n12336 = n857 ^ n429 ;
  assign n12337 = n12336 ^ n1738 ;
  assign n5246 = n1608 ^ n497 ;
  assign n12338 = n12337 ^ n5246 ;
  assign n12333 = n1001 ^ n151 ;
  assign n5631 = n500 ^ n178 ;
  assign n5632 = n5631 ^ n689 ;
  assign n12331 = n5632 ^ n772 ;
  assign n12332 = n12331 ^ n809 ;
  assign n12334 = n12333 ^ n12332 ;
  assign n12329 = n972 ^ n431 ;
  assign n3773 = n273 ^ n175 ;
  assign n12328 = n3773 ^ n3432 ;
  assign n12330 = n12329 ^ n12328 ;
  assign n12335 = n12334 ^ n12330 ;
  assign n12339 = n12338 ^ n12335 ;
  assign n5103 = n725 ^ n229 ;
  assign n12323 = n5103 ^ n2748 ;
  assign n12321 = n1148 ^ n745 ;
  assign n6333 = n677 ^ n155 ;
  assign n12322 = n12321 ^ n6333 ;
  assign n12324 = n12323 ^ n12322 ;
  assign n6419 = n2282 ^ n269 ;
  assign n12320 = n6419 ^ n495 ;
  assign n12325 = n12324 ^ n12320 ;
  assign n12316 = n1041 ^ n450 ;
  assign n12317 = n12316 ^ n201 ;
  assign n12314 = n2442 ^ n378 ;
  assign n12315 = n12314 ^ n261 ;
  assign n12318 = n12317 ^ n12315 ;
  assign n12319 = n12318 ^ n629 ;
  assign n12326 = n12325 ^ n12319 ;
  assign n12308 = n521 ^ n376 ;
  assign n12309 = n12308 ^ n285 ;
  assign n12310 = n12309 ^ n1280 ;
  assign n12307 = n1813 ^ n506 ;
  assign n12311 = n12310 ^ n12307 ;
  assign n12305 = n845 ^ n661 ;
  assign n3705 = n1389 ^ n804 ;
  assign n12303 = n3705 ^ n483 ;
  assign n12304 = n12303 ^ n303 ;
  assign n12306 = n12305 ^ n12304 ;
  assign n12312 = n12311 ^ n12306 ;
  assign n12313 = n12312 ^ n929 ;
  assign n12327 = n12326 ^ n12313 ;
  assign n12340 = n12339 ^ n12327 ;
  assign n12341 = ~n4196 & ~n12340 ;
  assign n12345 = n12344 ^ n12341 ;
  assign n3725 = n3724 ^ x31 ;
  assign n3726 = n3725 ^ n3513 ;
  assign n12300 = ~n445 & n3726 ;
  assign n12299 = ~n317 & ~n3724 ;
  assign n12301 = n12300 ^ n12299 ;
  assign n4072 = n3497 ^ n3494 ;
  assign n4073 = n4072 ^ n445 ;
  assign n12290 = n4073 ^ n649 ;
  assign n12289 = n4073 ^ n317 ;
  assign n12291 = n12290 ^ n12289 ;
  assign n12294 = ~x30 & n12291 ;
  assign n12295 = n12294 ^ n12290 ;
  assign n12296 = ~n3520 & ~n12295 ;
  assign n12297 = n12296 ^ n4073 ;
  assign n12298 = x31 & n12297 ;
  assign n12302 = n12301 ^ n12298 ;
  assign n12537 = n12344 ^ n12302 ;
  assign n12538 = ~n12345 & n12537 ;
  assign n12573 = n12572 ^ n12538 ;
  assign n12615 = n12582 ^ n12573 ;
  assign n12616 = n12585 & ~n12615 ;
  assign n12617 = n12616 ^ n12582 ;
  assign n12618 = n12572 ^ n12302 ;
  assign n12619 = n12538 & n12618 ;
  assign n12620 = n12619 ^ n12572 ;
  assign n12666 = n12617 & n12620 ;
  assign n12725 = n12701 ^ n12666 ;
  assign n12350 = ~n485 & n831 ;
  assign n3484 = n827 ^ n650 ;
  assign n12348 = n3484 & ~n3943 ;
  assign n12346 = n12345 ^ n12302 ;
  assign n12347 = n12346 ^ x29 ;
  assign n12349 = n12348 ^ n12347 ;
  assign n12351 = n12350 ^ n12349 ;
  assign n4536 = x29 ^ x28 ;
  assign n655 = n654 ^ n650 ;
  assign n3479 = n655 ^ x29 ;
  assign n3480 = n4536 ^ n3479 ;
  assign n651 = x29 & ~n650 ;
  assign n28635 = x29 & ~n651 ;
  assign n3477 = n28635 ^ x28 ;
  assign n3481 = n3480 ^ n3477 ;
  assign n12288 = n3481 & n4515 ;
  assign n12352 = n12351 ^ n12288 ;
  assign n12586 = n12585 ^ n12573 ;
  assign n12353 = n12061 ^ n11837 ;
  assign n12019 = ~n35 & ~n649 ;
  assign n12015 = x31 & ~n3520 ;
  assign n3955 = n3496 ^ n3493 ;
  assign n3956 = n3955 ^ n317 ;
  assign n12016 = n3956 ^ n649 ;
  assign n12017 = ~n12015 & ~n12016 ;
  assign n11938 = ~n35 & ~n3473 ;
  assign n12006 = n11938 ^ n3955 ;
  assign n12007 = n12006 ^ n317 ;
  assign n12008 = n12007 ^ n12006 ;
  assign n12009 = n12006 ^ n3726 ;
  assign n12010 = n12009 ^ n12006 ;
  assign n12011 = n12008 & ~n12010 ;
  assign n12012 = n12011 ^ n12006 ;
  assign n12013 = ~x31 & n12012 ;
  assign n12004 = n3726 ^ n649 ;
  assign n12005 = n12004 ^ n11938 ;
  assign n12014 = n12013 ^ n12005 ;
  assign n12018 = n12017 ^ n12014 ;
  assign n12020 = n12019 ^ n12018 ;
  assign n12354 = n12353 ^ n12020 ;
  assign n12355 = n12020 ^ n11837 ;
  assign n11940 = n11938 ^ n3475 ;
  assign n3476 = n3475 ^ n649 ;
  assign n11930 = n3476 ^ n3473 ;
  assign n11929 = n3476 ^ n824 ;
  assign n11931 = n11930 ^ n11929 ;
  assign n11934 = x30 & n11931 ;
  assign n11935 = n11934 ^ n11930 ;
  assign n11936 = ~n3520 & n11935 ;
  assign n11937 = n11936 ^ n3476 ;
  assign n11939 = n11938 ^ n11937 ;
  assign n11941 = n11940 ^ n11939 ;
  assign n11942 = n11940 ^ n3520 ;
  assign n11943 = n11942 ^ n11940 ;
  assign n11944 = ~n11941 & ~n11943 ;
  assign n11945 = n11944 ^ n11940 ;
  assign n11946 = ~x31 & n11945 ;
  assign n11947 = n11946 ^ n11937 ;
  assign n11884 = n1054 ^ n533 ;
  assign n3640 = n1085 ^ n414 ;
  assign n11883 = n3640 ^ n155 ;
  assign n11885 = n11884 ^ n11883 ;
  assign n5333 = n799 ^ n592 ;
  assign n11881 = n5333 ^ n3086 ;
  assign n11880 = n3066 ^ n1169 ;
  assign n11882 = n11881 ^ n11880 ;
  assign n11886 = n11885 ^ n11882 ;
  assign n11887 = n11886 ^ n1404 ;
  assign n11921 = n976 ^ n489 ;
  assign n11922 = n11921 ^ n2322 ;
  assign n11919 = n662 ^ n226 ;
  assign n4742 = n1028 ^ n520 ;
  assign n11920 = n11919 ^ n4742 ;
  assign n11923 = n11922 ^ n11920 ;
  assign n5016 = n577 ^ n497 ;
  assign n11915 = n5016 ^ n836 ;
  assign n11916 = n11915 ^ n397 ;
  assign n11914 = n1472 ^ n793 ;
  assign n11917 = n11916 ^ n11914 ;
  assign n11911 = n971 ^ n455 ;
  assign n11912 = n11911 ^ n2937 ;
  assign n3797 = n981 ^ n505 ;
  assign n11910 = n3797 ^ n3464 ;
  assign n11913 = n11912 ^ n11910 ;
  assign n11918 = n11917 ^ n11913 ;
  assign n11924 = n11923 ^ n11918 ;
  assign n4798 = n2610 ^ n1494 ;
  assign n4796 = n268 ^ n156 ;
  assign n4797 = n4796 ^ n540 ;
  assign n4799 = n4798 ^ n4797 ;
  assign n4793 = n790 ^ n161 ;
  assign n4794 = n4793 ^ n144 ;
  assign n4795 = n4794 ^ n570 ;
  assign n4800 = n4799 ^ n4795 ;
  assign n11925 = n11924 ^ n4800 ;
  assign n11906 = n1069 ^ n404 ;
  assign n11905 = n2627 ^ n561 ;
  assign n11907 = n11906 ^ n11905 ;
  assign n11902 = n1177 ^ n739 ;
  assign n11903 = n11902 ^ n628 ;
  assign n11900 = n1967 ^ n621 ;
  assign n5335 = n308 ^ n252 ;
  assign n11899 = n5335 ^ n2809 ;
  assign n11901 = n11900 ^ n11899 ;
  assign n11904 = n11903 ^ n11901 ;
  assign n11908 = n11907 ^ n11904 ;
  assign n11894 = n1093 ^ n321 ;
  assign n11895 = n11894 ^ n450 ;
  assign n11892 = n285 ^ n221 ;
  assign n11893 = n11892 ^ n362 ;
  assign n11896 = n11895 ^ n11893 ;
  assign n11890 = n1074 ^ n747 ;
  assign n11888 = n273 ^ n197 ;
  assign n11889 = n11888 ^ n2888 ;
  assign n11891 = n11890 ^ n11889 ;
  assign n11897 = n11896 ^ n11891 ;
  assign n11898 = n11897 ^ n2120 ;
  assign n11909 = n11908 ^ n11898 ;
  assign n11926 = n11925 ^ n11909 ;
  assign n11927 = ~n11887 & ~n11926 ;
  assign n11987 = n11947 ^ n11927 ;
  assign n12356 = n12355 ^ n11987 ;
  assign n12357 = n12356 ^ n12355 ;
  assign n12358 = n12020 ^ n11927 ;
  assign n12359 = n12358 ^ n12355 ;
  assign n12360 = ~n12357 & ~n12359 ;
  assign n12361 = n12360 ^ n12355 ;
  assign n12362 = n12354 & ~n12361 ;
  assign n12363 = n12362 ^ n12020 ;
  assign n12587 = n12586 ^ n12363 ;
  assign n12588 = n12587 ^ n12346 ;
  assign n12589 = n12588 ^ n12586 ;
  assign n12590 = n12352 & n12589 ;
  assign n12591 = n12590 ^ n12587 ;
  assign n12364 = n12363 ^ n12352 ;
  assign n3500 = n3499 ^ n485 ;
  assign n11963 = n3481 & n3500 ;
  assign n653 = n28635 ^ n650 ;
  assign n11960 = n826 ^ n653 ;
  assign n11961 = n445 & n11960 ;
  assign n11959 = n3484 ^ x29 ;
  assign n11962 = n11961 ^ n11959 ;
  assign n11964 = n11963 ^ n11962 ;
  assign n11958 = ~n317 & n831 ;
  assign n11965 = n11964 ^ n11958 ;
  assign n11966 = n11965 ^ x26 ;
  assign n12861 = n12860 ^ n80 ;
  assign n486 = n72 ^ n65 ;
  assign n487 = n486 ^ n55 ;
  assign n3501 = n487 ^ n64 ;
  assign n11955 = ~n3501 & ~n3920 ;
  assign n11956 = ~n12861 ^ n11955 ;
  assign n11957 = ~n3943 & ~n11956 ;
  assign n11967 = n11966 ^ n11957 ;
  assign n11928 = n11927 ^ n11837 ;
  assign n11948 = n11947 ^ n11928 ;
  assign n3858 = n2912 ^ n360 ;
  assign n3859 = n3858 ^ n273 ;
  assign n3857 = n2069 ^ n109 ;
  assign n3860 = n3859 ^ n3857 ;
  assign n3856 = n3855 ^ n2925 ;
  assign n3861 = n3860 ^ n3856 ;
  assign n3852 = n3851 ^ n1269 ;
  assign n3853 = n3852 ^ n2544 ;
  assign n3849 = n1171 ^ n621 ;
  assign n3850 = n3849 ^ n603 ;
  assign n3854 = n3853 ^ n3850 ;
  assign n3862 = n3861 ^ n3854 ;
  assign n3846 = n1839 ^ n380 ;
  assign n3844 = n1219 ^ n932 ;
  assign n3842 = n1197 ^ n238 ;
  assign n3843 = n3842 ^ n417 ;
  assign n3845 = n3844 ^ n3843 ;
  assign n3847 = n3846 ^ n3845 ;
  assign n3848 = n3847 ^ n1940 ;
  assign n3863 = n3862 ^ n3848 ;
  assign n3892 = n495 ^ n242 ;
  assign n3893 = n3892 ^ n954 ;
  assign n3889 = n607 ^ n249 ;
  assign n3890 = n3889 ^ n878 ;
  assign n3887 = n426 ^ n87 ;
  assign n3888 = n3887 ^ n1190 ;
  assign n3891 = n3890 ^ n3888 ;
  assign n3894 = n3893 ^ n3891 ;
  assign n3884 = n689 ^ n560 ;
  assign n3885 = n3884 ^ n662 ;
  assign n3882 = n520 ^ n407 ;
  assign n3881 = n2313 ^ n137 ;
  assign n3883 = n3882 ^ n3881 ;
  assign n3886 = n3885 ^ n3883 ;
  assign n3895 = n3894 ^ n3886 ;
  assign n3877 = n627 ^ n565 ;
  assign n3876 = n1283 ^ n521 ;
  assign n3878 = n3877 ^ n3876 ;
  assign n3874 = n1093 ^ n971 ;
  assign n3873 = n1509 ^ n1249 ;
  assign n3875 = n3874 ^ n3873 ;
  assign n3879 = n3878 ^ n3875 ;
  assign n3880 = n3879 ^ n3080 ;
  assign n3896 = n3895 ^ n3880 ;
  assign n3869 = n2060 ^ n172 ;
  assign n3870 = n3869 ^ n677 ;
  assign n3867 = n946 ^ n737 ;
  assign n3868 = n3867 ^ n1132 ;
  assign n3871 = n3870 ^ n3868 ;
  assign n3799 = n814 ^ n210 ;
  assign n3865 = n3799 ^ n3251 ;
  assign n3864 = n1009 ^ n693 ;
  assign n3866 = n3865 ^ n3864 ;
  assign n3872 = n3871 ^ n3866 ;
  assign n3897 = n3896 ^ n3872 ;
  assign n3898 = ~n3863 & ~n3897 ;
  assign n4039 = n3898 ^ x23 ;
  assign n3990 = n937 ^ n370 ;
  assign n3987 = n521 ^ n425 ;
  assign n3988 = n3987 ^ n284 ;
  assign n3989 = n3988 ^ n533 ;
  assign n3991 = n3990 ^ n3989 ;
  assign n3985 = n3041 ^ n518 ;
  assign n3983 = n2693 ^ n230 ;
  assign n3984 = n3983 ^ n592 ;
  assign n3986 = n3985 ^ n3984 ;
  assign n3992 = n3991 ^ n3986 ;
  assign n3993 = n3992 ^ n2157 ;
  assign n3978 = n1199 ^ n1129 ;
  assign n3977 = n2167 ^ n1266 ;
  assign n3979 = n3978 ^ n3977 ;
  assign n3975 = n129 ^ n97 ;
  assign n3973 = n1249 ^ n782 ;
  assign n3972 = n1088 ^ n90 ;
  assign n3974 = n3973 ^ n3972 ;
  assign n3976 = n3975 ^ n3974 ;
  assign n3980 = n3979 ^ n3976 ;
  assign n3981 = n3980 ^ n1815 ;
  assign n3968 = n765 ^ n417 ;
  assign n3638 = n542 ^ n153 ;
  assign n3967 = n3638 ^ n155 ;
  assign n3969 = n3968 ^ n3967 ;
  assign n3965 = n583 ^ n303 ;
  assign n3964 = n2161 ^ n526 ;
  assign n3966 = n3965 ^ n3964 ;
  assign n3970 = n3969 ^ n3966 ;
  assign n3673 = n625 ^ n87 ;
  assign n3961 = n3673 ^ n577 ;
  assign n3962 = n3961 ^ n2864 ;
  assign n3963 = n3962 ^ n2942 ;
  assign n3971 = n3970 ^ n3963 ;
  assign n3982 = n3981 ^ n3971 ;
  assign n3994 = n3993 ^ n3982 ;
  assign n4032 = n1518 ^ n774 ;
  assign n4030 = n1837 ^ n183 ;
  assign n4031 = n4030 ^ n672 ;
  assign n4033 = n4032 ^ n4031 ;
  assign n4027 = n1605 ^ n194 ;
  assign n4028 = n4027 ^ n450 ;
  assign n4024 = n1303 ^ n513 ;
  assign n4025 = n4024 ^ n2662 ;
  assign n4026 = n4025 ^ n212 ;
  assign n4029 = n4028 ^ n4026 ;
  assign n4034 = n4033 ^ n4029 ;
  assign n4021 = n1215 ^ n1001 ;
  assign n4022 = n4021 ^ n870 ;
  assign n4015 = n1152 ^ n877 ;
  assign n4016 = n4015 ^ n1986 ;
  assign n4020 = n4019 ^ n4016 ;
  assign n4023 = n4022 ^ n4020 ;
  assign n4035 = n4034 ^ n4023 ;
  assign n4011 = n1658 ^ n285 ;
  assign n4012 = n4011 ^ n392 ;
  assign n4007 = n400 ^ n144 ;
  assign n4006 = n621 ^ n268 ;
  assign n4008 = n4007 ^ n4006 ;
  assign n4009 = n4008 ^ n570 ;
  assign n4004 = n1197 ^ n378 ;
  assign n4005 = n4004 ^ n252 ;
  assign n4010 = n4009 ^ n4005 ;
  assign n4013 = n4012 ^ n4010 ;
  assign n4000 = n871 ^ n150 ;
  assign n3999 = n361 ^ n223 ;
  assign n4001 = n4000 ^ n3999 ;
  assign n3997 = n1899 ^ n1224 ;
  assign n3995 = n1956 ^ n641 ;
  assign n3996 = n3995 ^ n1437 ;
  assign n3998 = n3997 ^ n3996 ;
  assign n4002 = n4001 ^ n3998 ;
  assign n4003 = n4002 ^ n801 ;
  assign n4014 = n4013 ^ n4003 ;
  assign n4036 = n4035 ^ n4014 ;
  assign n4037 = n4036 ^ n2153 ;
  assign n4038 = ~n3994 & ~n4037 ;
  assign n11851 = n4038 ^ n3898 ;
  assign n11852 = n4039 & ~n11851 ;
  assign n11853 = n11852 ^ x23 ;
  assign n11876 = n11853 ^ n11837 ;
  assign n11845 = ~n649 & n831 ;
  assign n656 = n655 ^ n653 ;
  assign n11843 = ~n445 & n656 ;
  assign n11840 = ~n317 & n3484 ;
  assign n11839 = n3481 & n4073 ;
  assign n11841 = n11840 ^ n11839 ;
  assign n11842 = n11841 ^ x29 ;
  assign n11844 = n11843 ^ n11842 ;
  assign n11846 = n11845 ^ n11844 ;
  assign n11813 = ~n33 & n824 ;
  assign n3836 = ~n35 & n1109 ;
  assign n11812 = n3724 & ~n3836 ;
  assign n11814 = n11813 ^ n11812 ;
  assign n3508 = n3473 ^ n3388 ;
  assign n11810 = n3508 & n3520 ;
  assign n11808 = x31 & ~n824 ;
  assign n11807 = ~n3387 & n3726 ;
  assign n11809 = n11808 ^ n11807 ;
  assign n11811 = n11810 ^ n11809 ;
  assign n11815 = n11814 ^ n11811 ;
  assign n11873 = n11846 ^ n11815 ;
  assign n11877 = n11873 ^ n11853 ;
  assign n3613 = n1457 ^ n1123 ;
  assign n3614 = n3613 ^ n3302 ;
  assign n3610 = n2814 ^ n303 ;
  assign n3611 = n3610 ^ n1099 ;
  assign n3609 = n3440 ^ n230 ;
  assign n3612 = n3611 ^ n3609 ;
  assign n3615 = n3614 ^ n3612 ;
  assign n3606 = n331 ^ n201 ;
  assign n3602 = n512 ^ n197 ;
  assign n3604 = n3603 ^ n3602 ;
  assign n3601 = n1058 ^ n242 ;
  assign n3605 = n3604 ^ n3601 ;
  assign n3607 = n3606 ^ n3605 ;
  assign n3608 = n3607 ^ n1812 ;
  assign n3616 = n3615 ^ n3608 ;
  assign n3597 = n3596 ^ n667 ;
  assign n3598 = n3597 ^ n1269 ;
  assign n3592 = n483 ^ n429 ;
  assign n3593 = n3592 ^ n779 ;
  assign n3594 = n3593 ^ n725 ;
  assign n3590 = n970 ^ n219 ;
  assign n3589 = n1956 ^ n122 ;
  assign n3591 = n3590 ^ n3589 ;
  assign n3595 = n3594 ^ n3591 ;
  assign n3599 = n3598 ^ n3595 ;
  assign n3583 = n856 ^ n369 ;
  assign n3584 = n3583 ^ n151 ;
  assign n3582 = n3011 ^ n229 ;
  assign n3585 = n3584 ^ n3582 ;
  assign n3580 = n2377 ^ n181 ;
  assign n3581 = n3580 ^ n3086 ;
  assign n3586 = n3585 ^ n3581 ;
  assign n3578 = n1500 ^ n905 ;
  assign n3577 = n1366 ^ n365 ;
  assign n3579 = n3578 ^ n3577 ;
  assign n3587 = n3586 ^ n3579 ;
  assign n3588 = n3587 ^ n2457 ;
  assign n3600 = n3599 ^ n3588 ;
  assign n3617 = n3616 ^ n3600 ;
  assign n3630 = n2423 ^ n280 ;
  assign n3632 = n3631 ^ n3630 ;
  assign n3629 = n2765 ^ n629 ;
  assign n3633 = n3632 ^ n3629 ;
  assign n3626 = n804 ^ n417 ;
  assign n3624 = n2709 ^ n321 ;
  assign n3625 = n3624 ^ n838 ;
  assign n3627 = n3626 ^ n3625 ;
  assign n3621 = n1970 ^ n1728 ;
  assign n3620 = n3321 ^ n1921 ;
  assign n3622 = n3621 ^ n3620 ;
  assign n3618 = n3022 ^ n490 ;
  assign n3619 = n3618 ^ n381 ;
  assign n3623 = n3622 ^ n3619 ;
  assign n3628 = n3627 ^ n3623 ;
  assign n3634 = n3633 ^ n3628 ;
  assign n3635 = n3634 ^ n2145 ;
  assign n3636 = ~n3617 & ~n3635 ;
  assign n3637 = n3636 ^ x20 ;
  assign n3678 = n1311 ^ n1123 ;
  assign n3679 = n3678 ^ n272 ;
  assign n3677 = n836 ^ n298 ;
  assign n3680 = n3679 ^ n3677 ;
  assign n3675 = n1030 ^ n110 ;
  assign n3674 = n3673 ^ n130 ;
  assign n3676 = n3675 ^ n3674 ;
  assign n3681 = n3680 ^ n3676 ;
  assign n3670 = n3121 ^ n799 ;
  assign n3668 = n1641 ^ n497 ;
  assign n3669 = n3668 ^ n104 ;
  assign n3671 = n3670 ^ n3669 ;
  assign n3664 = n881 ^ n196 ;
  assign n3665 = n3664 ^ n1847 ;
  assign n3663 = n1739 ^ n1282 ;
  assign n3666 = n3665 ^ n3663 ;
  assign n3661 = n2433 ^ n218 ;
  assign n3660 = n2771 ^ n1721 ;
  assign n3662 = n3661 ^ n3660 ;
  assign n3667 = n3666 ^ n3662 ;
  assign n3672 = n3671 ^ n3667 ;
  assign n3682 = n3681 ^ n3672 ;
  assign n3655 = n677 ^ n642 ;
  assign n3656 = n3655 ^ n1982 ;
  assign n3654 = n1254 ^ n308 ;
  assign n3657 = n3656 ^ n3654 ;
  assign n3651 = n1512 ^ n245 ;
  assign n3650 = n1050 ^ n846 ;
  assign n3652 = n3651 ^ n3650 ;
  assign n3649 = n2818 ^ n915 ;
  assign n3653 = n3652 ^ n3649 ;
  assign n3658 = n3657 ^ n3653 ;
  assign n3645 = n1516 ^ n1130 ;
  assign n3643 = n1920 ^ n230 ;
  assign n3644 = n3643 ^ n672 ;
  assign n3646 = n3645 ^ n3644 ;
  assign n3641 = n3640 ^ n683 ;
  assign n3639 = n3638 ^ n1180 ;
  assign n3642 = n3641 ^ n3639 ;
  assign n3647 = n3646 ^ n3642 ;
  assign n3648 = n3647 ^ n2165 ;
  assign n3659 = n3658 ^ n3648 ;
  assign n3683 = n3682 ^ n3659 ;
  assign n3709 = n790 ^ n222 ;
  assign n3710 = n3709 ^ n794 ;
  assign n3711 = n3710 ^ n2495 ;
  assign n3707 = n2792 ^ n250 ;
  assign n3706 = n3705 ^ n1135 ;
  assign n3708 = n3707 ^ n3706 ;
  assign n3712 = n3711 ^ n3708 ;
  assign n3699 = n279 ^ n265 ;
  assign n3700 = n3699 ^ n1140 ;
  assign n3701 = n3700 ^ n2379 ;
  assign n3697 = n810 ^ n321 ;
  assign n3696 = n2850 ^ n1148 ;
  assign n3698 = n3697 ^ n3696 ;
  assign n3702 = n3701 ^ n3698 ;
  assign n3703 = n3702 ^ n3419 ;
  assign n3692 = n918 ^ n313 ;
  assign n3693 = n3692 ^ n1054 ;
  assign n3689 = n242 ^ n236 ;
  assign n3690 = n3689 ^ n1099 ;
  assign n3691 = n3690 ^ n1358 ;
  assign n3694 = n3693 ^ n3691 ;
  assign n3687 = n732 ^ n456 ;
  assign n3684 = n1542 ^ n728 ;
  assign n3685 = n3684 ^ n364 ;
  assign n3686 = n3685 ^ n622 ;
  assign n3688 = n3687 ^ n3686 ;
  assign n3695 = n3694 ^ n3688 ;
  assign n3704 = n3703 ^ n3695 ;
  assign n3713 = n3712 ^ n3704 ;
  assign n3714 = ~n3683 & ~n3713 ;
  assign n3715 = n3714 ^ n3636 ;
  assign n3716 = n3637 & ~n3715 ;
  assign n3717 = n3716 ^ x20 ;
  assign n3533 = n2834 ^ n218 ;
  assign n3569 = n597 ^ n177 ;
  assign n3567 = n2082 ^ n90 ;
  assign n3568 = n3567 ^ n305 ;
  assign n3570 = n3569 ^ n3568 ;
  assign n3571 = n3570 ^ n3261 ;
  assign n3564 = n3563 ^ n198 ;
  assign n3561 = n804 ^ n362 ;
  assign n3562 = n3561 ^ n537 ;
  assign n3565 = n3564 ^ n3562 ;
  assign n3558 = n853 ^ n492 ;
  assign n3559 = n3558 ^ n1184 ;
  assign n3556 = n2423 ^ n622 ;
  assign n3554 = n2276 ^ n259 ;
  assign n3555 = n3554 ^ n1249 ;
  assign n3557 = n3556 ^ n3555 ;
  assign n3560 = n3559 ^ n3557 ;
  assign n3566 = n3565 ^ n3560 ;
  assign n3572 = n3571 ^ n3566 ;
  assign n3551 = n2935 ^ n1743 ;
  assign n3549 = n905 ^ n244 ;
  assign n3550 = n3549 ^ n1921 ;
  assign n3552 = n3551 ^ n3550 ;
  assign n3544 = n672 ^ n255 ;
  assign n3545 = n3544 ^ n1088 ;
  assign n3542 = n1058 ^ n526 ;
  assign n3543 = n3542 ^ n2442 ;
  assign n3546 = n3545 ^ n3543 ;
  assign n3539 = n1956 ^ n584 ;
  assign n3540 = n3539 ^ n725 ;
  assign n3541 = n3540 ^ n1859 ;
  assign n3547 = n3546 ^ n3541 ;
  assign n3537 = n1037 ^ n897 ;
  assign n3534 = n1282 ^ n1014 ;
  assign n3535 = n3534 ^ n298 ;
  assign n3536 = n3535 ^ n636 ;
  assign n3538 = n3537 ^ n3536 ;
  assign n3548 = n3547 ^ n3538 ;
  assign n3553 = n3552 ^ n3548 ;
  assign n3573 = n3572 ^ n3553 ;
  assign n3574 = n3573 ^ n1681 ;
  assign n3575 = ~n3533 & ~n3574 ;
  assign n3840 = n3717 ^ n3575 ;
  assign n3521 = n3381 ^ n968 ;
  assign n3523 = n3521 ^ n1214 ;
  assign n3522 = n3521 ^ n1540 ;
  assign n3524 = n3523 ^ n3522 ;
  assign n3527 = x30 & n3524 ;
  assign n3528 = n3527 ^ n3523 ;
  assign n3529 = ~n3520 & ~n3528 ;
  assign n3530 = n3529 ^ n3521 ;
  assign n3531 = x31 & n3530 ;
  assign n3517 = ~n35 & n1214 ;
  assign n3515 = ~n35 & n968 ;
  assign n3516 = n3515 ^ n968 ;
  assign n3518 = n3517 ^ n3516 ;
  assign n3519 = ~n3514 & ~n3518 ;
  assign n3532 = n3531 ^ n3519 ;
  assign n4041 = n3717 ^ n3532 ;
  assign n4042 = ~n3840 & n4041 ;
  assign n4054 = ~n33 & n1109 ;
  assign n4053 = ~n3515 & n3724 ;
  assign n4055 = n4054 ^ n4053 ;
  assign n3903 = ~n968 & ~n3380 ;
  assign n3902 = n968 & ~n3379 ;
  assign n3904 = n3903 ^ n3902 ;
  assign n4043 = n1109 & n3904 ;
  assign n4044 = n4043 ^ n3902 ;
  assign n4050 = n4044 ^ n824 ;
  assign n4051 = n3520 & n4050 ;
  assign n4045 = n4044 ^ n1109 ;
  assign n4048 = n3726 & ~n4045 ;
  assign n4047 = x31 & ~n1109 ;
  assign n4049 = n4048 ^ n4047 ;
  assign n4052 = n4051 ^ n4049 ;
  assign n4056 = n4055 ^ n4052 ;
  assign n4058 = n4056 ^ n3898 ;
  assign n4057 = n4056 ^ n3532 ;
  assign n4059 = n4058 ^ n4057 ;
  assign n4060 = n4042 & n4059 ;
  assign n4061 = n4060 ^ n4058 ;
  assign n4040 = n4039 ^ n4038 ;
  assign n11848 = n4056 ^ n4040 ;
  assign n11849 = ~n4061 & n11848 ;
  assign n11850 = n11849 ^ n4056 ;
  assign n11878 = n11877 ^ n11850 ;
  assign n11879 = n11876 & ~n11878 ;
  assign n11949 = n11948 ^ n11879 ;
  assign n11874 = n11850 ^ n11815 ;
  assign n11875 = n11873 & ~n11874 ;
  assign n11950 = n11949 ^ n11875 ;
  assign n12082 = n11965 ^ n11950 ;
  assign n12083 = n11967 & ~n12082 ;
  assign n12084 = n12083 ^ n11965 ;
  assign n3944 = n3943 ^ n3924 ;
  assign n12077 = n3481 & n3944 ;
  assign n12065 = n3484 ^ n445 ;
  assign n12071 = ~n831 & ~n12065 ;
  assign n12069 = n831 ^ n485 ;
  assign n12070 = ~n3484 & ~n12069 ;
  assign n12072 = n12071 ^ n12070 ;
  assign n12073 = n3943 & n12072 ;
  assign n12074 = n12073 ^ n12071 ;
  assign n12075 = n12074 ^ n485 ;
  assign n12076 = n12075 ^ x29 ;
  assign n12079 = n12077 ^ n12076 ;
  assign n12279 = n12084 ^ n12079 ;
  assign n12278 = n12079 & ~n12084 ;
  assign n12280 = n12279 ^ n12278 ;
  assign n12592 = n12364 ^ n12280 ;
  assign n4062 = n4061 ^ n4040 ;
  assign n3959 = ~n649 & n3484 ;
  assign n3957 = n3481 & n3956 ;
  assign n3952 = ~n317 & n656 ;
  assign n3951 = n831 & ~n3473 ;
  assign n3953 = n3952 ^ n3951 ;
  assign n3954 = n3953 ^ x29 ;
  assign n3958 = n3957 ^ n3954 ;
  assign n3960 = n3959 ^ n3958 ;
  assign n4063 = n4062 ^ n3960 ;
  assign n3901 = x31 & ~n3517 ;
  assign n3910 = ~x30 & n968 ;
  assign n3905 = n3904 ^ n1109 ;
  assign n3911 = n3910 ^ n3905 ;
  assign n3912 = ~n3520 & ~n3911 ;
  assign n3913 = n3912 ^ n3905 ;
  assign n3914 = n3901 & n3913 ;
  assign n3576 = n3575 ^ n3532 ;
  assign n3841 = n3576 & ~n3840 ;
  assign n3899 = n3898 ^ n3841 ;
  assign n3837 = n3836 ^ n1109 ;
  assign n3838 = n3837 ^ n3515 ;
  assign n3839 = ~n3514 & ~n3838 ;
  assign n3900 = n3899 ^ n3839 ;
  assign n3915 = n3914 ^ n3900 ;
  assign n3718 = n3717 ^ n3576 ;
  assign n3511 = ~n824 & n3484 ;
  assign n3509 = n3481 & ~n3508 ;
  assign n3505 = n656 & ~n3473 ;
  assign n3504 = n831 & ~n1109 ;
  assign n3506 = n3505 ^ n3504 ;
  assign n3507 = n3506 ^ x29 ;
  assign n3510 = n3509 ^ n3507 ;
  assign n3512 = n3511 ^ n3510 ;
  assign n3719 = n3718 ^ n3512 ;
  assign n3738 = n3714 ^ x20 ;
  assign n3739 = n3738 ^ n3636 ;
  assign n3735 = ~n1433 & n24214 ;
  assign n3734 = ~n1540 & ~n3733 ;
  assign n3736 = n3735 ^ n3734 ;
  assign n4851 = n3514 ^ n33 ;
  assign n23912 = n24214 ^ n4851 ;
  assign n3730 = n3376 & n23912 ;
  assign n3729 = ~n1214 & n3520 ;
  assign n3731 = n3730 ^ n3729 ;
  assign n3737 = n3736 ^ n3731 ;
  assign n3740 = n3739 ^ n3737 ;
  assign n3821 = ~n1433 & ~n3733 ;
  assign n3820 = ~n1351 & n24214 ;
  assign n3822 = n3821 ^ n3820 ;
  assign n3809 = n1631 & n3368 ;
  assign n3813 = ~n1703 & ~n3809 ;
  assign n3814 = n1351 & ~n3813 ;
  assign n3808 = n3368 ^ n1631 ;
  assign n3810 = n3809 ^ n3808 ;
  assign n3811 = n1703 & n3810 ;
  assign n3812 = ~n1351 & ~n3811 ;
  assign n3815 = n3814 ^ n3812 ;
  assign n3816 = n1433 & n3815 ;
  assign n3817 = n3816 ^ n3814 ;
  assign n3818 = n3817 & n23912 ;
  assign n3807 = ~n1540 & n3520 ;
  assign n3819 = n3818 ^ n3807 ;
  assign n3823 = n3822 ^ n3819 ;
  assign n3763 = n3456 ^ n2276 ;
  assign n3762 = n2660 ^ n1222 ;
  assign n3764 = n3763 ^ n3762 ;
  assign n3760 = n1527 ^ n181 ;
  assign n3761 = n3760 ^ n1776 ;
  assign n3765 = n3764 ^ n3761 ;
  assign n3757 = n2085 ^ n836 ;
  assign n3758 = n3757 ^ n2274 ;
  assign n3755 = n1731 ^ n431 ;
  assign n3756 = n3755 ^ n622 ;
  assign n3759 = n3758 ^ n3756 ;
  assign n3766 = n3765 ^ n3759 ;
  assign n3751 = n838 ^ n689 ;
  assign n3750 = n1249 ^ n172 ;
  assign n3752 = n3751 ^ n3750 ;
  assign n3748 = n682 ^ n359 ;
  assign n3746 = n355 ^ n313 ;
  assign n3747 = n3746 ^ n100 ;
  assign n3749 = n3748 ^ n3747 ;
  assign n3753 = n3752 ^ n3749 ;
  assign n3743 = n914 ^ n913 ;
  assign n3744 = n3743 ^ n1444 ;
  assign n3741 = n1847 ^ n1014 ;
  assign n3742 = n3741 ^ n780 ;
  assign n3745 = n3744 ^ n3742 ;
  assign n3754 = n3753 ^ n3745 ;
  assign n3767 = n3766 ^ n3754 ;
  assign n3803 = n2676 ^ n1525 ;
  assign n3798 = n3797 ^ n3709 ;
  assign n3800 = n3799 ^ n3798 ;
  assign n3801 = n3800 ^ n2527 ;
  assign n3794 = n1494 ^ n976 ;
  assign n3795 = n3794 ^ n579 ;
  assign n3792 = n1282 ^ n617 ;
  assign n3793 = n3792 ^ n1837 ;
  assign n3796 = n3795 ^ n3793 ;
  assign n3802 = n3801 ^ n3796 ;
  assign n3804 = n3803 ^ n3802 ;
  assign n3787 = n624 ^ n379 ;
  assign n3788 = n3787 ^ n2611 ;
  assign n3785 = n2133 ^ n560 ;
  assign n3786 = n3785 ^ n2632 ;
  assign n3789 = n3788 ^ n3786 ;
  assign n3782 = n667 ^ n429 ;
  assign n3783 = n3782 ^ n155 ;
  assign n3780 = n1260 ^ n400 ;
  assign n3781 = n3780 ^ n567 ;
  assign n3784 = n3783 ^ n3781 ;
  assign n3790 = n3789 ^ n3784 ;
  assign n3775 = n971 ^ n518 ;
  assign n3776 = n3775 ^ n2111 ;
  assign n3774 = n3773 ^ n1450 ;
  assign n3777 = n3776 ^ n3774 ;
  assign n3778 = n3777 ^ n1695 ;
  assign n3771 = n1036 ^ n621 ;
  assign n3768 = n1254 ^ n592 ;
  assign n3769 = n3768 ^ n450 ;
  assign n3770 = n3769 ^ n227 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3779 = n3778 ^ n3772 ;
  assign n3791 = n3790 ^ n3779 ;
  assign n3805 = n3804 ^ n3791 ;
  assign n3806 = ~n3767 & ~n3805 ;
  assign n3824 = n3823 ^ n3806 ;
  assign n3827 = n3806 ^ n3737 ;
  assign n3828 = n3827 ^ n3738 ;
  assign n3829 = n3824 & ~n3828 ;
  assign n3830 = n3829 ^ n3738 ;
  assign n3831 = ~n3740 & n3830 ;
  assign n3832 = n3831 ^ n3737 ;
  assign n3833 = n3832 ^ n3512 ;
  assign n3834 = ~n3719 & n3833 ;
  assign n3835 = n3834 ^ n3512 ;
  assign n3948 = n3899 ^ n3835 ;
  assign n3949 = ~n3915 & ~n3948 ;
  assign n3950 = n3949 ^ n3899 ;
  assign n11857 = n3960 ^ n3950 ;
  assign n11858 = n4063 & ~n11857 ;
  assign n11859 = n11858 ^ n3960 ;
  assign n11864 = ~n3501 & n4515 ;
  assign n446 = n165 ^ n75 ;
  assign n11861 = n446 & ~n3943 ;
  assign n11860 = ~n485 & n12861 ;
  assign n11862 = n11861 ^ n11860 ;
  assign n11863 = n11862 ^ x26 ;
  assign n11865 = n11864 ^ n11863 ;
  assign n12086 = ~n11859 & ~n11865 ;
  assign n11968 = n11967 ^ n11950 ;
  assign n12087 = n12086 ^ n11968 ;
  assign n11854 = n11853 ^ n11850 ;
  assign n11838 = n11837 ^ n11815 ;
  assign n11847 = n11846 ^ n11838 ;
  assign n11855 = n11854 ^ n11847 ;
  assign n4068 = ~n487 & ~n3943 ;
  assign n4064 = n4063 ^ n3950 ;
  assign n4065 = n4064 ^ x26 ;
  assign n3947 = ~n445 & n12861 ;
  assign n4066 = n4065 ^ n3947 ;
  assign n3946 = n446 & ~n485 ;
  assign n4067 = n4066 ^ n3946 ;
  assign n4069 = n4068 ^ n4067 ;
  assign n3945 = ~n3501 & n3944 ;
  assign n4070 = n4069 ^ n3945 ;
  assign n3502 = n3500 & ~n3501 ;
  assign n3485 = ~n3473 & n3484 ;
  assign n3482 = ~n3476 & n3481 ;
  assign n832 = ~n824 & n831 ;
  assign n657 = ~n649 & n656 ;
  assign n833 = n832 ^ n657 ;
  assign n834 = n833 ^ x29 ;
  assign n3483 = n3482 ^ n834 ;
  assign n3486 = n3485 ^ n3483 ;
  assign n3487 = n3486 ^ x26 ;
  assign n488 = ~n485 & ~n487 ;
  assign n3488 = n3487 ^ n488 ;
  assign n447 = ~n445 & n446 ;
  assign n3489 = n3488 ^ n447 ;
  assign n319 = ~n317 & n12861 ;
  assign n3490 = n3489 ^ n319 ;
  assign n3503 = n3502 ^ n3490 ;
  assign n3916 = n3915 ^ n3835 ;
  assign n3917 = n3916 ^ n3486 ;
  assign n3918 = n3503 & ~n3917 ;
  assign n3919 = n3918 ^ n3486 ;
  assign n11867 = n4064 ^ n3919 ;
  assign n11868 = ~n4070 & ~n11867 ;
  assign n11869 = n11868 ^ n4064 ;
  assign n12089 = n11855 & n11869 ;
  assign n12088 = n11869 ^ n11855 ;
  assign n12090 = n12089 ^ n12088 ;
  assign n12091 = n12087 & n12090 ;
  assign n11866 = n11865 ^ n11859 ;
  assign n12092 = n12086 ^ n11866 ;
  assign n12093 = n12092 ^ n11968 ;
  assign n4071 = n4070 ^ n3919 ;
  assign n4488 = x21 ^ x20 ;
  assign n14005 = x23 & ~n4488 ;
  assign n14007 = n14005 ^ x23 ;
  assign n14008 = n14007 ^ n4488 ;
  assign n4490 = x22 & n4488 ;
  assign n4491 = n14008 ^ n4490 ;
  assign n4492 = n4491 ^ n4488 ;
  assign n4509 = ~n3920 & n4492 ;
  assign n4494 = ~x20 & ~x21 ;
  assign n4497 = ~x22 & n4494 ;
  assign n4498 = n4497 ^ n4488 ;
  assign n4495 = n4494 ^ n4488 ;
  assign n4493 = n4490 ^ x22 ;
  assign n4496 = n4495 ^ n4493 ;
  assign n4499 = n4498 ^ n4496 ;
  assign n4500 = n4499 ^ n4497 ;
  assign n4501 = n4497 ^ x23 ;
  assign n4502 = n4501 ^ n4499 ;
  assign n4503 = n4500 & n4502 ;
  assign n4504 = n4503 ^ n4497 ;
  assign n4510 = n4509 ^ n4504 ;
  assign n4511 = ~n3943 & n4510 ;
  assign n4512 = n4511 ^ x23 ;
  assign n4082 = n3832 ^ n3719 ;
  assign n4077 = ~n445 & ~n487 ;
  assign n4076 = ~n317 & n446 ;
  assign n4078 = n4077 ^ n4076 ;
  assign n4079 = n4078 ^ x26 ;
  assign n4075 = ~n649 & n12861 ;
  assign n4080 = n4079 ^ n4075 ;
  assign n4074 = ~n3501 & n4073 ;
  assign n4081 = n4080 ^ n4074 ;
  assign n4083 = n4082 ^ n4081 ;
  assign n4476 = ~n1109 & n3484 ;
  assign n4474 = n3481 & ~n4050 ;
  assign n4471 = n831 & ~n968 ;
  assign n4470 = n656 & ~n824 ;
  assign n4472 = n4471 ^ n4470 ;
  assign n4473 = n4472 ^ x29 ;
  assign n4475 = n4474 ^ n4473 ;
  assign n4477 = n4476 ^ n4475 ;
  assign n4084 = n3806 ^ n3636 ;
  assign n4085 = n4084 ^ n3823 ;
  assign n4255 = n1561 ^ n357 ;
  assign n4254 = n1028 ^ n769 ;
  assign n4256 = n4255 ^ n4254 ;
  assign n4251 = n478 ^ n250 ;
  assign n4250 = n2161 ^ n678 ;
  assign n4252 = n4251 ^ n4250 ;
  assign n4248 = n1458 ^ n660 ;
  assign n4249 = n4248 ^ n148 ;
  assign n4253 = n4252 ^ n4249 ;
  assign n4257 = n4256 ^ n4253 ;
  assign n4258 = n4257 ^ n3414 ;
  assign n4243 = n4242 ^ n198 ;
  assign n4245 = n4244 ^ n4243 ;
  assign n4239 = n2138 ^ n1355 ;
  assign n4240 = n4239 ^ n682 ;
  assign n4237 = n1641 ^ n360 ;
  assign n4238 = n4237 ^ n547 ;
  assign n4241 = n4240 ^ n4238 ;
  assign n4246 = n4245 ^ n4241 ;
  assign n4247 = n4246 ^ n3156 ;
  assign n4259 = n4258 ^ n4247 ;
  assign n4299 = n3784 ^ n2832 ;
  assign n4294 = n362 ^ n242 ;
  assign n4295 = n4294 ^ n118 ;
  assign n4292 = n760 ^ n677 ;
  assign n4293 = n4292 ^ n751 ;
  assign n4296 = n4295 ^ n4293 ;
  assign n4297 = n4296 ^ n1371 ;
  assign n4289 = n2774 ^ n99 ;
  assign n4290 = n4289 ^ n144 ;
  assign n4287 = n1509 ^ n359 ;
  assign n4288 = n4287 ^ n1074 ;
  assign n4291 = n4290 ^ n4288 ;
  assign n4298 = n4297 ^ n4291 ;
  assign n4300 = n4299 ^ n4298 ;
  assign n4282 = n867 ^ n739 ;
  assign n4283 = n4282 ^ n1608 ;
  assign n4284 = n4283 ^ n2167 ;
  assign n4279 = n3544 ^ n836 ;
  assign n4278 = n2789 ^ n541 ;
  assign n4280 = n4279 ^ n4278 ;
  assign n4281 = n4280 ^ n1744 ;
  assign n4285 = n4284 ^ n4281 ;
  assign n4275 = n4274 ^ n391 ;
  assign n4272 = n3539 ^ n932 ;
  assign n4276 = n4275 ^ n4272 ;
  assign n4267 = n897 ^ n175 ;
  assign n4268 = n4267 ^ n3011 ;
  assign n4266 = n1259 ^ n1184 ;
  assign n4269 = n4268 ^ n4266 ;
  assign n4270 = n4269 ^ n3684 ;
  assign n4263 = n1215 ^ n417 ;
  assign n4264 = n4263 ^ n1896 ;
  assign n4261 = n1495 ^ n230 ;
  assign n4260 = n3455 ^ n565 ;
  assign n4262 = n4261 ^ n4260 ;
  assign n4265 = n4264 ^ n4262 ;
  assign n4271 = n4270 ^ n4265 ;
  assign n4277 = n4276 ^ n4271 ;
  assign n4286 = n4285 ^ n4277 ;
  assign n4301 = n4300 ^ n4286 ;
  assign n4302 = ~n4259 & ~n4301 ;
  assign n4303 = n4302 ^ x14 ;
  assign n4311 = n762 ^ n212 ;
  assign n4312 = n4311 ^ n274 ;
  assign n4313 = n4312 ^ n2228 ;
  assign n4308 = n3746 ^ n370 ;
  assign n4307 = n3887 ^ n725 ;
  assign n4309 = n4308 ^ n4307 ;
  assign n4304 = n433 ^ n100 ;
  assign n4305 = n4304 ^ n116 ;
  assign n4306 = n4305 ^ n2465 ;
  assign n4310 = n4309 ^ n4306 ;
  assign n4314 = n4313 ^ n4310 ;
  assign n4331 = n1222 ^ n678 ;
  assign n4330 = n571 ^ n379 ;
  assign n4332 = n4331 ^ n4330 ;
  assign n4328 = n1906 ^ n1578 ;
  assign n4327 = n3321 ^ n949 ;
  assign n4329 = n4328 ^ n4327 ;
  assign n4333 = n4332 ^ n4329 ;
  assign n4324 = n1465 ^ n614 ;
  assign n4322 = n1586 ^ n364 ;
  assign n4323 = n4322 ^ n1201 ;
  assign n4325 = n4324 ^ n4323 ;
  assign n4318 = n774 ^ n229 ;
  assign n4319 = n4318 ^ n513 ;
  assign n4317 = n1614 ^ n375 ;
  assign n4320 = n4319 ^ n4317 ;
  assign n4127 = n848 ^ n403 ;
  assign n4315 = n4127 ^ n919 ;
  assign n4316 = n4315 ^ n2969 ;
  assign n4321 = n4320 ^ n4316 ;
  assign n4326 = n4325 ^ n4321 ;
  assign n4334 = n4333 ^ n4326 ;
  assign n4231 = n1597 ^ n178 ;
  assign n4229 = n4228 ^ n252 ;
  assign n4230 = n4229 ^ n722 ;
  assign n4232 = n4231 ^ n4230 ;
  assign n4233 = n4232 ^ n2895 ;
  assign n4335 = n4334 ^ n4233 ;
  assign n4371 = n259 ^ n175 ;
  assign n4372 = n4371 ^ n682 ;
  assign n4373 = n4372 ^ n1569 ;
  assign n4368 = n622 ^ n286 ;
  assign n4369 = n4368 ^ n2764 ;
  assign n4366 = n769 ^ n632 ;
  assign n4367 = n4366 ^ n202 ;
  assign n4370 = n4369 ^ n4367 ;
  assign n4374 = n4373 ^ n4370 ;
  assign n4362 = n1785 ^ n206 ;
  assign n4363 = n4362 ^ n1319 ;
  assign n4364 = n4363 ^ n894 ;
  assign n4358 = n583 ^ n176 ;
  assign n4359 = n4358 ^ n1414 ;
  assign n4356 = n540 ^ n483 ;
  assign n4357 = n4356 ^ n361 ;
  assign n4360 = n4359 ^ n4357 ;
  assign n4361 = n4360 ^ n2942 ;
  assign n4365 = n4364 ^ n4361 ;
  assign n4375 = n4374 ^ n4365 ;
  assign n4351 = n1122 ^ n242 ;
  assign n4352 = n4351 ^ n1129 ;
  assign n4348 = n3563 ^ n261 ;
  assign n4349 = n4348 ^ n109 ;
  assign n4347 = n559 ^ n219 ;
  assign n4350 = n4349 ^ n4347 ;
  assign n4353 = n4352 ^ n4350 ;
  assign n4354 = n4353 ^ n1034 ;
  assign n4342 = n1050 ^ n396 ;
  assign n4341 = n765 ^ n308 ;
  assign n4343 = n4342 ^ n4341 ;
  assign n4345 = n4344 ^ n4343 ;
  assign n4338 = n4183 ^ n1085 ;
  assign n4336 = n565 ^ n97 ;
  assign n4337 = n4336 ^ n2883 ;
  assign n4339 = n4338 ^ n4337 ;
  assign n4340 = n4339 ^ n3842 ;
  assign n4346 = n4345 ^ n4340 ;
  assign n4355 = n4354 ^ n4346 ;
  assign n4376 = n4375 ^ n4355 ;
  assign n4377 = ~n4335 & ~n4376 ;
  assign n4378 = ~n4314 & n4377 ;
  assign n4379 = n4378 ^ n4302 ;
  assign n4380 = n4303 & ~n4379 ;
  assign n4381 = n4380 ^ x14 ;
  assign n4197 = n4196 ^ n785 ;
  assign n4223 = n1014 ^ n512 ;
  assign n4224 = n4223 ^ n790 ;
  assign n4221 = n1828 ^ n489 ;
  assign n4222 = n4221 ^ n3398 ;
  assign n4225 = n4224 ^ n4222 ;
  assign n4219 = n225 ^ n88 ;
  assign n4217 = n571 ^ n505 ;
  assign n4218 = n4217 ^ n87 ;
  assign n4220 = n4219 ^ n4218 ;
  assign n4226 = n4225 ^ n4220 ;
  assign n4214 = n3433 ^ n888 ;
  assign n4213 = n658 ^ n590 ;
  assign n4215 = n4214 ^ n4213 ;
  assign n4216 = n4215 ^ n2563 ;
  assign n4227 = n4226 ^ n4216 ;
  assign n4234 = n4233 ^ n4227 ;
  assign n4209 = n2423 ^ n405 ;
  assign n4206 = n2308 ^ n1058 ;
  assign n4207 = n4206 ^ n932 ;
  assign n4205 = n2883 ^ n1513 ;
  assign n4208 = n4207 ^ n4205 ;
  assign n4210 = n4209 ^ n4208 ;
  assign n4211 = n4210 ^ n2976 ;
  assign n4202 = n2988 ^ n417 ;
  assign n4199 = n116 ^ n104 ;
  assign n4200 = n4199 ^ n731 ;
  assign n4201 = n4200 ^ n2495 ;
  assign n4203 = n4202 ^ n4201 ;
  assign n4198 = n3760 ^ n2784 ;
  assign n4204 = n4203 ^ n4198 ;
  assign n4212 = n4211 ^ n4204 ;
  assign n4235 = n4234 ^ n4212 ;
  assign n4236 = ~n4197 & ~n4235 ;
  assign n4382 = n4381 ^ n4236 ;
  assign n4404 = x31 & ~n1795 ;
  assign n4405 = n4404 ^ n1871 ;
  assign n4406 = ~n35 & ~n4405 ;
  assign n4400 = x31 & ~n1871 ;
  assign n4394 = ~n1631 & ~n23912 ;
  assign n4383 = n1994 & ~n3360 ;
  assign n4384 = n4383 ^ n3237 ;
  assign n4387 = n3237 ^ n1871 ;
  assign n4388 = n4387 ^ n3237 ;
  assign n4389 = n4384 & n4388 ;
  assign n4390 = n4389 ^ n3237 ;
  assign n4391 = n1872 & ~n4390 ;
  assign n4392 = n4391 ^ n1631 ;
  assign n4393 = x31 & ~n4392 ;
  assign n4395 = n4394 ^ n4393 ;
  assign n4401 = n4400 ^ n4395 ;
  assign n4402 = ~n3520 & n4401 ;
  assign n4403 = n4402 ^ n4395 ;
  assign n4407 = n4406 ^ n4403 ;
  assign n4408 = n4407 ^ n4381 ;
  assign n4409 = ~n4382 & n4408 ;
  assign n4132 = n971 ^ n579 ;
  assign n4133 = n4132 ^ n1201 ;
  assign n4130 = n1640 ^ n597 ;
  assign n4131 = n4130 ^ n737 ;
  assign n4134 = n4133 ^ n4131 ;
  assign n4128 = n4127 ^ n1783 ;
  assign n4129 = n4128 ^ n994 ;
  assign n4135 = n4134 ^ n4129 ;
  assign n4136 = n4135 ^ n891 ;
  assign n4137 = n4136 ^ n234 ;
  assign n4142 = n1512 ^ n489 ;
  assign n4140 = n2713 ^ n914 ;
  assign n4138 = n2647 ^ n245 ;
  assign n4139 = n4138 ^ n369 ;
  assign n4141 = n4140 ^ n4139 ;
  assign n4143 = n4142 ^ n4141 ;
  assign n4144 = n4143 ^ n2728 ;
  assign n4145 = n4144 ^ n2922 ;
  assign n4146 = n4145 ^ n3447 ;
  assign n4147 = ~n4137 & ~n4146 ;
  assign n4410 = n4407 ^ n4147 ;
  assign n4411 = n4409 & n4410 ;
  assign n4121 = n1355 ^ n848 ;
  assign n4122 = n4121 ^ n1767 ;
  assign n4119 = n2845 ^ n483 ;
  assign n4117 = n2432 ^ n417 ;
  assign n4118 = n4117 ^ n625 ;
  assign n4120 = n4119 ^ n4118 ;
  assign n4123 = n4122 ^ n4120 ;
  assign n4112 = n1494 ^ n1222 ;
  assign n4113 = n4112 ^ n660 ;
  assign n4110 = n505 ^ n192 ;
  assign n4111 = n4110 ^ n116 ;
  assign n4114 = n4113 ^ n4111 ;
  assign n4108 = n2085 ^ n1933 ;
  assign n4109 = n4108 ^ n1608 ;
  assign n4115 = n4114 ^ n4109 ;
  assign n4107 = n1648 ^ n367 ;
  assign n4116 = n4115 ^ n4107 ;
  assign n4124 = n4123 ^ n4116 ;
  assign n4101 = n1759 ^ n1219 ;
  assign n4102 = n4101 ^ n497 ;
  assign n4103 = n4102 ^ n1309 ;
  assign n4104 = n4103 ^ n3630 ;
  assign n4100 = n3144 ^ n1962 ;
  assign n4105 = n4104 ^ n4100 ;
  assign n4097 = n1480 ^ n835 ;
  assign n4095 = n2907 ^ n154 ;
  assign n4092 = n971 ^ n413 ;
  assign n4093 = n4092 ^ n614 ;
  assign n4094 = n4093 ^ n697 ;
  assign n4096 = n4095 ^ n4094 ;
  assign n4098 = n4097 ^ n4096 ;
  assign n4089 = n2334 ^ n403 ;
  assign n4090 = n4089 ^ n1602 ;
  assign n4087 = n810 ^ n512 ;
  assign n4086 = n1740 ^ n732 ;
  assign n4088 = n4087 ^ n4086 ;
  assign n4091 = n4090 ^ n4088 ;
  assign n4099 = n4098 ^ n4091 ;
  assign n4106 = n4105 ^ n4099 ;
  assign n4125 = n4124 ^ n4106 ;
  assign n4126 = ~n1108 & ~n4125 ;
  assign n4179 = n4126 ^ x17 ;
  assign n4412 = n4411 ^ n4179 ;
  assign n4430 = ~x30 & ~n1703 ;
  assign n4431 = n4430 ^ n1704 ;
  assign n4432 = ~n3520 & n4431 ;
  assign n4416 = n3813 ^ n3811 ;
  assign n4417 = n4416 ^ n1351 ;
  assign n4419 = n4417 ^ n1631 ;
  assign n4418 = n4417 ^ n1703 ;
  assign n4420 = n4419 ^ n4418 ;
  assign n4423 = ~x30 & n4420 ;
  assign n4424 = n4423 ^ n4419 ;
  assign n4425 = ~n3520 & ~n4424 ;
  assign n4426 = n4425 ^ n4417 ;
  assign n4427 = n4426 ^ n1351 ;
  assign n4433 = n4432 ^ n4427 ;
  assign n4434 = ~x31 & ~n4433 ;
  assign n4435 = n4434 ^ n4426 ;
  assign n4413 = n4179 ^ n4147 ;
  assign n4436 = n4435 ^ n4413 ;
  assign n4437 = n4412 & ~n4436 ;
  assign n4438 = n4437 ^ n4435 ;
  assign n4174 = ~n1214 & n3484 ;
  assign n4173 = n3481 & n3521 ;
  assign n4175 = n4174 ^ n4173 ;
  assign n4176 = n4175 ^ x29 ;
  assign n4172 = n656 & ~n968 ;
  assign n4177 = n4176 ^ n4172 ;
  assign n4171 = n831 & ~n1540 ;
  assign n4178 = n4177 ^ n4171 ;
  assign n4444 = n4438 ^ n4178 ;
  assign n4148 = n4147 ^ n4126 ;
  assign n4149 = n4147 ^ x17 ;
  assign n4150 = ~n4148 & n4149 ;
  assign n4151 = n4150 ^ x17 ;
  assign n4445 = n4444 ^ n4151 ;
  assign n4439 = ~n4178 & ~n4438 ;
  assign n4446 = n4445 ^ n4439 ;
  assign n4447 = n4446 ^ n4151 ;
  assign n4450 = n3636 & ~n4447 ;
  assign n4164 = ~n1433 & n3726 ;
  assign n4163 = ~n1351 & ~n3724 ;
  assign n4165 = n4164 ^ n4163 ;
  assign n4152 = n3815 ^ n1433 ;
  assign n4154 = n4152 ^ n1351 ;
  assign n4153 = n4152 ^ n1703 ;
  assign n4155 = n4154 ^ n4153 ;
  assign n4158 = x30 & n4155 ;
  assign n4159 = n4158 ^ n4154 ;
  assign n4160 = ~n3520 & ~n4159 ;
  assign n4161 = n4160 ^ n4152 ;
  assign n4162 = x31 & n4161 ;
  assign n4166 = n4165 ^ n4162 ;
  assign n4168 = ~n4151 & n4166 ;
  assign n4440 = ~n3636 & ~n4168 ;
  assign n4441 = n4439 & n4440 ;
  assign n4442 = n4441 ^ n4166 ;
  assign n4443 = n4442 ^ n4151 ;
  assign n4451 = n4450 ^ n4443 ;
  assign n4452 = n4451 ^ n4442 ;
  assign n4453 = n4441 ^ n4151 ;
  assign n4454 = n4453 ^ n4442 ;
  assign n4455 = n4452 & ~n4454 ;
  assign n4456 = n4455 ^ n4442 ;
  assign n4457 = n4085 & ~n4456 ;
  assign n4458 = n4457 ^ n4441 ;
  assign n4459 = n4178 ^ n3636 ;
  assign n4464 = ~n4444 & n4459 ;
  assign n4465 = n4464 ^ n3636 ;
  assign n4466 = ~n4458 & ~n4465 ;
  assign n4468 = n4466 ^ n4458 ;
  assign n4167 = n4166 ^ n4151 ;
  assign n4169 = n4168 ^ n4167 ;
  assign n4170 = ~n4085 & ~n4169 ;
  assign n4467 = n4170 & n4466 ;
  assign n4469 = n4468 ^ n4467 ;
  assign n4478 = n4477 ^ n4469 ;
  assign n4481 = n3824 & ~n4084 ;
  assign n4479 = n3738 ^ n3737 ;
  assign n4480 = n4479 ^ n4477 ;
  assign n4482 = n4481 ^ n4480 ;
  assign n4483 = ~n4478 & ~n4482 ;
  assign n4484 = n4483 ^ n4477 ;
  assign n4485 = n4484 ^ n4081 ;
  assign n4486 = ~n4083 & n4485 ;
  assign n4487 = n4486 ^ n4081 ;
  assign n4513 = n4512 ^ n4487 ;
  assign n4519 = n4484 ^ n4083 ;
  assign n4520 = n4519 ^ x23 ;
  assign n4518 = ~n3943 & ~n4496 ;
  assign n4521 = n4520 ^ n4518 ;
  assign n4517 = ~n485 & n4504 ;
  assign n4522 = n4521 ^ n4517 ;
  assign n4516 = n4492 & n4515 ;
  assign n4523 = n4522 ^ n4516 ;
  assign n4531 = n446 & ~n649 ;
  assign n4527 = n4482 ^ n4469 ;
  assign n4528 = n4527 ^ x26 ;
  assign n4526 = ~n3473 & n12861 ;
  assign n4529 = n4528 ^ n4526 ;
  assign n4525 = ~n317 & ~n487 ;
  assign n4530 = n4529 ^ n4525 ;
  assign n4532 = n4531 ^ n4530 ;
  assign n4524 = ~n3501 & n3956 ;
  assign n4533 = n4532 ^ n4524 ;
  assign n4552 = n831 & ~n1214 ;
  assign n4545 = ~n824 & n12861 ;
  assign n4544 = n446 & ~n3473 ;
  assign n4546 = n4545 ^ n4544 ;
  assign n4547 = n4546 ^ x26 ;
  assign n4543 = ~n487 & ~n649 ;
  assign n4548 = n4547 ^ n4543 ;
  assign n4542 = ~n3476 & ~n3501 ;
  assign n4549 = n4548 ^ n4542 ;
  assign n4550 = n4549 ^ x29 ;
  assign n4539 = ~n3904 & n4536 ;
  assign n4540 = n4539 ^ n1109 ;
  assign n4541 = n650 & ~n4540 ;
  assign n4551 = n4550 ^ n4541 ;
  assign n4553 = n4552 ^ n4551 ;
  assign n4534 = ~n968 & n3484 ;
  assign n4554 = n4553 ^ n4534 ;
  assign n4448 = n4151 ^ n3636 ;
  assign n4555 = n4438 ^ n4166 ;
  assign n4557 = n4555 ^ n4459 ;
  assign n4558 = n4448 & n4557 ;
  assign n4556 = ~n4444 & ~n4555 ;
  assign n4559 = n4558 ^ n4556 ;
  assign n4560 = n4559 ^ n4085 ;
  assign n4561 = n4560 ^ n4549 ;
  assign n4562 = n4554 & n4561 ;
  assign n4563 = n4562 ^ n4549 ;
  assign n4564 = n4563 ^ n4527 ;
  assign n4565 = n4533 & n4564 ;
  assign n4566 = n4565 ^ n4527 ;
  assign n4567 = n4566 ^ n4519 ;
  assign n4568 = ~n4523 & ~n4567 ;
  assign n4569 = n4568 ^ n4519 ;
  assign n4570 = n4569 ^ n4487 ;
  assign n4571 = ~n4513 & ~n4570 ;
  assign n4572 = n4571 ^ n4569 ;
  assign n4573 = n4071 & n4572 ;
  assign n11787 = n3916 ^ n3503 ;
  assign n11788 = n4572 ^ n4071 ;
  assign n11789 = n11788 ^ n4573 ;
  assign n11790 = n11787 & n11789 ;
  assign n4665 = ~n445 & n4504 ;
  assign n4700 = x23 ^ x22 ;
  assign n4661 = ~n3924 & n4700 ;
  assign n4662 = n4661 ^ n3943 ;
  assign n4663 = n4488 & ~n4662 ;
  assign n4664 = n4663 ^ x23 ;
  assign n4666 = n4665 ^ n4664 ;
  assign n4656 = ~n485 & ~n4496 ;
  assign n4667 = n4666 ^ n4656 ;
  assign n4655 = n4563 ^ n4533 ;
  assign n4668 = n4667 ^ n4655 ;
  assign n4582 = n4560 ^ n4554 ;
  assign n4579 = ~n485 & n4491 ;
  assign n4578 = ~n445 & ~n4496 ;
  assign n4580 = n4579 ^ n4578 ;
  assign n4575 = ~n317 & n4504 ;
  assign n4574 = n3500 & n4492 ;
  assign n4576 = n4575 ^ n4574 ;
  assign n4577 = n4576 ^ x23 ;
  assign n4581 = n4580 ^ n4577 ;
  assign n4583 = n4582 ^ n4581 ;
  assign n4587 = n4448 ^ n4166 ;
  assign n4588 = n4587 ^ n4178 ;
  assign n4589 = n4588 ^ n4438 ;
  assign n4651 = n4589 ^ n4581 ;
  assign n4593 = n446 & ~n824 ;
  assign n4590 = n4589 ^ x26 ;
  assign n4586 = ~n1109 & n12861 ;
  assign n4591 = n4590 ^ n4586 ;
  assign n4585 = ~n487 & ~n3473 ;
  assign n4592 = n4591 ^ n4585 ;
  assign n4594 = n4593 ^ n4592 ;
  assign n4584 = ~n3501 & ~n3508 ;
  assign n4595 = n4594 ^ n4584 ;
  assign n4603 = n3376 ^ n1214 ;
  assign n4604 = n3481 & ~n4603 ;
  assign n4601 = n831 & ~n1433 ;
  assign n4599 = n656 & ~n1214 ;
  assign n4597 = n4435 ^ n4412 ;
  assign n4598 = n4597 ^ x29 ;
  assign n4600 = n4599 ^ n4598 ;
  assign n4602 = n4601 ^ n4600 ;
  assign n4605 = n4604 ^ n4602 ;
  assign n4596 = ~n1540 & n3484 ;
  assign n4606 = n4605 ^ n4596 ;
  assign n4640 = n831 & ~n1351 ;
  assign n4631 = x30 & ~n1631 ;
  assign n4615 = n3808 ^ n1703 ;
  assign n4617 = n4615 ^ n1631 ;
  assign n4616 = n4615 ^ n1871 ;
  assign n4618 = n4617 ^ n4616 ;
  assign n4621 = x30 & n4618 ;
  assign n4622 = n4621 ^ n4617 ;
  assign n4623 = ~n3520 & n4622 ;
  assign n4624 = n4623 ^ n4615 ;
  assign n4625 = n4624 ^ n1703 ;
  assign n4626 = n4625 ^ n4624 ;
  assign n4632 = n4631 ^ n4626 ;
  assign n4633 = ~n3520 & ~n4632 ;
  assign n4634 = n4633 ^ n4625 ;
  assign n4635 = ~x31 & n4634 ;
  assign n4636 = n4635 ^ n4624 ;
  assign n4637 = n4636 ^ x29 ;
  assign n4612 = n3817 & n4536 ;
  assign n4613 = n4612 ^ n1540 ;
  assign n4614 = n650 & ~n4613 ;
  assign n4638 = n4637 ^ n4614 ;
  assign n4607 = ~n1433 & n3484 ;
  assign n4639 = n4638 ^ n4607 ;
  assign n4641 = n4640 ^ n4639 ;
  assign n4642 = n4409 ^ n4147 ;
  assign n4643 = n4642 ^ n4636 ;
  assign n4644 = ~n4641 & n4643 ;
  assign n4645 = n4644 ^ n4636 ;
  assign n4646 = n4645 ^ n4597 ;
  assign n4647 = ~n4606 & n4646 ;
  assign n4648 = n4647 ^ n4597 ;
  assign n4649 = n4648 ^ n4589 ;
  assign n4650 = ~n4595 & n4649 ;
  assign n4652 = n4651 ^ n4650 ;
  assign n4653 = n4583 & n4652 ;
  assign n4654 = n4653 ^ n4582 ;
  assign n11775 = n4668 ^ n4654 ;
  assign n4671 = n4566 ^ n4523 ;
  assign n11776 = n4671 ^ n4654 ;
  assign n11777 = n11776 ^ n4671 ;
  assign n11778 = n4671 ^ n4667 ;
  assign n11779 = n11778 ^ n4671 ;
  assign n11780 = n11777 & n11779 ;
  assign n11781 = n11780 ^ n4671 ;
  assign n11782 = n11775 & ~n11781 ;
  assign n4709 = n4648 ^ n4595 ;
  assign n4710 = n4709 ^ x23 ;
  assign n4706 = ~n4072 & n4700 ;
  assign n4707 = n4706 ^ n445 ;
  assign n4708 = n4488 & ~n4707 ;
  assign n4711 = n4710 ^ n4708 ;
  assign n4699 = ~n649 & n4504 ;
  assign n4712 = n4711 ^ n4699 ;
  assign n4698 = ~n317 & ~n4496 ;
  assign n4713 = n4712 ^ n4698 ;
  assign n4721 = ~n487 & ~n824 ;
  assign n4717 = n4645 ^ n4606 ;
  assign n4718 = n4717 ^ x26 ;
  assign n4716 = n446 & ~n1109 ;
  assign n4719 = n4718 ^ n4716 ;
  assign n4715 = ~n968 & n12861 ;
  assign n4720 = n4719 ^ n4715 ;
  assign n4722 = n4721 ^ n4720 ;
  assign n4714 = ~n3501 & ~n4050 ;
  assign n4723 = n4722 ^ n4714 ;
  assign n4732 = n4642 ^ n4641 ;
  assign n4727 = n446 & ~n968 ;
  assign n4726 = ~n1214 & n12861 ;
  assign n4728 = n4727 ^ n4726 ;
  assign n4729 = n4728 ^ x26 ;
  assign n4725 = ~n487 & ~n1109 ;
  assign n4730 = n4729 ^ n4725 ;
  assign n4724 = ~n3501 & n3905 ;
  assign n4731 = n4730 ^ n4724 ;
  assign n4733 = n4732 ^ n4731 ;
  assign n4838 = n1795 & n3520 ;
  assign n4817 = ~n1994 & n3520 ;
  assign n4834 = x31 & ~n3236 ;
  assign n4835 = n4817 & n4834 ;
  assign n4820 = n1994 ^ x31 ;
  assign n4832 = n4820 ^ n33 ;
  assign n4827 = ~n3236 & n3359 ;
  assign n4828 = ~n35 & n4827 ;
  assign n4829 = n4828 ^ n35 ;
  assign n4830 = n4829 ^ n4820 ;
  assign n4831 = n3720 & ~n4830 ;
  assign n4833 = n4832 ^ n4831 ;
  assign n4836 = n4835 ^ n4833 ;
  assign n4815 = x31 & n3360 ;
  assign n4816 = n33 & ~n2096 ;
  assign n4818 = n4817 ^ n4816 ;
  assign n4819 = n4815 & ~n4818 ;
  assign n4837 = n4836 ^ n4819 ;
  assign n4839 = n4838 ^ n4837 ;
  assign n4738 = n149 ^ n124 ;
  assign n4739 = n4738 ^ n483 ;
  assign n4736 = n624 ^ n197 ;
  assign n4735 = n1301 ^ n355 ;
  assign n4737 = n4736 ^ n4735 ;
  assign n4740 = n4739 ^ n4737 ;
  assign n4741 = n4740 ^ n2551 ;
  assign n4780 = n628 ^ n260 ;
  assign n4777 = n1088 ^ n104 ;
  assign n4778 = n4777 ^ n396 ;
  assign n4779 = n4778 ^ n97 ;
  assign n4781 = n4780 ^ n4779 ;
  assign n4775 = n1634 ^ n1355 ;
  assign n4773 = n3799 ^ n455 ;
  assign n4774 = n4773 ^ n2377 ;
  assign n4776 = n4775 ^ n4774 ;
  assign n4782 = n4781 ^ n4776 ;
  assign n4770 = n933 ^ n409 ;
  assign n4769 = n252 ^ n143 ;
  assign n4771 = n4770 ^ n4769 ;
  assign n4765 = n489 ^ n360 ;
  assign n4766 = n4765 ^ n4132 ;
  assign n4764 = n2745 ^ n1759 ;
  assign n4767 = n4766 ^ n4764 ;
  assign n4768 = n4767 ^ n1147 ;
  assign n4772 = n4771 ^ n4768 ;
  assign n4783 = n4782 ^ n4772 ;
  assign n4760 = n779 ^ n237 ;
  assign n4758 = n977 ^ n216 ;
  assign n4759 = n4758 ^ n413 ;
  assign n4761 = n4760 ^ n4759 ;
  assign n4756 = n3041 ^ n1677 ;
  assign n4753 = n661 ^ n559 ;
  assign n4751 = n797 ^ n264 ;
  assign n4752 = n4751 ^ n200 ;
  assign n4754 = n4753 ^ n4752 ;
  assign n4755 = n4754 ^ n1998 ;
  assign n4757 = n4756 ^ n4755 ;
  assign n4762 = n4761 ^ n4757 ;
  assign n4747 = n1970 ^ n845 ;
  assign n4748 = n4747 ^ n1451 ;
  assign n4749 = n4748 ^ n1244 ;
  assign n4745 = n987 ^ n635 ;
  assign n4743 = n4742 ^ n362 ;
  assign n4744 = n4743 ^ n2849 ;
  assign n4746 = n4745 ^ n4744 ;
  assign n4750 = n4749 ^ n4746 ;
  assign n4763 = n4762 ^ n4750 ;
  assign n4784 = n4783 ^ n4763 ;
  assign n4806 = n893 ^ n514 ;
  assign n4807 = n4806 ^ n1219 ;
  assign n4808 = n4807 ^ n4244 ;
  assign n4809 = n4808 ^ n2583 ;
  assign n4802 = n886 ^ n490 ;
  assign n4803 = n4802 ^ n643 ;
  assign n4805 = n4804 ^ n4803 ;
  assign n4810 = n4809 ^ n4805 ;
  assign n4790 = n1649 ^ n518 ;
  assign n4791 = n4790 ^ n3613 ;
  assign n4788 = n819 ^ n560 ;
  assign n4786 = n4785 ^ n2365 ;
  assign n4787 = n4786 ^ n313 ;
  assign n4789 = n4788 ^ n4787 ;
  assign n4792 = n4791 ^ n4789 ;
  assign n4801 = n4800 ^ n4792 ;
  assign n4811 = n4810 ^ n4801 ;
  assign n4812 = n4811 ^ n702 ;
  assign n4813 = ~n4784 & ~n4812 ;
  assign n4814 = ~n4741 & n4813 ;
  assign n4840 = n4839 ^ n4814 ;
  assign n4841 = n4839 ^ n4378 ;
  assign n4842 = ~n4840 & ~n4841 ;
  assign n4843 = n4842 ^ n4303 ;
  assign n4863 = n4842 ^ n4378 ;
  assign n4853 = n1994 & n24214 ;
  assign n4852 = ~n4404 & ~n4851 ;
  assign n4854 = n4853 ^ n4852 ;
  assign n4857 = ~n1795 & n4384 ;
  assign n4858 = n4857 ^ n3237 ;
  assign n4859 = n4858 ^ n1871 ;
  assign n4860 = n3520 & n4859 ;
  assign n4861 = ~n4854 & n4860 ;
  assign n4848 = ~n35 & n1872 ;
  assign n4849 = n4848 ^ n1871 ;
  assign n4850 = ~n3514 & ~n4849 ;
  assign n4855 = n4854 ^ n4850 ;
  assign n4862 = n4861 ^ n4855 ;
  assign n4864 = n4863 ^ n4862 ;
  assign n4865 = n4843 & ~n4864 ;
  assign n4866 = n4865 ^ n4862 ;
  assign n4878 = n4866 ^ n4731 ;
  assign n4734 = n4407 ^ n4382 ;
  assign n4867 = n4866 ^ n4734 ;
  assign n4871 = ~n1351 & n3484 ;
  assign n4870 = n3481 & n4152 ;
  assign n4872 = n4871 ^ n4870 ;
  assign n4873 = n4872 ^ x29 ;
  assign n4869 = n656 & ~n1433 ;
  assign n4874 = n4873 ^ n4869 ;
  assign n4868 = n831 & ~n1703 ;
  assign n4875 = n4874 ^ n4868 ;
  assign n4876 = n4875 ^ n4866 ;
  assign n4877 = n4867 & ~n4876 ;
  assign n4879 = n4878 ^ n4877 ;
  assign n4880 = n4733 & n4879 ;
  assign n4881 = n4880 ^ n4732 ;
  assign n4882 = n4881 ^ n4717 ;
  assign n4883 = n4723 & n4882 ;
  assign n4884 = n4883 ^ n4717 ;
  assign n4885 = n4884 ^ n4709 ;
  assign n4886 = n4713 & n4885 ;
  assign n4887 = n4886 ^ n4709 ;
  assign n4888 = n4887 ^ x20 ;
  assign n4675 = ~x17 & x18 ;
  assign n4677 = n4675 ^ x18 ;
  assign n4676 = n4675 ^ x17 ;
  assign n4678 = n4677 ^ n4676 ;
  assign n4681 = x19 & n4678 ;
  assign n14025 = n4681 ^ n4676 ;
  assign n4685 = x20 ^ x19 ;
  assign n4679 = x20 & ~n4678 ;
  assign n4686 = n4679 ^ n4676 ;
  assign n4687 = ~n4685 & n4686 ;
  assign n14026 = n14025 ^ n4687 ;
  assign n14027 = n14026 ^ x20 ;
  assign n4682 = n4681 ^ n4678 ;
  assign n4680 = n4679 ^ x20 ;
  assign n4683 = n4682 ^ n4680 ;
  assign n4684 = n4683 ^ n4678 ;
  assign n4695 = ~n3920 & n4684 ;
  assign n4696 = n14027 ^ n4695 ;
  assign n4697 = ~n3943 & n4696 ;
  assign n4889 = n4888 ^ n4697 ;
  assign n4890 = n4652 ^ n4582 ;
  assign n4891 = n4890 ^ n4887 ;
  assign n4892 = n4889 & ~n4891 ;
  assign n4893 = n4892 ^ n4887 ;
  assign n11783 = n11782 ^ n4893 ;
  assign n6023 = n4073 & n4684 ;
  assign n4915 = n4681 ^ x19 ;
  assign n4916 = n4915 ^ n4677 ;
  assign n6020 = ~n317 & n4916 ;
  assign n6018 = ~n445 & n4683 ;
  assign n6011 = ~n968 & n4504 ;
  assign n6009 = ~n824 & n4491 ;
  assign n6007 = ~n1109 & ~n4496 ;
  assign n6005 = ~n4050 & n4492 ;
  assign n5223 = n747 ^ n392 ;
  assign n5228 = n5227 ^ n5223 ;
  assign n5221 = n983 ^ n743 ;
  assign n5219 = n5218 ^ n155 ;
  assign n5217 = n2018 ^ n705 ;
  assign n5220 = n5219 ^ n5217 ;
  assign n5222 = n5221 ^ n5220 ;
  assign n5229 = n5228 ^ n5222 ;
  assign n5123 = n1399 ^ n1356 ;
  assign n5122 = n1906 ^ n818 ;
  assign n5124 = n5123 ^ n5122 ;
  assign n5119 = n742 ^ n193 ;
  assign n5120 = n5119 ^ n739 ;
  assign n5115 = n1093 ^ n149 ;
  assign n5116 = n5115 ^ n897 ;
  assign n5117 = n5116 ^ n396 ;
  assign n5113 = n2307 ^ n106 ;
  assign n5114 = n5113 ^ n413 ;
  assign n5118 = n5117 ^ n5114 ;
  assign n5121 = n5120 ^ n5118 ;
  assign n5125 = n5124 ^ n5121 ;
  assign n5230 = n5229 ^ n5125 ;
  assign n5232 = n4221 ^ n2062 ;
  assign n5231 = n4024 ^ n2628 ;
  assign n5233 = n5232 ^ n5231 ;
  assign n5234 = n5233 ^ n3599 ;
  assign n5235 = n5234 ^ n3872 ;
  assign n5258 = n5257 ^ n360 ;
  assign n5255 = n2348 ^ n124 ;
  assign n5256 = n5255 ^ n535 ;
  assign n5259 = n5258 ^ n5256 ;
  assign n5251 = n265 ^ n194 ;
  assign n5250 = n2320 ^ n222 ;
  assign n5252 = n5251 ^ n5250 ;
  assign n5248 = n1116 ^ n567 ;
  assign n5249 = n5248 ^ n156 ;
  assign n5253 = n5252 ^ n5249 ;
  assign n5245 = n1159 ^ n682 ;
  assign n5247 = n5246 ^ n5245 ;
  assign n5254 = n5253 ^ n5247 ;
  assign n5260 = n5259 ^ n5254 ;
  assign n5242 = n2920 ^ n1426 ;
  assign n5240 = n1590 ^ n197 ;
  assign n5237 = n584 ^ n272 ;
  assign n5236 = n540 ^ n226 ;
  assign n5238 = n5237 ^ n5236 ;
  assign n5239 = n5238 ^ n261 ;
  assign n5241 = n5240 ^ n5239 ;
  assign n5243 = n5242 ^ n5241 ;
  assign n5244 = n5243 ^ n1420 ;
  assign n5261 = n5260 ^ n5244 ;
  assign n5262 = ~n5235 & ~n5261 ;
  assign n5263 = ~n5230 & n5262 ;
  assign n5264 = n5263 ^ x11 ;
  assign n5018 = n732 ^ n660 ;
  assign n5136 = n5018 ^ n3448 ;
  assign n5134 = n364 ^ n265 ;
  assign n5135 = n5134 ^ n1308 ;
  assign n5137 = n5136 ^ n5135 ;
  assign n5132 = n1834 ^ n172 ;
  assign n5129 = n1122 ^ n272 ;
  assign n5130 = n5129 ^ n4185 ;
  assign n5128 = n3103 ^ n1549 ;
  assign n5131 = n5130 ^ n5128 ;
  assign n5133 = n5132 ^ n5131 ;
  assign n5138 = n5137 ^ n5133 ;
  assign n5127 = n4361 ^ n2247 ;
  assign n5139 = n5138 ^ n5127 ;
  assign n5107 = n222 ^ n196 ;
  assign n5108 = n5107 ^ n394 ;
  assign n5109 = n5108 ^ n2910 ;
  assign n5106 = n2358 ^ n607 ;
  assign n5110 = n5109 ^ n5106 ;
  assign n5104 = n5103 ^ n637 ;
  assign n5102 = n5101 ^ n1586 ;
  assign n5105 = n5104 ^ n5102 ;
  assign n5111 = n5110 ^ n5105 ;
  assign n5097 = n1128 ^ n279 ;
  assign n5098 = n5097 ^ n702 ;
  assign n5099 = n5098 ^ n751 ;
  assign n5095 = n1943 ^ n592 ;
  assign n5094 = n3674 ^ n1197 ;
  assign n5096 = n5095 ^ n5094 ;
  assign n5100 = n5099 ^ n5096 ;
  assign n5112 = n5111 ^ n5100 ;
  assign n5126 = n5125 ^ n5112 ;
  assign n5140 = n5139 ^ n5126 ;
  assign n5141 = ~n876 & ~n5140 ;
  assign n5265 = n5264 ^ n5141 ;
  assign n4980 = n799 ^ n210 ;
  assign n4981 = n4980 ^ n274 ;
  assign n4982 = n4981 ^ n3423 ;
  assign n4979 = n1002 ^ n153 ;
  assign n4983 = n4982 ^ n4979 ;
  assign n4984 = n4983 ^ n1572 ;
  assign n4976 = n4199 ^ n764 ;
  assign n4977 = n4976 ^ n3390 ;
  assign n4973 = n739 ^ n429 ;
  assign n4974 = n4973 ^ n230 ;
  assign n4975 = n4974 ^ n2677 ;
  assign n4978 = n4977 ^ n4975 ;
  assign n4985 = n4984 ^ n4978 ;
  assign n4969 = n528 ^ n258 ;
  assign n4968 = n2117 ^ n137 ;
  assign n4970 = n4969 ^ n4968 ;
  assign n4971 = n4970 ^ n2827 ;
  assign n4964 = n689 ^ n255 ;
  assign n4965 = n4964 ^ n728 ;
  assign n4962 = n520 ^ n226 ;
  assign n4961 = n2982 ^ n505 ;
  assign n4963 = n4962 ^ n4961 ;
  assign n4966 = n4965 ^ n4963 ;
  assign n4967 = n4966 ^ n4005 ;
  assign n4972 = n4971 ^ n4967 ;
  assign n4986 = n4985 ^ n4972 ;
  assign n5028 = n2864 ^ n914 ;
  assign n5027 = n4765 ^ n322 ;
  assign n5029 = n5028 ^ n5027 ;
  assign n5030 = n5029 ^ n2421 ;
  assign n5023 = n863 ^ n194 ;
  assign n5024 = n5023 ^ n292 ;
  assign n5021 = n961 ^ n355 ;
  assign n5022 = n5021 ^ n641 ;
  assign n5025 = n5024 ^ n5022 ;
  assign n5019 = n5018 ^ n2240 ;
  assign n5017 = n5016 ^ n1359 ;
  assign n5020 = n5019 ^ n5017 ;
  assign n5026 = n5025 ^ n5020 ;
  assign n5031 = n5030 ^ n5026 ;
  assign n5003 = n3787 ^ n737 ;
  assign n5004 = n5003 ^ n2963 ;
  assign n5002 = n3448 ^ n2702 ;
  assign n5005 = n5004 ^ n5002 ;
  assign n5015 = n5014 ^ n5005 ;
  assign n5032 = n5031 ^ n5015 ;
  assign n4997 = n117 ^ n100 ;
  assign n4998 = n4997 ^ n762 ;
  assign n4995 = n1159 ^ n239 ;
  assign n4996 = n4995 ^ n814 ;
  assign n4999 = n4998 ^ n4996 ;
  assign n5000 = n4999 ^ n2092 ;
  assign n4991 = n2408 ^ n1339 ;
  assign n4990 = n3673 ^ n3601 ;
  assign n4992 = n4991 ^ n4990 ;
  assign n4988 = n3972 ^ n2693 ;
  assign n4987 = n4356 ^ n1534 ;
  assign n4989 = n4988 ^ n4987 ;
  assign n4993 = n4992 ^ n4989 ;
  assign n4994 = n4993 ^ n4276 ;
  assign n5001 = n5000 ^ n4994 ;
  assign n5033 = n5032 ^ n5001 ;
  assign n5034 = ~n4986 & ~n5033 ;
  assign n5035 = n5034 ^ x8 ;
  assign n5058 = n970 ^ n559 ;
  assign n5056 = n352 ^ n178 ;
  assign n5054 = n5016 ^ n418 ;
  assign n5055 = n5054 ^ n883 ;
  assign n5057 = n5056 ^ n5055 ;
  assign n5059 = n5058 ^ n5057 ;
  assign n5051 = n1819 ^ n356 ;
  assign n5049 = n5048 ^ n217 ;
  assign n5050 = n5049 ^ n192 ;
  assign n5052 = n5051 ^ n5050 ;
  assign n5046 = n3427 ^ n1836 ;
  assign n5047 = n5046 ^ n2243 ;
  assign n5053 = n5052 ^ n5047 ;
  assign n5060 = n5059 ^ n5053 ;
  assign n5042 = n4121 ^ n219 ;
  assign n5040 = n4294 ^ n1029 ;
  assign n5041 = n5040 ^ n97 ;
  assign n5043 = n5042 ^ n5041 ;
  assign n5044 = n5043 ^ n1971 ;
  assign n5037 = n1042 ^ n478 ;
  assign n5036 = n1188 ^ n183 ;
  assign n5038 = n5037 ^ n5036 ;
  assign n5039 = n5038 ^ n3761 ;
  assign n5045 = n5044 ^ n5039 ;
  assign n5061 = n5060 ^ n5045 ;
  assign n5062 = n5061 ^ n3791 ;
  assign n5083 = n4804 ^ n897 ;
  assign n5084 = n5083 ^ n507 ;
  assign n5082 = n961 ^ n622 ;
  assign n5085 = n5084 ^ n5082 ;
  assign n5086 = n5085 ^ n793 ;
  assign n5087 = n5086 ^ n1389 ;
  assign n5078 = n635 ^ n252 ;
  assign n5079 = n5078 ^ n557 ;
  assign n5076 = n772 ^ n571 ;
  assign n5077 = n5076 ^ n872 ;
  assign n5080 = n5079 ^ n5077 ;
  assign n5074 = n4292 ^ n403 ;
  assign n5075 = n5074 ^ n492 ;
  assign n5081 = n5080 ^ n5075 ;
  assign n5088 = n5087 ^ n5081 ;
  assign n5071 = n1731 ^ n396 ;
  assign n5069 = n662 ^ n414 ;
  assign n5070 = n5069 ^ n4017 ;
  assign n5072 = n5071 ^ n5070 ;
  assign n5065 = n2208 ^ n1002 ;
  assign n5066 = n5065 ^ n1847 ;
  assign n5063 = n2132 ^ n1658 ;
  assign n5064 = n5063 ^ n742 ;
  assign n5067 = n5066 ^ n5064 ;
  assign n5068 = n5067 ^ n619 ;
  assign n5073 = n5072 ^ n5068 ;
  assign n5089 = n5088 ^ n5073 ;
  assign n5090 = ~n5062 & ~n5089 ;
  assign n5091 = n5090 ^ n5034 ;
  assign n5092 = n5035 & ~n5091 ;
  assign n5093 = n5092 ^ x8 ;
  assign n5142 = n5141 ^ n5093 ;
  assign n5154 = ~n35 & ~n2268 ;
  assign n5143 = n3357 ^ n3233 ;
  assign n5144 = n5143 ^ n2268 ;
  assign n5146 = n5144 ^ n2364 ;
  assign n5145 = n5144 ^ n2449 ;
  assign n5147 = n5146 ^ n5145 ;
  assign n5150 = x30 & n5147 ;
  assign n5151 = n5150 ^ n5146 ;
  assign n5152 = ~n3520 & ~n5151 ;
  assign n5153 = n5152 ^ n5144 ;
  assign n5155 = n5154 ^ n5153 ;
  assign n4936 = ~n35 & ~n2364 ;
  assign n4937 = n4936 ^ n2268 ;
  assign n5156 = n5155 ^ n4937 ;
  assign n5157 = n5156 ^ n5153 ;
  assign n5160 = ~n33 & ~n5157 ;
  assign n5161 = n5160 ^ n5153 ;
  assign n5162 = ~x31 & n5161 ;
  assign n5163 = n5162 ^ n5153 ;
  assign n5164 = n5163 ^ n5093 ;
  assign n5165 = ~n5142 & n5164 ;
  assign n5208 = n4851 ^ x31 ;
  assign n5209 = ~n2185 & n5208 ;
  assign n5204 = ~n2096 & n3520 ;
  assign n5198 = ~n35 & ~n2185 ;
  assign n5199 = n5198 ^ n5154 ;
  assign n5205 = n5204 ^ n5199 ;
  assign n5206 = ~x31 & n5205 ;
  assign n5207 = n5206 ^ n5154 ;
  assign n5210 = n5209 ^ n5207 ;
  assign n5195 = n3359 ^ n3235 ;
  assign n5196 = n5195 ^ n2096 ;
  assign n5197 = n5196 & n23912 ;
  assign n5211 = n5210 ^ n5197 ;
  assign n5212 = n5211 ^ n5141 ;
  assign n5213 = n5212 ^ n5211 ;
  assign n4955 = n2586 ^ n798 ;
  assign n4954 = n885 ^ n768 ;
  assign n4956 = n4955 ^ n4954 ;
  assign n4950 = n2111 ^ n612 ;
  assign n4951 = n4950 ^ n841 ;
  assign n4948 = n2912 ^ n751 ;
  assign n4947 = n2890 ^ n780 ;
  assign n4949 = n4948 ^ n4947 ;
  assign n4952 = n4951 ^ n4949 ;
  assign n4944 = n739 ^ n196 ;
  assign n4945 = n4944 ^ n1839 ;
  assign n4941 = n945 ^ n97 ;
  assign n4942 = n4941 ^ n518 ;
  assign n4940 = n1783 ^ n571 ;
  assign n4943 = n4942 ^ n4940 ;
  assign n4946 = n4945 ^ n4943 ;
  assign n4953 = n4952 ^ n4946 ;
  assign n4957 = n4956 ^ n4953 ;
  assign n4958 = n4957 ^ n3886 ;
  assign n4959 = ~n1277 & ~n2267 ;
  assign n4960 = ~n4958 & n4959 ;
  assign n5214 = n5213 ^ n4960 ;
  assign n5215 = n5165 & ~n5214 ;
  assign n5216 = n5215 ^ n5212 ;
  assign n5266 = n5265 ^ n5216 ;
  assign n5192 = ~n1795 & n3484 ;
  assign n5184 = n4859 ^ n1871 ;
  assign n5188 = n4536 & n5184 ;
  assign n5189 = n5188 ^ n1871 ;
  assign n5190 = n650 & ~n5189 ;
  assign n5191 = n5190 ^ x29 ;
  assign n5193 = n5192 ^ n5191 ;
  assign n5183 = n831 & ~n1994 ;
  assign n5194 = n5193 ^ n5183 ;
  assign n5267 = n5266 ^ n5194 ;
  assign n5448 = ~n1871 & n3484 ;
  assign n5444 = n4391 & n4536 ;
  assign n5445 = n5444 ^ n1631 ;
  assign n5446 = n650 & ~n5445 ;
  assign n5447 = n5446 ^ x29 ;
  assign n5449 = n5448 ^ n5447 ;
  assign n5439 = n831 & ~n1795 ;
  assign n5450 = n5449 ^ n5439 ;
  assign n5436 = n5265 ^ n5211 ;
  assign n5437 = ~n5216 & ~n5436 ;
  assign n5438 = n5437 ^ n5265 ;
  assign n5451 = n5450 ^ n5438 ;
  assign n5430 = n5141 ^ x11 ;
  assign n5431 = n5263 ^ n5141 ;
  assign n5432 = n5430 & ~n5431 ;
  assign n5433 = n5432 ^ x11 ;
  assign n5425 = n5198 ^ n4816 ;
  assign n5423 = ~n35 & ~n2096 ;
  assign n5424 = n5423 ^ n4817 ;
  assign n5426 = n5425 ^ n5424 ;
  assign n5408 = n3360 ^ n3236 ;
  assign n5409 = n5408 ^ n1994 ;
  assign n5422 = n3520 & n5409 ;
  assign n5427 = n5426 ^ n5422 ;
  assign n5428 = x31 & n5427 ;
  assign n5429 = n5428 ^ n5424 ;
  assign n5434 = n5433 ^ n5429 ;
  assign n5435 = n5434 ^ n4378 ;
  assign n5452 = n5451 ^ n5435 ;
  assign n5453 = n5452 ^ n5194 ;
  assign n5454 = n5453 ^ n5452 ;
  assign n5166 = n5165 ^ n4960 ;
  assign n4938 = n3720 & ~n4937 ;
  assign n4933 = ~n2185 & n3520 ;
  assign n4930 = n3358 ^ n3234 ;
  assign n4931 = n4930 ^ n2268 ;
  assign n4932 = n4931 & n23912 ;
  assign n4934 = n4933 ^ n4932 ;
  assign n4935 = n4934 ^ n2268 ;
  assign n4939 = n4938 ^ n4935 ;
  assign n5167 = n5166 ^ n4939 ;
  assign n5179 = n831 & ~n2096 ;
  assign n5177 = ~n1994 & n3484 ;
  assign n5175 = n4939 ^ x29 ;
  assign n5172 = ~n4384 & n4536 ;
  assign n5173 = n5172 ^ n1795 ;
  assign n5174 = n650 & ~n5173 ;
  assign n5176 = n5175 ^ n5174 ;
  assign n5178 = n5177 ^ n5176 ;
  assign n5180 = n5179 ^ n5178 ;
  assign n5181 = n5167 & n5180 ;
  assign n5182 = n5181 ^ n5166 ;
  assign n5455 = n5454 ^ n5182 ;
  assign n5456 = ~n5267 & ~n5455 ;
  assign n5457 = n5456 ^ n5453 ;
  assign n5740 = ~n968 & ~n4496 ;
  assign n5739 = ~n1214 & n4504 ;
  assign n5741 = n5740 ^ n5739 ;
  assign n5732 = n1109 ^ x23 ;
  assign n5733 = n5732 ^ x22 ;
  assign n5734 = n5733 ^ n1109 ;
  assign n5735 = ~n3904 & n5734 ;
  assign n5736 = n5735 ^ n1109 ;
  assign n5737 = n4488 & ~n5736 ;
  assign n5738 = n5737 ^ x23 ;
  assign n5742 = n5741 ^ n5738 ;
  assign n5744 = n5742 ^ n5452 ;
  assign n5461 = ~n487 & ~n1433 ;
  assign n5460 = ~n1703 & n12861 ;
  assign n5462 = n5461 ^ n5460 ;
  assign n5463 = n5462 ^ x26 ;
  assign n5459 = n446 & ~n1351 ;
  assign n5464 = n5463 ^ n5459 ;
  assign n5458 = ~n3501 & n4152 ;
  assign n5465 = n5464 ^ n5458 ;
  assign n5743 = n5742 ^ n5465 ;
  assign n5745 = n5744 ^ n5743 ;
  assign n5746 = n5457 & n5745 ;
  assign n5747 = n5746 ^ n5744 ;
  assign n5772 = n656 & ~n1703 ;
  assign n5764 = n446 & ~n1433 ;
  assign n5763 = ~n487 & ~n1540 ;
  assign n5765 = n5764 ^ n5763 ;
  assign n5766 = n5765 ^ x26 ;
  assign n5762 = ~n1351 & n12861 ;
  assign n5767 = n5766 ^ n5762 ;
  assign n4610 = n3817 ^ n1540 ;
  assign n5761 = ~n3501 & ~n4610 ;
  assign n5768 = n5767 ^ n5761 ;
  assign n5769 = n5768 ^ x29 ;
  assign n5760 = n3481 & ~n4615 ;
  assign n5770 = n5769 ^ n5760 ;
  assign n5759 = ~n1631 & n3484 ;
  assign n5771 = n5770 ^ n5759 ;
  assign n5773 = n5772 ^ n5771 ;
  assign n5758 = n831 & ~n1871 ;
  assign n5774 = n5773 ^ n5758 ;
  assign n5748 = n5450 ^ n5429 ;
  assign n5756 = n5451 & ~n5748 ;
  assign n5749 = n5748 ^ n5433 ;
  assign n5750 = n5749 ^ n5438 ;
  assign n5752 = n4840 ^ n4378 ;
  assign n5751 = n5433 ^ n4840 ;
  assign n5753 = n5752 ^ n5751 ;
  assign n5754 = n5750 & n5753 ;
  assign n5755 = n5754 ^ n5752 ;
  assign n5757 = n5756 ^ n5755 ;
  assign n5775 = n5774 ^ n5757 ;
  assign n6001 = n5775 ^ n5742 ;
  assign n6002 = n5747 & ~n6001 ;
  assign n6003 = n6002 ^ n5742 ;
  assign n6004 = n6003 ^ x23 ;
  assign n6006 = n6005 ^ n6004 ;
  assign n6008 = n6007 ^ n6006 ;
  assign n6010 = n6009 ^ n6008 ;
  assign n6012 = n6011 ^ n6010 ;
  assign n5970 = n5768 ^ n5757 ;
  assign n5971 = n5774 & ~n5970 ;
  assign n5972 = n5971 ^ n5768 ;
  assign n5967 = ~n1433 & n12861 ;
  assign n5960 = ~n1703 & n3484 ;
  assign n5956 = n4862 ^ n4303 ;
  assign n5957 = n5956 ^ n4842 ;
  assign n5958 = n5957 ^ x29 ;
  assign n5953 = ~n4416 & n4536 ;
  assign n5954 = n5953 ^ n1351 ;
  assign n5955 = n650 & ~n5954 ;
  assign n5959 = n5958 ^ n5955 ;
  assign n5961 = n5960 ^ n5959 ;
  assign n5947 = n831 & ~n1631 ;
  assign n5962 = n5961 ^ n5947 ;
  assign n5903 = ~n5438 & n5450 ;
  assign n5904 = ~n5433 & n5903 ;
  assign n5905 = ~n4378 & n5429 ;
  assign n5906 = n5904 & n5905 ;
  assign n5907 = n5906 ^ n4378 ;
  assign n5908 = n5438 ^ n5433 ;
  assign n5909 = ~n5749 & n5908 ;
  assign n5910 = n5909 ^ n5433 ;
  assign n5911 = ~n5907 & n5910 ;
  assign n5912 = n5911 ^ n5907 ;
  assign n5913 = n5912 ^ n5429 ;
  assign n5914 = n5913 ^ n5912 ;
  assign n5917 = n5912 ^ n5450 ;
  assign n5918 = n5917 ^ n5912 ;
  assign n5919 = n5911 & n5918 ;
  assign n5920 = n5914 & n5919 ;
  assign n5921 = n5920 ^ n5914 ;
  assign n5922 = n5921 ^ n5913 ;
  assign n5923 = n4840 & ~n5922 ;
  assign n5924 = n5923 ^ n5907 ;
  assign n5925 = n4378 & n4840 ;
  assign n5926 = n5925 ^ n5450 ;
  assign n5927 = n5926 ^ n5925 ;
  assign n5928 = n5925 ^ n5433 ;
  assign n5929 = n5928 ^ n5925 ;
  assign n5930 = ~n5927 & n5929 ;
  assign n5931 = n5930 ^ n5925 ;
  assign n5939 = n5929 ^ n5927 ;
  assign n5940 = n5939 ^ n5925 ;
  assign n5933 = n5925 ^ n5429 ;
  assign n5932 = n5925 ^ n5438 ;
  assign n5934 = n5933 ^ n5932 ;
  assign n5935 = n5932 ^ n5928 ;
  assign n5936 = n5935 ^ n5926 ;
  assign n5937 = n5936 ^ n5925 ;
  assign n5938 = n5934 & ~n5937 ;
  assign n5941 = n5940 ^ n5938 ;
  assign n5942 = n5931 & ~n5941 ;
  assign n5943 = n5942 ^ n5925 ;
  assign n5946 = n5924 & ~n5943 ;
  assign n5963 = n5962 ^ n5946 ;
  assign n5964 = n5963 ^ x26 ;
  assign n5902 = n446 & ~n1540 ;
  assign n5965 = n5964 ^ n5902 ;
  assign n5901 = ~n487 & ~n1214 ;
  assign n5966 = n5965 ^ n5901 ;
  assign n5968 = n5967 ^ n5966 ;
  assign n5900 = ~n3501 & ~n4603 ;
  assign n5969 = n5968 ^ n5900 ;
  assign n6013 = n5972 ^ n5969 ;
  assign n6014 = n6013 ^ n6003 ;
  assign n6015 = ~n6012 & n6014 ;
  assign n6016 = n6015 ^ n6013 ;
  assign n6017 = n6016 ^ x20 ;
  assign n6019 = n6018 ^ n6017 ;
  assign n6021 = n6020 ^ n6019 ;
  assign n6000 = ~n649 & n14027 ;
  assign n6022 = n6021 ^ n6000 ;
  assign n6024 = n6023 ^ n6022 ;
  assign n5996 = ~n1109 & n4504 ;
  assign n5989 = n5957 ^ n5946 ;
  assign n5990 = n5962 & n5989 ;
  assign n5991 = n5990 ^ n5957 ;
  assign n5986 = ~n1540 & n12861 ;
  assign n5982 = n4875 ^ n4867 ;
  assign n5983 = n5982 ^ x26 ;
  assign n5981 = n446 & ~n1214 ;
  assign n5984 = n5983 ^ n5981 ;
  assign n5980 = ~n487 & ~n968 ;
  assign n5985 = n5984 ^ n5980 ;
  assign n5987 = n5986 ^ n5985 ;
  assign n5979 = ~n3501 & n3521 ;
  assign n5988 = n5987 ^ n5979 ;
  assign n5992 = n5991 ^ n5988 ;
  assign n5993 = n5992 ^ x23 ;
  assign n5978 = ~n3508 & n4492 ;
  assign n5994 = n5993 ^ n5978 ;
  assign n5977 = ~n824 & ~n4496 ;
  assign n5995 = n5994 ^ n5977 ;
  assign n5997 = n5996 ^ n5995 ;
  assign n5976 = ~n3473 & n4491 ;
  assign n5998 = n5997 ^ n5976 ;
  assign n5973 = n5972 ^ n5963 ;
  assign n5974 = n5969 & n5973 ;
  assign n5975 = n5974 ^ n5963 ;
  assign n5999 = n5998 ^ n5975 ;
  assign n11640 = n6016 ^ n5999 ;
  assign n11641 = n6024 & n11640 ;
  assign n11642 = n11641 ^ n6016 ;
  assign n4897 = x12 ^ x11 ;
  assign n4896 = ~x11 & ~x12 ;
  assign n4898 = n4897 ^ n4896 ;
  assign n4906 = n4896 ^ x14 ;
  assign n4907 = n4896 ^ x13 ;
  assign n4908 = ~n4906 & n4907 ;
  assign n4909 = ~n3943 & n4908 ;
  assign n4903 = ~x13 & ~n3943 ;
  assign n4904 = n4903 ^ x14 ;
  assign n4905 = ~n3920 & ~n4904 ;
  assign n4910 = n4909 ^ n4905 ;
  assign n4911 = n4898 & n4910 ;
  assign n5780 = n4909 ^ x14 ;
  assign n5783 = n4911 & n5780 ;
  assign n5776 = n5775 ^ n5747 ;
  assign n5725 = ~n824 & n14027 ;
  assign n5724 = ~n3473 & n4916 ;
  assign n5726 = n5725 ^ n5724 ;
  assign n5727 = n5726 ^ x20 ;
  assign n5723 = ~n649 & n4683 ;
  assign n5728 = n5727 ^ n5723 ;
  assign n5722 = ~n3476 & n4684 ;
  assign n5729 = n5728 ^ n5722 ;
  assign n5472 = ~n968 & n4491 ;
  assign n5471 = ~n1214 & ~n4496 ;
  assign n5473 = n5472 ^ n5471 ;
  assign n5468 = ~n1540 & n4504 ;
  assign n5467 = n3521 & n4492 ;
  assign n5469 = n5468 ^ n5467 ;
  assign n5470 = n5469 ^ x23 ;
  assign n5474 = n5473 ^ n5470 ;
  assign n5730 = n5729 ^ n5474 ;
  assign n5466 = n5465 ^ n5457 ;
  assign n5475 = n5474 ^ n5466 ;
  assign n5268 = n5267 ^ n5182 ;
  assign n4925 = ~n1631 & n12861 ;
  assign n4924 = n446 & ~n1703 ;
  assign n4926 = n4925 ^ n4924 ;
  assign n4927 = n4926 ^ x26 ;
  assign n4923 = ~n487 & ~n1351 ;
  assign n4928 = n4927 ^ n4923 ;
  assign n4922 = ~n3501 & n4417 ;
  assign n4929 = n4928 ^ n4922 ;
  assign n5269 = n5268 ^ n4929 ;
  assign n5274 = n446 & ~n1631 ;
  assign n5273 = ~n487 & ~n1703 ;
  assign n5275 = n5274 ^ n5273 ;
  assign n5276 = n5275 ^ x26 ;
  assign n5272 = ~n1871 & n12861 ;
  assign n5277 = n5276 ^ n5272 ;
  assign n5271 = ~n3501 & ~n4615 ;
  assign n5278 = n5277 ^ n5271 ;
  assign n5270 = n5180 ^ n5166 ;
  assign n5279 = n5278 ^ n5270 ;
  assign n5402 = n5163 ^ n5142 ;
  assign n5281 = x31 ^ x30 ;
  assign n5294 = ~n2449 & n5281 ;
  assign n5287 = ~x31 & ~n2364 ;
  assign n5295 = n5294 ^ n5287 ;
  assign n5296 = ~n3520 & n5295 ;
  assign n5285 = ~n2486 & n24214 ;
  assign n5282 = n3356 ^ n3232 ;
  assign n5283 = n5282 ^ n2364 ;
  assign n5284 = n5283 & n23912 ;
  assign n5286 = n5285 ^ n5284 ;
  assign n5288 = n5287 ^ n5286 ;
  assign n5297 = n5296 ^ n5288 ;
  assign n5280 = n5090 ^ n5035 ;
  assign n5298 = n5297 ^ n5280 ;
  assign n5323 = n5085 ^ n5005 ;
  assign n5319 = n977 ^ n401 ;
  assign n5320 = n5319 ^ n918 ;
  assign n5317 = n809 ^ n218 ;
  assign n5318 = n5317 ^ n274 ;
  assign n5321 = n5320 ^ n5318 ;
  assign n5315 = n3583 ^ n1247 ;
  assign n5314 = n5076 ^ n1075 ;
  assign n5316 = n5315 ^ n5314 ;
  assign n5322 = n5321 ^ n5316 ;
  assign n5324 = n5323 ^ n5322 ;
  assign n5309 = n1987 ^ n853 ;
  assign n5310 = n5309 ^ n1021 ;
  assign n5307 = n5078 ^ n3408 ;
  assign n5308 = n5307 ^ n1597 ;
  assign n5311 = n5310 ^ n5308 ;
  assign n5304 = n797 ^ n417 ;
  assign n5301 = n3664 ^ n249 ;
  assign n5302 = n5301 ^ n697 ;
  assign n5303 = n5302 ^ n391 ;
  assign n5305 = n5304 ^ n5303 ;
  assign n5299 = n2208 ^ n2069 ;
  assign n5300 = n5299 ^ n766 ;
  assign n5306 = n5305 ^ n5300 ;
  assign n5312 = n5311 ^ n5306 ;
  assign n5313 = n5312 ^ n1315 ;
  assign n5325 = n5324 ^ n5313 ;
  assign n5326 = ~n3659 & ~n5325 ;
  assign n5327 = n5326 ^ n5034 ;
  assign n5328 = x5 ^ x2 ;
  assign n5347 = n917 ^ n804 ;
  assign n5343 = n1020 ^ n867 ;
  assign n5341 = n2474 ^ n181 ;
  assign n5342 = n5341 ^ n3046 ;
  assign n5344 = n5343 ^ n5342 ;
  assign n5345 = n5344 ^ n728 ;
  assign n5339 = n3263 ^ n963 ;
  assign n5336 = n5335 ^ n330 ;
  assign n5332 = n621 ^ n156 ;
  assign n5334 = n5333 ^ n5332 ;
  assign n5337 = n5336 ^ n5334 ;
  assign n5330 = n627 ^ n237 ;
  assign n5329 = n1373 ^ n258 ;
  assign n5331 = n5330 ^ n5329 ;
  assign n5338 = n5337 ^ n5331 ;
  assign n5340 = n5339 ^ n5338 ;
  assign n5346 = n5345 ^ n5340 ;
  assign n5348 = n5347 ^ n5346 ;
  assign n5374 = n5373 ^ n5348 ;
  assign n5375 = ~n4259 & ~n5374 ;
  assign n5376 = n5375 ^ x5 ;
  assign n5377 = n5328 & ~n5376 ;
  assign n5378 = n5377 ^ x2 ;
  assign n5379 = n5378 ^ n5034 ;
  assign n5391 = ~n2554 & ~n3733 ;
  assign n5390 = ~n2609 & n24214 ;
  assign n5392 = n5391 ^ n5390 ;
  assign n5380 = n3354 ^ n3230 ;
  assign n5387 = x31 & ~n5380 ;
  assign n5388 = n5387 ^ n2486 ;
  assign n5389 = n3520 & ~n5388 ;
  assign n5393 = n5392 ^ n5389 ;
  assign n5394 = n5393 ^ n5378 ;
  assign n5395 = ~n5379 & n5394 ;
  assign n5396 = ~n5327 & n5395 ;
  assign n5397 = n5396 ^ n5034 ;
  assign n5398 = n5397 ^ n5297 ;
  assign n5399 = ~n5298 & n5398 ;
  assign n5400 = n5399 ^ n5297 ;
  assign n5403 = n5402 ^ n5400 ;
  assign n5412 = ~n2096 & n3484 ;
  assign n5410 = n3481 & n5409 ;
  assign n5405 = n831 & ~n2185 ;
  assign n5404 = n656 & ~n1994 ;
  assign n5406 = n5405 ^ n5404 ;
  assign n5407 = n5406 ^ x29 ;
  assign n5411 = n5410 ^ n5407 ;
  assign n5413 = n5412 ^ n5411 ;
  assign n5414 = n5413 ^ n5400 ;
  assign n5415 = ~n5403 & n5414 ;
  assign n5401 = n5400 ^ n5270 ;
  assign n5416 = n5415 ^ n5401 ;
  assign n5417 = n5279 & ~n5416 ;
  assign n5418 = n5417 ^ n5278 ;
  assign n5419 = n5418 ^ n4929 ;
  assign n5420 = n5269 & n5419 ;
  assign n5421 = n5420 ^ n4929 ;
  assign n5720 = n5474 ^ n5421 ;
  assign n5721 = n5475 & n5720 ;
  assign n5731 = n5730 ^ n5721 ;
  assign n5777 = n5776 ^ n5731 ;
  assign n5693 = x15 ^ x14 ;
  assign n24304 = x16 & n5693 ;
  assign n17163 = x17 & n5693 ;
  assign n5696 = n17163 ^ n5693 ;
  assign n5702 = n24304 ^ n5696 ;
  assign n5715 = ~n485 & n5702 ;
  assign n5699 = x16 ^ x15 ;
  assign n5700 = ~n5693 & n5699 ;
  assign n5714 = ~n445 & n5700 ;
  assign n5716 = n5715 ^ n5714 ;
  assign n5717 = n5716 ^ x17 ;
  assign n5705 = n5700 ^ n5693 ;
  assign n5697 = x14 & x15 ;
  assign n5706 = x16 & n5697 ;
  assign n20726 = n5706 ^ x17 ;
  assign n5707 = n5706 ^ n5705 ;
  assign n20727 = n20726 ^ n5707 ;
  assign n20730 = ~n5705 & n20727 ;
  assign n20731 = n20730 ^ n5706 ;
  assign n5713 = ~n317 & n20731 ;
  assign n5718 = n5717 ^ n5713 ;
  assign n5703 = n5702 ^ n5693 ;
  assign n5704 = n3500 & n5703 ;
  assign n5719 = n5718 ^ n5704 ;
  assign n5778 = n5777 ^ n5719 ;
  assign n5476 = n5475 ^ n5421 ;
  assign n4917 = ~n824 & n4916 ;
  assign n4914 = ~n3473 & n4683 ;
  assign n4918 = n4917 ^ n4914 ;
  assign n4919 = n4918 ^ x20 ;
  assign n4913 = ~n1109 & n14027 ;
  assign n4920 = n4919 ^ n4913 ;
  assign n4912 = ~n3508 & n4684 ;
  assign n4921 = n4920 ^ n4912 ;
  assign n5477 = n5476 ^ n4921 ;
  assign n5481 = n5418 ^ n5269 ;
  assign n5689 = n5481 ^ n4921 ;
  assign n5485 = ~n1214 & n4491 ;
  assign n5482 = n5481 ^ x23 ;
  assign n5480 = n4492 & ~n4603 ;
  assign n5483 = n5482 ^ n5480 ;
  assign n5479 = ~n1540 & ~n4496 ;
  assign n5484 = n5483 ^ n5479 ;
  assign n5486 = n5485 ^ n5484 ;
  assign n5478 = ~n1433 & n4504 ;
  assign n5487 = n5486 ^ n5478 ;
  assign n5494 = ~n1433 & ~n4496 ;
  assign n5493 = ~n1540 & n4491 ;
  assign n5495 = n5494 ^ n5493 ;
  assign n5490 = ~n1351 & n4504 ;
  assign n5489 = n4492 & ~n4610 ;
  assign n5491 = n5490 ^ n5489 ;
  assign n5492 = n5491 ^ x23 ;
  assign n5496 = n5495 ^ n5492 ;
  assign n5488 = n5416 ^ n5278 ;
  assign n5497 = n5496 ^ n5488 ;
  assign n5506 = n5413 ^ n5403 ;
  assign n5501 = n446 & ~n1871 ;
  assign n5500 = ~n1795 & n12861 ;
  assign n5502 = n5501 ^ n5500 ;
  assign n5503 = n5502 ^ x26 ;
  assign n5499 = ~n487 & ~n1631 ;
  assign n5504 = n5503 ^ n5499 ;
  assign n5498 = ~n3501 & ~n4392 ;
  assign n5505 = n5504 ^ n5498 ;
  assign n5507 = n5506 ^ n5505 ;
  assign n5516 = n5397 ^ n5298 ;
  assign n5514 = ~n2185 & n3484 ;
  assign n5512 = n3481 & n5196 ;
  assign n5509 = n831 & ~n2268 ;
  assign n5508 = n656 & ~n2096 ;
  assign n5510 = n5509 ^ n5508 ;
  assign n5511 = n5510 ^ x29 ;
  assign n5513 = n5512 ^ n5511 ;
  assign n5515 = n5514 ^ n5513 ;
  assign n5517 = n5516 ^ n5515 ;
  assign n5525 = ~n2486 & ~n3733 ;
  assign n5524 = ~n2449 & n3726 ;
  assign n5526 = n5525 ^ n5524 ;
  assign n5522 = ~n2554 & n24214 ;
  assign n5519 = n3355 ^ n3231 ;
  assign n5520 = n5519 ^ n2449 ;
  assign n5521 = n5520 & n23912 ;
  assign n5523 = n5522 ^ n5521 ;
  assign n5527 = n5526 ^ n5523 ;
  assign n5518 = n5395 ^ n5326 ;
  assign n5528 = n5527 ^ n5518 ;
  assign n5536 = ~n2364 & n3484 ;
  assign n5534 = n3481 & n5144 ;
  assign n5531 = n656 & ~n2268 ;
  assign n5530 = n831 & ~n2449 ;
  assign n5532 = n5531 ^ n5530 ;
  assign n5533 = n5532 ^ x29 ;
  assign n5535 = n5534 ^ n5533 ;
  assign n5537 = n5536 ^ n5535 ;
  assign n5674 = n5537 ^ n5527 ;
  assign n5529 = n5393 ^ n5379 ;
  assign n5538 = n5537 ^ n5529 ;
  assign n5551 = ~n2609 & ~n3733 ;
  assign n5550 = ~n3227 & n24214 ;
  assign n5552 = n5551 ^ n5550 ;
  assign n5540 = n3353 ^ n3229 ;
  assign n5547 = x31 & ~n5540 ;
  assign n5548 = n5547 ^ n2554 ;
  assign n5549 = n3520 & ~n5548 ;
  assign n5553 = n5552 ^ n5549 ;
  assign n5671 = n5553 ^ n5537 ;
  assign n5539 = n5375 ^ n5328 ;
  assign n5554 = n5553 ^ n5539 ;
  assign n5613 = n3799 ^ n1387 ;
  assign n5614 = n5613 ^ n3602 ;
  assign n5615 = n5614 ^ n870 ;
  assign n5610 = n5078 ^ n393 ;
  assign n5611 = n5610 ^ n2072 ;
  assign n5612 = n5611 ^ n4325 ;
  assign n5616 = n5615 ^ n5612 ;
  assign n5597 = n1450 ^ n662 ;
  assign n5596 = n5595 ^ n3596 ;
  assign n5598 = n5597 ^ n5596 ;
  assign n5593 = n456 ^ n104 ;
  assign n5591 = n1254 ^ n940 ;
  assign n5592 = n5591 ^ n237 ;
  assign n5594 = n5593 ^ n5592 ;
  assign n5599 = n5598 ^ n5594 ;
  assign n5609 = n5608 ^ n5599 ;
  assign n5617 = n5616 ^ n5609 ;
  assign n5618 = n5617 ^ n1187 ;
  assign n5619 = ~n3062 & ~n5618 ;
  assign n5585 = n4950 ^ n2964 ;
  assign n5586 = n5585 ^ n2354 ;
  assign n5587 = n5586 ^ n5029 ;
  assign n5582 = n2536 ^ n1054 ;
  assign n5583 = n5582 ^ n940 ;
  assign n5580 = n1180 ^ n1039 ;
  assign n5578 = n974 ^ n814 ;
  assign n5579 = n5578 ^ n3431 ;
  assign n5581 = n5580 ^ n5579 ;
  assign n5584 = n5583 ^ n5581 ;
  assign n5588 = n5587 ^ n5584 ;
  assign n5566 = n5565 ^ n3318 ;
  assign n5568 = n5567 ^ n5566 ;
  assign n5562 = n2474 ^ n589 ;
  assign n5560 = n4941 ^ n175 ;
  assign n5561 = n5560 ^ n408 ;
  assign n5563 = n5562 ^ n5561 ;
  assign n5557 = n512 ^ n109 ;
  assign n5558 = n5557 ^ n785 ;
  assign n5555 = n623 ^ n130 ;
  assign n5556 = n5555 ^ n161 ;
  assign n5559 = n5558 ^ n5556 ;
  assign n5564 = n5563 ^ n5559 ;
  assign n5569 = n5568 ^ n5564 ;
  assign n5576 = n5575 ^ n5569 ;
  assign n5577 = n5576 ^ n3281 ;
  assign n5589 = n5588 ^ n5577 ;
  assign n5590 = ~n1993 & ~n5589 ;
  assign n5620 = n5619 ^ n5590 ;
  assign n5621 = n2881 ^ n723 ;
  assign n5640 = n1039 ^ n455 ;
  assign n5641 = n5640 ^ n625 ;
  assign n5639 = n790 ^ n190 ;
  assign n5642 = n5641 ^ n5639 ;
  assign n5637 = n1387 ^ n522 ;
  assign n5638 = n5637 ^ n5238 ;
  assign n5643 = n5642 ^ n5638 ;
  assign n5635 = n978 ^ n786 ;
  assign n5633 = n5632 ^ n181 ;
  assign n5630 = n1180 ^ n541 ;
  assign n5634 = n5633 ^ n5630 ;
  assign n5636 = n5635 ^ n5634 ;
  assign n5644 = n5643 ^ n5636 ;
  assign n5625 = n627 ^ n279 ;
  assign n5626 = n5625 ^ n751 ;
  assign n5627 = n5626 ^ n2436 ;
  assign n5622 = n1471 ^ n197 ;
  assign n5623 = n5622 ^ n3390 ;
  assign n5624 = n5623 ^ n525 ;
  assign n5628 = n5627 ^ n5624 ;
  assign n5629 = n5628 ^ n1854 ;
  assign n5645 = n5644 ^ n5629 ;
  assign n5646 = n5645 ^ n3211 ;
  assign n5647 = ~n5621 & ~n5646 ;
  assign n5648 = n5647 ^ n5619 ;
  assign n5649 = n5590 ^ x2 ;
  assign n5660 = ~n35 & ~n2646 ;
  assign n5661 = n5660 ^ n2836 ;
  assign n5662 = ~n5661 & ~n24214 ;
  assign n5656 = ~n35 & ~n2738 ;
  assign n5657 = n5656 ^ n2646 ;
  assign n5658 = ~n3514 & ~n5657 ;
  assign n5653 = ~n2738 & n5208 ;
  assign n5650 = n3350 ^ n3154 ;
  assign n5651 = n5650 ^ n2646 ;
  assign n5652 = ~n5651 & n23912 ;
  assign n5654 = n5653 ^ n5652 ;
  assign n5655 = n5654 ^ n2836 ;
  assign n5659 = n5658 ^ n5655 ;
  assign n5663 = n5662 ^ n5659 ;
  assign n5664 = n5663 ^ n5590 ;
  assign n5665 = ~n5649 & ~n5664 ;
  assign n5666 = ~n5648 & n5665 ;
  assign n5667 = ~n5620 & n5666 ;
  assign n5668 = n5667 ^ x2 ;
  assign n5669 = n5668 ^ n5553 ;
  assign n5670 = ~n5554 & n5669 ;
  assign n5672 = n5671 ^ n5670 ;
  assign n5673 = ~n5538 & n5672 ;
  assign n5675 = n5674 ^ n5673 ;
  assign n5676 = ~n5528 & n5675 ;
  assign n5677 = n5676 ^ n5527 ;
  assign n5678 = n5677 ^ n5515 ;
  assign n5679 = ~n5517 & n5678 ;
  assign n5680 = n5679 ^ n5515 ;
  assign n5681 = n5680 ^ n5505 ;
  assign n5682 = ~n5507 & n5681 ;
  assign n5683 = n5682 ^ n5505 ;
  assign n5684 = n5683 ^ n5496 ;
  assign n5685 = n5497 & n5684 ;
  assign n5686 = n5685 ^ n5496 ;
  assign n5687 = n5686 ^ n5481 ;
  assign n5688 = n5487 & n5687 ;
  assign n5690 = n5689 ^ n5688 ;
  assign n5691 = n5477 & ~n5690 ;
  assign n5692 = n5691 ^ n5476 ;
  assign n5779 = n5778 ^ n5692 ;
  assign n5781 = n5780 ^ n5779 ;
  assign n5784 = n5783 ^ n5781 ;
  assign n5793 = ~n968 & n14027 ;
  assign n5789 = n5686 ^ n5487 ;
  assign n5790 = n5789 ^ x20 ;
  assign n5788 = ~n1109 & n4916 ;
  assign n5791 = n5790 ^ n5788 ;
  assign n5787 = ~n824 & n4683 ;
  assign n5792 = n5791 ^ n5787 ;
  assign n5794 = n5793 ^ n5792 ;
  assign n5786 = ~n4050 & n4684 ;
  assign n5795 = n5794 ^ n5786 ;
  assign n5804 = n5683 ^ n5497 ;
  assign n5799 = ~n1109 & n4683 ;
  assign n5798 = ~n1214 & n14027 ;
  assign n5800 = n5799 ^ n5798 ;
  assign n5801 = n5800 ^ x20 ;
  assign n5797 = ~n968 & n4916 ;
  assign n5802 = n5801 ^ n5797 ;
  assign n5796 = n3905 & n4684 ;
  assign n5803 = n5802 ^ n5796 ;
  assign n5805 = n5804 ^ n5803 ;
  assign n5818 = n5680 ^ n5507 ;
  assign n5857 = n5818 ^ n5804 ;
  assign n5815 = ~n1703 & n4504 ;
  assign n5814 = ~n1351 & ~n4496 ;
  assign n5816 = n5815 ^ n5814 ;
  assign n5807 = n1433 ^ x22 ;
  assign n5808 = n5807 ^ x23 ;
  assign n5809 = n5808 ^ n1433 ;
  assign n5810 = ~n3815 & n5809 ;
  assign n5811 = n5810 ^ n1433 ;
  assign n5812 = n4488 & ~n5811 ;
  assign n5813 = n5812 ^ x23 ;
  assign n5817 = n5816 ^ n5813 ;
  assign n5819 = n5818 ^ n5817 ;
  assign n5842 = n5677 ^ n5517 ;
  assign n5854 = n5842 ^ n5817 ;
  assign n5835 = ~n2268 & n3484 ;
  assign n5832 = n4930 ^ n2185 ;
  assign n5833 = n3481 & n5832 ;
  assign n5829 = n656 & ~n2185 ;
  assign n5828 = n831 & ~n2364 ;
  assign n5830 = n5829 ^ n5828 ;
  assign n5831 = n5830 ^ x29 ;
  assign n5834 = n5833 ^ n5831 ;
  assign n5836 = n5835 ^ n5834 ;
  assign n5823 = ~n2096 & n12861 ;
  assign n5822 = n446 & ~n1994 ;
  assign n5824 = n5823 ^ n5822 ;
  assign n5825 = n5824 ^ x26 ;
  assign n5821 = ~n487 & ~n1795 ;
  assign n5826 = n5825 ^ n5821 ;
  assign n5168 = n4384 ^ n1795 ;
  assign n5820 = ~n3501 & n5168 ;
  assign n5827 = n5826 ^ n5820 ;
  assign n5837 = n5836 ^ n5827 ;
  assign n5838 = n5675 ^ n5518 ;
  assign n5839 = n5838 ^ n5836 ;
  assign n5840 = n5837 & ~n5839 ;
  assign n5841 = n5840 ^ n5836 ;
  assign n5843 = n5842 ^ n5841 ;
  assign n5850 = ~n1994 & n12861 ;
  assign n5848 = ~n487 & ~n1871 ;
  assign n5846 = n446 & ~n1795 ;
  assign n5845 = n5842 ^ x26 ;
  assign n5847 = n5846 ^ n5845 ;
  assign n5849 = n5848 ^ n5847 ;
  assign n5851 = n5850 ^ n5849 ;
  assign n5844 = ~n3501 & ~n4859 ;
  assign n5852 = n5851 ^ n5844 ;
  assign n5853 = ~n5843 & ~n5852 ;
  assign n5855 = n5854 ^ n5853 ;
  assign n5856 = ~n5819 & n5855 ;
  assign n5858 = n5857 ^ n5856 ;
  assign n5859 = n5805 & ~n5858 ;
  assign n5860 = n5859 ^ n5804 ;
  assign n5861 = n5860 ^ n5789 ;
  assign n5862 = n5795 & n5861 ;
  assign n5863 = n5862 ^ n5789 ;
  assign n5785 = n5690 ^ n5476 ;
  assign n5864 = n5863 ^ n5785 ;
  assign n5866 = ~n317 & n5700 ;
  assign n5865 = ~n649 & n20731 ;
  assign n5867 = n5866 ^ n5865 ;
  assign n5694 = x17 & ~n5693 ;
  assign n5875 = n5867 ^ n5694 ;
  assign n5881 = n5875 ^ n5785 ;
  assign n5868 = n5867 ^ x17 ;
  assign n5876 = n5868 ^ n445 ;
  assign n5869 = n5868 ^ x16 ;
  assign n5870 = ~n4072 & n5869 ;
  assign n5877 = n5876 ^ n5870 ;
  assign n5871 = n5870 ^ n445 ;
  assign n5872 = n5868 ^ n5696 ;
  assign n5873 = ~n5871 & ~n5872 ;
  assign n5878 = n5877 ^ n5873 ;
  assign n5879 = ~n5875 & ~n5878 ;
  assign n5882 = n5881 ^ n5879 ;
  assign n5884 = n5864 & ~n5882 ;
  assign n5885 = n5884 ^ n5863 ;
  assign n5886 = n5885 ^ n5779 ;
  assign n5887 = ~n5784 & ~n5886 ;
  assign n5888 = n5887 ^ n5779 ;
  assign n5895 = n3944 & n5693 ;
  assign n5893 = ~n485 & n5700 ;
  assign n5891 = ~n445 & n20731 ;
  assign n5890 = n5888 ^ x17 ;
  assign n5892 = n5891 ^ n5890 ;
  assign n5894 = n5893 ^ n5892 ;
  assign n5896 = n5895 ^ n5894 ;
  assign n5889 = ~n3924 & n5702 ;
  assign n5897 = n5896 ^ n5889 ;
  assign n5898 = ~n5888 & n5897 ;
  assign n5899 = n5898 ^ n5897 ;
  assign n6046 = ~n485 & n20731 ;
  assign n6044 = ~n3943 & n5700 ;
  assign n6031 = n5776 ^ n5729 ;
  assign n6032 = ~n5731 & ~n6031 ;
  assign n6033 = n6032 ^ n5776 ;
  assign n6034 = n6033 ^ x20 ;
  assign n6030 = ~n3473 & n14027 ;
  assign n6035 = n6034 ^ n6030 ;
  assign n6029 = ~n317 & n4683 ;
  assign n6036 = n6035 ^ n6029 ;
  assign n6028 = ~n649 & n4916 ;
  assign n6037 = n6036 ^ n6028 ;
  assign n6027 = n3956 & n4684 ;
  assign n6038 = n6037 ^ n6027 ;
  assign n6039 = n6013 ^ n6012 ;
  assign n6040 = n6039 ^ n6033 ;
  assign n6041 = n6038 & ~n6040 ;
  assign n6042 = n6041 ^ n6039 ;
  assign n6043 = n6042 ^ x17 ;
  assign n6045 = n6044 ^ n6043 ;
  assign n6047 = n6046 ^ n6045 ;
  assign n6026 = n4515 & n5703 ;
  assign n6048 = n6047 ^ n6026 ;
  assign n6025 = n6024 ^ n5999 ;
  assign n6049 = n6048 ^ n6025 ;
  assign n6053 = n6039 ^ n6038 ;
  assign n6050 = n5719 ^ n5692 ;
  assign n6051 = ~n5778 & n6050 ;
  assign n6052 = n6051 ^ n5719 ;
  assign n6054 = n6053 ^ n6052 ;
  assign n11611 = n5885 ^ n5784 ;
  assign n6648 = x9 ^ x8 ;
  assign n6656 = x11 & n6648 ;
  assign n6645 = x8 & x9 ;
  assign n6647 = n6645 ^ x10 ;
  assign n15412 = n6656 ^ n6647 ;
  assign n6649 = x10 & n6648 ;
  assign n6650 = n6649 ^ n6647 ;
  assign n15413 = n15412 ^ n6650 ;
  assign n6664 = ~n3920 & n15413 ;
  assign n16288 = x10 ^ x9 ;
  assign n16289 = ~n6648 & ~n16288 ;
  assign n16290 = n16289 ^ x11 ;
  assign n6652 = ~x11 & ~n16289 ;
  assign n6646 = x10 & n6645 ;
  assign n6653 = n6652 ^ n6646 ;
  assign n6655 = ~n16290 ^ n6653 ;
  assign n6665 = n6664 ^ n6655 ;
  assign n6666 = ~n3943 & n6665 ;
  assign n6667 = n6666 ^ x11 ;
  assign n6565 = ~n824 & n5700 ;
  assign n6121 = ~n1703 & ~n4496 ;
  assign n6118 = n5852 ^ n5841 ;
  assign n6119 = n6118 ^ x23 ;
  assign n6115 = ~n4416 & n4700 ;
  assign n6116 = n6115 ^ n1351 ;
  assign n6117 = n4488 & ~n6116 ;
  assign n6120 = n6119 ^ n6117 ;
  assign n6122 = n6121 ^ n6120 ;
  assign n6112 = ~n1631 & n4504 ;
  assign n6123 = n6122 ^ n6112 ;
  assign n6131 = ~n1703 & n4491 ;
  assign n6127 = n5839 ^ n5827 ;
  assign n6128 = n6127 ^ x23 ;
  assign n6126 = n4492 & ~n4615 ;
  assign n6129 = n6128 ^ n6126 ;
  assign n6125 = ~n1871 & n4504 ;
  assign n6130 = n6129 ^ n6125 ;
  assign n6132 = n6131 ^ n6130 ;
  assign n6124 = ~n1631 & ~n4496 ;
  assign n6133 = n6132 ^ n6124 ;
  assign n6145 = n5672 ^ n5529 ;
  assign n6141 = ~n2185 & n12861 ;
  assign n6140 = n446 & ~n2096 ;
  assign n6142 = n6141 ^ n6140 ;
  assign n6143 = n6142 ^ x26 ;
  assign n6137 = n467 & ~n5408 ;
  assign n6138 = n6137 ^ n1994 ;
  assign n6139 = n64 & ~n6138 ;
  assign n6144 = n6143 ^ n6139 ;
  assign n6146 = n6145 ^ n6144 ;
  assign n6155 = n5668 ^ n5554 ;
  assign n6153 = ~n2449 & n3484 ;
  assign n6151 = n3481 & n5283 ;
  assign n6148 = n831 & ~n2486 ;
  assign n6147 = n656 & ~n2364 ;
  assign n6149 = n6148 ^ n6147 ;
  assign n6150 = n6149 ^ x29 ;
  assign n6152 = n6151 ^ n6150 ;
  assign n6154 = n6153 ^ n6152 ;
  assign n6156 = n6155 ^ n6154 ;
  assign n6171 = n3352 ^ n3228 ;
  assign n6172 = ~n6171 & n23912 ;
  assign n6170 = ~n2609 & n3520 ;
  assign n6173 = n6172 ^ n6170 ;
  assign n6166 = ~n3227 & ~n3725 ;
  assign n6167 = n6166 ^ n5660 ;
  assign n6168 = ~n3732 & n6167 ;
  assign n6157 = n5663 ^ n5619 ;
  assign n6158 = n5665 & ~n6157 ;
  assign n6159 = n6158 ^ n5647 ;
  assign n6160 = n6159 ^ n5660 ;
  assign n6169 = n6168 ^ n6160 ;
  assign n6174 = n6173 ^ n6169 ;
  assign n6183 = n5665 ^ n5619 ;
  assign n6181 = n3720 & ~n5657 ;
  assign n6176 = n3351 ^ n3155 ;
  assign n6177 = n6176 ^ n2646 ;
  assign n6178 = n6177 & n23912 ;
  assign n6175 = ~n3227 & n3520 ;
  assign n6179 = n6178 ^ n6175 ;
  assign n6180 = n6179 ^ n2646 ;
  assign n6182 = n6181 ^ n6180 ;
  assign n6184 = n6183 ^ n6182 ;
  assign n6192 = ~n2609 & n3484 ;
  assign n5541 = n5540 ^ n2554 ;
  assign n6190 = n3481 & n5541 ;
  assign n6187 = n656 & ~n2554 ;
  assign n6186 = n831 & ~n3227 ;
  assign n6188 = n6187 ^ n6186 ;
  assign n6189 = n6188 ^ x29 ;
  assign n6191 = n6190 ^ n6189 ;
  assign n6193 = n6192 ^ n6191 ;
  assign n6519 = n6193 ^ n6182 ;
  assign n6185 = n5663 ^ n5649 ;
  assign n6194 = n6193 ^ n6185 ;
  assign n6215 = n2358 ^ n1099 ;
  assign n6216 = n6215 ^ n5365 ;
  assign n6217 = n6216 ^ n5591 ;
  assign n6212 = n911 ^ n804 ;
  assign n6213 = n6212 ^ n2301 ;
  assign n6206 = n396 ^ n325 ;
  assign n6207 = n6206 ^ n841 ;
  assign n6210 = n6209 ^ n6207 ;
  assign n6204 = n2466 ^ n1219 ;
  assign n6202 = n1806 ^ n203 ;
  assign n6203 = n6202 ^ n1272 ;
  assign n6205 = n6204 ^ n6203 ;
  assign n6211 = n6210 ^ n6205 ;
  assign n6214 = n6213 ^ n6211 ;
  assign n6218 = n6217 ^ n6214 ;
  assign n6219 = n6218 ^ n4247 ;
  assign n6229 = n4282 ^ n2077 ;
  assign n6230 = n6229 ^ n1634 ;
  assign n6231 = n6230 ^ n4320 ;
  assign n6225 = n1130 ^ n261 ;
  assign n6226 = n6225 ^ n1739 ;
  assign n6224 = n1331 ^ n371 ;
  assign n6227 = n6226 ^ n6224 ;
  assign n6222 = n932 ^ n225 ;
  assign n6220 = n744 ^ n635 ;
  assign n6221 = n6220 ^ n613 ;
  assign n6223 = n6222 ^ n6221 ;
  assign n6228 = n6227 ^ n6223 ;
  assign n6232 = n6231 ^ n6228 ;
  assign n6233 = n6232 ^ n2407 ;
  assign n6234 = n6233 ^ n4300 ;
  assign n6235 = ~n6219 & ~n6234 ;
  assign n6199 = ~n2836 & ~n3733 ;
  assign n6198 = ~n3151 & n24214 ;
  assign n6200 = n6199 ^ n6198 ;
  assign n6196 = n3347 & n23912 ;
  assign n6195 = ~n2738 & n3520 ;
  assign n6197 = n6196 ^ n6195 ;
  assign n6201 = n6200 ^ n6197 ;
  assign n6236 = n6235 ^ n6201 ;
  assign n6257 = n5056 ^ n4189 ;
  assign n6255 = n1023 ^ n602 ;
  assign n6254 = n2962 ^ n848 ;
  assign n6256 = n6255 ^ n6254 ;
  assign n6258 = n6257 ^ n6256 ;
  assign n6251 = n5625 ^ n4311 ;
  assign n6250 = n4941 ^ n231 ;
  assign n6252 = n6251 ^ n6250 ;
  assign n6253 = n6252 ^ n4096 ;
  assign n6259 = n6258 ^ n6253 ;
  assign n6260 = n6259 ^ n1211 ;
  assign n6274 = n3316 ^ n2310 ;
  assign n6271 = n1450 ^ n433 ;
  assign n6270 = n3215 ^ n1093 ;
  assign n6272 = n6271 ^ n6270 ;
  assign n6273 = n6272 ^ n2092 ;
  assign n6275 = n6274 ^ n6273 ;
  assign n6267 = n2507 ^ n1428 ;
  assign n6268 = n6267 ^ n1086 ;
  assign n6264 = n4244 ^ n514 ;
  assign n6263 = n4980 ^ n2334 ;
  assign n6265 = n6264 ^ n6263 ;
  assign n6261 = n3455 ^ n380 ;
  assign n6262 = n6261 ^ n326 ;
  assign n6266 = n6265 ^ n6262 ;
  assign n6269 = n6268 ^ n6266 ;
  assign n6276 = n6275 ^ n6269 ;
  assign n6277 = n6276 ^ n5243 ;
  assign n6278 = ~n6260 & ~n6277 ;
  assign n6247 = ~n2836 & n3726 ;
  assign n6246 = ~n3151 & ~n3733 ;
  assign n6248 = n6247 ^ n6246 ;
  assign n6237 = n3345 ^ n2836 ;
  assign n6243 = n3520 & n6237 ;
  assign n6238 = ~n35 & ~n2924 ;
  assign n6244 = n6243 ^ n6238 ;
  assign n6245 = x31 & n6244 ;
  assign n6249 = n6248 ^ n6245 ;
  assign n6279 = n6278 ^ n6249 ;
  assign n6338 = n4943 ^ n4119 ;
  assign n6334 = n6333 ^ n6225 ;
  assign n6332 = n5134 ^ n4311 ;
  assign n6335 = n6334 ^ n6332 ;
  assign n6336 = n6335 ^ n3296 ;
  assign n6330 = n1809 ^ n1521 ;
  assign n6327 = n3041 ^ n1029 ;
  assign n6328 = n6327 ^ n697 ;
  assign n6325 = n416 ^ n223 ;
  assign n6326 = n6325 ^ n264 ;
  assign n6329 = n6328 ^ n6326 ;
  assign n6331 = n6330 ^ n6329 ;
  assign n6337 = n6336 ^ n6331 ;
  assign n6339 = n6338 ^ n6337 ;
  assign n6320 = n526 ^ n237 ;
  assign n6321 = n6320 ^ n5631 ;
  assign n6319 = n4342 ^ n4242 ;
  assign n6322 = n6321 ^ n6319 ;
  assign n6317 = n881 ^ n200 ;
  assign n6316 = n1667 ^ n642 ;
  assign n6318 = n6317 ^ n6316 ;
  assign n6323 = n6322 ^ n6318 ;
  assign n6310 = n867 ^ n203 ;
  assign n6311 = n6310 ^ n490 ;
  assign n6308 = n521 ^ n284 ;
  assign n6309 = n6308 ^ n414 ;
  assign n6312 = n6311 ^ n6309 ;
  assign n6306 = n2805 ^ n351 ;
  assign n6307 = n6306 ^ n229 ;
  assign n6313 = n6312 ^ n6307 ;
  assign n6314 = n6313 ^ n634 ;
  assign n6303 = n1937 ^ n914 ;
  assign n6302 = n2569 ^ n291 ;
  assign n6304 = n6303 ^ n6302 ;
  assign n6305 = n6304 ^ n2747 ;
  assign n6315 = n6314 ^ n6305 ;
  assign n6324 = n6323 ^ n6315 ;
  assign n6340 = n6339 ^ n6324 ;
  assign n6341 = ~n4986 & ~n6340 ;
  assign n6280 = n3342 ^ n3102 ;
  assign n6281 = n6280 ^ n3343 ;
  assign n6282 = n6281 ^ n3342 ;
  assign n6283 = n6282 ^ n6238 ;
  assign n6284 = n6283 ^ n3520 ;
  assign n6285 = n6284 ^ n6283 ;
  assign n6286 = n6282 ^ n3151 ;
  assign n6288 = n6286 ^ n2924 ;
  assign n6287 = n6286 ^ n2958 ;
  assign n6289 = n6288 ^ n6287 ;
  assign n6292 = x30 & n6289 ;
  assign n6293 = n6292 ^ n6288 ;
  assign n6294 = ~n3520 & ~n6293 ;
  assign n6295 = n6294 ^ n6286 ;
  assign n6296 = n6295 ^ n6238 ;
  assign n6297 = n6296 ^ n6283 ;
  assign n6298 = ~n6285 & ~n6297 ;
  assign n6299 = n6298 ^ n6283 ;
  assign n6300 = ~x31 & ~n6299 ;
  assign n6301 = n6300 ^ n6295 ;
  assign n6342 = n6341 ^ n6301 ;
  assign n6391 = n2111 ^ n206 ;
  assign n6392 = n6391 ^ n1828 ;
  assign n6393 = n6392 ^ n3797 ;
  assign n6388 = n217 ^ n180 ;
  assign n6387 = n1058 ^ n815 ;
  assign n6389 = n6388 ^ n6387 ;
  assign n6385 = n1495 ^ n497 ;
  assign n6384 = n3253 ^ n1116 ;
  assign n6386 = n6385 ^ n6384 ;
  assign n6390 = n6389 ^ n6386 ;
  assign n6394 = n6393 ^ n6390 ;
  assign n6380 = n1076 ^ n568 ;
  assign n6378 = n3086 ^ n264 ;
  assign n6377 = n2805 ^ n1379 ;
  assign n6379 = n6378 ^ n6377 ;
  assign n6381 = n6380 ^ n6379 ;
  assign n6373 = n495 ^ n143 ;
  assign n6375 = n6374 ^ n6373 ;
  assign n6372 = n4008 ^ n2249 ;
  assign n6376 = n6375 ^ n6372 ;
  assign n6382 = n6381 ^ n6376 ;
  assign n6368 = n612 ^ n88 ;
  assign n6366 = n2744 ^ n99 ;
  assign n6367 = n6366 ^ n222 ;
  assign n6369 = n6368 ^ n6367 ;
  assign n6370 = n6369 ^ n3397 ;
  assign n6371 = n6370 ^ n1297 ;
  assign n6383 = n6382 ^ n6371 ;
  assign n6395 = n6394 ^ n6383 ;
  assign n6396 = n2688 & ~n6395 ;
  assign n6360 = x30 & ~n2958 ;
  assign n6361 = n6360 ^ n2924 ;
  assign n6362 = ~n3520 & ~n6361 ;
  assign n6343 = n3342 ^ n3101 ;
  assign n6344 = n6343 ^ n2924 ;
  assign n6346 = n6344 ^ n2958 ;
  assign n6345 = n6344 ^ n3099 ;
  assign n6347 = n6346 ^ n6345 ;
  assign n6350 = x30 & n6347 ;
  assign n6351 = n6350 ^ n6346 ;
  assign n6352 = ~n3520 & ~n6351 ;
  assign n6353 = n6352 ^ n6344 ;
  assign n6354 = n6353 ^ n2924 ;
  assign n6363 = n6362 ^ n6354 ;
  assign n6364 = ~x31 & ~n6363 ;
  assign n6365 = n6364 ^ n6353 ;
  assign n6397 = n6396 ^ n6365 ;
  assign n6453 = x30 & ~n3099 ;
  assign n6454 = n6453 ^ n2958 ;
  assign n6455 = ~n3520 & ~n6454 ;
  assign n6456 = n6455 ^ n2958 ;
  assign n6439 = n3341 ^ n3100 ;
  assign n6440 = n6439 ^ n2958 ;
  assign n6457 = n6456 ^ n6440 ;
  assign n6442 = n6440 ^ n3027 ;
  assign n6441 = n6440 ^ n3099 ;
  assign n6443 = n6442 ^ n6441 ;
  assign n6446 = ~x30 & n6443 ;
  assign n6447 = n6446 ^ n6442 ;
  assign n6448 = ~n3520 & ~n6447 ;
  assign n6458 = n6457 ^ n6448 ;
  assign n6459 = x31 & ~n6458 ;
  assign n6460 = n6459 ^ n6456 ;
  assign n6414 = n255 ^ n218 ;
  assign n6415 = n6414 ^ n193 ;
  assign n6416 = n6415 ^ n2060 ;
  assign n6412 = n2234 ^ n1015 ;
  assign n6413 = n6412 ^ n1305 ;
  assign n6417 = n6416 ^ n6413 ;
  assign n6408 = n3601 ^ n3129 ;
  assign n6409 = n6408 ^ n850 ;
  assign n6405 = n1280 ^ n155 ;
  assign n6406 = n6405 ^ n2726 ;
  assign n6403 = n732 ^ n130 ;
  assign n6402 = n3213 ^ n1206 ;
  assign n6404 = n6403 ^ n6402 ;
  assign n6407 = n6406 ^ n6404 ;
  assign n6410 = n6409 ^ n6407 ;
  assign n6398 = n761 ^ n407 ;
  assign n6399 = n6398 ^ n660 ;
  assign n6400 = n6399 ^ n2864 ;
  assign n6401 = n6400 ^ n6373 ;
  assign n6411 = n6410 ^ n6401 ;
  assign n6418 = n6417 ^ n6411 ;
  assign n6433 = n1181 ^ n782 ;
  assign n6431 = n3192 ^ n116 ;
  assign n6432 = n6431 ^ n636 ;
  assign n6434 = n6433 ^ n6432 ;
  assign n6428 = n3889 ^ n2195 ;
  assign n6427 = n1721 ^ n872 ;
  assign n6429 = n6428 ^ n6427 ;
  assign n6430 = n6429 ^ n2265 ;
  assign n6435 = n6434 ^ n6430 ;
  assign n6423 = n6422 ^ n416 ;
  assign n6424 = n6423 ^ n790 ;
  assign n6420 = n6419 ^ n450 ;
  assign n6421 = n6420 ^ n584 ;
  assign n6425 = n6424 ^ n6421 ;
  assign n6426 = n6425 ^ n3074 ;
  assign n6436 = n6435 ^ n6426 ;
  assign n6437 = n6436 ^ n2028 ;
  assign n6438 = ~n6418 & ~n6437 ;
  assign n6461 = n6460 ^ n6438 ;
  assign n6472 = ~n3337 & n24214 ;
  assign n6470 = n3027 & ~n3733 ;
  assign n6466 = ~n3339 & ~n3720 ;
  assign n6467 = n6466 ^ n3099 ;
  assign n6468 = n3520 & ~n6467 ;
  assign n6469 = n6468 ^ n3720 ;
  assign n6471 = n6470 ^ n6469 ;
  assign n6473 = n6472 ^ n6471 ;
  assign n6474 = n4014 ^ n1516 ;
  assign n6491 = n672 ^ n269 ;
  assign n6492 = n6491 ^ n1208 ;
  assign n6493 = n6492 ^ n2488 ;
  assign n6488 = n2234 ^ n405 ;
  assign n6489 = n6488 ^ n704 ;
  assign n6486 = n2200 ^ n409 ;
  assign n6487 = n6486 ^ n1181 ;
  assign n6490 = n6489 ^ n6487 ;
  assign n6494 = n6493 ^ n6490 ;
  assign n6483 = n3415 ^ n426 ;
  assign n6484 = n6483 ^ n550 ;
  assign n6480 = n1311 ^ n728 ;
  assign n6478 = n857 ^ n212 ;
  assign n6479 = n6478 ^ n613 ;
  assign n6481 = n6480 ^ n6479 ;
  assign n6476 = n2348 ^ n1414 ;
  assign n6475 = n6320 ^ n837 ;
  assign n6477 = n6476 ^ n6475 ;
  assign n6482 = n6481 ^ n6477 ;
  assign n6485 = n6484 ^ n6482 ;
  assign n6495 = n6494 ^ n6485 ;
  assign n6496 = n6495 ^ n3224 ;
  assign n6497 = n6496 ^ n4106 ;
  assign n6498 = ~n6474 & ~n6497 ;
  assign n6500 = n6473 & n6498 ;
  assign n6499 = n6498 ^ n6473 ;
  assign n6501 = n6500 ^ n6499 ;
  assign n6502 = n6501 ^ n6460 ;
  assign n6503 = n6461 & n6502 ;
  assign n6504 = n6503 ^ n6460 ;
  assign n6505 = n6504 ^ n6365 ;
  assign n6506 = ~n6397 & ~n6505 ;
  assign n6507 = n6506 ^ n6365 ;
  assign n6508 = n6507 ^ n6301 ;
  assign n6509 = n6342 & n6508 ;
  assign n6510 = n6509 ^ n6507 ;
  assign n6511 = n6510 ^ n6249 ;
  assign n6512 = ~n6279 & n6511 ;
  assign n6513 = n6512 ^ n6249 ;
  assign n6514 = n6513 ^ n6201 ;
  assign n6515 = ~n6236 & n6514 ;
  assign n6516 = n6515 ^ n6201 ;
  assign n6517 = n6516 ^ n6193 ;
  assign n6518 = n6194 & n6517 ;
  assign n6520 = n6519 ^ n6518 ;
  assign n6521 = n6184 & n6520 ;
  assign n6522 = n6521 ^ n6183 ;
  assign n6523 = n6522 ^ n6159 ;
  assign n6524 = ~n6174 & n6523 ;
  assign n6525 = n6524 ^ n6159 ;
  assign n6526 = n6525 ^ n6154 ;
  assign n6527 = ~n6156 & ~n6526 ;
  assign n6528 = n6527 ^ n6154 ;
  assign n6529 = n6528 ^ n6144 ;
  assign n6530 = n6146 & n6529 ;
  assign n6531 = n6530 ^ n6528 ;
  assign n6532 = n6531 ^ n6127 ;
  assign n6533 = ~n6133 & ~n6532 ;
  assign n6534 = n6533 ^ n6127 ;
  assign n6535 = n6534 ^ n6118 ;
  assign n6536 = ~n6123 & n6535 ;
  assign n6537 = n6536 ^ n6118 ;
  assign n6109 = ~n1540 & n14027 ;
  assign n6105 = n5855 ^ n5818 ;
  assign n6106 = n6105 ^ x20 ;
  assign n6104 = ~n1214 & n4916 ;
  assign n6107 = n6106 ^ n6104 ;
  assign n6103 = ~n968 & n4683 ;
  assign n6108 = n6107 ^ n6103 ;
  assign n6110 = n6109 ^ n6108 ;
  assign n6102 = n3521 & n4684 ;
  assign n6111 = n6110 ^ n6102 ;
  assign n6561 = n6537 ^ n6111 ;
  assign n6562 = n6561 ^ x17 ;
  assign n6560 = ~n1109 & n20731 ;
  assign n6563 = n6562 ^ n6560 ;
  assign n6559 = ~n3473 & n5702 ;
  assign n6564 = n6563 ^ n6559 ;
  assign n6566 = n6565 ^ n6564 ;
  assign n6558 = ~n3508 & n5703 ;
  assign n6567 = n6566 ^ n6558 ;
  assign n6575 = ~n1540 & n4916 ;
  assign n6573 = ~n1433 & n14027 ;
  assign n6571 = ~n1214 & n4683 ;
  assign n6569 = n6534 ^ n6123 ;
  assign n6570 = n6569 ^ x20 ;
  assign n6572 = n6571 ^ n6570 ;
  assign n6574 = n6573 ^ n6572 ;
  assign n6576 = n6575 ^ n6574 ;
  assign n6568 = ~n4603 & n4684 ;
  assign n6577 = n6576 ^ n6568 ;
  assign n6585 = ~n1540 & n4683 ;
  assign n6581 = n6531 ^ n6133 ;
  assign n6582 = n6581 ^ x20 ;
  assign n6580 = ~n1351 & n14027 ;
  assign n6583 = n6582 ^ n6580 ;
  assign n6579 = ~n1433 & n4916 ;
  assign n6584 = n6583 ^ n6579 ;
  assign n6586 = n6585 ^ n6584 ;
  assign n6578 = ~n4610 & n4684 ;
  assign n6587 = n6586 ^ n6578 ;
  assign n6594 = ~n1631 & n4491 ;
  assign n6593 = ~n1871 & ~n4496 ;
  assign n6595 = n6594 ^ n6593 ;
  assign n6590 = ~n1795 & n4504 ;
  assign n6589 = ~n4392 & n4492 ;
  assign n6591 = n6590 ^ n6589 ;
  assign n6592 = n6591 ^ x23 ;
  assign n6596 = n6595 ^ n6592 ;
  assign n6588 = n6528 ^ n6146 ;
  assign n6597 = n6596 ^ n6588 ;
  assign n6602 = ~n2268 & n12861 ;
  assign n6601 = ~n487 & ~n2096 ;
  assign n6603 = n6602 ^ n6601 ;
  assign n6604 = n6603 ^ x26 ;
  assign n6600 = n446 & ~n2185 ;
  assign n6605 = n6604 ^ n6600 ;
  assign n6599 = ~n3501 & n5196 ;
  assign n6606 = n6605 ^ n6599 ;
  assign n6631 = n6606 ^ n6588 ;
  assign n6598 = n6525 ^ n6156 ;
  assign n6607 = n6606 ^ n6598 ;
  assign n6623 = n3481 & n5520 ;
  assign n6621 = n831 & ~n2554 ;
  assign n6619 = n656 & ~n2449 ;
  assign n6611 = n446 & ~n2268 ;
  assign n6610 = ~n487 & ~n2185 ;
  assign n6612 = n6611 ^ n6610 ;
  assign n6613 = n6612 ^ x26 ;
  assign n6609 = ~n2364 & n12861 ;
  assign n6614 = n6613 ^ n6609 ;
  assign n6608 = ~n3501 & n5832 ;
  assign n6615 = n6614 ^ n6608 ;
  assign n6618 = n6615 ^ x29 ;
  assign n6620 = n6619 ^ n6618 ;
  assign n6622 = n6621 ^ n6620 ;
  assign n6624 = n6623 ^ n6622 ;
  assign n6617 = ~n2486 & n3484 ;
  assign n6625 = n6624 ^ n6617 ;
  assign n6626 = n6522 ^ n6174 ;
  assign n6627 = n6626 ^ n6615 ;
  assign n6628 = n6625 & n6627 ;
  assign n6616 = n6615 ^ n6598 ;
  assign n6629 = n6628 ^ n6616 ;
  assign n6630 = n6607 & ~n6629 ;
  assign n6632 = n6631 ^ n6630 ;
  assign n6633 = ~n6597 & n6632 ;
  assign n6634 = n6633 ^ n6596 ;
  assign n6635 = n6634 ^ n6581 ;
  assign n6636 = ~n6587 & ~n6635 ;
  assign n6637 = n6636 ^ n6581 ;
  assign n6638 = n6637 ^ n6569 ;
  assign n6639 = n6577 & ~n6638 ;
  assign n6640 = n6639 ^ n6569 ;
  assign n6641 = n6640 ^ n6561 ;
  assign n6642 = ~n6567 & ~n6641 ;
  assign n6643 = n6642 ^ n6561 ;
  assign n6057 = ~x13 & n4897 ;
  assign n6078 = ~x14 & n6057 ;
  assign n6079 = ~n485 & n6078 ;
  assign n6074 = n6057 ^ n4907 ;
  assign n6075 = ~n445 & ~n6074 ;
  assign n6066 = x13 ^ x12 ;
  assign n15382 = ~n4897 & ~n6066 ;
  assign n15385 = n15382 ^ x14 ;
  assign n6055 = x13 & ~n4898 ;
  assign n6059 = n15382 ^ n6055 ;
  assign n6061 = n4897 ^ x14 ;
  assign n6060 = x14 & n4897 ;
  assign n6062 = n6061 ^ n6060 ;
  assign n6065 = ~x12 & ~x13 ;
  assign n6067 = n6066 ^ n6065 ;
  assign n6068 = ~n6062 & n6067 ;
  assign n6063 = n6062 ^ x14 ;
  assign n6064 = n6063 ^ n6055 ;
  assign n6069 = n6068 ^ n6064 ;
  assign n6070 = ~n6059 & n6069 ;
  assign n6072 = n15385 ^ n6070 ;
  assign n6073 = ~n317 & ~n6072 ;
  assign n6076 = n6075 ^ n6073 ;
  assign n6077 = n6076 ^ x14 ;
  assign n6080 = n6079 ^ n6077 ;
  assign n6081 = n6080 ^ x14 ;
  assign n6087 = ~x13 & ~n3499 ;
  assign n6088 = n6087 ^ n485 ;
  assign n6089 = n4897 & ~n6088 ;
  assign n6091 = n6089 ^ n6079 ;
  assign n6092 = n6091 ^ n3500 ;
  assign n6093 = n6092 ^ n6091 ;
  assign n8434 = n6057 ^ n4897 ;
  assign n6098 = n6093 & n8434 ;
  assign n6099 = n6098 ^ n6091 ;
  assign n6100 = ~n6080 & ~n6099 ;
  assign n6101 = n6081 & ~n6100 ;
  assign n6548 = ~n3473 & n5700 ;
  assign n6544 = n5858 ^ n5803 ;
  assign n6545 = n6544 ^ x17 ;
  assign n6543 = ~n649 & n5702 ;
  assign n6546 = n6545 ^ n6543 ;
  assign n6542 = ~n824 & n20731 ;
  assign n6547 = n6546 ^ n6542 ;
  assign n6549 = n6548 ^ n6547 ;
  assign n6541 = ~n3476 & n5703 ;
  assign n6550 = n6549 ^ n6541 ;
  assign n6538 = n6537 ^ n6105 ;
  assign n6539 = n6111 & ~n6538 ;
  assign n6540 = n6539 ^ n6105 ;
  assign n6551 = n6550 ^ n6540 ;
  assign n6552 = n6551 ^ n6091 ;
  assign n6553 = n6552 ^ n6100 ;
  assign n6554 = n6553 ^ x14 ;
  assign n6555 = n6554 ^ n6551 ;
  assign n6556 = n6101 & n6555 ;
  assign n6557 = n6556 ^ n6553 ;
  assign n6644 = n6643 ^ n6557 ;
  assign n6668 = n6667 ^ n6644 ;
  assign n6675 = ~n445 & n6078 ;
  assign n6672 = ~n317 & ~n6074 ;
  assign n6671 = ~n649 & ~n6072 ;
  assign n6673 = n6672 ^ n6671 ;
  assign n6674 = n6673 ^ x14 ;
  assign n6676 = n6675 ^ n6674 ;
  assign n6679 = ~x13 & ~n4072 ;
  assign n6680 = n6679 ^ n445 ;
  assign n6681 = n4897 & ~n6680 ;
  assign n6683 = n6681 ^ n6675 ;
  assign n6686 = n6683 ^ n4073 ;
  assign n6687 = n6686 ^ n6683 ;
  assign n6688 = n6687 & n8434 ;
  assign n6689 = n6688 ^ n6683 ;
  assign n6690 = ~n6676 & ~n6689 ;
  assign n6691 = n6690 ^ n6683 ;
  assign n6692 = n6691 ^ x14 ;
  assign n6693 = n6691 ^ n6676 ;
  assign n6694 = ~n6690 & ~n6693 ;
  assign n6695 = n6692 & n6694 ;
  assign n6696 = n6695 ^ n6691 ;
  assign n6669 = n6640 ^ n6567 ;
  assign n6697 = n6696 ^ n6669 ;
  assign n6782 = ~n968 & n20731 ;
  assign n6781 = ~n824 & n5702 ;
  assign n6783 = n6782 ^ n6781 ;
  assign n6784 = n6783 ^ x17 ;
  assign n6780 = ~n1109 & n5700 ;
  assign n6785 = n6784 ^ n6780 ;
  assign n6779 = ~n4050 & n5703 ;
  assign n6786 = n6785 ^ n6779 ;
  assign n6705 = ~n968 & n5700 ;
  assign n6701 = n6634 ^ n6587 ;
  assign n6702 = n6701 ^ x17 ;
  assign n6700 = ~n1214 & n20731 ;
  assign n6703 = n6702 ^ n6700 ;
  assign n6699 = ~n1109 & n5702 ;
  assign n6704 = n6703 ^ n6699 ;
  assign n6706 = n6705 ^ n6704 ;
  assign n6698 = n3905 & n5703 ;
  assign n6707 = n6706 ^ n6698 ;
  assign n6716 = n6632 ^ n6596 ;
  assign n6711 = ~n1433 & n4683 ;
  assign n6710 = ~n1703 & n14027 ;
  assign n6712 = n6711 ^ n6710 ;
  assign n6713 = n6712 ^ x20 ;
  assign n6709 = ~n1351 & n4916 ;
  assign n6714 = n6713 ^ n6709 ;
  assign n6708 = n4152 & n4684 ;
  assign n6715 = n6714 ^ n6708 ;
  assign n6717 = n6716 ^ n6715 ;
  assign n6748 = n6626 ^ n6625 ;
  assign n6735 = n6520 ^ n6183 ;
  assign n6730 = ~n487 & ~n2268 ;
  assign n6729 = n446 & ~n2364 ;
  assign n6731 = n6730 ^ n6729 ;
  assign n6732 = n6731 ^ x26 ;
  assign n6728 = ~n2449 & n12861 ;
  assign n6733 = n6732 ^ n6728 ;
  assign n6727 = ~n3501 & n5144 ;
  assign n6734 = n6733 ^ n6727 ;
  assign n6736 = n6735 ^ n6734 ;
  assign n5381 = n5380 ^ n2486 ;
  assign n6743 = n3481 & n5381 ;
  assign n6741 = n656 & ~n2486 ;
  assign n6739 = n831 & ~n2609 ;
  assign n6738 = n6734 ^ x29 ;
  assign n6740 = n6739 ^ n6738 ;
  assign n6742 = n6741 ^ n6740 ;
  assign n6744 = n6743 ^ n6742 ;
  assign n6737 = ~n2554 & n3484 ;
  assign n6745 = n6744 ^ n6737 ;
  assign n6746 = n6736 & ~n6745 ;
  assign n6747 = n6746 ^ n6735 ;
  assign n6749 = n6748 ^ n6747 ;
  assign n6760 = ~n1994 & ~n4496 ;
  assign n6758 = n6747 ^ x23 ;
  assign n6755 = ~n4384 & n4700 ;
  assign n6756 = n6755 ^ n1795 ;
  assign n6757 = n4488 & ~n6756 ;
  assign n6759 = n6758 ^ n6757 ;
  assign n6761 = n6760 ^ n6759 ;
  assign n6750 = ~n2096 & n4504 ;
  assign n6762 = n6761 ^ n6750 ;
  assign n6763 = n6749 & ~n6762 ;
  assign n6764 = n6763 ^ n6748 ;
  assign n6772 = n6764 ^ n6716 ;
  assign n6765 = n6764 ^ x23 ;
  assign n6724 = n4700 & n5184 ;
  assign n6725 = n6724 ^ n1871 ;
  assign n6726 = n4488 & ~n6725 ;
  assign n6766 = n6765 ^ n6726 ;
  assign n6719 = ~n1795 & ~n4496 ;
  assign n6767 = n6766 ^ n6719 ;
  assign n6718 = ~n1994 & n4504 ;
  assign n6768 = n6767 ^ n6718 ;
  assign n6769 = n6629 ^ n6606 ;
  assign n6770 = n6769 ^ n6764 ;
  assign n6771 = n6768 & n6770 ;
  assign n6773 = n6772 ^ n6771 ;
  assign n6774 = ~n6717 & ~n6773 ;
  assign n6775 = n6774 ^ n6716 ;
  assign n6776 = n6775 ^ n6701 ;
  assign n6777 = ~n6707 & n6776 ;
  assign n6778 = n6777 ^ n6701 ;
  assign n6787 = n6786 ^ n6778 ;
  assign n6788 = n6637 ^ n6577 ;
  assign n6789 = n6788 ^ n6696 ;
  assign n6790 = n6789 ^ n6778 ;
  assign n6791 = n6790 ^ n6696 ;
  assign n6792 = n6787 & n6791 ;
  assign n6793 = n6792 ^ n6789 ;
  assign n6794 = n6697 & ~n6793 ;
  assign n6670 = n6669 ^ n6667 ;
  assign n6795 = n6794 ^ n6670 ;
  assign n6796 = ~n6668 & ~n6795 ;
  assign n6797 = n6796 ^ n6667 ;
  assign n6798 = n6643 ^ n6551 ;
  assign n6799 = n6557 & n6798 ;
  assign n6800 = n6799 ^ n6551 ;
  assign n6801 = n6800 ^ n6797 ;
  assign n6812 = n6544 ^ n6540 ;
  assign n6813 = ~n6550 & ~n6812 ;
  assign n6814 = n6813 ^ n6544 ;
  assign n6809 = ~n649 & n5700 ;
  assign n6805 = n5860 ^ n5795 ;
  assign n6806 = n6805 ^ x17 ;
  assign n6804 = ~n3473 & n20731 ;
  assign n6807 = n6806 ^ n6804 ;
  assign n6803 = ~n317 & n5702 ;
  assign n6808 = n6807 ^ n6803 ;
  assign n6810 = n6809 ^ n6808 ;
  assign n6802 = n3956 & n5703 ;
  assign n6811 = n6810 ^ n6802 ;
  assign n6815 = n6814 ^ n6811 ;
  assign n6816 = n6815 ^ n6800 ;
  assign n6817 = n6801 & ~n6816 ;
  assign n6818 = ~n6797 & n6817 ;
  assign n6824 = n3944 ^ x13 ;
  assign n6825 = n6824 ^ n3944 ;
  assign n6826 = ~n3924 & n6825 ;
  assign n6827 = n6826 ^ n3944 ;
  assign n6828 = n6060 & n6827 ;
  assign n6820 = ~n485 & ~n6074 ;
  assign n6819 = ~n445 & ~n6072 ;
  assign n6821 = n6820 ^ n6819 ;
  assign n6822 = n6821 ^ x14 ;
  assign n6829 = n6828 ^ n6822 ;
  assign n6832 = x13 & ~n3924 ;
  assign n6833 = n6832 ^ n3943 ;
  assign n6834 = n4897 & ~n6833 ;
  assign n6835 = n6834 ^ n6821 ;
  assign n6836 = ~x14 & n6835 ;
  assign n6837 = ~n6829 & n6836 ;
  assign n6838 = n6837 ^ n6829 ;
  assign n7110 = n6795 ^ n6644 ;
  assign n6844 = ~n485 & n6655 ;
  assign n6842 = ~n3943 & n6650 ;
  assign n6840 = n6793 ^ n6669 ;
  assign n6841 = n6840 ^ x11 ;
  assign n6843 = n6842 ^ n6841 ;
  assign n6845 = n6844 ^ n6843 ;
  assign n6839 = n4515 & n15413 ;
  assign n6846 = n6845 ^ n6839 ;
  assign n7073 = n6788 ^ n6778 ;
  assign n7074 = n7073 ^ n6786 ;
  assign n6850 = ~n824 & ~n6072 ;
  assign n6849 = ~n3473 & ~n6074 ;
  assign n6851 = n6850 ^ n6849 ;
  assign n6860 = n6851 ^ x14 ;
  assign n6859 = n6775 ^ n6707 ;
  assign n6861 = n6860 ^ n6859 ;
  assign n6852 = n6851 ^ n649 ;
  assign n4899 = x14 ^ x13 ;
  assign n6847 = n4899 ^ n649 ;
  assign n6853 = n6852 ^ n6847 ;
  assign n6856 = ~n3475 & n6853 ;
  assign n6857 = n6856 ^ n6847 ;
  assign n6858 = n4897 & ~n6857 ;
  assign n6862 = n6861 ^ n6858 ;
  assign n7057 = n6773 ^ n6715 ;
  assign n6870 = ~n1351 & n4683 ;
  assign n6866 = n6769 ^ n6768 ;
  assign n6867 = n6866 ^ x20 ;
  assign n6865 = ~n1703 & n4916 ;
  assign n6868 = n6867 ^ n6865 ;
  assign n6864 = ~n1631 & n14027 ;
  assign n6869 = n6868 ^ n6864 ;
  assign n6871 = n6870 ^ n6869 ;
  assign n6863 = n4417 & n4684 ;
  assign n6872 = n6871 ^ n6863 ;
  assign n6880 = ~n1871 & n14027 ;
  assign n6876 = n6762 ^ n6748 ;
  assign n6877 = n6876 ^ x20 ;
  assign n6875 = ~n1703 & n4683 ;
  assign n6878 = n6877 ^ n6875 ;
  assign n6874 = ~n1631 & n4916 ;
  assign n6879 = n6878 ^ n6874 ;
  assign n6881 = n6880 ^ n6879 ;
  assign n6873 = ~n4615 & n4684 ;
  assign n6882 = n6881 ^ n6873 ;
  assign n6890 = ~n1994 & n4491 ;
  assign n6886 = n6745 ^ n6735 ;
  assign n6887 = n6886 ^ x23 ;
  assign n6885 = n4492 & n5409 ;
  assign n6888 = n6887 ^ n6885 ;
  assign n6884 = ~n2096 & ~n4496 ;
  assign n6889 = n6888 ^ n6884 ;
  assign n6891 = n6890 ^ n6889 ;
  assign n6883 = ~n2185 & n4504 ;
  assign n6892 = n6891 ^ n6883 ;
  assign n7035 = n6516 ^ n6194 ;
  assign n7021 = n6513 ^ n6236 ;
  assign n6900 = n6176 ^ n3227 ;
  assign n6901 = n3481 & n6900 ;
  assign n6896 = n6510 ^ n6279 ;
  assign n6897 = n6896 ^ x29 ;
  assign n6895 = n656 & ~n3227 ;
  assign n6898 = n6897 ^ n6895 ;
  assign n6894 = n831 & ~n2738 ;
  assign n6899 = n6898 ^ n6894 ;
  assign n6902 = n6901 ^ n6899 ;
  assign n6893 = ~n2646 & n3484 ;
  assign n6903 = n6902 ^ n6893 ;
  assign n7005 = n6507 ^ n6342 ;
  assign n6912 = n656 & ~n2738 ;
  assign n6910 = ~n2836 & n3484 ;
  assign n6907 = n3347 ^ n2738 ;
  assign n6908 = n3481 & ~n6907 ;
  assign n6905 = n6504 ^ n6397 ;
  assign n6906 = n6905 ^ x29 ;
  assign n6909 = n6908 ^ n6906 ;
  assign n6911 = n6910 ^ n6909 ;
  assign n6913 = n6912 ^ n6911 ;
  assign n6904 = n831 & ~n3151 ;
  assign n6914 = n6913 ^ n6904 ;
  assign n6922 = ~n3151 & n3484 ;
  assign n6920 = n3481 & n6237 ;
  assign n6917 = n656 & ~n2836 ;
  assign n6916 = n831 & ~n2924 ;
  assign n6918 = n6917 ^ n6916 ;
  assign n6919 = n6918 ^ x29 ;
  assign n6921 = n6920 ^ n6919 ;
  assign n6923 = n6922 ^ n6921 ;
  assign n6915 = n6501 ^ n6461 ;
  assign n6924 = n6923 ^ n6915 ;
  assign n6934 = ~n2924 & n3484 ;
  assign n6930 = n4536 & ~n6282 ;
  assign n6931 = n6930 ^ n3151 ;
  assign n6932 = n650 & ~n6931 ;
  assign n6933 = n6932 ^ x29 ;
  assign n6935 = n6934 ^ n6933 ;
  assign n6925 = n831 & ~n2958 ;
  assign n6936 = n6935 ^ n6925 ;
  assign n6988 = n6936 ^ n6500 ;
  assign n6978 = ~n2958 & n3484 ;
  assign n6976 = n3481 & n6344 ;
  assign n6973 = n831 & ~n3099 ;
  assign n6972 = n656 & ~n2924 ;
  assign n6974 = n6973 ^ n6972 ;
  assign n6975 = n6974 ^ x29 ;
  assign n6977 = n6976 ^ n6975 ;
  assign n6979 = n6978 ^ n6977 ;
  assign n6941 = n650 & ~n2958 ;
  assign n6940 = n3481 & ~n6439 ;
  assign n6942 = n6941 ^ n6940 ;
  assign n6938 = n831 & ~n3027 ;
  assign n6937 = ~n3099 & n3484 ;
  assign n6939 = n6938 ^ n6937 ;
  assign n6943 = n6942 ^ n6939 ;
  assign n6947 = ~x30 & ~n3337 ;
  assign n6956 = ~n3027 & n3484 ;
  assign n6955 = n831 & ~n3337 ;
  assign n6957 = n6956 ^ n6955 ;
  assign n6952 = n3339 & n4536 ;
  assign n6953 = n6952 ^ n3099 ;
  assign n6954 = n650 & ~n6953 ;
  assign n6958 = n6957 ^ n6954 ;
  assign n6959 = n650 & ~n3027 ;
  assign n6960 = n827 & ~n3337 ;
  assign n6961 = ~n6959 & n6960 ;
  assign n6962 = n6961 ^ n6959 ;
  assign n6963 = ~n6958 & ~n6962 ;
  assign n6966 = ~n6947 & ~n6963 ;
  assign n6967 = x29 & n6966 ;
  assign n6968 = n6967 ^ x29 ;
  assign n6944 = ~n34 & ~n3337 ;
  assign n6969 = n6968 ^ n6944 ;
  assign n6970 = ~n6943 & n6969 ;
  assign n6971 = n6970 ^ n6944 ;
  assign n6980 = n6979 ^ n6971 ;
  assign n6982 = ~n3337 & ~n3720 ;
  assign n6981 = ~n3027 & n3520 ;
  assign n6983 = n6982 ^ n6981 ;
  assign n6984 = n6983 ^ n6979 ;
  assign n6985 = n6980 & n6984 ;
  assign n6986 = n6985 ^ n6979 ;
  assign n6989 = n6986 ^ n6936 ;
  assign n6990 = ~n6988 & ~n6989 ;
  assign n6991 = n6990 ^ n6500 ;
  assign n6993 = n6991 ^ n6923 ;
  assign n6987 = n6936 & n6986 ;
  assign n6992 = n6991 ^ n6987 ;
  assign n6994 = n6993 ^ n6992 ;
  assign n6995 = n6994 ^ n6993 ;
  assign n6996 = n6993 ^ n6501 ;
  assign n6997 = n6996 ^ n6993 ;
  assign n6998 = ~n6995 & ~n6997 ;
  assign n6999 = n6998 ^ n6993 ;
  assign n7000 = ~n6924 & ~n6999 ;
  assign n7001 = n7000 ^ n6923 ;
  assign n7002 = n7001 ^ n6905 ;
  assign n7003 = n6914 & n7002 ;
  assign n7004 = n7003 ^ n6905 ;
  assign n7006 = n7005 ^ n7004 ;
  assign n7013 = n3481 & ~n5651 ;
  assign n7011 = n831 & ~n2836 ;
  assign n7009 = n656 & ~n2646 ;
  assign n7008 = n7005 ^ x29 ;
  assign n7010 = n7009 ^ n7008 ;
  assign n7012 = n7011 ^ n7010 ;
  assign n7014 = n7013 ^ n7012 ;
  assign n7007 = ~n2738 & n3484 ;
  assign n7015 = n7014 ^ n7007 ;
  assign n7016 = ~n7006 & ~n7015 ;
  assign n7017 = n7016 ^ n7005 ;
  assign n7018 = n7017 ^ n6896 ;
  assign n7019 = ~n6903 & n7018 ;
  assign n7020 = n7019 ^ n6896 ;
  assign n7022 = n7021 ^ n7020 ;
  assign n7029 = n6171 ^ n2609 ;
  assign n7030 = n3481 & n7029 ;
  assign n7027 = n656 & ~n2609 ;
  assign n7025 = n831 & ~n2646 ;
  assign n7024 = n7021 ^ x29 ;
  assign n7026 = n7025 ^ n7024 ;
  assign n7028 = n7027 ^ n7026 ;
  assign n7031 = n7030 ^ n7028 ;
  assign n7023 = ~n3227 & n3484 ;
  assign n7032 = n7031 ^ n7023 ;
  assign n7033 = n7022 & ~n7032 ;
  assign n7034 = n7033 ^ n7021 ;
  assign n7036 = n7035 ^ n7034 ;
  assign n7043 = ~n487 & ~n2364 ;
  assign n7041 = ~n2486 & n12861 ;
  assign n7039 = n446 & ~n2449 ;
  assign n7038 = n7035 ^ x26 ;
  assign n7040 = n7039 ^ n7038 ;
  assign n7042 = n7041 ^ n7040 ;
  assign n7044 = n7043 ^ n7042 ;
  assign n7037 = ~n3501 & n5283 ;
  assign n7045 = n7044 ^ n7037 ;
  assign n7046 = ~n7036 & n7045 ;
  assign n7047 = n7046 ^ n7035 ;
  assign n7048 = n7047 ^ n6886 ;
  assign n7049 = n6892 & n7048 ;
  assign n7050 = n7049 ^ n6886 ;
  assign n7051 = n7050 ^ n6876 ;
  assign n7052 = n6882 & n7051 ;
  assign n7053 = n7052 ^ n6876 ;
  assign n7054 = n7053 ^ n6866 ;
  assign n7055 = n6872 & n7054 ;
  assign n7056 = n7055 ^ n6866 ;
  assign n7058 = n7057 ^ n7056 ;
  assign n7065 = ~n1214 & n5700 ;
  assign n7063 = ~n968 & n5702 ;
  assign n7061 = ~n1540 & n20731 ;
  assign n7060 = n7057 ^ x17 ;
  assign n7062 = n7061 ^ n7060 ;
  assign n7064 = n7063 ^ n7062 ;
  assign n7066 = n7065 ^ n7064 ;
  assign n7059 = n3521 & n5703 ;
  assign n7067 = n7066 ^ n7059 ;
  assign n7068 = ~n7058 & ~n7067 ;
  assign n7069 = n7068 ^ n7057 ;
  assign n7070 = n7069 ^ n6859 ;
  assign n7071 = n6862 & ~n7070 ;
  assign n7072 = n7071 ^ n6859 ;
  assign n7075 = n7074 ^ n7072 ;
  assign n7086 = ~n317 & n6078 ;
  assign n7078 = n3956 ^ n317 ;
  assign n7079 = ~x13 & ~n7078 ;
  assign n7080 = n7079 ^ n317 ;
  assign n7081 = n4897 & ~n7080 ;
  assign n7090 = n7086 ^ n7081 ;
  assign n7102 = n7090 ^ n7074 ;
  assign n7083 = ~n3473 & ~n6072 ;
  assign n7082 = ~n649 & ~n6074 ;
  assign n7084 = n7083 ^ n7082 ;
  assign n7085 = n7084 ^ x14 ;
  assign n7087 = n7086 ^ n7085 ;
  assign n7097 = n3956 & n8434 ;
  assign n7098 = n7097 ^ n7090 ;
  assign n7099 = ~n7087 & ~n7098 ;
  assign n7103 = n7102 ^ n7099 ;
  assign n7091 = n7090 ^ x14 ;
  assign n7092 = n7090 ^ n7087 ;
  assign n7100 = ~n7092 & ~n7099 ;
  assign n7101 = n7091 & n7100 ;
  assign n7104 = n7103 ^ n7101 ;
  assign n7105 = n7075 & ~n7104 ;
  assign n7106 = n7105 ^ n7074 ;
  assign n7107 = n7106 ^ n6840 ;
  assign n7108 = ~n6846 & ~n7107 ;
  assign n7109 = n7108 ^ n6840 ;
  assign n7111 = n7110 ^ n7109 ;
  assign n7113 = n7104 ^ n7072 ;
  assign n7122 = ~n445 & n6655 ;
  assign n9154 = x11 ^ x10 ;
  assign n7118 = ~n3924 & n9154 ;
  assign n7119 = n7118 ^ n3943 ;
  assign n7120 = n6648 & ~n7119 ;
  assign n7121 = n7120 ^ x11 ;
  assign n7123 = n7122 ^ n7121 ;
  assign n7114 = ~n485 & n6650 ;
  assign n7124 = n7123 ^ n7114 ;
  assign n7125 = ~n7113 & n7124 ;
  assign n7112 = n7106 ^ n6846 ;
  assign n7126 = n7125 ^ n7112 ;
  assign n7128 = x6 ^ x5 ;
  assign n7132 = x7 & n7128 ;
  assign n7129 = x8 & n7128 ;
  assign n7130 = n7129 ^ n7128 ;
  assign n7131 = n7130 ^ x7 ;
  assign n7133 = n7132 ^ n7131 ;
  assign n7134 = n7133 ^ n7129 ;
  assign n7135 = n7134 ^ n7131 ;
  assign n8044 = ~n3920 & n7135 ;
  assign n7137 = x5 & x6 ;
  assign n7138 = x7 & n7137 ;
  assign n7145 = n7138 ^ x8 ;
  assign n18155 = x7 ^ x6 ;
  assign n18156 = ~n7128 & ~n18155 ;
  assign n7144 = x8 & ~n18156 ;
  assign n7146 = n7145 ^ n7144 ;
  assign n8045 = n8044 ^ n7146 ;
  assign n8046 = ~n3943 & n8045 ;
  assign n8047 = n8046 ^ x8 ;
  assign n8034 = ~n317 & n6655 ;
  assign n8030 = n7069 ^ n6862 ;
  assign n8031 = n8030 ^ x11 ;
  assign n8029 = ~n445 & n6650 ;
  assign n8032 = n8031 ^ n8029 ;
  assign n6657 = n6656 ^ n6648 ;
  assign n6658 = n6657 ^ n6649 ;
  assign n8028 = ~n485 & n6658 ;
  assign n8033 = n8032 ^ n8028 ;
  assign n8035 = n8034 ^ n8033 ;
  assign n8027 = n3500 & n15413 ;
  assign n8036 = n8035 ^ n8027 ;
  assign n7698 = n7067 ^ n7056 ;
  assign n7699 = n7698 ^ x14 ;
  assign n7688 = ~n3473 & n4897 ;
  assign n7694 = x14 & ~n3388 ;
  assign n7696 = n7688 & n7694 ;
  assign n7691 = ~n824 & ~n6074 ;
  assign n7690 = ~n1109 & ~n6072 ;
  assign n7692 = n7691 ^ n7690 ;
  assign n8435 = n8434 ^ n6060 ;
  assign n7689 = n8435 ^ n7688 ;
  assign n7693 = n7692 ^ n7689 ;
  assign n7697 = n7696 ^ n7693 ;
  assign n7700 = n7699 ^ n7697 ;
  assign n7685 = n3473 & n6060 ;
  assign n7686 = n8434 ^ n7685 ;
  assign n7687 = ~n3388 & n7686 ;
  assign n7701 = n7700 ^ n7687 ;
  assign n7672 = ~n1540 & n5700 ;
  assign n7668 = n7053 ^ n6872 ;
  assign n7669 = n7668 ^ x17 ;
  assign n7667 = ~n1214 & n5702 ;
  assign n7670 = n7669 ^ n7667 ;
  assign n7666 = ~n1433 & n20731 ;
  assign n7671 = n7670 ^ n7666 ;
  assign n7673 = n7672 ^ n7671 ;
  assign n7665 = ~n4603 & n5703 ;
  assign n7674 = n7673 ^ n7665 ;
  assign n7594 = ~n1351 & n20731 ;
  assign n7590 = n7050 ^ n6882 ;
  assign n7591 = n7590 ^ x17 ;
  assign n7589 = ~n1540 & n5702 ;
  assign n7592 = n7591 ^ n7589 ;
  assign n7588 = ~n1433 & n5700 ;
  assign n7593 = n7592 ^ n7588 ;
  assign n7595 = n7594 ^ n7593 ;
  assign n7587 = ~n4610 & n5703 ;
  assign n7596 = n7595 ^ n7587 ;
  assign n7355 = ~n1631 & n4683 ;
  assign n7351 = n7047 ^ n6892 ;
  assign n7352 = n7351 ^ x20 ;
  assign n7350 = ~n1795 & n14027 ;
  assign n7353 = n7352 ^ n7350 ;
  assign n7349 = ~n1871 & n4916 ;
  assign n7354 = n7353 ^ n7349 ;
  assign n7356 = n7355 ^ n7354 ;
  assign n7348 = ~n4392 & n4684 ;
  assign n7357 = n7356 ^ n7348 ;
  assign n7167 = ~n2096 & n4491 ;
  assign n7165 = ~n2185 & ~n4496 ;
  assign n7163 = n4492 & n5196 ;
  assign n7161 = n7045 ^ n7034 ;
  assign n7162 = n7161 ^ x23 ;
  assign n7164 = n7163 ^ n7162 ;
  assign n7166 = n7165 ^ n7164 ;
  assign n7168 = n7167 ^ n7166 ;
  assign n7160 = ~n2268 & n4504 ;
  assign n7169 = n7168 ^ n7160 ;
  assign n7332 = n7032 ^ n7020 ;
  assign n7177 = ~n487 & ~n2486 ;
  assign n7173 = n7017 ^ n6903 ;
  assign n7174 = n7173 ^ x26 ;
  assign n7172 = ~n2609 & n12861 ;
  assign n7175 = n7174 ^ n7172 ;
  assign n7171 = n446 & ~n2554 ;
  assign n7176 = n7175 ^ n7171 ;
  assign n7178 = n7177 ^ n7176 ;
  assign n7170 = ~n3501 & n5381 ;
  assign n7179 = n7178 ^ n7170 ;
  assign n7316 = n7015 ^ n7004 ;
  assign n7187 = ~n2646 & n12861 ;
  assign n7183 = n7001 ^ n6914 ;
  assign n7184 = n7183 ^ x26 ;
  assign n7182 = n446 & ~n3227 ;
  assign n7185 = n7184 ^ n7182 ;
  assign n7181 = ~n487 & ~n2609 ;
  assign n7186 = n7185 ^ n7181 ;
  assign n7188 = n7187 ^ n7186 ;
  assign n7180 = ~n3501 & n7029 ;
  assign n7189 = n7188 ^ n7180 ;
  assign n7199 = ~n487 & ~n3227 ;
  assign n7194 = ~n6501 & n6992 ;
  assign n7193 = n6993 ^ n6461 ;
  assign n7195 = n7194 ^ n7193 ;
  assign n7196 = n7195 ^ x26 ;
  assign n7192 = n446 & ~n2646 ;
  assign n7197 = n7196 ^ n7192 ;
  assign n7191 = ~n2738 & n12861 ;
  assign n7198 = n7197 ^ n7191 ;
  assign n7200 = n7199 ^ n7198 ;
  assign n7190 = ~n3501 & n6900 ;
  assign n7201 = n7200 ^ n7190 ;
  assign n7295 = n6936 ^ n6473 ;
  assign n7296 = n7295 ^ n6498 ;
  assign n7297 = n7296 ^ n6986 ;
  assign n7282 = n6984 ^ n6971 ;
  assign n7268 = n6944 ^ n6943 ;
  assign n7265 = n6963 ^ n6944 ;
  assign n7266 = n7265 ^ n6947 ;
  assign n7267 = x29 & ~n7266 ;
  assign n7269 = n7268 ^ n7267 ;
  assign n7254 = ~n487 & ~n3151 ;
  assign n7253 = n446 & ~n2924 ;
  assign n7255 = n7254 ^ n7253 ;
  assign n7256 = n7255 ^ x26 ;
  assign n7252 = ~n2958 & n12861 ;
  assign n7257 = n7256 ^ n7252 ;
  assign n7251 = ~n3501 & n6286 ;
  assign n7258 = n7257 ^ n7251 ;
  assign n7210 = n826 & ~n3337 ;
  assign n7211 = n7210 ^ n6959 ;
  assign n7205 = n446 & ~n2958 ;
  assign n7204 = ~n3099 & n12861 ;
  assign n7206 = n7205 ^ n7204 ;
  assign n7207 = n7206 ^ x26 ;
  assign n7203 = ~n487 & ~n2924 ;
  assign n7208 = n7207 ^ n7203 ;
  assign n7202 = ~n3501 & n6344 ;
  assign n7209 = n7208 ^ n7202 ;
  assign n7212 = n7211 ^ n7209 ;
  assign n7213 = n650 & ~n3337 ;
  assign n7214 = n446 ^ n64 ;
  assign n7215 = n64 & ~n3027 ;
  assign n7216 = x26 & ~n7215 ;
  assign n7217 = n7214 & n7216 ;
  assign n7218 = ~n3337 & n7217 ;
  assign n7219 = n7218 ^ n7216 ;
  assign n7233 = ~n3337 & n12861 ;
  assign n7230 = n64 & ~n3099 ;
  assign n7231 = n467 & n3339 ;
  assign n7232 = n7230 & ~n7231 ;
  assign n7234 = n7233 ^ n7232 ;
  assign n7224 = n3099 & n3337 ;
  assign n7227 = ~n3501 & n7224 ;
  assign n7228 = n7227 ^ n446 ;
  assign n7229 = ~n3027 & n7228 ;
  assign n7235 = n7234 ^ n7229 ;
  assign n7236 = n7219 & ~n7235 ;
  assign n7237 = ~n7213 & ~n7236 ;
  assign n7241 = ~n487 & ~n2958 ;
  assign n7240 = n446 & ~n3099 ;
  assign n7242 = n7241 ^ n7240 ;
  assign n7243 = n7242 ^ x26 ;
  assign n7239 = ~n3027 & n12861 ;
  assign n7244 = n7243 ^ n7239 ;
  assign n7238 = ~n3501 & n6440 ;
  assign n7245 = n7244 ^ n7238 ;
  assign n7246 = n7237 & n7245 ;
  assign n7247 = n7246 ^ n7245 ;
  assign n7248 = n7247 ^ n7209 ;
  assign n7249 = n7212 & ~n7248 ;
  assign n7250 = n7249 ^ n7211 ;
  assign n7259 = n7258 ^ n7250 ;
  assign n7261 = x29 & n6962 ;
  assign n7260 = n7258 ^ n6958 ;
  assign n7262 = n7261 ^ n7260 ;
  assign n7263 = n7259 & n7262 ;
  assign n7264 = n7263 ^ n7258 ;
  assign n7270 = n7269 ^ n7264 ;
  assign n7277 = ~n487 & ~n2836 ;
  assign n7275 = n446 & ~n3151 ;
  assign n7273 = ~n2924 & n12861 ;
  assign n7272 = n7269 ^ x26 ;
  assign n7274 = n7273 ^ n7272 ;
  assign n7276 = n7275 ^ n7274 ;
  assign n7278 = n7277 ^ n7276 ;
  assign n7271 = ~n3501 & n6237 ;
  assign n7279 = n7278 ^ n7271 ;
  assign n7280 = n7270 & n7279 ;
  assign n7281 = n7280 ^ n7269 ;
  assign n7283 = n7282 ^ n7281 ;
  assign n7290 = ~n487 & ~n2738 ;
  assign n7288 = n446 & ~n2836 ;
  assign n7286 = ~n3151 & n12861 ;
  assign n7285 = n7282 ^ x26 ;
  assign n7287 = n7286 ^ n7285 ;
  assign n7289 = n7288 ^ n7287 ;
  assign n7291 = n7290 ^ n7289 ;
  assign n7284 = ~n3501 & ~n6907 ;
  assign n7292 = n7291 ^ n7284 ;
  assign n7293 = n7283 & n7292 ;
  assign n7294 = n7293 ^ n7282 ;
  assign n7298 = n7297 ^ n7294 ;
  assign n7305 = n446 & ~n2738 ;
  assign n7303 = ~n2836 & n12861 ;
  assign n7301 = ~n487 & ~n2646 ;
  assign n7300 = n7297 ^ x26 ;
  assign n7302 = n7301 ^ n7300 ;
  assign n7304 = n7303 ^ n7302 ;
  assign n7306 = n7305 ^ n7304 ;
  assign n7299 = ~n3501 & ~n5651 ;
  assign n7307 = n7306 ^ n7299 ;
  assign n7308 = n7298 & n7307 ;
  assign n7309 = n7308 ^ n7297 ;
  assign n7310 = n7309 ^ n7195 ;
  assign n7311 = ~n7201 & ~n7310 ;
  assign n7312 = n7311 ^ n7195 ;
  assign n7313 = n7312 ^ n7183 ;
  assign n7314 = n7189 & ~n7313 ;
  assign n7315 = n7314 ^ n7183 ;
  assign n7317 = n7316 ^ n7315 ;
  assign n7324 = ~n3227 & n12861 ;
  assign n7322 = ~n487 & ~n2554 ;
  assign n7320 = n446 & ~n2609 ;
  assign n7319 = n7316 ^ x26 ;
  assign n7321 = n7320 ^ n7319 ;
  assign n7323 = n7322 ^ n7321 ;
  assign n7325 = n7324 ^ n7323 ;
  assign n7318 = ~n3501 & n5541 ;
  assign n7326 = n7325 ^ n7318 ;
  assign n7327 = ~n7317 & ~n7326 ;
  assign n7328 = n7327 ^ n7316 ;
  assign n7329 = n7328 ^ n7173 ;
  assign n7330 = n7179 & ~n7329 ;
  assign n7331 = n7330 ^ n7173 ;
  assign n7333 = n7332 ^ n7331 ;
  assign n7340 = ~n487 & ~n2449 ;
  assign n7338 = ~n2554 & n12861 ;
  assign n7336 = n446 & ~n2486 ;
  assign n7335 = n7332 ^ x26 ;
  assign n7337 = n7336 ^ n7335 ;
  assign n7339 = n7338 ^ n7337 ;
  assign n7341 = n7340 ^ n7339 ;
  assign n7334 = ~n3501 & n5520 ;
  assign n7342 = n7341 ^ n7334 ;
  assign n7343 = n7333 & n7342 ;
  assign n7344 = n7343 ^ n7332 ;
  assign n7345 = n7344 ^ n7161 ;
  assign n7346 = ~n7169 & ~n7345 ;
  assign n7347 = n7346 ^ n7161 ;
  assign n7584 = n7351 ^ n7347 ;
  assign n7585 = n7357 & ~n7584 ;
  assign n7586 = n7585 ^ n7351 ;
  assign n7662 = n7590 ^ n7586 ;
  assign n7663 = n7596 & n7662 ;
  assign n7664 = n7663 ^ n7590 ;
  assign n7678 = n7668 ^ n7664 ;
  assign n7679 = n7674 & n7678 ;
  assign n7680 = n7679 ^ n7668 ;
  assign n8024 = n7698 ^ n7680 ;
  assign n8025 = ~n7701 & ~n8024 ;
  assign n8026 = n8025 ^ n7698 ;
  assign n8037 = n8036 ^ n8026 ;
  assign n7702 = n7701 ^ n7680 ;
  assign n8038 = n8037 ^ n7702 ;
  assign n7675 = n7674 ^ n7664 ;
  assign n7703 = n7702 ^ n7675 ;
  assign n7603 = x14 & n8434 ;
  assign n7636 = ~n824 & n7603 ;
  assign n7633 = ~n968 & ~n6072 ;
  assign n7632 = ~n1109 & ~n6074 ;
  assign n7634 = n7633 ^ n7632 ;
  assign n7635 = n7634 ^ x14 ;
  assign n7637 = n7636 ^ n7635 ;
  assign n7640 = ~n4050 & ~n7634 ;
  assign n7641 = n7640 ^ n824 ;
  assign n7642 = x13 & ~n7641 ;
  assign n7643 = n7642 ^ n824 ;
  assign n7644 = n4897 & ~n7643 ;
  assign n7647 = n7644 ^ n7636 ;
  assign n7648 = n7647 ^ n6057 ;
  assign n7649 = n7648 ^ n7647 ;
  assign n7652 = ~n4050 & n7649 ;
  assign n7653 = n7652 ^ n7647 ;
  assign n7654 = n7637 & ~n7653 ;
  assign n7655 = n7654 ^ n7647 ;
  assign n7656 = n7655 ^ x14 ;
  assign n7657 = n7655 ^ n7637 ;
  assign n7658 = ~n7654 & n7657 ;
  assign n7659 = ~n7656 & n7658 ;
  assign n7660 = n7659 ^ n7655 ;
  assign n7597 = n7596 ^ n7586 ;
  assign n7362 = ~n1351 & n5700 ;
  assign n7358 = n7357 ^ n7347 ;
  assign n7359 = n7358 ^ x17 ;
  assign n7159 = ~n1703 & n20731 ;
  assign n7360 = n7359 ^ n7159 ;
  assign n7158 = ~n1433 & n5702 ;
  assign n7361 = n7360 ^ n7158 ;
  assign n7363 = n7362 ^ n7361 ;
  assign n7157 = n4152 & n5703 ;
  assign n7364 = n7363 ^ n7157 ;
  assign n7372 = ~n1795 & n4916 ;
  assign n7368 = n7344 ^ n7169 ;
  assign n7369 = n7368 ^ x20 ;
  assign n7367 = ~n1994 & n14027 ;
  assign n7370 = n7369 ^ n7367 ;
  assign n7366 = ~n1871 & n4683 ;
  assign n7371 = n7370 ^ n7366 ;
  assign n7373 = n7372 ^ n7371 ;
  assign n7365 = n4684 & ~n4859 ;
  assign n7374 = n7373 ^ n7365 ;
  assign n7565 = n7342 ^ n7331 ;
  assign n7382 = ~n2449 & n4504 ;
  assign n7378 = n7328 ^ n7179 ;
  assign n7379 = n7378 ^ x23 ;
  assign n7377 = n4492 & n5144 ;
  assign n7380 = n7379 ^ n7377 ;
  assign n7376 = ~n2364 & ~n4496 ;
  assign n7381 = n7380 ^ n7376 ;
  assign n7383 = n7382 ^ n7381 ;
  assign n7375 = ~n2268 & n4491 ;
  assign n7384 = n7383 ^ n7375 ;
  assign n7549 = n7326 ^ n7315 ;
  assign n7392 = ~n2449 & n4491 ;
  assign n7388 = n7312 ^ n7189 ;
  assign n7389 = n7388 ^ x23 ;
  assign n7387 = n4492 & n5520 ;
  assign n7390 = n7389 ^ n7387 ;
  assign n7386 = ~n2486 & ~n4496 ;
  assign n7391 = n7390 ^ n7386 ;
  assign n7393 = n7392 ^ n7391 ;
  assign n7385 = ~n2554 & n4504 ;
  assign n7394 = n7393 ^ n7385 ;
  assign n7533 = n7309 ^ n7201 ;
  assign n7520 = n7307 ^ n7294 ;
  assign n7507 = n7292 ^ n7281 ;
  assign n7494 = n7279 ^ n7264 ;
  assign n7481 = n7262 ^ n7250 ;
  assign n7403 = n7247 ^ n7212 ;
  assign n7400 = ~n2738 & n4491 ;
  assign n7399 = ~n3151 & n4504 ;
  assign n7401 = n7400 ^ n7399 ;
  assign n7396 = ~n2836 & ~n4496 ;
  assign n7395 = n4492 & ~n6907 ;
  assign n7397 = n7396 ^ n7395 ;
  assign n7398 = n7397 ^ x23 ;
  assign n7402 = n7401 ^ n7398 ;
  assign n7404 = n7403 ^ n7402 ;
  assign n7413 = n7236 ^ n7213 ;
  assign n7414 = n7413 ^ n7245 ;
  assign n7410 = ~n2836 & n4491 ;
  assign n7409 = ~n2924 & n4504 ;
  assign n7411 = n7410 ^ n7409 ;
  assign n7406 = ~n3151 & ~n4496 ;
  assign n7405 = n4492 & n6237 ;
  assign n7407 = n7406 ^ n7405 ;
  assign n7408 = n7407 ^ x23 ;
  assign n7412 = n7411 ^ n7408 ;
  assign n7415 = n7414 ^ n7412 ;
  assign n7422 = ~n2958 & n4504 ;
  assign n7421 = ~n3151 & n4491 ;
  assign n7423 = n7422 ^ n7421 ;
  assign n7418 = ~n2924 & ~n4496 ;
  assign n7417 = n4492 & n6286 ;
  assign n7419 = n7418 ^ n7417 ;
  assign n7420 = n7419 ^ x23 ;
  assign n7424 = n7423 ^ n7420 ;
  assign n7474 = n7424 ^ n7414 ;
  assign n7220 = n7219 ^ x26 ;
  assign n7416 = n7235 ^ n7220 ;
  assign n7425 = n7424 ^ n7416 ;
  assign n7434 = n112 ^ n75 ;
  assign n7435 = ~n3337 & ~n7434 ;
  assign n7436 = n7435 ^ n7215 ;
  assign n7431 = ~n3099 & n4504 ;
  assign n7430 = ~n2924 & n4491 ;
  assign n7432 = n7431 ^ n7430 ;
  assign n7427 = ~n2958 & ~n4496 ;
  assign n7426 = n4492 & n6344 ;
  assign n7428 = n7427 ^ n7426 ;
  assign n7429 = n7428 ^ x23 ;
  assign n7433 = n7432 ^ n7429 ;
  assign n7437 = n7436 ^ n7433 ;
  assign n7438 = n64 & ~n3337 ;
  assign n7439 = ~n3027 & n4488 ;
  assign n7440 = x23 & ~n7439 ;
  assign n7441 = ~n4500 & n7440 ;
  assign n7442 = ~n3337 & n7441 ;
  assign n7443 = n7442 ^ n7440 ;
  assign n7454 = ~n3099 & n4488 ;
  assign n7453 = ~n3337 & n4504 ;
  assign n7455 = n7454 ^ n7453 ;
  assign n7450 = n3337 & n4492 ;
  assign n7451 = n7450 ^ n4496 ;
  assign n7452 = ~n3027 & ~n7451 ;
  assign n7456 = n7455 ^ n7452 ;
  assign n7457 = n7443 & ~n7456 ;
  assign n7458 = ~n7438 & ~n7457 ;
  assign n7464 = ~n2958 & n4491 ;
  assign n7463 = ~n3027 & n4504 ;
  assign n7465 = n7464 ^ n7463 ;
  assign n7460 = ~n3099 & ~n4496 ;
  assign n7459 = n4492 & n6440 ;
  assign n7461 = n7460 ^ n7459 ;
  assign n7462 = n7461 ^ x23 ;
  assign n7466 = n7465 ^ n7462 ;
  assign n7467 = n7458 & n7466 ;
  assign n7468 = n7467 ^ n7466 ;
  assign n7469 = n7468 ^ n7433 ;
  assign n7470 = n7437 & ~n7469 ;
  assign n7471 = n7470 ^ n7436 ;
  assign n7472 = n7471 ^ n7424 ;
  assign n7473 = n7425 & n7472 ;
  assign n7475 = n7474 ^ n7473 ;
  assign n7476 = n7415 & n7475 ;
  assign n7477 = n7476 ^ n7414 ;
  assign n7478 = n7477 ^ n7402 ;
  assign n7479 = n7404 & n7478 ;
  assign n7480 = n7479 ^ n7402 ;
  assign n7482 = n7481 ^ n7480 ;
  assign n7489 = ~n2646 & n4491 ;
  assign n7487 = ~n2738 & ~n4496 ;
  assign n7485 = n4492 & ~n5651 ;
  assign n7484 = n7481 ^ x23 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7488 = n7487 ^ n7486 ;
  assign n7490 = n7489 ^ n7488 ;
  assign n7483 = ~n2836 & n4504 ;
  assign n7491 = n7490 ^ n7483 ;
  assign n7492 = n7482 & n7491 ;
  assign n7493 = n7492 ^ n7481 ;
  assign n7495 = n7494 ^ n7493 ;
  assign n7502 = ~n2646 & ~n4496 ;
  assign n7500 = ~n2738 & n4504 ;
  assign n7498 = n4492 & n6900 ;
  assign n7497 = n7494 ^ x23 ;
  assign n7499 = n7498 ^ n7497 ;
  assign n7501 = n7500 ^ n7499 ;
  assign n7503 = n7502 ^ n7501 ;
  assign n7496 = ~n3227 & n4491 ;
  assign n7504 = n7503 ^ n7496 ;
  assign n7505 = n7495 & n7504 ;
  assign n7506 = n7505 ^ n7494 ;
  assign n7508 = n7507 ^ n7506 ;
  assign n7515 = ~n2646 & n4504 ;
  assign n7513 = ~n3227 & ~n4496 ;
  assign n7511 = n4492 & n7029 ;
  assign n7510 = n7507 ^ x23 ;
  assign n7512 = n7511 ^ n7510 ;
  assign n7514 = n7513 ^ n7512 ;
  assign n7516 = n7515 ^ n7514 ;
  assign n7509 = ~n2609 & n4491 ;
  assign n7517 = n7516 ^ n7509 ;
  assign n7518 = n7508 & n7517 ;
  assign n7519 = n7518 ^ n7507 ;
  assign n7521 = n7520 ^ n7519 ;
  assign n7528 = ~n3227 & n4504 ;
  assign n7526 = ~n2609 & ~n4496 ;
  assign n7524 = n4492 & n5541 ;
  assign n7523 = n7520 ^ x23 ;
  assign n7525 = n7524 ^ n7523 ;
  assign n7527 = n7526 ^ n7525 ;
  assign n7529 = n7528 ^ n7527 ;
  assign n7522 = ~n2554 & n4491 ;
  assign n7530 = n7529 ^ n7522 ;
  assign n7531 = n7521 & n7530 ;
  assign n7532 = n7531 ^ n7520 ;
  assign n7534 = n7533 ^ n7532 ;
  assign n7541 = ~n2609 & n4504 ;
  assign n7539 = ~n2554 & ~n4496 ;
  assign n7537 = n4492 & n5381 ;
  assign n7536 = n7533 ^ x23 ;
  assign n7538 = n7537 ^ n7536 ;
  assign n7540 = n7539 ^ n7538 ;
  assign n7542 = n7541 ^ n7540 ;
  assign n7535 = ~n2486 & n4491 ;
  assign n7543 = n7542 ^ n7535 ;
  assign n7544 = ~n7534 & ~n7543 ;
  assign n7545 = n7544 ^ n7533 ;
  assign n7546 = n7545 ^ n7388 ;
  assign n7547 = ~n7394 & n7546 ;
  assign n7548 = n7547 ^ n7388 ;
  assign n7550 = n7549 ^ n7548 ;
  assign n7557 = ~n2364 & n4491 ;
  assign n7555 = ~n2449 & ~n4496 ;
  assign n7553 = n4492 & n5283 ;
  assign n7552 = n7549 ^ x23 ;
  assign n7554 = n7553 ^ n7552 ;
  assign n7556 = n7555 ^ n7554 ;
  assign n7558 = n7557 ^ n7556 ;
  assign n7551 = ~n2486 & n4504 ;
  assign n7559 = n7558 ^ n7551 ;
  assign n7560 = n7550 & ~n7559 ;
  assign n7561 = n7560 ^ n7549 ;
  assign n7562 = n7561 ^ n7378 ;
  assign n7563 = ~n7384 & n7562 ;
  assign n7564 = n7563 ^ n7378 ;
  assign n7566 = n7565 ^ n7564 ;
  assign n7573 = ~n2364 & n4504 ;
  assign n7571 = ~n2268 & ~n4496 ;
  assign n7569 = n4492 & n5832 ;
  assign n7568 = n7565 ^ x23 ;
  assign n7570 = n7569 ^ n7568 ;
  assign n7572 = n7571 ^ n7570 ;
  assign n7574 = n7573 ^ n7572 ;
  assign n7567 = ~n2185 & n4491 ;
  assign n7575 = n7574 ^ n7567 ;
  assign n7576 = ~n7566 & n7575 ;
  assign n7577 = n7576 ^ n7565 ;
  assign n7578 = n7577 ^ n7368 ;
  assign n7579 = ~n7374 & ~n7578 ;
  assign n7580 = n7579 ^ n7368 ;
  assign n7581 = n7580 ^ n7358 ;
  assign n7582 = ~n7364 & n7581 ;
  assign n7583 = n7582 ^ n7358 ;
  assign n7598 = n7597 ^ n7583 ;
  assign n7604 = ~n1109 & n7603 ;
  assign n7600 = ~n968 & ~n6074 ;
  assign n7599 = ~n1214 & ~n6072 ;
  assign n7601 = n7600 ^ n7599 ;
  assign n7602 = n7601 ^ x14 ;
  assign n7605 = n7604 ^ n7602 ;
  assign n7606 = n7605 ^ x14 ;
  assign n7611 = x13 & ~n3904 ;
  assign n7612 = n7611 ^ n1109 ;
  assign n7613 = n4897 & ~n7612 ;
  assign n7615 = n7613 ^ n7604 ;
  assign n7616 = n7615 ^ n6057 ;
  assign n7617 = n7616 ^ n7615 ;
  assign n7618 = n7615 ^ n3905 ;
  assign n7619 = n7618 ^ n7615 ;
  assign n7620 = n7617 & n7619 ;
  assign n7621 = n7620 ^ n7615 ;
  assign n7622 = n7605 & ~n7621 ;
  assign n7623 = n7606 & ~n7622 ;
  assign n7624 = n7615 ^ n7597 ;
  assign n7625 = n7624 ^ n7622 ;
  assign n7626 = n7625 ^ x14 ;
  assign n7627 = n7626 ^ n7597 ;
  assign n7628 = n7623 & ~n7627 ;
  assign n7629 = n7628 ^ n7625 ;
  assign n7630 = ~n7598 & n7629 ;
  assign n7631 = n7630 ^ n7597 ;
  assign n7661 = n7660 ^ n7631 ;
  assign n7676 = n7675 ^ n7660 ;
  assign n7677 = ~n7661 & n7676 ;
  assign n7704 = n7703 ^ n7677 ;
  assign n7152 = ~n445 & n6658 ;
  assign n7151 = ~n317 & n6650 ;
  assign n7153 = n7152 ^ n7151 ;
  assign n7154 = n7153 ^ x11 ;
  assign n7150 = ~n649 & n6655 ;
  assign n7155 = n7154 ^ n7150 ;
  assign n7149 = n4073 & n15413 ;
  assign n7156 = n7155 ^ n7149 ;
  assign n8022 = n7702 ^ n7156 ;
  assign n8023 = ~n7704 & ~n8022 ;
  assign n8039 = n8038 ^ n8023 ;
  assign n8048 = n8047 ^ n8039 ;
  assign n7705 = n7704 ^ n7156 ;
  assign n7706 = n7705 ^ x8 ;
  assign n7140 = n7137 ^ x7 ;
  assign n7141 = n7140 ^ n7132 ;
  assign n7148 = ~n3943 & n7141 ;
  assign n7707 = n7706 ^ n7148 ;
  assign n7147 = ~n485 & n7146 ;
  assign n7708 = n7707 ^ n7147 ;
  assign n7136 = n4515 & n7135 ;
  assign n7709 = n7708 ^ n7136 ;
  assign n8006 = n7676 ^ n7631 ;
  assign n7717 = ~n3473 & n6650 ;
  assign n7713 = n7629 ^ n7583 ;
  assign n7714 = n7713 ^ x11 ;
  assign n7712 = ~n649 & n6658 ;
  assign n7715 = n7714 ^ n7712 ;
  assign n7711 = ~n824 & n6655 ;
  assign n7716 = n7715 ^ n7711 ;
  assign n7718 = n7717 ^ n7716 ;
  assign n7710 = ~n3476 & n15413 ;
  assign n7719 = n7718 ^ n7710 ;
  assign n7968 = n7580 ^ n7364 ;
  assign n7727 = ~n1351 & n5702 ;
  assign n7723 = n7577 ^ n7374 ;
  assign n7724 = n7723 ^ x17 ;
  assign n7722 = ~n1703 & n5700 ;
  assign n7725 = n7724 ^ n7722 ;
  assign n7721 = ~n1631 & n20731 ;
  assign n7726 = n7725 ^ n7721 ;
  assign n7728 = n7727 ^ n7726 ;
  assign n7720 = n4417 & n5703 ;
  assign n7729 = n7728 ^ n7720 ;
  assign n7950 = n7575 ^ n7564 ;
  assign n7737 = ~n2185 & n14027 ;
  assign n7733 = n7561 ^ n7384 ;
  assign n7734 = n7733 ^ x20 ;
  assign n7732 = ~n1994 & n4683 ;
  assign n7735 = n7734 ^ n7732 ;
  assign n7731 = ~n2096 & n4916 ;
  assign n7736 = n7735 ^ n7731 ;
  assign n7738 = n7737 ^ n7736 ;
  assign n7730 = n4684 & n5409 ;
  assign n7739 = n7738 ^ n7730 ;
  assign n7934 = n7559 ^ n7548 ;
  assign n7747 = ~n2268 & n4916 ;
  assign n7743 = n7545 ^ n7394 ;
  assign n7744 = n7743 ^ x20 ;
  assign n7742 = ~n2364 & n14027 ;
  assign n7745 = n7744 ^ n7742 ;
  assign n7741 = ~n2185 & n4683 ;
  assign n7746 = n7745 ^ n7741 ;
  assign n7748 = n7747 ^ n7746 ;
  assign n7740 = n4684 & n5832 ;
  assign n7749 = n7748 ^ n7740 ;
  assign n7918 = n7543 ^ n7532 ;
  assign n7758 = n7530 ^ n7519 ;
  assign n7753 = ~n2449 & n4916 ;
  assign n7752 = ~n2364 & n4683 ;
  assign n7754 = n7753 ^ n7752 ;
  assign n7755 = n7754 ^ x20 ;
  assign n7751 = ~n2486 & n14027 ;
  assign n7756 = n7755 ^ n7751 ;
  assign n7750 = n4684 & n5283 ;
  assign n7757 = n7756 ^ n7750 ;
  assign n7759 = n7758 ^ n7757 ;
  assign n7890 = n7504 ^ n7493 ;
  assign n7877 = n7491 ^ n7480 ;
  assign n7864 = n7477 ^ n7404 ;
  assign n7851 = n7475 ^ n7412 ;
  assign n7769 = n7471 ^ n7425 ;
  assign n7764 = ~n2738 & n4916 ;
  assign n7763 = ~n2836 & n14027 ;
  assign n7765 = n7764 ^ n7763 ;
  assign n7766 = n7765 ^ x20 ;
  assign n7762 = ~n2646 & n4683 ;
  assign n7767 = n7766 ^ n7762 ;
  assign n7761 = n4684 & ~n5651 ;
  assign n7768 = n7767 ^ n7761 ;
  assign n7770 = n7769 ^ n7768 ;
  assign n7779 = n7468 ^ n7437 ;
  assign n7774 = ~n2738 & n4683 ;
  assign n7773 = ~n2836 & n4916 ;
  assign n7775 = n7774 ^ n7773 ;
  assign n7776 = n7775 ^ x20 ;
  assign n7772 = ~n3151 & n14027 ;
  assign n7777 = n7776 ^ n7772 ;
  assign n7771 = n4684 & ~n6907 ;
  assign n7778 = n7777 ^ n7771 ;
  assign n7780 = n7779 ^ n7778 ;
  assign n7789 = n7457 ^ n7438 ;
  assign n7790 = n7789 ^ n7466 ;
  assign n7784 = ~n3151 & n4916 ;
  assign n7783 = ~n2924 & n14027 ;
  assign n7785 = n7784 ^ n7783 ;
  assign n7786 = n7785 ^ x20 ;
  assign n7782 = ~n2836 & n4683 ;
  assign n7787 = n7786 ^ n7782 ;
  assign n7781 = n4684 & n6237 ;
  assign n7788 = n7787 ^ n7781 ;
  assign n7791 = n7790 ^ n7788 ;
  assign n7444 = n7443 ^ x23 ;
  assign n7800 = n7456 ^ n7444 ;
  assign n7795 = ~n3151 & n4683 ;
  assign n7794 = ~n2924 & n4916 ;
  assign n7796 = n7795 ^ n7794 ;
  assign n7797 = n7796 ^ x20 ;
  assign n7793 = ~n2958 & n14027 ;
  assign n7798 = n7797 ^ n7793 ;
  assign n7792 = n4684 & n6286 ;
  assign n7799 = n7798 ^ n7792 ;
  assign n7801 = n7800 ^ n7799 ;
  assign n7810 = n4495 ^ x22 ;
  assign n7811 = ~n3337 & ~n7810 ;
  assign n7812 = n7811 ^ n7439 ;
  assign n7805 = ~n2958 & n4916 ;
  assign n7804 = ~n3099 & n14027 ;
  assign n7806 = n7805 ^ n7804 ;
  assign n7807 = n7806 ^ x20 ;
  assign n7803 = ~n2924 & n4683 ;
  assign n7808 = n7807 ^ n7803 ;
  assign n7802 = n4684 & n6344 ;
  assign n7809 = n7808 ^ n7802 ;
  assign n7813 = n7812 ^ n7809 ;
  assign n7814 = ~n3337 & n4488 ;
  assign n7818 = ~n2958 & n4683 ;
  assign n7817 = ~n3027 & n14027 ;
  assign n7819 = n7818 ^ n7817 ;
  assign n7820 = n7819 ^ x20 ;
  assign n7816 = ~n3099 & n4916 ;
  assign n7821 = n7820 ^ n7816 ;
  assign n7815 = n4684 & n6440 ;
  assign n7822 = n7821 ^ n7815 ;
  assign n7823 = ~n7814 & n7822 ;
  assign n7824 = n4916 ^ n4678 ;
  assign n7828 = ~n3337 & n14027 ;
  assign n7825 = ~n3099 & n4678 ;
  assign n7826 = n3339 & n4685 ;
  assign n7827 = n7825 & ~n7826 ;
  assign n7829 = n7828 ^ n7827 ;
  assign n7830 = x20 & ~n7829 ;
  assign n7831 = ~n3338 & n7830 ;
  assign n7832 = n7824 & n7831 ;
  assign n7833 = n7832 ^ n7830 ;
  assign n7834 = n7823 & ~n7833 ;
  assign n7835 = n7834 ^ n7822 ;
  assign n7836 = n7835 ^ n7809 ;
  assign n7837 = n7813 & ~n7836 ;
  assign n7838 = n7837 ^ n7812 ;
  assign n7839 = n7838 ^ n7799 ;
  assign n7840 = n7801 & n7839 ;
  assign n7841 = n7840 ^ n7799 ;
  assign n7842 = n7841 ^ n7788 ;
  assign n7843 = n7791 & n7842 ;
  assign n7844 = n7843 ^ n7788 ;
  assign n7845 = n7844 ^ n7778 ;
  assign n7846 = n7780 & n7845 ;
  assign n7847 = n7846 ^ n7778 ;
  assign n7848 = n7847 ^ n7768 ;
  assign n7849 = n7770 & n7848 ;
  assign n7850 = n7849 ^ n7768 ;
  assign n7852 = n7851 ^ n7850 ;
  assign n7859 = ~n3227 & n4683 ;
  assign n7857 = ~n2738 & n14027 ;
  assign n7855 = ~n2646 & n4916 ;
  assign n7854 = n7851 ^ x20 ;
  assign n7856 = n7855 ^ n7854 ;
  assign n7858 = n7857 ^ n7856 ;
  assign n7860 = n7859 ^ n7858 ;
  assign n7853 = n4684 & n6900 ;
  assign n7861 = n7860 ^ n7853 ;
  assign n7862 = n7852 & n7861 ;
  assign n7863 = n7862 ^ n7851 ;
  assign n7865 = n7864 ^ n7863 ;
  assign n7872 = ~n2609 & n4683 ;
  assign n7870 = ~n3227 & n4916 ;
  assign n7868 = ~n2646 & n14027 ;
  assign n7867 = n7864 ^ x20 ;
  assign n7869 = n7868 ^ n7867 ;
  assign n7871 = n7870 ^ n7869 ;
  assign n7873 = n7872 ^ n7871 ;
  assign n7866 = n4684 & n7029 ;
  assign n7874 = n7873 ^ n7866 ;
  assign n7875 = n7865 & n7874 ;
  assign n7876 = n7875 ^ n7864 ;
  assign n7878 = n7877 ^ n7876 ;
  assign n7885 = ~n2554 & n4683 ;
  assign n7883 = ~n2609 & n4916 ;
  assign n7881 = ~n3227 & n14027 ;
  assign n7880 = n7877 ^ x20 ;
  assign n7882 = n7881 ^ n7880 ;
  assign n7884 = n7883 ^ n7882 ;
  assign n7886 = n7885 ^ n7884 ;
  assign n7879 = n4684 & n5541 ;
  assign n7887 = n7886 ^ n7879 ;
  assign n7888 = n7878 & n7887 ;
  assign n7889 = n7888 ^ n7877 ;
  assign n7891 = n7890 ^ n7889 ;
  assign n7898 = ~n2486 & n4683 ;
  assign n7896 = ~n2554 & n4916 ;
  assign n7894 = ~n2609 & n14027 ;
  assign n7893 = n7890 ^ x20 ;
  assign n7895 = n7894 ^ n7893 ;
  assign n7897 = n7896 ^ n7895 ;
  assign n7899 = n7898 ^ n7897 ;
  assign n7892 = n4684 & n5381 ;
  assign n7900 = n7899 ^ n7892 ;
  assign n7901 = n7891 & n7900 ;
  assign n7902 = n7901 ^ n7890 ;
  assign n7914 = n7902 ^ n7757 ;
  assign n7760 = n7517 ^ n7506 ;
  assign n7903 = n7902 ^ n7760 ;
  assign n7910 = ~n2449 & n4683 ;
  assign n7908 = ~n2554 & n14027 ;
  assign n7906 = ~n2486 & n4916 ;
  assign n7905 = n7760 ^ x20 ;
  assign n7907 = n7906 ^ n7905 ;
  assign n7909 = n7908 ^ n7907 ;
  assign n7911 = n7910 ^ n7909 ;
  assign n7904 = n4684 & n5520 ;
  assign n7912 = n7911 ^ n7904 ;
  assign n7913 = n7903 & ~n7912 ;
  assign n7915 = n7914 ^ n7913 ;
  assign n7916 = n7759 & ~n7915 ;
  assign n7917 = n7916 ^ n7758 ;
  assign n7919 = n7918 ^ n7917 ;
  assign n7926 = ~n2268 & n4683 ;
  assign n7924 = ~n2449 & n14027 ;
  assign n7922 = ~n2364 & n4916 ;
  assign n7921 = n7918 ^ x20 ;
  assign n7923 = n7922 ^ n7921 ;
  assign n7925 = n7924 ^ n7923 ;
  assign n7927 = n7926 ^ n7925 ;
  assign n7920 = n4684 & n5144 ;
  assign n7928 = n7927 ^ n7920 ;
  assign n7929 = ~n7919 & ~n7928 ;
  assign n7930 = n7929 ^ n7918 ;
  assign n7931 = n7930 ^ n7743 ;
  assign n7932 = n7749 & ~n7931 ;
  assign n7933 = n7932 ^ n7743 ;
  assign n7935 = n7934 ^ n7933 ;
  assign n7942 = ~n2096 & n4683 ;
  assign n7940 = ~n2268 & n14027 ;
  assign n7938 = ~n2185 & n4916 ;
  assign n7937 = n7934 ^ x20 ;
  assign n7939 = n7938 ^ n7937 ;
  assign n7941 = n7940 ^ n7939 ;
  assign n7943 = n7942 ^ n7941 ;
  assign n7936 = n4684 & n5196 ;
  assign n7944 = n7943 ^ n7936 ;
  assign n7945 = n7935 & n7944 ;
  assign n7946 = n7945 ^ n7934 ;
  assign n7947 = n7946 ^ n7733 ;
  assign n7948 = n7739 & n7947 ;
  assign n7949 = n7948 ^ n7733 ;
  assign n7951 = n7950 ^ n7949 ;
  assign n7959 = n7950 ^ x20 ;
  assign n7958 = ~n2096 & n14027 ;
  assign n7960 = n7959 ^ n7958 ;
  assign n7957 = ~n1994 & n4916 ;
  assign n7961 = n7960 ^ n7957 ;
  assign n7954 = ~n4384 & n4685 ;
  assign n7955 = n7954 ^ n1795 ;
  assign n7956 = n4678 & ~n7955 ;
  assign n7962 = n7961 ^ n7956 ;
  assign n7963 = ~n7951 & ~n7962 ;
  assign n7964 = n7963 ^ n7950 ;
  assign n7965 = n7964 ^ n7723 ;
  assign n7966 = ~n7729 & n7965 ;
  assign n7967 = n7966 ^ n7723 ;
  assign n7969 = n7968 ^ n7967 ;
  assign n7974 = ~n968 & n7603 ;
  assign n7971 = ~n1214 & ~n6074 ;
  assign n7970 = ~n1540 & ~n6072 ;
  assign n7972 = n7971 ^ n7970 ;
  assign n7973 = n7972 ^ x14 ;
  assign n7975 = n7974 ^ n7973 ;
  assign n7976 = n7975 ^ x14 ;
  assign n7982 = x13 & ~n3381 ;
  assign n7983 = n7982 ^ n968 ;
  assign n7984 = n4897 & ~n7983 ;
  assign n7986 = n7984 ^ n7974 ;
  assign n7987 = n7986 ^ n6057 ;
  assign n7988 = n7987 ^ n7986 ;
  assign n7989 = n7986 ^ n3521 ;
  assign n7990 = n7989 ^ n7986 ;
  assign n7991 = n7988 & n7990 ;
  assign n7992 = n7991 ^ n7986 ;
  assign n7993 = n7975 & ~n7992 ;
  assign n7994 = n7976 & ~n7993 ;
  assign n7995 = n7986 ^ n7968 ;
  assign n7996 = n7995 ^ n7993 ;
  assign n7997 = n7996 ^ x14 ;
  assign n7998 = n7997 ^ n7968 ;
  assign n7999 = n7994 & ~n7998 ;
  assign n8000 = n7999 ^ n7996 ;
  assign n8001 = ~n7969 & n8000 ;
  assign n8002 = n8001 ^ n7968 ;
  assign n8003 = n8002 ^ n7713 ;
  assign n8004 = ~n7719 & ~n8003 ;
  assign n8005 = n8004 ^ n7713 ;
  assign n8007 = n8006 ^ n8005 ;
  assign n8014 = ~n649 & n6650 ;
  assign n8012 = ~n317 & n6658 ;
  assign n8010 = ~n3473 & n6655 ;
  assign n8009 = n8006 ^ x11 ;
  assign n8011 = n8010 ^ n8009 ;
  assign n8013 = n8012 ^ n8011 ;
  assign n8015 = n8014 ^ n8013 ;
  assign n8008 = n3956 & n15413 ;
  assign n8016 = n8015 ^ n8008 ;
  assign n8017 = ~n8007 & n8016 ;
  assign n8018 = n8017 ^ n8006 ;
  assign n8019 = n8018 ^ n7705 ;
  assign n8020 = ~n7709 & ~n8019 ;
  assign n8021 = n8020 ^ n7705 ;
  assign n8049 = n8048 ^ n8021 ;
  assign n11522 = n8018 ^ n7709 ;
  assign n11519 = n8016 ^ n8005 ;
  assign n11534 = n11522 ^ n11519 ;
  assign n8069 = ~n824 & n6650 ;
  assign n8065 = n8000 ^ n7967 ;
  assign n8066 = n8065 ^ x11 ;
  assign n8064 = ~n1109 & n6655 ;
  assign n8067 = n8066 ^ n8064 ;
  assign n8063 = ~n3473 & n6658 ;
  assign n8068 = n8067 ^ n8063 ;
  assign n8070 = n8069 ^ n8068 ;
  assign n8062 = ~n3508 & n15413 ;
  assign n8071 = n8070 ^ n8062 ;
  assign n8075 = ~n1433 & ~n6072 ;
  assign n8074 = ~n1540 & ~n6074 ;
  assign n8076 = n8075 ^ n8074 ;
  assign n8085 = n8076 ^ x14 ;
  assign n8084 = n7964 ^ n7729 ;
  assign n8086 = n8085 ^ n8084 ;
  assign n8077 = n8076 ^ n1214 ;
  assign n8072 = n4899 ^ n1214 ;
  assign n8078 = n8077 ^ n8072 ;
  assign n8081 = ~n3376 & n8078 ;
  assign n8082 = n8081 ^ n8072 ;
  assign n8083 = n4897 & ~n8082 ;
  assign n8087 = n8086 ^ n8083 ;
  assign n8376 = n7962 ^ n7949 ;
  assign n8095 = ~n1795 & n20731 ;
  assign n8091 = n7946 ^ n7739 ;
  assign n8092 = n8091 ^ x17 ;
  assign n8090 = ~n1871 & n5700 ;
  assign n8093 = n8092 ^ n8090 ;
  assign n8089 = ~n1631 & n5702 ;
  assign n8094 = n8093 ^ n8089 ;
  assign n8096 = n8095 ^ n8094 ;
  assign n8088 = ~n4392 & n5703 ;
  assign n8097 = n8096 ^ n8088 ;
  assign n8360 = n7944 ^ n7933 ;
  assign n8105 = ~n1795 & n5702 ;
  assign n8101 = n7930 ^ n7749 ;
  assign n8102 = n8101 ^ x17 ;
  assign n8100 = ~n1994 & n5700 ;
  assign n8103 = n8102 ^ n8100 ;
  assign n8099 = ~n2096 & n20731 ;
  assign n8104 = n8103 ^ n8099 ;
  assign n8106 = n8105 ^ n8104 ;
  assign n8098 = n5168 & n5703 ;
  assign n8107 = n8106 ^ n8098 ;
  assign n8344 = n7928 ^ n7917 ;
  assign n8331 = n7915 ^ n7758 ;
  assign n8112 = ~n2364 & n5700 ;
  assign n8110 = ~n2268 & n5702 ;
  assign n8109 = ~n2449 & n20731 ;
  assign n8111 = n8110 ^ n8109 ;
  assign n8113 = n8112 ^ n8111 ;
  assign n8108 = n5144 & n5703 ;
  assign n8114 = n8113 ^ n8108 ;
  assign n8115 = n8114 ^ x17 ;
  assign n8121 = ~n2364 & n20731 ;
  assign n8119 = ~n2268 & n5700 ;
  assign n8118 = ~n2185 & n5702 ;
  assign n8120 = n8119 ^ n8118 ;
  assign n8122 = n8121 ^ n8120 ;
  assign n8117 = n5703 & n5832 ;
  assign n8123 = n8122 ^ n8117 ;
  assign n8124 = n8123 ^ n8114 ;
  assign n8116 = n7912 ^ n7902 ;
  assign n8125 = n8124 ^ n8116 ;
  assign n8126 = ~n8115 & n8125 ;
  assign n8306 = n7887 ^ n7876 ;
  assign n8293 = n7874 ^ n7863 ;
  assign n8280 = n7861 ^ n7850 ;
  assign n8267 = n7847 ^ n7770 ;
  assign n8254 = n7844 ^ n7780 ;
  assign n8241 = n7841 ^ n7791 ;
  assign n8228 = n7838 ^ n7801 ;
  assign n8135 = n7835 ^ n7813 ;
  assign n8130 = ~n2738 & n5702 ;
  assign n8129 = ~n2836 & n5700 ;
  assign n8131 = n8130 ^ n8129 ;
  assign n8132 = n8131 ^ x17 ;
  assign n8128 = ~n3151 & n20731 ;
  assign n8133 = n8132 ^ n8128 ;
  assign n8127 = n5703 & ~n6907 ;
  assign n8134 = n8133 ^ n8127 ;
  assign n8136 = n8135 ^ n8134 ;
  assign n8145 = n7833 ^ n7814 ;
  assign n8146 = n8145 ^ n7822 ;
  assign n8140 = ~n2836 & n5702 ;
  assign n8139 = ~n2924 & n20731 ;
  assign n8141 = n8140 ^ n8139 ;
  assign n8142 = n8141 ^ x17 ;
  assign n8138 = ~n3151 & n5700 ;
  assign n8143 = n8142 ^ n8138 ;
  assign n8137 = n5703 & n6237 ;
  assign n8144 = n8143 ^ n8137 ;
  assign n8147 = n8146 ^ n8144 ;
  assign n8198 = ~n2958 & n20731 ;
  assign n8197 = ~n3151 & n5702 ;
  assign n8199 = n8198 ^ n8197 ;
  assign n8200 = n8199 ^ x17 ;
  assign n8196 = ~n2924 & n5700 ;
  assign n8201 = n8200 ^ n8196 ;
  assign n8195 = n5703 & n6286 ;
  assign n8202 = n8201 ^ n8195 ;
  assign n8158 = ~n3027 & n4678 ;
  assign n8156 = n4677 ^ x19 ;
  assign n8157 = ~n3337 & n8156 ;
  assign n8159 = n8158 ^ n8157 ;
  assign n8151 = ~n3099 & n20731 ;
  assign n8150 = ~n2924 & n5702 ;
  assign n8152 = n8151 ^ n8150 ;
  assign n8153 = n8152 ^ x17 ;
  assign n8149 = ~n2958 & n5700 ;
  assign n8154 = n8153 ^ n8149 ;
  assign n8148 = n5703 & n6344 ;
  assign n8155 = n8154 ^ n8148 ;
  assign n8160 = n8159 ^ n8155 ;
  assign n8161 = ~n3337 & n4678 ;
  assign n8162 = ~n3027 & n5693 ;
  assign n8163 = x17 & ~n8162 ;
  assign n8164 = n5705 & n8163 ;
  assign n8165 = ~n3337 & n8164 ;
  assign n8166 = n8165 ^ n8163 ;
  assign n8178 = ~n3099 & n5693 ;
  assign n8176 = ~n3337 & n20731 ;
  assign n8173 = n3337 & n5703 ;
  assign n8174 = n8173 ^ n5700 ;
  assign n8175 = ~n3027 & n8174 ;
  assign n8177 = n8176 ^ n8175 ;
  assign n8179 = n8178 ^ n8177 ;
  assign n8180 = n8166 & ~n8179 ;
  assign n8181 = ~n8161 & ~n8180 ;
  assign n8185 = ~n2958 & n5702 ;
  assign n8184 = ~n3099 & n5700 ;
  assign n8186 = n8185 ^ n8184 ;
  assign n8187 = n8186 ^ x17 ;
  assign n8183 = ~n3027 & n20731 ;
  assign n8188 = n8187 ^ n8183 ;
  assign n8182 = n5703 & n6440 ;
  assign n8189 = n8188 ^ n8182 ;
  assign n8190 = n8181 & n8189 ;
  assign n8191 = n8190 ^ n8189 ;
  assign n8192 = n8191 ^ n8155 ;
  assign n8193 = n8160 & ~n8192 ;
  assign n8194 = n8193 ^ n8159 ;
  assign n8203 = n8202 ^ n8194 ;
  assign n8213 = ~x19 & ~n4676 ;
  assign n8212 = n4687 ^ x19 ;
  assign n8214 = n8213 ^ n8212 ;
  assign n8217 = n3337 & ~n8158 ;
  assign n8218 = ~n8214 & n8217 ;
  assign n8211 = n8202 ^ n7829 ;
  assign n8215 = n8214 ^ n8211 ;
  assign n8208 = n4684 & n7224 ;
  assign n8209 = n8208 ^ n4916 ;
  assign n8210 = ~n3027 & n8209 ;
  assign n8216 = n8215 ^ n8210 ;
  assign n8219 = n8218 ^ n8216 ;
  assign n8220 = n8203 & ~n8219 ;
  assign n8221 = n8220 ^ n8202 ;
  assign n8222 = n8221 ^ n8144 ;
  assign n8223 = n8147 & n8222 ;
  assign n8224 = n8223 ^ n8144 ;
  assign n8225 = n8224 ^ n8134 ;
  assign n8226 = n8136 & n8225 ;
  assign n8227 = n8226 ^ n8134 ;
  assign n8229 = n8228 ^ n8227 ;
  assign n8236 = ~n2836 & n20731 ;
  assign n8234 = ~n2738 & n5700 ;
  assign n8232 = ~n2646 & n5702 ;
  assign n8231 = n8228 ^ x17 ;
  assign n8233 = n8232 ^ n8231 ;
  assign n8235 = n8234 ^ n8233 ;
  assign n8237 = n8236 ^ n8235 ;
  assign n8230 = ~n5651 & n5703 ;
  assign n8238 = n8237 ^ n8230 ;
  assign n8239 = n8229 & n8238 ;
  assign n8240 = n8239 ^ n8228 ;
  assign n8242 = n8241 ^ n8240 ;
  assign n8249 = ~n2646 & n5700 ;
  assign n8247 = ~n2738 & n20731 ;
  assign n8245 = ~n3227 & n5702 ;
  assign n8244 = n8241 ^ x17 ;
  assign n8246 = n8245 ^ n8244 ;
  assign n8248 = n8247 ^ n8246 ;
  assign n8250 = n8249 ^ n8248 ;
  assign n8243 = n5703 & n6900 ;
  assign n8251 = n8250 ^ n8243 ;
  assign n8252 = n8242 & n8251 ;
  assign n8253 = n8252 ^ n8241 ;
  assign n8255 = n8254 ^ n8253 ;
  assign n8262 = ~n2646 & n20731 ;
  assign n8260 = ~n2609 & n5702 ;
  assign n8258 = ~n3227 & n5700 ;
  assign n8257 = n8254 ^ x17 ;
  assign n8259 = n8258 ^ n8257 ;
  assign n8261 = n8260 ^ n8259 ;
  assign n8263 = n8262 ^ n8261 ;
  assign n8256 = n5703 & n7029 ;
  assign n8264 = n8263 ^ n8256 ;
  assign n8265 = n8255 & n8264 ;
  assign n8266 = n8265 ^ n8254 ;
  assign n8268 = n8267 ^ n8266 ;
  assign n8275 = ~n2609 & n5700 ;
  assign n8273 = ~n2554 & n5702 ;
  assign n8271 = ~n3227 & n20731 ;
  assign n8270 = n8267 ^ x17 ;
  assign n8272 = n8271 ^ n8270 ;
  assign n8274 = n8273 ^ n8272 ;
  assign n8276 = n8275 ^ n8274 ;
  assign n8269 = n5541 & n5703 ;
  assign n8277 = n8276 ^ n8269 ;
  assign n8278 = n8268 & n8277 ;
  assign n8279 = n8278 ^ n8267 ;
  assign n8281 = n8280 ^ n8279 ;
  assign n8288 = ~n2554 & n5700 ;
  assign n8286 = ~n2486 & n5702 ;
  assign n8284 = ~n2609 & n20731 ;
  assign n8283 = n8280 ^ x17 ;
  assign n8285 = n8284 ^ n8283 ;
  assign n8287 = n8286 ^ n8285 ;
  assign n8289 = n8288 ^ n8287 ;
  assign n8282 = n5381 & n5703 ;
  assign n8290 = n8289 ^ n8282 ;
  assign n8291 = n8281 & n8290 ;
  assign n8292 = n8291 ^ n8280 ;
  assign n8294 = n8293 ^ n8292 ;
  assign n8301 = ~n2486 & n5700 ;
  assign n8299 = ~n2554 & n20731 ;
  assign n8297 = ~n2449 & n5702 ;
  assign n8296 = n8293 ^ x17 ;
  assign n8298 = n8297 ^ n8296 ;
  assign n8300 = n8299 ^ n8298 ;
  assign n8302 = n8301 ^ n8300 ;
  assign n8295 = n5520 & n5703 ;
  assign n8303 = n8302 ^ n8295 ;
  assign n8304 = n8294 & n8303 ;
  assign n8305 = n8304 ^ n8293 ;
  assign n8307 = n8306 ^ n8305 ;
  assign n8314 = ~n2449 & n5700 ;
  assign n8312 = ~n2486 & n20731 ;
  assign n8310 = ~n2364 & n5702 ;
  assign n8309 = n8306 ^ x17 ;
  assign n8311 = n8310 ^ n8309 ;
  assign n8313 = n8312 ^ n8311 ;
  assign n8315 = n8314 ^ n8313 ;
  assign n8308 = n5283 & n5703 ;
  assign n8316 = n8315 ^ n8308 ;
  assign n8317 = n8307 & n8316 ;
  assign n8318 = n8317 ^ n8306 ;
  assign n8319 = n7900 ^ n7889 ;
  assign n8321 = ~n8318 & ~n8319 ;
  assign n8320 = n8319 ^ n8318 ;
  assign n8322 = n8321 ^ n8320 ;
  assign n8323 = n8321 ^ n8116 ;
  assign n8324 = n8123 ^ x17 ;
  assign n8325 = n8324 ^ n8321 ;
  assign n8326 = ~n8323 & n8325 ;
  assign n8327 = n8326 ^ n8116 ;
  assign n8328 = n8322 & n8327 ;
  assign n8329 = n8126 & n8328 ;
  assign n8330 = n8329 ^ n8327 ;
  assign n8332 = n8331 ^ n8330 ;
  assign n8339 = ~n2268 & n20731 ;
  assign n8337 = ~n2185 & n5700 ;
  assign n8335 = ~n2096 & n5702 ;
  assign n8334 = n8331 ^ x17 ;
  assign n8336 = n8335 ^ n8334 ;
  assign n8338 = n8337 ^ n8336 ;
  assign n8340 = n8339 ^ n8338 ;
  assign n8333 = n5196 & n5703 ;
  assign n8341 = n8340 ^ n8333 ;
  assign n8342 = n8332 & n8341 ;
  assign n8343 = n8342 ^ n8331 ;
  assign n8345 = n8344 ^ n8343 ;
  assign n8352 = ~n2096 & n5700 ;
  assign n8350 = ~n2185 & n20731 ;
  assign n8348 = ~n1994 & n5702 ;
  assign n8347 = n8344 ^ x17 ;
  assign n8349 = n8348 ^ n8347 ;
  assign n8351 = n8350 ^ n8349 ;
  assign n8353 = n8352 ^ n8351 ;
  assign n8346 = n5409 & n5703 ;
  assign n8354 = n8353 ^ n8346 ;
  assign n8355 = ~n8345 & ~n8354 ;
  assign n8356 = n8355 ^ n8344 ;
  assign n8357 = n8356 ^ n8101 ;
  assign n8358 = ~n8107 & n8357 ;
  assign n8359 = n8358 ^ n8101 ;
  assign n8361 = n8360 ^ n8359 ;
  assign n8368 = ~n1795 & n5700 ;
  assign n8366 = ~n1871 & n5702 ;
  assign n8364 = ~n1994 & n20731 ;
  assign n8363 = n8360 ^ x17 ;
  assign n8365 = n8364 ^ n8363 ;
  assign n8367 = n8366 ^ n8365 ;
  assign n8369 = n8368 ^ n8367 ;
  assign n8362 = ~n4859 & n5703 ;
  assign n8370 = n8369 ^ n8362 ;
  assign n8371 = ~n8361 & n8370 ;
  assign n8372 = n8371 ^ n8360 ;
  assign n8373 = n8372 ^ n8091 ;
  assign n8374 = n8097 & n8373 ;
  assign n8375 = n8374 ^ n8091 ;
  assign n8377 = n8376 ^ n8375 ;
  assign n8384 = ~n1871 & n20731 ;
  assign n8382 = ~n1631 & n5700 ;
  assign n8380 = ~n1703 & n5702 ;
  assign n8379 = n8376 ^ x17 ;
  assign n8381 = n8380 ^ n8379 ;
  assign n8383 = n8382 ^ n8381 ;
  assign n8385 = n8384 ^ n8383 ;
  assign n8378 = ~n4615 & n5703 ;
  assign n8386 = n8385 ^ n8378 ;
  assign n8387 = ~n8377 & ~n8386 ;
  assign n8388 = n8387 ^ n8376 ;
  assign n8389 = n8388 ^ n8084 ;
  assign n8390 = n8087 & ~n8389 ;
  assign n8391 = n8390 ^ n8084 ;
  assign n8392 = n8391 ^ n8065 ;
  assign n8393 = ~n8071 & ~n8392 ;
  assign n8394 = n8393 ^ n8065 ;
  assign n8060 = ~n317 & n7146 ;
  assign n8057 = ~n445 & n7141 ;
  assign n8054 = n7133 ^ x7 ;
  assign n8055 = ~n485 & n8054 ;
  assign n8051 = n8002 ^ n7719 ;
  assign n8052 = n8051 ^ x8 ;
  assign n8056 = n8055 ^ n8052 ;
  assign n8058 = n8057 ^ n8056 ;
  assign n8050 = n3500 & n7135 ;
  assign n8059 = n8058 ^ n8050 ;
  assign n8061 = n8060 ^ n8059 ;
  assign n10106 = n8394 ^ n8061 ;
  assign n10107 = n10106 ^ x5 ;
  assign n9077 = x3 ^ x2 ;
  assign n25052 = x5 & n9077 ;
  assign n9078 = x4 & n9077 ;
  assign n9081 = n25052 ^ n9078 ;
  assign n10103 = ~n3920 & n9081 ;
  assign n9088 = x4 ^ x3 ;
  assign n18627 = ~n9077 & ~n9088 ;
  assign n9089 = x5 ^ x4 ;
  assign n9090 = ~n9088 & ~n9089 ;
  assign n9091 = ~n9077 & n9090 ;
  assign n9092 = ~n18627 ^ n9091 ;
  assign n10104 = n10103 ^ n9092 ;
  assign n10105 = ~n3943 & ~n10104 ;
  assign n10108 = n10107 ^ n10105 ;
  assign n9073 = n4073 & n7135 ;
  assign n9071 = ~n445 & n8054 ;
  assign n9069 = ~n649 & n7146 ;
  assign n9067 = n8391 ^ n8071 ;
  assign n9068 = n9067 ^ x8 ;
  assign n9070 = n9069 ^ n9068 ;
  assign n9072 = n9071 ^ n9070 ;
  assign n9074 = n9073 ^ n9072 ;
  assign n9066 = ~n317 & n7141 ;
  assign n9075 = n9074 ^ n9066 ;
  assign n8409 = ~n968 & n6655 ;
  assign n8408 = ~n1109 & n6650 ;
  assign n8410 = n8409 ^ n8408 ;
  assign n8411 = n8410 ^ n6656 ;
  assign n8412 = n8411 ^ x11 ;
  assign n8413 = n8410 ^ x11 ;
  assign n8420 = n4044 & n8413 ;
  assign n8414 = n8413 ^ n6657 ;
  assign n8421 = n8420 ^ n8414 ;
  assign n8415 = n8414 ^ n824 ;
  assign n8416 = n8415 ^ x10 ;
  assign n8417 = n8416 ^ n8413 ;
  assign n8424 = n8417 ^ n8415 ;
  assign n8425 = n4044 & n8424 ;
  assign n8426 = n8425 ^ n8415 ;
  assign n8427 = ~n8414 & ~n8426 ;
  assign n8428 = ~n8421 & n8427 ;
  assign n8429 = n8428 ^ n8425 ;
  assign n8430 = n8429 ^ n6657 ;
  assign n8431 = n8430 ^ n8415 ;
  assign n8432 = ~n8412 & n8431 ;
  assign n8407 = n8388 ^ n8087 ;
  assign n8433 = n8432 ^ n8407 ;
  assign n8447 = ~x14 & ~n3817 ;
  assign n8444 = n1540 & n4897 ;
  assign n8448 = n8444 ^ n4897 ;
  assign n8453 = n8447 & n8448 ;
  assign n8450 = ~n1433 & ~n6074 ;
  assign n8449 = ~n1351 & ~n6072 ;
  assign n8451 = n8450 ^ n8449 ;
  assign n8454 = n8453 ^ n8451 ;
  assign n8445 = n8444 ^ n6060 ;
  assign n8446 = n8445 ^ n6057 ;
  assign n8455 = n8454 ^ n8446 ;
  assign n8442 = n8386 ^ n8375 ;
  assign n8443 = n8442 ^ x14 ;
  assign n8456 = n8455 ^ n8443 ;
  assign n8439 = n1540 & n6063 ;
  assign n8440 = n8439 ^ n6057 ;
  assign n8441 = ~n3817 & n8440 ;
  assign n8457 = n8456 ^ n8441 ;
  assign n8460 = ~n1703 & ~n6072 ;
  assign n8459 = ~n1351 & ~n6074 ;
  assign n8461 = n8460 ^ n8459 ;
  assign n8462 = n8461 ^ n6060 ;
  assign n8463 = n8462 ^ x14 ;
  assign n8472 = n8461 ^ x14 ;
  assign n8475 = ~x13 & ~n3815 ;
  assign n8476 = n8475 ^ n1433 ;
  assign n8477 = ~n8472 & n8476 ;
  assign n8478 = n8477 ^ n1433 ;
  assign n8464 = n4908 ^ x13 ;
  assign n8465 = n8464 ^ n6072 ;
  assign n8466 = n4152 ^ n3815 ;
  assign n8469 = ~n6063 & ~n8466 ;
  assign n8470 = n8469 ^ n4152 ;
  assign n8471 = n8465 & n8470 ;
  assign n8479 = n8478 ^ n8471 ;
  assign n8480 = ~n8463 & ~n8479 ;
  assign n8458 = n8372 ^ n8097 ;
  assign n8481 = n8480 ^ n8458 ;
  assign n9032 = n8370 ^ n8359 ;
  assign n9016 = n8356 ^ n8107 ;
  assign n8982 = n8354 ^ n8343 ;
  assign n8967 = n8341 ^ n8330 ;
  assign n8500 = n8319 ^ n8115 ;
  assign n8501 = ~n8320 & n8500 ;
  assign n8502 = n8501 ^ n8125 ;
  assign n8491 = ~n1795 & n4897 ;
  assign n8492 = n4384 & n8491 ;
  assign n8494 = ~n2096 & ~n6072 ;
  assign n8493 = ~n1994 & ~n6074 ;
  assign n8495 = n8494 ^ n8493 ;
  assign n8496 = x14 & ~n8495 ;
  assign n8497 = n8492 & n8496 ;
  assign n8498 = n8497 ^ n8495 ;
  assign n8499 = n8498 ^ x14 ;
  assign n8503 = n8502 ^ n8499 ;
  assign n8486 = ~x14 & ~n1795 ;
  assign n8482 = n4899 ^ n1795 ;
  assign n8487 = n8486 ^ n8482 ;
  assign n8488 = n4384 & ~n8487 ;
  assign n8489 = n8488 ^ n8482 ;
  assign n8490 = n4897 & ~n8489 ;
  assign n8504 = n8503 ^ n8490 ;
  assign n8930 = n8320 ^ n8115 ;
  assign n8897 = n8316 ^ n8305 ;
  assign n8868 = n8303 ^ n8292 ;
  assign n8519 = n8277 ^ n8266 ;
  assign n8509 = ~n2486 & ~n6072 ;
  assign n8508 = ~n2449 & ~n6074 ;
  assign n8510 = n8509 ^ n8508 ;
  assign n8518 = n8510 ^ x14 ;
  assign n8520 = n8519 ^ n8518 ;
  assign n8511 = n8510 ^ n2364 ;
  assign n8506 = n4899 ^ n2364 ;
  assign n8512 = n8511 ^ n8506 ;
  assign n8515 = n5282 & n8512 ;
  assign n8516 = n8515 ^ n8506 ;
  assign n8517 = n4897 & ~n8516 ;
  assign n8521 = n8520 ^ n8517 ;
  assign n8817 = n8264 ^ n8253 ;
  assign n8785 = n8251 ^ n8240 ;
  assign n17542 = n6063 ^ x13 ;
  assign n8528 = n4899 ^ n2554 ;
  assign n8523 = ~n2609 & ~n6074 ;
  assign n8522 = ~n3227 & ~n6072 ;
  assign n8524 = n8523 ^ n8522 ;
  assign n8529 = n8528 ^ n8524 ;
  assign n8531 = n17542 ^ n8529 ;
  assign n8532 = n8524 ^ n4899 ;
  assign n8533 = n17542 ^ n8532 ;
  assign n8534 = n8531 & ~n8533 ;
  assign n8535 = n17542 ^ n8534 ;
  assign n8536 = n5540 & ~n8535 ;
  assign n8537 = n8536 ^ n8528 ;
  assign n8538 = n4897 & ~n8537 ;
  assign n8526 = n8238 ^ n8227 ;
  assign n8525 = n8524 ^ x14 ;
  assign n8527 = n8526 ^ n8525 ;
  assign n8539 = n8538 ^ n8527 ;
  assign n8563 = n8221 ^ n8147 ;
  assign n8542 = ~n2738 & ~n6072 ;
  assign n8541 = ~n2646 & ~n6074 ;
  assign n8543 = n8542 ^ n8541 ;
  assign n8544 = n8543 ^ n6060 ;
  assign n8545 = n8544 ^ x14 ;
  assign n8558 = ~n3227 & n8465 ;
  assign n8557 = x13 & ~n6900 ;
  assign n8559 = n8558 ^ n8557 ;
  assign n8560 = ~n6063 & n8559 ;
  assign n8546 = n8543 ^ x14 ;
  assign n8553 = ~x13 & ~n6176 ;
  assign n8554 = n8553 ^ n3227 ;
  assign n8555 = ~n8546 & n8554 ;
  assign n8550 = n8465 ^ n6176 ;
  assign n8556 = n8555 ^ n8550 ;
  assign n8561 = n8560 ^ n8556 ;
  assign n8562 = ~n8545 & n8561 ;
  assign n8564 = n8563 ^ n8562 ;
  assign n8593 = n8219 ^ n8194 ;
  assign n8569 = ~n2646 & n6078 ;
  assign n8566 = ~n2738 & ~n6074 ;
  assign n8565 = ~n2836 & ~n6072 ;
  assign n8567 = n8566 ^ n8565 ;
  assign n8568 = n8567 ^ x14 ;
  assign n8570 = n8569 ^ n8568 ;
  assign n8574 = ~x13 & n5650 ;
  assign n8575 = n8574 ^ n2646 ;
  assign n8576 = n4897 & ~n8575 ;
  assign n8579 = n8576 ^ n8569 ;
  assign n8580 = n8579 ^ n8434 ;
  assign n8581 = n8580 ^ n8579 ;
  assign n8582 = n8579 ^ n5651 ;
  assign n8583 = n8582 ^ n8579 ;
  assign n8584 = n8581 & ~n8583 ;
  assign n8585 = n8584 ^ n8579 ;
  assign n8586 = ~n8570 & ~n8585 ;
  assign n8587 = n8586 ^ n8579 ;
  assign n8588 = n8587 ^ x14 ;
  assign n8589 = n8587 ^ n8570 ;
  assign n8590 = ~n8586 & ~n8589 ;
  assign n8591 = n8588 & n8590 ;
  assign n8592 = n8591 ^ n8587 ;
  assign n8594 = n8593 ^ n8592 ;
  assign n8598 = ~n2836 & ~n6074 ;
  assign n8597 = ~n3151 & ~n6072 ;
  assign n8599 = n8598 ^ n8597 ;
  assign n8609 = n8599 ^ x14 ;
  assign n8601 = n4899 ^ n2738 ;
  assign n8603 = n8601 ^ x13 ;
  assign n8604 = ~n2738 & ~n8603 ;
  assign n8605 = n8604 ^ n8601 ;
  assign n8606 = ~n3347 & ~n8605 ;
  assign n8607 = n8606 ^ n8601 ;
  assign n8608 = n4897 & ~n8607 ;
  assign n8610 = n8609 ^ n8608 ;
  assign n8596 = n3348 & n6060 ;
  assign n8611 = n8610 ^ n8596 ;
  assign n8595 = n8191 ^ n8160 ;
  assign n8612 = n8611 ^ n8595 ;
  assign n8641 = n8180 ^ n8161 ;
  assign n8642 = n8641 ^ n8189 ;
  assign n8617 = ~n2836 & n7603 ;
  assign n8614 = ~n3151 & ~n6074 ;
  assign n8613 = ~n2924 & ~n6072 ;
  assign n8615 = n8614 ^ n8613 ;
  assign n8616 = n8615 ^ x14 ;
  assign n8618 = n8617 ^ n8616 ;
  assign n8622 = x13 & ~n3345 ;
  assign n8623 = n8622 ^ n2836 ;
  assign n8624 = n4897 & ~n8623 ;
  assign n8627 = n8624 ^ n8617 ;
  assign n8628 = n8627 ^ n6057 ;
  assign n8629 = n8628 ^ n8627 ;
  assign n8630 = n8627 ^ n6237 ;
  assign n8631 = n8630 ^ n8627 ;
  assign n8632 = n8629 & n8631 ;
  assign n8633 = n8632 ^ n8627 ;
  assign n8634 = n8618 & ~n8633 ;
  assign n8635 = n8634 ^ n8627 ;
  assign n8636 = n8635 ^ x14 ;
  assign n8637 = n8635 ^ n8618 ;
  assign n8638 = ~n8634 & n8637 ;
  assign n8639 = ~n8636 & n8638 ;
  assign n8640 = n8639 ^ n8635 ;
  assign n8643 = n8642 ^ n8640 ;
  assign n8167 = n8166 ^ x17 ;
  assign n8673 = n8179 ^ n8167 ;
  assign n8648 = ~n3151 & n7603 ;
  assign n8645 = ~n2958 & ~n6072 ;
  assign n8644 = ~n2924 & ~n6074 ;
  assign n8646 = n8645 ^ n8644 ;
  assign n8647 = n8646 ^ x14 ;
  assign n8649 = n8648 ^ n8647 ;
  assign n8654 = x13 & ~n6282 ;
  assign n8655 = n8654 ^ n3151 ;
  assign n8656 = n4897 & ~n8655 ;
  assign n8659 = n8656 ^ n8648 ;
  assign n8660 = n8659 ^ n6057 ;
  assign n8661 = n8660 ^ n8659 ;
  assign n8662 = n8659 ^ n6286 ;
  assign n8663 = n8662 ^ n8659 ;
  assign n8664 = n8661 & n8663 ;
  assign n8665 = n8664 ^ n8659 ;
  assign n8666 = n8649 & ~n8665 ;
  assign n8667 = n8666 ^ n8659 ;
  assign n8668 = n8667 ^ x14 ;
  assign n8669 = n8667 ^ n8649 ;
  assign n8670 = ~n8666 & n8669 ;
  assign n8671 = ~n8668 & n8670 ;
  assign n8672 = n8671 ^ n8667 ;
  assign n8674 = n8673 ^ n8672 ;
  assign n5698 = n5697 ^ x16 ;
  assign n8726 = ~n3337 & n5698 ;
  assign n8727 = n8726 ^ n8162 ;
  assign n8679 = ~n2958 & n6078 ;
  assign n8676 = ~n3027 & ~n6072 ;
  assign n8675 = ~n3099 & ~n6074 ;
  assign n8677 = n8676 ^ n8675 ;
  assign n8678 = n8677 ^ x14 ;
  assign n8680 = n8679 ^ n8678 ;
  assign n8694 = n6440 & n8434 ;
  assign n8684 = ~x13 & ~n6439 ;
  assign n8685 = n8684 ^ n2958 ;
  assign n8686 = n4897 & ~n8685 ;
  assign n8689 = n8686 ^ n8679 ;
  assign n8695 = n8694 ^ n8689 ;
  assign n8696 = ~n8680 & ~n8695 ;
  assign n8697 = n8696 ^ n8689 ;
  assign n8698 = n8697 ^ x14 ;
  assign n8699 = n8697 ^ n8680 ;
  assign n8700 = ~n8696 & ~n8699 ;
  assign n8701 = n8698 & n8700 ;
  assign n8702 = n8701 ^ n8697 ;
  assign n8703 = ~n3337 & n5693 ;
  assign n8704 = n4897 ^ n3337 ;
  assign n8706 = ~n3027 & n4897 ;
  assign n8705 = n15382 ^ n3337 ;
  assign n8707 = n8706 ^ n8705 ;
  assign n8708 = n8707 ^ n3337 ;
  assign n8709 = ~n8704 & n8708 ;
  assign n8710 = n8709 ^ n3337 ;
  assign n8711 = x14 & ~n8710 ;
  assign n8712 = n8711 ^ x14 ;
  assign n8719 = ~n3027 & ~n6074 ;
  assign n8718 = ~n3337 & ~n6072 ;
  assign n8720 = n8719 ^ n8718 ;
  assign n8715 = n3339 & n4899 ;
  assign n8716 = n8715 ^ n3099 ;
  assign n8717 = n4897 & ~n8716 ;
  assign n8721 = n8720 ^ n8717 ;
  assign n8722 = n8712 & ~n8721 ;
  assign n8723 = ~n8703 & ~n8722 ;
  assign n8724 = ~n8702 & n8723 ;
  assign n8725 = n8724 ^ n8702 ;
  assign n8728 = n8727 ^ n8725 ;
  assign n8741 = ~n2958 & ~n6074 ;
  assign n8740 = ~n3099 & ~n6072 ;
  assign n8742 = n8741 ^ n8740 ;
  assign n8735 = ~x14 & ~n2924 ;
  assign n8731 = n4899 ^ n2924 ;
  assign n8736 = n8735 ^ n8731 ;
  assign n8737 = n6343 & ~n8736 ;
  assign n8738 = n8737 ^ n8731 ;
  assign n8739 = n4897 & ~n8738 ;
  assign n8743 = n8742 ^ n8739 ;
  assign n8747 = n8743 ^ x14 ;
  assign n8729 = ~n2924 & n4897 ;
  assign n8730 = n6344 & n8729 ;
  assign n8745 = x14 & ~n8742 ;
  assign n8746 = n8730 & n8745 ;
  assign n8748 = n8747 ^ n8746 ;
  assign n8749 = n8748 ^ n8725 ;
  assign n8750 = ~n8728 & n8749 ;
  assign n8751 = n8750 ^ n8727 ;
  assign n8752 = n8751 ^ n8672 ;
  assign n8753 = n8674 & ~n8752 ;
  assign n8754 = n8753 ^ n8673 ;
  assign n8755 = n8754 ^ n8640 ;
  assign n8756 = ~n8643 & n8755 ;
  assign n8757 = n8756 ^ n8754 ;
  assign n8758 = n8757 ^ n8611 ;
  assign n8759 = n8612 & n8758 ;
  assign n8760 = n8759 ^ n8611 ;
  assign n8761 = n8760 ^ n8592 ;
  assign n8762 = ~n8594 & ~n8761 ;
  assign n8763 = n8762 ^ n8760 ;
  assign n8764 = n8763 ^ n8563 ;
  assign n8765 = ~n8564 & n8764 ;
  assign n8766 = n8765 ^ n8563 ;
  assign n8540 = n8224 ^ n8136 ;
  assign n8767 = n8766 ^ n8540 ;
  assign n8777 = ~n2646 & ~n6072 ;
  assign n8775 = ~n3227 & ~n6074 ;
  assign n8774 = n8540 ^ x14 ;
  assign n8776 = n8775 ^ n8774 ;
  assign n8778 = n8777 ^ n8776 ;
  assign n8768 = n7029 ^ n2609 ;
  assign n8771 = n4899 & ~n8768 ;
  assign n8772 = n8771 ^ n2609 ;
  assign n8773 = n4897 & ~n8772 ;
  assign n8779 = n8778 ^ n8773 ;
  assign n8780 = n8767 & ~n8779 ;
  assign n8781 = n8780 ^ n8766 ;
  assign n8782 = n8781 ^ n8526 ;
  assign n8783 = n8539 & n8782 ;
  assign n8784 = n8783 ^ n8526 ;
  assign n8786 = n8785 ^ n8784 ;
  assign n8791 = ~n2486 & n7603 ;
  assign n8788 = ~n2554 & ~n6074 ;
  assign n8787 = ~n2609 & ~n6072 ;
  assign n8789 = n8788 ^ n8787 ;
  assign n8790 = n8789 ^ x14 ;
  assign n8792 = n8791 ^ n8790 ;
  assign n8793 = n8792 ^ x14 ;
  assign n8796 = x13 & ~n5380 ;
  assign n8797 = n8796 ^ n2486 ;
  assign n8798 = n4897 & ~n8797 ;
  assign n8800 = n8798 ^ n8791 ;
  assign n8801 = n8800 ^ n6057 ;
  assign n8802 = n8801 ^ n8800 ;
  assign n8803 = n8800 ^ n5381 ;
  assign n8804 = n8803 ^ n8800 ;
  assign n8805 = n8802 & n8804 ;
  assign n8806 = n8805 ^ n8800 ;
  assign n8807 = n8792 & ~n8806 ;
  assign n8808 = n8793 & ~n8807 ;
  assign n8809 = n8800 ^ n8785 ;
  assign n8810 = n8809 ^ n8807 ;
  assign n8811 = n8810 ^ x14 ;
  assign n8812 = n8811 ^ n8785 ;
  assign n8813 = n8808 & ~n8812 ;
  assign n8814 = n8813 ^ n8810 ;
  assign n8815 = n8786 & n8814 ;
  assign n8816 = n8815 ^ n8785 ;
  assign n8818 = n8817 ^ n8816 ;
  assign n8823 = ~n2449 & n6078 ;
  assign n8820 = ~n2554 & ~n6072 ;
  assign n8819 = ~n2486 & ~n6074 ;
  assign n8821 = n8820 ^ n8819 ;
  assign n8822 = n8821 ^ x14 ;
  assign n8824 = n8823 ^ n8822 ;
  assign n8825 = n8824 ^ x14 ;
  assign n8829 = ~x13 & ~n5519 ;
  assign n8830 = n8829 ^ n2449 ;
  assign n8831 = n4897 & ~n8830 ;
  assign n8833 = n8831 ^ n8823 ;
  assign n8834 = n8833 ^ n8434 ;
  assign n8835 = n8834 ^ n8833 ;
  assign n8836 = n8833 ^ n5520 ;
  assign n8837 = n8836 ^ n8833 ;
  assign n8838 = n8835 & n8837 ;
  assign n8839 = n8838 ^ n8833 ;
  assign n8840 = ~n8824 & ~n8839 ;
  assign n8841 = n8825 & ~n8840 ;
  assign n8842 = n8833 ^ n8817 ;
  assign n8843 = n8842 ^ n8840 ;
  assign n8844 = n8843 ^ x14 ;
  assign n8845 = n8844 ^ n8817 ;
  assign n8846 = n8841 & n8845 ;
  assign n8847 = n8846 ^ n8843 ;
  assign n8848 = n8818 & ~n8847 ;
  assign n8849 = n8848 ^ n8817 ;
  assign n8850 = n8849 ^ n8519 ;
  assign n8851 = n8521 & n8850 ;
  assign n8852 = n8851 ^ n8519 ;
  assign n8505 = n8290 ^ n8279 ;
  assign n8853 = n8852 ^ n8505 ;
  assign n8863 = ~n2364 & ~n6074 ;
  assign n8861 = ~n2449 & ~n6072 ;
  assign n8860 = n8505 ^ x14 ;
  assign n8862 = n8861 ^ n8860 ;
  assign n8864 = n8863 ^ n8862 ;
  assign n8855 = n5144 ^ n4899 ;
  assign n8856 = n8855 ^ n5144 ;
  assign n8857 = ~n5143 & ~n8856 ;
  assign n8858 = n8857 ^ n5144 ;
  assign n8859 = n4897 & n8858 ;
  assign n8865 = n8864 ^ n8859 ;
  assign n8866 = n8853 & ~n8865 ;
  assign n8867 = n8866 ^ n8852 ;
  assign n8869 = n8868 ^ n8867 ;
  assign n8870 = n5195 ^ n3234 ;
  assign n8871 = x14 & ~n8870 ;
  assign n8883 = ~n2268 & ~n6074 ;
  assign n8882 = ~n2364 & ~n6072 ;
  assign n8884 = n8883 ^ n8882 ;
  assign n8891 = n8884 ^ n8868 ;
  assign n8880 = ~n2185 & n4897 ;
  assign n8881 = n4930 & n8880 ;
  assign n8885 = ~x14 & ~n8884 ;
  assign n8886 = n8881 & n8885 ;
  assign n8887 = n8886 ^ n8884 ;
  assign n8888 = n8887 ^ x14 ;
  assign n8889 = n8888 ^ n8868 ;
  assign n8872 = n2185 ^ x14 ;
  assign n8873 = n8872 ^ x13 ;
  assign n8874 = n8873 ^ x14 ;
  assign n8877 = ~n4930 & ~n8874 ;
  assign n8878 = n8877 ^ x14 ;
  assign n8879 = n4897 & n8878 ;
  assign n8890 = n8889 ^ n8879 ;
  assign n8892 = n8891 ^ n8890 ;
  assign n8893 = n8871 & ~n8892 ;
  assign n8894 = n8893 ^ n8890 ;
  assign n8895 = n8869 & n8894 ;
  assign n8896 = n8895 ^ n8868 ;
  assign n8898 = n8897 ^ n8896 ;
  assign n8903 = ~n2096 & n7603 ;
  assign n8900 = ~n2268 & ~n6072 ;
  assign n8899 = ~n2185 & ~n6074 ;
  assign n8901 = n8900 ^ n8899 ;
  assign n8902 = n8901 ^ x14 ;
  assign n8904 = n8903 ^ n8902 ;
  assign n8905 = n8904 ^ x14 ;
  assign n8909 = x13 & ~n5195 ;
  assign n8910 = n8909 ^ n2096 ;
  assign n8911 = n4897 & ~n8910 ;
  assign n8913 = n8911 ^ n8903 ;
  assign n8914 = n8913 ^ n6057 ;
  assign n8915 = n8914 ^ n8913 ;
  assign n8916 = n8913 ^ n5196 ;
  assign n8917 = n8916 ^ n8913 ;
  assign n8918 = n8915 & n8917 ;
  assign n8919 = n8918 ^ n8913 ;
  assign n8920 = n8904 & ~n8919 ;
  assign n8921 = n8905 & ~n8920 ;
  assign n8922 = n8913 ^ n8897 ;
  assign n8923 = n8922 ^ n8920 ;
  assign n8924 = n8923 ^ x14 ;
  assign n8925 = n8924 ^ n8897 ;
  assign n8926 = n8921 & ~n8925 ;
  assign n8927 = n8926 ^ n8923 ;
  assign n8928 = n8898 & n8927 ;
  assign n8929 = n8928 ^ n8897 ;
  assign n8931 = n8930 ^ n8929 ;
  assign n8936 = ~n1994 & n7603 ;
  assign n8933 = ~n2185 & ~n6072 ;
  assign n8932 = ~n2096 & ~n6074 ;
  assign n8934 = n8933 ^ n8932 ;
  assign n8935 = n8934 ^ x14 ;
  assign n8937 = n8936 ^ n8935 ;
  assign n8938 = n8937 ^ x14 ;
  assign n8943 = x13 & ~n5408 ;
  assign n8944 = n8943 ^ n1994 ;
  assign n8945 = n4897 & ~n8944 ;
  assign n8947 = n8945 ^ n8936 ;
  assign n8948 = n8947 ^ n6057 ;
  assign n8949 = n8948 ^ n8947 ;
  assign n8950 = n8947 ^ n5409 ;
  assign n8951 = n8950 ^ n8947 ;
  assign n8952 = n8949 & n8951 ;
  assign n8953 = n8952 ^ n8947 ;
  assign n8954 = n8937 & ~n8953 ;
  assign n8955 = n8938 & ~n8954 ;
  assign n8956 = n8947 ^ n8930 ;
  assign n8957 = n8956 ^ n8954 ;
  assign n8958 = n8957 ^ x14 ;
  assign n8959 = n8958 ^ n8930 ;
  assign n8960 = n8955 & ~n8959 ;
  assign n8961 = n8960 ^ n8957 ;
  assign n8962 = n8931 & n8961 ;
  assign n8963 = n8962 ^ n8930 ;
  assign n8964 = n8963 ^ n8502 ;
  assign n8965 = n8504 & n8964 ;
  assign n8966 = n8965 ^ n8502 ;
  assign n8968 = n8967 ^ n8966 ;
  assign n8977 = ~n1795 & ~n6074 ;
  assign n8975 = ~n1994 & ~n6072 ;
  assign n8974 = n8967 ^ x14 ;
  assign n8976 = n8975 ^ n8974 ;
  assign n8978 = n8977 ^ n8976 ;
  assign n8971 = ~n4899 & n5184 ;
  assign n8972 = n8971 ^ n4859 ;
  assign n8973 = n4897 & ~n8972 ;
  assign n8979 = n8978 ^ n8973 ;
  assign n8980 = n8968 & n8979 ;
  assign n8981 = n8980 ^ n8967 ;
  assign n8983 = n8982 ^ n8981 ;
  assign n8988 = ~n1631 & n6078 ;
  assign n8985 = ~n1871 & ~n6074 ;
  assign n8984 = ~n1795 & ~n6072 ;
  assign n8986 = n8985 ^ n8984 ;
  assign n8987 = n8986 ^ x14 ;
  assign n8989 = n8988 ^ n8987 ;
  assign n8990 = n8989 ^ x14 ;
  assign n8995 = ~x13 & n4391 ;
  assign n8996 = n8995 ^ n1631 ;
  assign n8997 = n4897 & ~n8996 ;
  assign n8999 = n8997 ^ n8988 ;
  assign n9000 = n8999 ^ n8434 ;
  assign n9001 = n9000 ^ n8999 ;
  assign n9002 = n8999 ^ n4392 ;
  assign n9003 = n9002 ^ n8999 ;
  assign n9004 = n9001 & ~n9003 ;
  assign n9005 = n9004 ^ n8999 ;
  assign n9006 = ~n8989 & ~n9005 ;
  assign n9007 = n8990 & ~n9006 ;
  assign n9008 = n8999 ^ n8982 ;
  assign n9009 = n9008 ^ n9006 ;
  assign n9010 = n9009 ^ x14 ;
  assign n9011 = n9010 ^ n8982 ;
  assign n9012 = n9007 & n9011 ;
  assign n9013 = n9012 ^ n9009 ;
  assign n9014 = ~n8983 & n9013 ;
  assign n9015 = n9014 ^ n8982 ;
  assign n9017 = n9016 ^ n9015 ;
  assign n9026 = n9016 ^ x14 ;
  assign n9025 = ~n1631 & ~n6074 ;
  assign n9027 = n9026 ^ n9025 ;
  assign n9024 = ~n1871 & ~n6072 ;
  assign n9028 = n9027 ^ n9024 ;
  assign n9021 = n3808 & ~n4899 ;
  assign n9022 = n9021 ^ n4615 ;
  assign n9023 = n4897 & ~n9022 ;
  assign n9029 = n9028 ^ n9023 ;
  assign n9030 = ~n9017 & n9029 ;
  assign n9031 = n9030 ^ n9016 ;
  assign n9033 = n9032 ^ n9031 ;
  assign n9039 = n4417 ^ x13 ;
  assign n9040 = n9039 ^ n4417 ;
  assign n9041 = ~n4416 & n9040 ;
  assign n9042 = n9041 ^ n4417 ;
  assign n9043 = n6060 & n9042 ;
  assign n9035 = ~n1631 & ~n6072 ;
  assign n9034 = ~n1703 & ~n6074 ;
  assign n9036 = n9035 ^ n9034 ;
  assign n9037 = n9036 ^ x14 ;
  assign n9044 = n9043 ^ n9037 ;
  assign n9053 = n9044 ^ n9032 ;
  assign n9047 = x13 & ~n4416 ;
  assign n9048 = n9047 ^ n1351 ;
  assign n9049 = n4897 & ~n9048 ;
  assign n9050 = n9049 ^ n9036 ;
  assign n9051 = ~x14 & n9050 ;
  assign n9052 = ~n9044 & n9051 ;
  assign n9054 = n9053 ^ n9052 ;
  assign n9055 = ~n9033 & ~n9054 ;
  assign n9056 = n9055 ^ n9032 ;
  assign n9057 = n9056 ^ n8458 ;
  assign n9058 = ~n8481 & ~n9057 ;
  assign n9059 = n9058 ^ n8458 ;
  assign n9060 = n9059 ^ n8442 ;
  assign n9061 = ~n8457 & ~n9060 ;
  assign n9062 = n9061 ^ n8442 ;
  assign n9063 = n9062 ^ n8407 ;
  assign n9064 = n8433 & n9063 ;
  assign n9065 = n9064 ^ n8407 ;
  assign n10096 = n9067 ^ n9065 ;
  assign n10097 = ~n9075 & n10096 ;
  assign n10098 = n10097 ^ n9067 ;
  assign n11516 = n10106 ^ n10098 ;
  assign n11517 = n10108 & ~n11516 ;
  assign n11518 = n11517 ^ n10106 ;
  assign n11520 = n11519 ^ n11518 ;
  assign n9076 = n9075 ^ n9065 ;
  assign n9573 = ~n3943 & n9077 ;
  assign n9566 = n3956 & n7135 ;
  assign n9562 = n9062 ^ n8433 ;
  assign n9563 = n9562 ^ x8 ;
  assign n9561 = ~n3473 & n7146 ;
  assign n9564 = n9563 ^ n9561 ;
  assign n9560 = ~n317 & n8054 ;
  assign n9565 = n9564 ^ n9560 ;
  assign n9567 = n9566 ^ n9565 ;
  assign n9559 = ~n649 & n7141 ;
  assign n9568 = n9567 ^ n9559 ;
  assign n9101 = ~n1109 & n6658 ;
  assign n9097 = n9059 ^ n8457 ;
  assign n9098 = n9097 ^ x11 ;
  assign n9096 = ~n1214 & n6655 ;
  assign n9099 = n9098 ^ n9096 ;
  assign n9095 = ~n968 & n6650 ;
  assign n9100 = n9099 ^ n9095 ;
  assign n9102 = n9101 ^ n9100 ;
  assign n9094 = n3905 & n15413 ;
  assign n9103 = n9102 ^ n9094 ;
  assign n9111 = ~n1540 & n6655 ;
  assign n9107 = n9056 ^ n8481 ;
  assign n9108 = n9107 ^ x11 ;
  assign n9106 = ~n1214 & n6650 ;
  assign n9109 = n9108 ^ n9106 ;
  assign n9105 = ~n968 & n6658 ;
  assign n9110 = n9109 ^ n9105 ;
  assign n9112 = n9111 ^ n9110 ;
  assign n9104 = n3521 & n15413 ;
  assign n9113 = n9112 ^ n9104 ;
  assign n9540 = n9054 ^ n9031 ;
  assign n9121 = ~n1351 & n6655 ;
  assign n9117 = n9029 ^ n9015 ;
  assign n9118 = n9117 ^ x11 ;
  assign n9116 = ~n1540 & n6658 ;
  assign n9119 = n9118 ^ n9116 ;
  assign n9115 = ~n1433 & n6650 ;
  assign n9120 = n9119 ^ n9115 ;
  assign n9122 = n9121 ^ n9120 ;
  assign n9114 = ~n4610 & n15413 ;
  assign n9123 = n9122 ^ n9114 ;
  assign n9524 = n9013 ^ n8981 ;
  assign n9511 = n8979 ^ n8966 ;
  assign n9131 = ~n1871 & n6655 ;
  assign n9127 = n8963 ^ n8504 ;
  assign n9128 = n9127 ^ x11 ;
  assign n9126 = ~n1703 & n6658 ;
  assign n9129 = n9128 ^ n9126 ;
  assign n9125 = ~n1631 & n6650 ;
  assign n9130 = n9129 ^ n9125 ;
  assign n9132 = n9131 ^ n9130 ;
  assign n9124 = ~n4615 & n15413 ;
  assign n9133 = n9132 ^ n9124 ;
  assign n9141 = ~n1795 & n6655 ;
  assign n9137 = n8961 ^ n8929 ;
  assign n9138 = n9137 ^ x11 ;
  assign n9136 = ~n1871 & n6650 ;
  assign n9139 = n9138 ^ n9136 ;
  assign n9135 = ~n1631 & n6658 ;
  assign n9140 = n9139 ^ n9135 ;
  assign n9142 = n9141 ^ n9140 ;
  assign n9134 = ~n4392 & n15413 ;
  assign n9143 = n9142 ^ n9134 ;
  assign n9151 = ~n1871 & n6658 ;
  assign n9147 = n8927 ^ n8896 ;
  assign n9148 = n9147 ^ x11 ;
  assign n9146 = ~n1795 & n6650 ;
  assign n9149 = n9148 ^ n9146 ;
  assign n9145 = ~n1994 & n6655 ;
  assign n9150 = n9149 ^ n9145 ;
  assign n9152 = n9151 ^ n9150 ;
  assign n9144 = ~n4859 & n15413 ;
  assign n9153 = n9152 ^ n9144 ;
  assign n9489 = n8894 ^ n8867 ;
  assign n9162 = n8865 ^ n8852 ;
  assign n9163 = n9162 ^ x11 ;
  assign n9161 = ~n2185 & n6655 ;
  assign n9164 = n9163 ^ n9161 ;
  assign n9160 = ~n2096 & n6650 ;
  assign n9165 = n9164 ^ n9160 ;
  assign n9155 = n9154 ^ n5409 ;
  assign n9156 = n9155 ^ n5409 ;
  assign n9157 = ~n5408 & ~n9156 ;
  assign n9158 = n9157 ^ n5409 ;
  assign n9159 = n6648 & n9158 ;
  assign n9166 = n9165 ^ n9159 ;
  assign n9473 = n8849 ^ n8521 ;
  assign n9447 = n8781 ^ n8539 ;
  assign n9197 = n8779 ^ n8766 ;
  assign n9192 = ~n2554 & n6655 ;
  assign n9191 = ~n2449 & n6658 ;
  assign n9193 = n9192 ^ n9191 ;
  assign n9194 = n9193 ^ x11 ;
  assign n9190 = ~n2486 & n6650 ;
  assign n9195 = n9194 ^ n9190 ;
  assign n9189 = n5520 & n15413 ;
  assign n9196 = n9195 ^ n9189 ;
  assign n9198 = n9197 ^ n9196 ;
  assign n9431 = n8763 ^ n8564 ;
  assign n9443 = n9431 ^ n9196 ;
  assign n9416 = n8760 ^ n8594 ;
  assign n9203 = ~n2738 & n6655 ;
  assign n9201 = ~n3227 & n6658 ;
  assign n9200 = ~n2646 & n6650 ;
  assign n9202 = n9201 ^ n9200 ;
  assign n9204 = n9203 ^ n9202 ;
  assign n9199 = n6900 & n15413 ;
  assign n9205 = n9204 ^ n9199 ;
  assign n9206 = n9205 ^ x11 ;
  assign n9216 = ~n3227 & n6650 ;
  assign n9215 = ~n2646 & n6655 ;
  assign n9217 = n9216 ^ n9215 ;
  assign n9212 = ~n8768 & n9154 ;
  assign n9213 = n9212 ^ n2609 ;
  assign n9214 = n6648 & ~n9213 ;
  assign n9218 = n9217 ^ n9214 ;
  assign n9219 = n9218 ^ n9205 ;
  assign n9207 = n8757 ^ n8612 ;
  assign n9220 = n9219 ^ n9207 ;
  assign n9221 = n9206 & ~n9220 ;
  assign n9238 = n8749 ^ n8727 ;
  assign n9233 = ~n2738 & n6658 ;
  assign n9232 = ~n2836 & n6650 ;
  assign n9234 = n9233 ^ n9232 ;
  assign n9235 = n9234 ^ x11 ;
  assign n9231 = ~n3151 & n6655 ;
  assign n9236 = n9235 ^ n9231 ;
  assign n9230 = ~n6907 & n15413 ;
  assign n9237 = n9236 ^ n9230 ;
  assign n9239 = n9238 ^ n9237 ;
  assign n9248 = ~n3151 & n6650 ;
  assign n9243 = n8722 ^ n8703 ;
  assign n9244 = n9243 ^ n8702 ;
  assign n9245 = n9244 ^ x11 ;
  assign n9242 = ~n2924 & n6655 ;
  assign n9246 = n9245 ^ n9242 ;
  assign n9241 = ~n2836 & n6658 ;
  assign n9247 = n9246 ^ n9241 ;
  assign n9249 = n9248 ^ n9247 ;
  assign n9240 = n6237 & n15413 ;
  assign n9250 = n9249 ^ n9240 ;
  assign n9259 = n8721 ^ n8711 ;
  assign n9254 = ~n2958 & n6655 ;
  assign n9253 = ~n3151 & n6658 ;
  assign n9255 = n9254 ^ n9253 ;
  assign n9256 = n9255 ^ x11 ;
  assign n9252 = ~n2924 & n6650 ;
  assign n9257 = n9256 ^ n9252 ;
  assign n9251 = n6286 & n15413 ;
  assign n9258 = n9257 ^ n9251 ;
  assign n9260 = n9259 ^ n9258 ;
  assign n9379 = ~n3099 & n6655 ;
  assign n9378 = ~n2924 & n6658 ;
  assign n9380 = n9379 ^ n9378 ;
  assign n9381 = n9380 ^ x11 ;
  assign n9377 = ~n2958 & n6650 ;
  assign n9382 = n9381 ^ n9377 ;
  assign n9376 = n6344 & n15413 ;
  assign n9383 = n9382 ^ n9376 ;
  assign n9302 = n3337 ^ x11 ;
  assign n9268 = ~n3027 & n6648 ;
  assign n9269 = x11 & ~n16289 ;
  assign n9270 = n3337 & n9269 ;
  assign n9271 = ~n9268 & n9270 ;
  assign n9272 = n9271 ^ n9269 ;
  assign n9273 = n9272 ^ x11 ;
  assign n9282 = ~n3099 & n6648 ;
  assign n9281 = ~n3337 & n6655 ;
  assign n9283 = n9282 ^ n9281 ;
  assign n9278 = n3337 & n15413 ;
  assign n9279 = n9278 ^ n6650 ;
  assign n9280 = ~n3027 & n9279 ;
  assign n9284 = n9283 ^ n9280 ;
  assign n9285 = n9273 & ~n9284 ;
  assign n9265 = ~n2958 & n6658 ;
  assign n9263 = ~n3027 & n6655 ;
  assign n9262 = ~n3099 & n6650 ;
  assign n9264 = n9263 ^ n9262 ;
  assign n9266 = n9265 ^ n9264 ;
  assign n9261 = n6440 & n15413 ;
  assign n9267 = n9266 ^ n9261 ;
  assign n9286 = n9285 ^ n9267 ;
  assign n9287 = n9286 ^ x12 ;
  assign n9303 = n9302 ^ n9287 ;
  assign n9337 = n9303 ^ n9267 ;
  assign n9288 = n9287 ^ n3337 ;
  assign n9289 = n9288 ^ n9286 ;
  assign n9365 = n9337 ^ n9289 ;
  assign n9366 = n9365 ^ x12 ;
  assign n9367 = n9366 ^ n9267 ;
  assign n9319 = n9267 & ~n9286 ;
  assign n9320 = n9319 ^ n9288 ;
  assign n9304 = n9303 ^ n9289 ;
  assign n9321 = n9320 ^ n9304 ;
  assign n9322 = n9321 ^ n9285 ;
  assign n9323 = n9304 ^ n3337 ;
  assign n9324 = n9323 ^ n9285 ;
  assign n9325 = n9322 & n9324 ;
  assign n9301 = n9288 ^ n9267 ;
  assign n9308 = n9301 ^ n9287 ;
  assign n9310 = n9308 ^ n9304 ;
  assign n9326 = n9310 ^ n9287 ;
  assign n9327 = n9326 ^ n9302 ;
  assign n9328 = n9310 ^ n9288 ;
  assign n9329 = n9328 ^ n9302 ;
  assign n9330 = ~n9327 & ~n9329 ;
  assign n9331 = n9325 & n9330 ;
  assign n9332 = n9331 ^ n9319 ;
  assign n9333 = n9332 ^ n3337 ;
  assign n9372 = n9367 ^ n9333 ;
  assign n9293 = n9288 ^ x11 ;
  assign n9295 = n9293 ^ x12 ;
  assign n9297 = n9295 ^ n9267 ;
  assign n9298 = n9297 ^ n9293 ;
  assign n9373 = n9372 ^ n9298 ;
  assign n9374 = n9373 ^ n9285 ;
  assign n9375 = n9374 ^ n9297 ;
  assign n9384 = n9383 ^ n9375 ;
  assign n6056 = n4898 ^ x13 ;
  assign n9386 = ~n3337 & ~n6056 ;
  assign n9385 = n9383 ^ n8706 ;
  assign n9387 = n9386 ^ n9385 ;
  assign n9388 = n9384 & n9387 ;
  assign n9389 = n9388 ^ n9383 ;
  assign n9390 = n9389 ^ n9258 ;
  assign n9391 = n9260 & n9390 ;
  assign n9392 = n9391 ^ n9258 ;
  assign n9393 = n9392 ^ n9244 ;
  assign n9394 = ~n9250 & ~n9393 ;
  assign n9395 = n9394 ^ n9244 ;
  assign n9396 = n9395 ^ n9237 ;
  assign n9397 = ~n9239 & ~n9396 ;
  assign n9398 = n9397 ^ n9237 ;
  assign n9225 = ~n2836 & n6655 ;
  assign n9224 = ~n2646 & n6658 ;
  assign n9226 = n9225 ^ n9224 ;
  assign n9227 = n9226 ^ x11 ;
  assign n9223 = ~n2738 & n6650 ;
  assign n9228 = n9227 ^ n9223 ;
  assign n9222 = ~n5651 & n15413 ;
  assign n9229 = n9228 ^ n9222 ;
  assign n9399 = n9398 ^ n9229 ;
  assign n9400 = n9229 ^ n8674 ;
  assign n9401 = n9400 ^ n8751 ;
  assign n9402 = n9399 & ~n9401 ;
  assign n9403 = n9402 ^ n9398 ;
  assign n9404 = n8754 ^ n8643 ;
  assign n9406 = n9403 & n9404 ;
  assign n9405 = n9404 ^ n9403 ;
  assign n9407 = n9406 ^ n9405 ;
  assign n9408 = n9406 ^ n9207 ;
  assign n9409 = n9218 ^ x11 ;
  assign n9410 = n9409 ^ n9406 ;
  assign n9411 = n9408 & ~n9410 ;
  assign n9412 = n9411 ^ n9207 ;
  assign n9413 = n9407 & ~n9412 ;
  assign n9414 = n9221 & n9413 ;
  assign n9415 = n9414 ^ n9412 ;
  assign n9417 = n9416 ^ n9415 ;
  assign n9425 = n9416 ^ x11 ;
  assign n9424 = ~n2609 & n6650 ;
  assign n9426 = n9425 ^ n9424 ;
  assign n9423 = ~n3227 & n6655 ;
  assign n9427 = n9426 ^ n9423 ;
  assign n9418 = n9154 ^ n5541 ;
  assign n9419 = n9418 ^ n5541 ;
  assign n9420 = ~n5540 & ~n9419 ;
  assign n9421 = n9420 ^ n5541 ;
  assign n9422 = n6648 & n9421 ;
  assign n9428 = n9427 ^ n9422 ;
  assign n9429 = n9417 & n9428 ;
  assign n9430 = n9429 ^ n9416 ;
  assign n9432 = n9431 ^ n9430 ;
  assign n9439 = ~n2609 & n6655 ;
  assign n9437 = ~n2554 & n6650 ;
  assign n9435 = ~n2486 & n6658 ;
  assign n9434 = n9431 ^ x11 ;
  assign n9436 = n9435 ^ n9434 ;
  assign n9438 = n9437 ^ n9436 ;
  assign n9440 = n9439 ^ n9438 ;
  assign n9433 = n5381 & n15413 ;
  assign n9441 = n9440 ^ n9433 ;
  assign n9442 = ~n9432 & ~n9441 ;
  assign n9444 = n9443 ^ n9442 ;
  assign n9445 = n9198 & n9444 ;
  assign n9446 = n9445 ^ n9197 ;
  assign n9448 = n9447 ^ n9446 ;
  assign n9455 = ~n2449 & n6650 ;
  assign n9453 = ~n2486 & n6655 ;
  assign n9451 = ~n2364 & n6658 ;
  assign n9450 = n9447 ^ x11 ;
  assign n9452 = n9451 ^ n9450 ;
  assign n9454 = n9453 ^ n9452 ;
  assign n9456 = n9455 ^ n9454 ;
  assign n9449 = n5283 & n15413 ;
  assign n9457 = n9456 ^ n9449 ;
  assign n9458 = n9448 & n9457 ;
  assign n9459 = n9458 ^ n9447 ;
  assign n9184 = n8814 ^ n8784 ;
  assign n9181 = ~n2364 & n6650 ;
  assign n9179 = ~n2268 & n6658 ;
  assign n9178 = ~n2449 & n6655 ;
  assign n9180 = n9179 ^ n9178 ;
  assign n9182 = n9181 ^ n9180 ;
  assign n9177 = n5144 & n15413 ;
  assign n9183 = n9182 ^ n9177 ;
  assign n9460 = n9183 ^ x11 ;
  assign n9461 = n9184 & n9460 ;
  assign n9462 = ~n9459 & n9461 ;
  assign n9463 = n9462 ^ n9459 ;
  assign n9171 = ~n2364 & n6655 ;
  assign n9169 = ~n2268 & n6650 ;
  assign n9168 = ~n2185 & n6658 ;
  assign n9170 = n9169 ^ n9168 ;
  assign n9172 = n9171 ^ n9170 ;
  assign n9167 = n5832 & n15413 ;
  assign n9173 = n9172 ^ n9167 ;
  assign n9174 = n8847 ^ n8816 ;
  assign n9175 = ~n9173 & ~n9174 ;
  assign n9186 = n9175 ^ n9173 ;
  assign n9185 = n9183 & ~n9184 ;
  assign n9466 = n9185 ^ n9184 ;
  assign n9467 = n9186 & n9466 ;
  assign n9468 = n9463 & n9467 ;
  assign n9187 = n9186 ^ n9174 ;
  assign n9469 = n9187 ^ n9173 ;
  assign n9470 = ~x11 & n9469 ;
  assign n9471 = ~n9468 & n9470 ;
  assign n9176 = x11 & ~n9175 ;
  assign n9188 = ~n9185 & n9187 ;
  assign n9464 = n9188 & n9463 ;
  assign n9465 = n9176 & ~n9464 ;
  assign n9472 = n9471 ^ n9465 ;
  assign n9474 = n9473 ^ n9472 ;
  assign n9478 = ~n2268 & n6655 ;
  assign n9477 = ~n2096 & n6658 ;
  assign n9479 = n9478 ^ n9477 ;
  assign n9480 = n9479 ^ x11 ;
  assign n9476 = ~n2185 & n6650 ;
  assign n9481 = n9480 ^ n9476 ;
  assign n9475 = n5196 & n15413 ;
  assign n9482 = n9481 ^ n9475 ;
  assign n9483 = n9482 ^ n9472 ;
  assign n9484 = ~n9474 & n9483 ;
  assign n9485 = n9484 ^ n9473 ;
  assign n9486 = n9485 ^ n9162 ;
  assign n9487 = n9166 & n9486 ;
  assign n9488 = n9487 ^ n9162 ;
  assign n9490 = n9489 ^ n9488 ;
  assign n9497 = ~n1795 & n6658 ;
  assign n9495 = ~n2096 & n6655 ;
  assign n9493 = ~n1994 & n6650 ;
  assign n9492 = n9489 ^ x11 ;
  assign n9494 = n9493 ^ n9492 ;
  assign n9496 = n9495 ^ n9494 ;
  assign n9498 = n9497 ^ n9496 ;
  assign n9491 = n5168 & n15413 ;
  assign n9499 = n9498 ^ n9491 ;
  assign n9500 = n9490 & n9499 ;
  assign n9501 = n9500 ^ n9489 ;
  assign n9502 = n9501 ^ n9147 ;
  assign n9503 = n9153 & n9502 ;
  assign n9504 = n9503 ^ n9147 ;
  assign n9505 = n9504 ^ n9137 ;
  assign n9506 = n9143 & n9505 ;
  assign n9507 = n9506 ^ n9137 ;
  assign n9508 = n9507 ^ n9127 ;
  assign n9509 = n9133 & n9508 ;
  assign n9510 = n9509 ^ n9127 ;
  assign n9512 = n9511 ^ n9510 ;
  assign n9519 = ~n1351 & n6658 ;
  assign n9517 = ~n1631 & n6655 ;
  assign n9515 = ~n1703 & n6650 ;
  assign n9514 = n9511 ^ x11 ;
  assign n9516 = n9515 ^ n9514 ;
  assign n9518 = n9517 ^ n9516 ;
  assign n9520 = n9519 ^ n9518 ;
  assign n9513 = n4417 & n15413 ;
  assign n9521 = n9520 ^ n9513 ;
  assign n9522 = n9512 & n9521 ;
  assign n9523 = n9522 ^ n9511 ;
  assign n9525 = n9524 ^ n9523 ;
  assign n9532 = ~n1351 & n6650 ;
  assign n9530 = ~n1433 & n6658 ;
  assign n9528 = ~n1703 & n6655 ;
  assign n9527 = n9524 ^ x11 ;
  assign n9529 = n9528 ^ n9527 ;
  assign n9531 = n9530 ^ n9529 ;
  assign n9533 = n9532 ^ n9531 ;
  assign n9526 = n4152 & n15413 ;
  assign n9534 = n9533 ^ n9526 ;
  assign n9535 = n9525 & n9534 ;
  assign n9536 = n9535 ^ n9524 ;
  assign n9537 = n9536 ^ n9117 ;
  assign n9538 = ~n9123 & ~n9537 ;
  assign n9539 = n9538 ^ n9117 ;
  assign n9541 = n9540 ^ n9539 ;
  assign n9548 = ~n1540 & n6650 ;
  assign n9546 = ~n1433 & n6655 ;
  assign n9544 = ~n1214 & n6658 ;
  assign n9543 = n9540 ^ x11 ;
  assign n9545 = n9544 ^ n9543 ;
  assign n9547 = n9546 ^ n9545 ;
  assign n9549 = n9548 ^ n9547 ;
  assign n9542 = ~n4603 & n15413 ;
  assign n9550 = n9549 ^ n9542 ;
  assign n9551 = n9541 & ~n9550 ;
  assign n9552 = n9551 ^ n9540 ;
  assign n9553 = n9552 ^ n9107 ;
  assign n9554 = n9113 & ~n9553 ;
  assign n9555 = n9554 ^ n9107 ;
  assign n9556 = n9555 ^ n9097 ;
  assign n9557 = ~n9103 & ~n9556 ;
  assign n9558 = n9557 ^ n9097 ;
  assign n9569 = n9568 ^ n9558 ;
  assign n9570 = n9569 ^ x5 ;
  assign n9093 = ~n445 & ~n9092 ;
  assign n9571 = n9570 ^ n9093 ;
  assign n9084 = x2 & x3 ;
  assign n9083 = n9078 ^ x4 ;
  assign n9085 = n9084 ^ n9083 ;
  assign n9086 = ~n485 & n9085 ;
  assign n9572 = n9571 ^ n9086 ;
  assign n9574 = n9573 ^ n9572 ;
  assign n9082 = ~n3924 & n9081 ;
  assign n9575 = n9574 ^ n9082 ;
  assign n9588 = n9555 ^ n9103 ;
  assign n9584 = ~n824 & n7146 ;
  assign n9583 = ~n3473 & n7141 ;
  assign n9585 = n9584 ^ n9583 ;
  assign n9586 = n9585 ^ x8 ;
  assign n9577 = x8 ^ x7 ;
  assign n9580 = n3475 & ~n9577 ;
  assign n9581 = n9580 ^ n3476 ;
  assign n9582 = n7128 & ~n9581 ;
  assign n9587 = n9586 ^ n9582 ;
  assign n9589 = n9588 ^ n9587 ;
  assign n9597 = ~n3508 & n7135 ;
  assign n9595 = ~n3473 & n8054 ;
  assign n9593 = ~n1109 & n7146 ;
  assign n9591 = n9552 ^ n9113 ;
  assign n9592 = n9591 ^ x8 ;
  assign n9594 = n9593 ^ n9592 ;
  assign n9596 = n9595 ^ n9594 ;
  assign n9598 = n9597 ^ n9596 ;
  assign n9590 = ~n824 & n7141 ;
  assign n9599 = n9598 ^ n9590 ;
  assign n9607 = ~n4050 & n7135 ;
  assign n9603 = n9550 ^ n9539 ;
  assign n9604 = n9603 ^ x8 ;
  assign n9602 = ~n824 & n8054 ;
  assign n9605 = n9604 ^ n9602 ;
  assign n9601 = ~n968 & n7146 ;
  assign n9606 = n9605 ^ n9601 ;
  assign n9608 = n9607 ^ n9606 ;
  assign n9600 = ~n1109 & n7141 ;
  assign n9609 = n9608 ^ n9600 ;
  assign n9621 = n9536 ^ n9123 ;
  assign n9618 = ~n1214 & n7146 ;
  assign n9611 = n1109 ^ x8 ;
  assign n9612 = n9611 ^ x7 ;
  assign n9613 = n9612 ^ n1109 ;
  assign n9614 = ~n3904 & n9613 ;
  assign n9615 = n9614 ^ n1109 ;
  assign n9616 = n7128 & ~n9615 ;
  assign n9617 = n9616 ^ x8 ;
  assign n9619 = n9618 ^ n9617 ;
  assign n9610 = ~n968 & n7141 ;
  assign n9620 = n9619 ^ n9610 ;
  assign n9622 = n9621 ^ n9620 ;
  assign n10056 = n9534 ^ n9523 ;
  assign n10068 = n10056 ^ n9621 ;
  assign n10043 = n9521 ^ n9510 ;
  assign n9630 = ~n4610 & n7135 ;
  assign n9628 = ~n1433 & n7141 ;
  assign n9626 = ~n1540 & n8054 ;
  assign n9624 = n9507 ^ n9133 ;
  assign n9625 = n9624 ^ x8 ;
  assign n9627 = n9626 ^ n9625 ;
  assign n9629 = n9628 ^ n9627 ;
  assign n9631 = n9630 ^ n9629 ;
  assign n9623 = ~n1351 & n7146 ;
  assign n9632 = n9631 ^ n9623 ;
  assign n9640 = n4152 & n7135 ;
  assign n9638 = ~n1433 & n8054 ;
  assign n9636 = ~n1351 & n7141 ;
  assign n9634 = n9504 ^ n9143 ;
  assign n9635 = n9634 ^ x8 ;
  assign n9637 = n9636 ^ n9635 ;
  assign n9639 = n9638 ^ n9637 ;
  assign n9641 = n9640 ^ n9639 ;
  assign n9633 = ~n1703 & n7146 ;
  assign n9642 = n9641 ^ n9633 ;
  assign n10022 = n9501 ^ n9153 ;
  assign n9651 = n9499 ^ n9488 ;
  assign n9649 = ~n1871 & n7146 ;
  assign n9647 = ~n4615 & n7135 ;
  assign n9644 = ~n1631 & n7141 ;
  assign n9643 = ~n1703 & n8054 ;
  assign n9645 = n9644 ^ n9643 ;
  assign n9646 = n9645 ^ x8 ;
  assign n9648 = n9647 ^ n9646 ;
  assign n9650 = n9649 ^ n9648 ;
  assign n9652 = n9651 ^ n9650 ;
  assign n10006 = n9485 ^ n9166 ;
  assign n9662 = ~n1795 & n7141 ;
  assign n9659 = n9482 ^ n9474 ;
  assign n9660 = n9659 ^ x8 ;
  assign n9656 = n5184 & ~n9577 ;
  assign n9657 = n9656 ^ n4859 ;
  assign n9658 = n7128 & ~n9657 ;
  assign n9661 = n9660 ^ n9658 ;
  assign n9663 = n9662 ^ n9661 ;
  assign n9653 = ~n1994 & n7146 ;
  assign n9664 = n9663 ^ n9653 ;
  assign n9679 = ~n1994 & n7141 ;
  assign n9674 = n9183 ^ n9173 ;
  assign n9675 = n9674 ^ n9174 ;
  assign n9671 = n9460 ^ n9459 ;
  assign n9672 = n9460 ^ n9184 ;
  assign n9673 = n9671 & n9672 ;
  assign n9676 = n9675 ^ n9673 ;
  assign n9677 = n9676 ^ x8 ;
  assign n9668 = ~n4384 & ~n9577 ;
  assign n9669 = n9668 ^ n5168 ;
  assign n9670 = n7128 & n9669 ;
  assign n9678 = n9677 ^ n9670 ;
  assign n9680 = n9679 ^ n9678 ;
  assign n9665 = ~n2096 & n7146 ;
  assign n9681 = n9680 ^ n9665 ;
  assign n9986 = n9459 ^ n9184 ;
  assign n9987 = n9986 ^ n9460 ;
  assign n9686 = ~n2185 & n7141 ;
  assign n9685 = n5196 & n7135 ;
  assign n9687 = n9686 ^ n9685 ;
  assign n9688 = n9687 ^ x8 ;
  assign n9684 = ~n2268 & n7146 ;
  assign n9689 = n9688 ^ n9684 ;
  assign n9683 = ~n2096 & n8054 ;
  assign n9690 = n9689 ^ n9683 ;
  assign n9682 = n9457 ^ n9446 ;
  assign n9691 = n9690 ^ n9682 ;
  assign n9700 = n5144 & n7135 ;
  assign n9698 = ~n2268 & n8054 ;
  assign n9696 = ~n2449 & n7146 ;
  assign n9694 = n9441 ^ n9430 ;
  assign n9695 = n9694 ^ x8 ;
  assign n9697 = n9696 ^ n9695 ;
  assign n9699 = n9698 ^ n9697 ;
  assign n9701 = n9700 ^ n9699 ;
  assign n9693 = ~n2364 & n7141 ;
  assign n9702 = n9701 ^ n9693 ;
  assign n9711 = n9428 ^ n9415 ;
  assign n9709 = ~n2449 & n7141 ;
  assign n9707 = n5283 & n7135 ;
  assign n9704 = ~n2486 & n7146 ;
  assign n9703 = ~n2364 & n8054 ;
  assign n9705 = n9704 ^ n9703 ;
  assign n9706 = n9705 ^ x8 ;
  assign n9708 = n9707 ^ n9706 ;
  assign n9710 = n9709 ^ n9708 ;
  assign n9712 = n9711 ^ n9710 ;
  assign n9722 = n5520 & n7135 ;
  assign n9720 = ~n2554 & n7146 ;
  assign n9718 = ~n2449 & n8054 ;
  assign n9714 = n9404 ^ n9206 ;
  assign n9715 = ~n9405 & n9714 ;
  assign n9716 = n9715 ^ n9220 ;
  assign n9717 = n9716 ^ x8 ;
  assign n9719 = n9718 ^ n9717 ;
  assign n9721 = n9720 ^ n9719 ;
  assign n9723 = n9722 ^ n9721 ;
  assign n9713 = ~n2486 & n7141 ;
  assign n9724 = n9723 ^ n9713 ;
  assign n9949 = n9405 ^ n9206 ;
  assign n9733 = n5541 & n7135 ;
  assign n9731 = ~n2554 & n8054 ;
  assign n9729 = ~n3227 & n7146 ;
  assign n9726 = n9398 ^ n8751 ;
  assign n9727 = n9726 ^ n9400 ;
  assign n9728 = n9727 ^ x8 ;
  assign n9730 = n9729 ^ n9728 ;
  assign n9732 = n9731 ^ n9730 ;
  assign n9734 = n9733 ^ n9732 ;
  assign n9725 = ~n2609 & n7141 ;
  assign n9735 = n9734 ^ n9725 ;
  assign n9744 = n9395 ^ n9239 ;
  assign n9742 = ~n3227 & n7141 ;
  assign n9740 = n7029 & n7135 ;
  assign n9737 = ~n2609 & n8054 ;
  assign n9736 = ~n2646 & n7146 ;
  assign n9738 = n9737 ^ n9736 ;
  assign n9739 = n9738 ^ x8 ;
  assign n9741 = n9740 ^ n9739 ;
  assign n9743 = n9742 ^ n9741 ;
  assign n9745 = n9744 ^ n9743 ;
  assign n9753 = n6900 & n7135 ;
  assign n9749 = n9392 ^ n9250 ;
  assign n9750 = n9749 ^ x8 ;
  assign n9748 = ~n3227 & n8054 ;
  assign n9751 = n9750 ^ n9748 ;
  assign n9747 = ~n2738 & n7146 ;
  assign n9752 = n9751 ^ n9747 ;
  assign n9754 = n9753 ^ n9752 ;
  assign n9746 = ~n2646 & n7141 ;
  assign n9755 = n9754 ^ n9746 ;
  assign n9927 = n9389 ^ n9260 ;
  assign n9763 = ~n6907 & n7135 ;
  assign n9761 = ~n2738 & n8054 ;
  assign n9759 = ~n2836 & n7141 ;
  assign n9757 = n9387 ^ n9375 ;
  assign n9758 = n9757 ^ x8 ;
  assign n9760 = n9759 ^ n9758 ;
  assign n9762 = n9761 ^ n9760 ;
  assign n9764 = n9763 ^ n9762 ;
  assign n9756 = ~n3151 & n7146 ;
  assign n9765 = n9764 ^ n9756 ;
  assign n9775 = n9285 ^ x11 ;
  assign n9776 = n9775 ^ n9267 ;
  assign n9773 = ~n3151 & n7141 ;
  assign n9771 = n6237 & n7135 ;
  assign n9768 = ~n2836 & n8054 ;
  assign n9767 = ~n2924 & n7146 ;
  assign n9769 = n9768 ^ n9767 ;
  assign n9770 = n9769 ^ x8 ;
  assign n9772 = n9771 ^ n9770 ;
  assign n9774 = n9773 ^ n9772 ;
  assign n9777 = n9776 ^ n9774 ;
  assign n9766 = ~n3337 & n4897 ;
  assign n9778 = n9777 ^ n9766 ;
  assign n9787 = n9284 ^ n9272 ;
  assign n9785 = ~n2958 & n7146 ;
  assign n9783 = n6286 & n7135 ;
  assign n9780 = ~n3151 & n8054 ;
  assign n9779 = ~n2924 & n7141 ;
  assign n9781 = n9780 ^ n9779 ;
  assign n9782 = n9781 ^ x8 ;
  assign n9784 = n9783 ^ n9782 ;
  assign n9786 = n9785 ^ n9784 ;
  assign n9788 = n9787 ^ n9786 ;
  assign n9910 = ~n2958 & n7141 ;
  assign n9908 = n6344 & n7135 ;
  assign n9905 = ~n3099 & n7146 ;
  assign n9904 = ~n2924 & n8054 ;
  assign n9906 = n9905 ^ n9904 ;
  assign n9907 = n9906 ^ x8 ;
  assign n9909 = n9908 ^ n9907 ;
  assign n9911 = n9910 ^ n9909 ;
  assign n9830 = n3337 ^ x8 ;
  assign n9796 = ~n3337 & ~n18156 ;
  assign n9797 = ~n3027 & n7128 ;
  assign n9798 = x8 & ~n9797 ;
  assign n9799 = ~n9796 & n9798 ;
  assign n9810 = ~n3099 & n7128 ;
  assign n9809 = ~n3337 & n7146 ;
  assign n9811 = n9810 ^ n9809 ;
  assign n9806 = n3337 & n7135 ;
  assign n9807 = n9806 ^ n7141 ;
  assign n9808 = ~n3027 & n9807 ;
  assign n9812 = n9811 ^ n9808 ;
  assign n9813 = n9799 & ~n9812 ;
  assign n9793 = ~n2958 & n7128 ;
  assign n9792 = ~n6439 & n7135 ;
  assign n9794 = n9793 ^ n9792 ;
  assign n9790 = ~n3027 & n7146 ;
  assign n9789 = ~n3099 & n7141 ;
  assign n9791 = n9790 ^ n9789 ;
  assign n9795 = n9794 ^ n9791 ;
  assign n9814 = n9813 ^ n9795 ;
  assign n9815 = n9814 ^ x9 ;
  assign n9831 = n9830 ^ n9815 ;
  assign n9865 = n9831 ^ n9795 ;
  assign n9816 = n9815 ^ n3337 ;
  assign n9817 = n9816 ^ n9814 ;
  assign n9893 = n9865 ^ n9817 ;
  assign n9894 = n9893 ^ x9 ;
  assign n9895 = n9894 ^ n9795 ;
  assign n9847 = n9795 & ~n9814 ;
  assign n9848 = n9847 ^ n9816 ;
  assign n9832 = n9831 ^ n9817 ;
  assign n9849 = n9848 ^ n9832 ;
  assign n9850 = n9849 ^ n9813 ;
  assign n9851 = n9832 ^ n3337 ;
  assign n9852 = n9851 ^ n9813 ;
  assign n9853 = n9850 & n9852 ;
  assign n9829 = n9816 ^ n9795 ;
  assign n9836 = n9829 ^ n9815 ;
  assign n9838 = n9836 ^ n9832 ;
  assign n9854 = n9838 ^ n9815 ;
  assign n9855 = n9854 ^ n9830 ;
  assign n9856 = n9838 ^ n9816 ;
  assign n9857 = n9856 ^ n9830 ;
  assign n9858 = ~n9855 & ~n9857 ;
  assign n9859 = n9853 & n9858 ;
  assign n9860 = n9859 ^ n9847 ;
  assign n9861 = n9860 ^ n3337 ;
  assign n9900 = n9895 ^ n9861 ;
  assign n9821 = n9816 ^ x8 ;
  assign n9823 = n9821 ^ x9 ;
  assign n9825 = n9823 ^ n9795 ;
  assign n9826 = n9825 ^ n9821 ;
  assign n9901 = n9900 ^ n9826 ;
  assign n9902 = n9901 ^ n9813 ;
  assign n9903 = n9902 ^ n9825 ;
  assign n9912 = n9911 ^ n9903 ;
  assign n9914 = ~n3337 & n6647 ;
  assign n9913 = n9911 ^ n9268 ;
  assign n9915 = n9914 ^ n9913 ;
  assign n9916 = n9912 & n9915 ;
  assign n9917 = n9916 ^ n9911 ;
  assign n9918 = n9917 ^ n9786 ;
  assign n9919 = n9788 & n9918 ;
  assign n9920 = n9919 ^ n9786 ;
  assign n9921 = n9920 ^ n9774 ;
  assign n9922 = n9778 & n9921 ;
  assign n9923 = n9922 ^ n9774 ;
  assign n9924 = n9923 ^ n9757 ;
  assign n9925 = n9765 & n9924 ;
  assign n9926 = n9925 ^ n9757 ;
  assign n9928 = n9927 ^ n9926 ;
  assign n9935 = ~n5651 & n7135 ;
  assign n9933 = ~n2836 & n7146 ;
  assign n9931 = ~n2646 & n8054 ;
  assign n9930 = n9927 ^ x8 ;
  assign n9932 = n9931 ^ n9930 ;
  assign n9934 = n9933 ^ n9932 ;
  assign n9936 = n9935 ^ n9934 ;
  assign n9929 = ~n2738 & n7141 ;
  assign n9937 = n9936 ^ n9929 ;
  assign n9938 = n9928 & n9937 ;
  assign n9939 = n9938 ^ n9927 ;
  assign n9940 = n9939 ^ n9749 ;
  assign n9941 = ~n9755 & ~n9940 ;
  assign n9942 = n9941 ^ n9749 ;
  assign n9943 = n9942 ^ n9743 ;
  assign n9944 = n9745 & ~n9943 ;
  assign n9945 = n9944 ^ n9743 ;
  assign n9946 = n9945 ^ n9727 ;
  assign n9947 = n9735 & n9946 ;
  assign n9948 = n9947 ^ n9727 ;
  assign n9950 = n9949 ^ n9948 ;
  assign n9957 = n5381 & n7135 ;
  assign n9955 = ~n2486 & n8054 ;
  assign n9953 = ~n2609 & n7146 ;
  assign n9952 = n9949 ^ x8 ;
  assign n9954 = n9953 ^ n9952 ;
  assign n9956 = n9955 ^ n9954 ;
  assign n9958 = n9957 ^ n9956 ;
  assign n9951 = ~n2554 & n7141 ;
  assign n9959 = n9958 ^ n9951 ;
  assign n9960 = n9950 & n9959 ;
  assign n9961 = n9960 ^ n9949 ;
  assign n9962 = n9961 ^ n9716 ;
  assign n9963 = n9724 & n9962 ;
  assign n9964 = n9963 ^ n9716 ;
  assign n9965 = n9964 ^ n9710 ;
  assign n9966 = n9712 & n9965 ;
  assign n9967 = n9966 ^ n9710 ;
  assign n9968 = n9967 ^ n9694 ;
  assign n9969 = ~n9702 & ~n9968 ;
  assign n9970 = n9969 ^ n9694 ;
  assign n9692 = n9444 ^ n9197 ;
  assign n9971 = n9970 ^ n9692 ;
  assign n9978 = ~n2185 & n8054 ;
  assign n9976 = ~n2268 & n7141 ;
  assign n9974 = n5832 & n7135 ;
  assign n9973 = n9692 ^ x8 ;
  assign n9975 = n9974 ^ n9973 ;
  assign n9977 = n9976 ^ n9975 ;
  assign n9979 = n9978 ^ n9977 ;
  assign n9972 = ~n2364 & n7146 ;
  assign n9980 = n9979 ^ n9972 ;
  assign n9981 = n9971 & n9980 ;
  assign n9982 = n9981 ^ n9970 ;
  assign n9983 = n9982 ^ n9682 ;
  assign n9984 = n9691 & n9983 ;
  assign n9985 = n9984 ^ n9690 ;
  assign n9988 = n9987 ^ n9985 ;
  assign n9995 = n5409 & n7135 ;
  assign n9993 = ~n2185 & n7146 ;
  assign n9991 = ~n1994 & n8054 ;
  assign n9990 = n9987 ^ x8 ;
  assign n9992 = n9991 ^ n9990 ;
  assign n9994 = n9993 ^ n9992 ;
  assign n9996 = n9995 ^ n9994 ;
  assign n9989 = ~n2096 & n7141 ;
  assign n9997 = n9996 ^ n9989 ;
  assign n9998 = n9988 & n9997 ;
  assign n9999 = n9998 ^ n9987 ;
  assign n10000 = n9999 ^ n9676 ;
  assign n10001 = n9681 & ~n10000 ;
  assign n10002 = n10001 ^ n9999 ;
  assign n10003 = n10002 ^ n9659 ;
  assign n10004 = ~n9664 & ~n10003 ;
  assign n10005 = n10004 ^ n9659 ;
  assign n10007 = n10006 ^ n10005 ;
  assign n10014 = ~n4392 & n7135 ;
  assign n10012 = ~n1631 & n8054 ;
  assign n10010 = ~n1871 & n7141 ;
  assign n10009 = n10006 ^ x8 ;
  assign n10011 = n10010 ^ n10009 ;
  assign n10013 = n10012 ^ n10011 ;
  assign n10015 = n10014 ^ n10013 ;
  assign n10008 = ~n1795 & n7146 ;
  assign n10016 = n10015 ^ n10008 ;
  assign n10017 = ~n10007 & n10016 ;
  assign n10018 = n10017 ^ n10006 ;
  assign n10019 = n10018 ^ n9650 ;
  assign n10020 = n9652 & n10019 ;
  assign n10021 = n10020 ^ n9650 ;
  assign n10023 = n10022 ^ n10021 ;
  assign n10032 = ~n1703 & n7141 ;
  assign n10030 = n10022 ^ x8 ;
  assign n10025 = n9577 ^ n4417 ;
  assign n10026 = n10025 ^ n4417 ;
  assign n10027 = ~n4416 & ~n10026 ;
  assign n10028 = n10027 ^ n4417 ;
  assign n10029 = n7128 & n10028 ;
  assign n10031 = n10030 ^ n10029 ;
  assign n10033 = n10032 ^ n10031 ;
  assign n10024 = ~n1631 & n7146 ;
  assign n10034 = n10033 ^ n10024 ;
  assign n10035 = n10023 & n10034 ;
  assign n10036 = n10035 ^ n10022 ;
  assign n10037 = n10036 ^ n9634 ;
  assign n10038 = n9642 & n10037 ;
  assign n10039 = n10038 ^ n9634 ;
  assign n10040 = n10039 ^ n9624 ;
  assign n10041 = n9632 & n10040 ;
  assign n10042 = n10041 ^ n9624 ;
  assign n10044 = n10043 ^ n10042 ;
  assign n10051 = ~n4603 & n7135 ;
  assign n10049 = ~n1433 & n7146 ;
  assign n10047 = ~n1214 & n8054 ;
  assign n10046 = n10043 ^ x8 ;
  assign n10048 = n10047 ^ n10046 ;
  assign n10050 = n10049 ^ n10048 ;
  assign n10052 = n10051 ^ n10050 ;
  assign n10045 = ~n1540 & n7141 ;
  assign n10053 = n10052 ^ n10045 ;
  assign n10054 = n10044 & n10053 ;
  assign n10055 = n10054 ^ n10043 ;
  assign n10057 = n10056 ^ n10055 ;
  assign n10064 = n3521 & n7135 ;
  assign n10062 = ~n968 & n8054 ;
  assign n10060 = ~n1214 & n7141 ;
  assign n10059 = n10056 ^ x8 ;
  assign n10061 = n10060 ^ n10059 ;
  assign n10063 = n10062 ^ n10061 ;
  assign n10065 = n10064 ^ n10063 ;
  assign n10058 = ~n1540 & n7146 ;
  assign n10066 = n10065 ^ n10058 ;
  assign n10067 = n10057 & n10066 ;
  assign n10069 = n10068 ^ n10067 ;
  assign n10070 = ~n9622 & ~n10069 ;
  assign n10071 = n10070 ^ n9621 ;
  assign n10072 = n10071 ^ n9603 ;
  assign n10073 = n9609 & ~n10072 ;
  assign n10074 = n10073 ^ n9603 ;
  assign n10075 = n10074 ^ n9591 ;
  assign n10076 = ~n9599 & ~n10075 ;
  assign n10077 = n10076 ^ n9591 ;
  assign n10078 = n10077 ^ n9587 ;
  assign n10079 = n9589 & ~n10078 ;
  assign n10080 = n10079 ^ n10077 ;
  assign n10081 = n10080 ^ n9569 ;
  assign n10082 = n9575 & ~n10081 ;
  assign n10083 = n10082 ^ n9569 ;
  assign n10084 = n9562 ^ n9558 ;
  assign n10085 = ~n9568 & n10084 ;
  assign n10086 = n10085 ^ n9562 ;
  assign n10087 = ~n10083 & n10086 ;
  assign n10088 = ~n9076 & n10087 ;
  assign n10093 = n4515 & n9081 ;
  assign n10090 = ~n3943 & n9085 ;
  assign n10089 = ~n485 & ~n9092 ;
  assign n10091 = n10090 ^ n10089 ;
  assign n10092 = n10091 ^ x5 ;
  assign n10094 = n10093 ^ n10092 ;
  assign n10095 = n10088 & ~n10094 ;
  assign n10109 = n10108 ^ n10098 ;
  assign n10110 = ~n10095 & n10109 ;
  assign n10121 = n10094 ^ n9076 ;
  assign n10122 = n10121 ^ n10086 ;
  assign n10123 = n10122 ^ n10083 ;
  assign n10111 = n10086 ^ n9076 ;
  assign n10113 = n10086 ^ n10083 ;
  assign n10114 = n10111 & ~n10113 ;
  assign n10117 = n10114 ^ n10083 ;
  assign n10118 = n10094 ^ n10088 ;
  assign n10119 = n10118 ^ n10095 ;
  assign n10120 = ~n10117 & ~n10119 ;
  assign n10124 = n10123 ^ n10120 ;
  assign n10112 = n10111 ^ n10088 ;
  assign n10115 = n10114 ^ n10112 ;
  assign n10116 = n10094 & n10115 ;
  assign n10125 = n10124 ^ n10116 ;
  assign n10126 = n10110 & n10125 ;
  assign n10127 = n10126 ^ n10095 ;
  assign n11496 = n10080 ^ n9575 ;
  assign n10131 = n9081 ^ n9077 ;
  assign n10132 = ~n445 & n10131 ;
  assign n10130 = ~n317 & n9085 ;
  assign n10133 = n10132 ^ n10130 ;
  assign n10134 = n10133 ^ x5 ;
  assign n10129 = ~n649 & ~n9092 ;
  assign n10135 = n10134 ^ n10129 ;
  assign n10128 = n4073 & n9081 ;
  assign n10136 = n10135 ^ n10128 ;
  assign n10145 = n10071 ^ n9609 ;
  assign n10140 = ~n317 & n10131 ;
  assign n10139 = ~n3473 & ~n9092 ;
  assign n10141 = n10140 ^ n10139 ;
  assign n10142 = n10141 ^ x5 ;
  assign n10138 = ~n649 & n9085 ;
  assign n10143 = n10142 ^ n10138 ;
  assign n10137 = n3956 & n9081 ;
  assign n10144 = n10143 ^ n10137 ;
  assign n10146 = n10145 ^ n10144 ;
  assign n10158 = ~n1109 & ~n9092 ;
  assign n10155 = n10066 ^ n10055 ;
  assign n10156 = n10155 ^ x5 ;
  assign n10152 = n3388 & n9089 ;
  assign n10153 = n10152 ^ n3473 ;
  assign n10154 = n9077 & ~n10153 ;
  assign n10157 = n10156 ^ n10154 ;
  assign n10159 = n10158 ^ n10157 ;
  assign n10148 = ~n824 & n9085 ;
  assign n10160 = n10159 ^ n10148 ;
  assign n10171 = ~n1109 & n9085 ;
  assign n10168 = n10053 ^ n10042 ;
  assign n10169 = n10168 ^ x5 ;
  assign n10165 = n4044 & n9089 ;
  assign n10166 = n10165 ^ n824 ;
  assign n10167 = n9077 & ~n10166 ;
  assign n10170 = n10169 ^ n10167 ;
  assign n10172 = n10171 ^ n10170 ;
  assign n10161 = ~n968 & ~n9092 ;
  assign n10173 = n10172 ^ n10161 ;
  assign n10666 = n10039 ^ n9632 ;
  assign n10651 = n10036 ^ n9642 ;
  assign n10194 = ~n1351 & n9085 ;
  assign n10191 = n10016 ^ n10005 ;
  assign n10192 = n10191 ^ x5 ;
  assign n10188 = ~n3815 & n9089 ;
  assign n10189 = n10188 ^ n1433 ;
  assign n10190 = n9077 & ~n10189 ;
  assign n10193 = n10192 ^ n10190 ;
  assign n10195 = n10194 ^ n10193 ;
  assign n10183 = ~n1703 & ~n9092 ;
  assign n10196 = n10195 ^ n10183 ;
  assign n10205 = n10002 ^ n9664 ;
  assign n10200 = ~n1703 & n9085 ;
  assign n10199 = n4417 & n9081 ;
  assign n10201 = n10200 ^ n10199 ;
  assign n10202 = n10201 ^ x5 ;
  assign n10198 = ~n1631 & ~n9092 ;
  assign n10203 = n10202 ^ n10198 ;
  assign n10197 = ~n1351 & n10131 ;
  assign n10204 = n10203 ^ n10197 ;
  assign n10206 = n10205 ^ n10204 ;
  assign n10216 = ~n1631 & n9085 ;
  assign n10215 = ~n1871 & ~n9092 ;
  assign n10217 = n10216 ^ n10215 ;
  assign n10208 = n1703 ^ x5 ;
  assign n10209 = n10208 ^ x4 ;
  assign n10210 = n10209 ^ n1703 ;
  assign n10211 = n3808 & n10210 ;
  assign n10212 = n10211 ^ n1703 ;
  assign n10213 = n9077 & ~n10212 ;
  assign n10214 = n10213 ^ x5 ;
  assign n10218 = n10217 ^ n10214 ;
  assign n10207 = n9999 ^ n9681 ;
  assign n10219 = n10218 ^ n10207 ;
  assign n10230 = n9997 ^ n9985 ;
  assign n10226 = ~n1871 & n9085 ;
  assign n10225 = ~n1795 & ~n9092 ;
  assign n10227 = n10226 ^ n10225 ;
  assign n10228 = n10227 ^ x5 ;
  assign n10222 = n4391 & ~n9089 ;
  assign n10223 = n10222 ^ n4392 ;
  assign n10224 = n9077 & ~n10223 ;
  assign n10229 = n10228 ^ n10224 ;
  assign n10231 = n10230 ^ n10229 ;
  assign n10240 = n9982 ^ n9691 ;
  assign n10235 = ~n1994 & ~n9092 ;
  assign n10234 = ~n4859 & n9081 ;
  assign n10236 = n10235 ^ n10234 ;
  assign n10237 = n10236 ^ x5 ;
  assign n10233 = ~n1795 & n9085 ;
  assign n10238 = n10237 ^ n10233 ;
  assign n10232 = ~n1871 & n10131 ;
  assign n10239 = n10238 ^ n10232 ;
  assign n10241 = n10240 ^ n10239 ;
  assign n10250 = ~n1795 & n10131 ;
  assign n10245 = n9980 ^ n9970 ;
  assign n10246 = n10245 ^ x5 ;
  assign n10244 = ~n2096 & ~n9092 ;
  assign n10247 = n10246 ^ n10244 ;
  assign n10243 = ~n1994 & n9085 ;
  assign n10248 = n10247 ^ n10243 ;
  assign n10242 = n5168 & n9081 ;
  assign n10249 = n10248 ^ n10242 ;
  assign n10251 = n10250 ^ n10249 ;
  assign n10260 = n9967 ^ n9702 ;
  assign n10255 = ~n2185 & ~n9092 ;
  assign n10254 = ~n2096 & n9085 ;
  assign n10256 = n10255 ^ n10254 ;
  assign n10257 = n10256 ^ x5 ;
  assign n10253 = n5409 & n9081 ;
  assign n10258 = n10257 ^ n10253 ;
  assign n10252 = ~n1994 & n10131 ;
  assign n10259 = n10258 ^ n10252 ;
  assign n10261 = n10260 ^ n10259 ;
  assign n10593 = n9964 ^ n9712 ;
  assign n10269 = n5832 & n9081 ;
  assign n10265 = n9961 ^ n9724 ;
  assign n10266 = n10265 ^ x5 ;
  assign n10264 = ~n2364 & ~n9092 ;
  assign n10267 = n10266 ^ n10264 ;
  assign n10263 = ~n2268 & n9085 ;
  assign n10268 = n10267 ^ n10263 ;
  assign n10270 = n10269 ^ n10268 ;
  assign n10262 = ~n2185 & n10131 ;
  assign n10271 = n10270 ^ n10262 ;
  assign n10577 = n9959 ^ n9948 ;
  assign n10279 = n5283 & n9081 ;
  assign n10277 = ~n2486 & ~n9092 ;
  assign n10275 = ~n2449 & n9085 ;
  assign n10273 = n9945 ^ n9735 ;
  assign n10274 = n10273 ^ x5 ;
  assign n10276 = n10275 ^ n10274 ;
  assign n10278 = n10277 ^ n10276 ;
  assign n10280 = n10279 ^ n10278 ;
  assign n10272 = ~n2364 & n10131 ;
  assign n10281 = n10280 ^ n10272 ;
  assign n10561 = n9942 ^ n9745 ;
  assign n10289 = n5381 & n9081 ;
  assign n10287 = ~n2554 & n9085 ;
  assign n10285 = ~n2609 & ~n9092 ;
  assign n10283 = n9939 ^ n9755 ;
  assign n10284 = n10283 ^ x5 ;
  assign n10286 = n10285 ^ n10284 ;
  assign n10288 = n10287 ^ n10286 ;
  assign n10290 = n10289 ^ n10288 ;
  assign n10282 = ~n2486 & n10131 ;
  assign n10291 = n10290 ^ n10282 ;
  assign n10545 = n9937 ^ n9926 ;
  assign n10299 = n7029 & n9081 ;
  assign n10295 = n9923 ^ n9765 ;
  assign n10296 = n10295 ^ x5 ;
  assign n10294 = ~n2646 & ~n9092 ;
  assign n10297 = n10296 ^ n10294 ;
  assign n10293 = ~n3227 & n9085 ;
  assign n10298 = n10297 ^ n10293 ;
  assign n10300 = n10299 ^ n10298 ;
  assign n10292 = ~n2609 & n10131 ;
  assign n10301 = n10300 ^ n10292 ;
  assign n10312 = ~n2646 & n9085 ;
  assign n10309 = n9920 ^ n9778 ;
  assign n10310 = n10309 ^ x5 ;
  assign n10306 = ~n6176 & n9089 ;
  assign n10307 = n10306 ^ n3227 ;
  assign n10308 = n9077 & ~n10307 ;
  assign n10311 = n10310 ^ n10308 ;
  assign n10313 = n10312 ^ n10311 ;
  assign n10302 = ~n2738 & ~n9092 ;
  assign n10314 = n10313 ^ n10302 ;
  assign n10526 = n9917 ^ n9788 ;
  assign n10323 = n9915 ^ n9903 ;
  assign n10319 = ~n2836 & n9085 ;
  assign n10318 = ~n3151 & ~n9092 ;
  assign n10320 = n10319 ^ n10318 ;
  assign n10321 = n10320 ^ x5 ;
  assign n10316 = n3347 & n9081 ;
  assign n10315 = ~n2738 & n9077 ;
  assign n10317 = n10316 ^ n10315 ;
  assign n10322 = n10321 ^ n10317 ;
  assign n10324 = n10323 ^ n10322 ;
  assign n10510 = ~n2924 & ~n9092 ;
  assign n10509 = n6237 & n9081 ;
  assign n10511 = n10510 ^ n10509 ;
  assign n10512 = n10511 ^ x5 ;
  assign n10508 = ~n3151 & n9085 ;
  assign n10513 = n10512 ^ n10508 ;
  assign n10507 = ~n2836 & n10131 ;
  assign n10514 = n10513 ^ n10507 ;
  assign n9800 = n9799 ^ x8 ;
  assign n10333 = n9812 ^ n9800 ;
  assign n10329 = ~n2958 & ~n9092 ;
  assign n10328 = ~n2924 & n9085 ;
  assign n10330 = n10329 ^ n10328 ;
  assign n10331 = n10330 ^ x5 ;
  assign n10326 = ~n6282 & n9081 ;
  assign n10325 = ~n3151 & n9077 ;
  assign n10327 = n10326 ^ n10325 ;
  assign n10332 = n10331 ^ n10327 ;
  assign n10334 = n10333 ^ n10332 ;
  assign n10490 = n7140 & n9796 ;
  assign n10491 = n10490 ^ n9797 ;
  assign n10335 = ~n3027 & n9077 ;
  assign n10336 = x5 & ~n18627 ;
  assign n10337 = n3337 & n10336 ;
  assign n10338 = ~n10335 & n10337 ;
  assign n10339 = n10338 ^ n10336 ;
  assign n10340 = n10339 ^ x5 ;
  assign n10349 = ~n3099 & n9077 ;
  assign n10348 = ~n3337 & ~n9092 ;
  assign n10350 = n10349 ^ n10348 ;
  assign n10345 = n3337 & n9081 ;
  assign n10346 = n10345 ^ n9085 ;
  assign n10347 = ~n3027 & n10346 ;
  assign n10351 = n10350 ^ n10347 ;
  assign n10352 = n10340 & ~n10351 ;
  assign n10357 = ~n3027 & ~n9092 ;
  assign n10355 = ~n2958 & n10131 ;
  assign n10354 = ~n3099 & n9085 ;
  assign n10356 = n10355 ^ n10354 ;
  assign n10358 = n10357 ^ n10356 ;
  assign n10353 = n6440 & n9081 ;
  assign n10359 = n10358 ^ n10353 ;
  assign n10428 = ~n10352 & n10359 ;
  assign n10411 = n3337 ^ x5 ;
  assign n10408 = n10411 ^ n10352 ;
  assign n10429 = n10428 ^ n10408 ;
  assign n10418 = n10352 ^ x5 ;
  assign n10430 = n10429 ^ n10418 ;
  assign n10360 = n10359 ^ n10352 ;
  assign n10431 = n10430 ^ n10360 ;
  assign n10375 = n3337 ^ x6 ;
  assign n10414 = n10375 ^ n10359 ;
  assign n10415 = n10414 ^ x5 ;
  assign n10416 = n10415 ^ n10352 ;
  assign n10424 = n10416 ^ n10408 ;
  assign n10432 = n10424 ^ n10418 ;
  assign n10433 = n10432 ^ n10360 ;
  assign n10434 = ~n10431 & n10433 ;
  assign n10417 = n10416 ^ n10411 ;
  assign n10419 = n10418 ^ n10417 ;
  assign n10435 = n10419 ^ n10416 ;
  assign n10421 = n10419 ^ n10360 ;
  assign n10436 = n10435 ^ n10421 ;
  assign n10437 = n10419 ^ n10408 ;
  assign n10438 = n10437 ^ n10421 ;
  assign n10439 = n10436 & n10438 ;
  assign n10440 = n10434 & n10439 ;
  assign n10441 = n10440 ^ n10428 ;
  assign n10442 = n10441 ^ n10424 ;
  assign n10422 = n10421 ^ n10417 ;
  assign n10443 = n10442 ^ n10422 ;
  assign n10444 = n10443 ^ n10414 ;
  assign n10364 = n10360 ^ x6 ;
  assign n10365 = n10364 ^ n3337 ;
  assign n10366 = n10365 ^ n10360 ;
  assign n10361 = n10360 ^ x5 ;
  assign n10367 = n10366 ^ n10361 ;
  assign n10369 = n10367 ^ x6 ;
  assign n10370 = n10369 ^ n10359 ;
  assign n10489 = n10444 ^ n10370 ;
  assign n10492 = n10491 ^ n10489 ;
  assign n10500 = ~n2924 & n10131 ;
  assign n10496 = n10491 ^ x5 ;
  assign n10495 = ~n3099 & ~n9092 ;
  assign n10497 = n10496 ^ n10495 ;
  assign n10494 = n6344 & n9081 ;
  assign n10498 = n10497 ^ n10494 ;
  assign n10493 = ~n2958 & n9085 ;
  assign n10499 = n10498 ^ n10493 ;
  assign n10501 = n10500 ^ n10499 ;
  assign n10502 = n10492 & n10501 ;
  assign n10503 = n10502 ^ n10491 ;
  assign n10504 = n10503 ^ n10332 ;
  assign n10505 = n10334 & n10504 ;
  assign n10506 = n10505 ^ n10332 ;
  assign n10515 = n10514 ^ n10506 ;
  assign n10519 = ~n3337 & n6648 ;
  assign n10516 = n9813 ^ x8 ;
  assign n10517 = n10516 ^ n9795 ;
  assign n10518 = n10517 ^ n10514 ;
  assign n10520 = n10519 ^ n10518 ;
  assign n10521 = n10515 & n10520 ;
  assign n10522 = n10521 ^ n10514 ;
  assign n10523 = n10522 ^ n10322 ;
  assign n10524 = n10324 & n10523 ;
  assign n10525 = n10524 ^ n10322 ;
  assign n10527 = n10526 ^ n10525 ;
  assign n10535 = n5650 & n9081 ;
  assign n10531 = n10526 ^ x5 ;
  assign n10530 = ~n2738 & n9085 ;
  assign n10532 = n10531 ^ n10530 ;
  assign n10529 = ~n2836 & ~n9092 ;
  assign n10533 = n10532 ^ n10529 ;
  assign n10528 = ~n2646 & n9077 ;
  assign n10534 = n10533 ^ n10528 ;
  assign n10536 = n10535 ^ n10534 ;
  assign n10537 = n10527 & n10536 ;
  assign n10538 = n10537 ^ n10526 ;
  assign n10539 = n10538 ^ n10309 ;
  assign n10540 = n10314 & n10539 ;
  assign n10541 = n10540 ^ n10309 ;
  assign n10542 = n10541 ^ n10295 ;
  assign n10543 = n10301 & n10542 ;
  assign n10544 = n10543 ^ n10295 ;
  assign n10546 = n10545 ^ n10544 ;
  assign n10553 = n5541 & n9081 ;
  assign n10551 = ~n2609 & n9085 ;
  assign n10549 = ~n3227 & ~n9092 ;
  assign n10548 = n10545 ^ x5 ;
  assign n10550 = n10549 ^ n10548 ;
  assign n10552 = n10551 ^ n10550 ;
  assign n10554 = n10553 ^ n10552 ;
  assign n10547 = ~n2554 & n10131 ;
  assign n10555 = n10554 ^ n10547 ;
  assign n10556 = n10546 & n10555 ;
  assign n10557 = n10556 ^ n10545 ;
  assign n10558 = n10557 ^ n10283 ;
  assign n10559 = ~n10291 & ~n10558 ;
  assign n10560 = n10559 ^ n10283 ;
  assign n10562 = n10561 ^ n10560 ;
  assign n10569 = n5520 & n9081 ;
  assign n10567 = ~n2554 & ~n9092 ;
  assign n10565 = ~n2486 & n9085 ;
  assign n10564 = n10561 ^ x5 ;
  assign n10566 = n10565 ^ n10564 ;
  assign n10568 = n10567 ^ n10566 ;
  assign n10570 = n10569 ^ n10568 ;
  assign n10563 = ~n2449 & n10131 ;
  assign n10571 = n10570 ^ n10563 ;
  assign n10572 = n10562 & ~n10571 ;
  assign n10573 = n10572 ^ n10561 ;
  assign n10574 = n10573 ^ n10273 ;
  assign n10575 = n10281 & ~n10574 ;
  assign n10576 = n10575 ^ n10273 ;
  assign n10578 = n10577 ^ n10576 ;
  assign n10585 = n5144 & n9081 ;
  assign n10583 = ~n2268 & n10131 ;
  assign n10581 = ~n2364 & n9085 ;
  assign n10580 = n10577 ^ x5 ;
  assign n10582 = n10581 ^ n10580 ;
  assign n10584 = n10583 ^ n10582 ;
  assign n10586 = n10585 ^ n10584 ;
  assign n10579 = ~n2449 & ~n9092 ;
  assign n10587 = n10586 ^ n10579 ;
  assign n10588 = n10578 & n10587 ;
  assign n10589 = n10588 ^ n10577 ;
  assign n10590 = n10589 ^ n10265 ;
  assign n10591 = n10271 & n10590 ;
  assign n10592 = n10591 ^ n10265 ;
  assign n10594 = n10593 ^ n10592 ;
  assign n10601 = n5196 & n9081 ;
  assign n10599 = ~n2268 & ~n9092 ;
  assign n10597 = ~n2185 & n9085 ;
  assign n10596 = n10593 ^ x5 ;
  assign n10598 = n10597 ^ n10596 ;
  assign n10600 = n10599 ^ n10598 ;
  assign n10602 = n10601 ^ n10600 ;
  assign n10595 = ~n2096 & n10131 ;
  assign n10603 = n10602 ^ n10595 ;
  assign n10604 = n10594 & n10603 ;
  assign n10605 = n10604 ^ n10593 ;
  assign n10606 = n10605 ^ n10259 ;
  assign n10607 = ~n10261 & ~n10606 ;
  assign n10608 = n10607 ^ n10260 ;
  assign n10609 = n10608 ^ n10245 ;
  assign n10610 = n10251 & ~n10609 ;
  assign n10611 = n10610 ^ n10245 ;
  assign n10612 = n10611 ^ n10239 ;
  assign n10613 = ~n10241 & ~n10612 ;
  assign n10614 = n10613 ^ n10240 ;
  assign n10615 = n10614 ^ n10229 ;
  assign n10616 = n10231 & n10615 ;
  assign n10617 = n10616 ^ n10230 ;
  assign n10618 = n10617 ^ n10207 ;
  assign n10619 = ~n10219 & n10618 ;
  assign n10620 = n10619 ^ n10218 ;
  assign n10621 = n10620 ^ n10204 ;
  assign n10622 = ~n10206 & n10621 ;
  assign n10623 = n10622 ^ n10204 ;
  assign n10624 = n10623 ^ n10191 ;
  assign n10625 = ~n10196 & ~n10624 ;
  assign n10626 = n10625 ^ n10191 ;
  assign n10627 = n10018 ^ n9652 ;
  assign n10632 = ~n10626 & n10627 ;
  assign n10633 = n10632 ^ n10627 ;
  assign n10178 = ~n1433 & n9085 ;
  assign n10177 = ~n4610 & n9081 ;
  assign n10179 = n10178 ^ n10177 ;
  assign n10180 = n10179 ^ x5 ;
  assign n10176 = ~n1351 & ~n9092 ;
  assign n10181 = n10180 ^ n10176 ;
  assign n10175 = ~n1540 & n10131 ;
  assign n10182 = n10181 ^ n10175 ;
  assign n10628 = n10627 ^ n10626 ;
  assign n10630 = ~n10182 & n10628 ;
  assign n10629 = n10628 ^ n10182 ;
  assign n10631 = n10630 ^ n10629 ;
  assign n10634 = n10633 ^ n10631 ;
  assign n10635 = n10634 ^ n10627 ;
  assign n10174 = n10034 ^ n10021 ;
  assign n10636 = n10635 ^ n10174 ;
  assign n10645 = n10174 ^ x5 ;
  assign n10644 = ~n1433 & ~n9092 ;
  assign n10646 = n10645 ^ n10644 ;
  assign n10643 = ~n1540 & n9085 ;
  assign n10647 = n10646 ^ n10643 ;
  assign n10637 = n4603 ^ n1214 ;
  assign n10640 = ~n9089 & n10637 ;
  assign n10641 = n10640 ^ n4603 ;
  assign n10642 = n9077 & ~n10641 ;
  assign n10648 = n10647 ^ n10642 ;
  assign n10649 = n10636 & ~n10648 ;
  assign n10650 = n10649 ^ n10635 ;
  assign n10652 = n10651 ^ n10650 ;
  assign n10661 = ~n1540 & ~n9092 ;
  assign n10659 = n10651 ^ x5 ;
  assign n10656 = ~n3381 & n9089 ;
  assign n10657 = n10656 ^ n968 ;
  assign n10658 = n9077 & ~n10657 ;
  assign n10660 = n10659 ^ n10658 ;
  assign n10662 = n10661 ^ n10660 ;
  assign n10653 = ~n1214 & n9085 ;
  assign n10663 = n10662 ^ n10653 ;
  assign n10664 = n10652 & n10663 ;
  assign n10665 = n10664 ^ n10651 ;
  assign n10667 = n10666 ^ n10665 ;
  assign n10674 = n3905 & n9081 ;
  assign n10672 = ~n968 & n9085 ;
  assign n10670 = ~n1214 & ~n9092 ;
  assign n10669 = n10666 ^ x5 ;
  assign n10671 = n10670 ^ n10669 ;
  assign n10673 = n10672 ^ n10671 ;
  assign n10675 = n10674 ^ n10673 ;
  assign n10668 = ~n1109 & n10131 ;
  assign n10676 = n10675 ^ n10668 ;
  assign n10677 = n10667 & n10676 ;
  assign n10678 = n10677 ^ n10666 ;
  assign n10679 = n10678 ^ n10168 ;
  assign n10680 = n10173 & n10679 ;
  assign n10681 = n10680 ^ n10168 ;
  assign n10682 = n10681 ^ n10155 ;
  assign n10683 = n10160 & n10682 ;
  assign n10684 = n10683 ^ n10155 ;
  assign n10696 = n10684 ^ n10144 ;
  assign n10147 = n10069 ^ n9620 ;
  assign n10685 = n10684 ^ n10147 ;
  assign n10692 = ~n3473 & n9085 ;
  assign n10690 = ~n824 & ~n9092 ;
  assign n10688 = ~n3476 & n9081 ;
  assign n10687 = n10147 ^ x5 ;
  assign n10689 = n10688 ^ n10687 ;
  assign n10691 = n10690 ^ n10689 ;
  assign n10693 = n10692 ^ n10691 ;
  assign n10686 = ~n649 & n10131 ;
  assign n10694 = n10693 ^ n10686 ;
  assign n10695 = ~n10685 & n10694 ;
  assign n10697 = n10696 ^ n10695 ;
  assign n10698 = ~n10146 & ~n10697 ;
  assign n10699 = n10698 ^ n10145 ;
  assign n10700 = n10136 & ~n10699 ;
  assign n10702 = x0 & x2 ;
  assign n10726 = n3923 & n3943 ;
  assign n10727 = x1 & x2 ;
  assign n10728 = x0 & x1 ;
  assign n10729 = ~n10727 & n10728 ;
  assign n10730 = n10726 & n10729 ;
  assign n10703 = n3943 ^ x2 ;
  assign n10704 = n10703 ^ x1 ;
  assign n10705 = n10704 ^ x0 ;
  assign n10712 = n10705 ^ n10703 ;
  assign n10713 = x2 ^ x0 ;
  assign n10716 = ~n10712 & ~n10713 ;
  assign n10717 = n10716 ^ x0 ;
  assign n10718 = n10703 ^ n485 ;
  assign n10719 = n10716 ^ n10712 ;
  assign n10720 = ~n10718 & ~n10719 ;
  assign n10721 = n10720 ^ n485 ;
  assign n10722 = n10721 ^ n10718 ;
  assign n10723 = n10717 & ~n10722 ;
  assign n10724 = n10723 ^ n10720 ;
  assign n10725 = n10724 ^ n10703 ;
  assign n10731 = n10730 ^ n10725 ;
  assign n10732 = n10702 & n10731 ;
  assign n10735 = n3922 & ~n3943 ;
  assign n10736 = n10735 ^ n3921 ;
  assign n10737 = n10732 & ~n10736 ;
  assign n10738 = n10737 ^ n10731 ;
  assign n10739 = n485 & n10738 ;
  assign n10743 = ~n3943 & n10728 ;
  assign n10746 = ~n3921 & n10743 ;
  assign n10740 = x2 & n3943 ;
  assign n10747 = n10746 ^ n10740 ;
  assign n10748 = n10739 & n10747 ;
  assign n10749 = n10748 ^ n10738 ;
  assign n10701 = n10074 ^ n9599 ;
  assign n10768 = n10749 ^ n10701 ;
  assign n10760 = ~n10727 & ~n10740 ;
  assign n10761 = n10743 ^ n10702 ;
  assign n10762 = ~n3920 & n10761 ;
  assign n10763 = n10762 ^ n10702 ;
  assign n10764 = n10760 & ~n10763 ;
  assign n10758 = ~n445 & n9085 ;
  assign n10756 = n3500 & n9081 ;
  assign n10753 = ~n485 & n10131 ;
  assign n10752 = ~n317 & ~n9092 ;
  assign n10754 = n10753 ^ n10752 ;
  assign n10755 = n10754 ^ x5 ;
  assign n10757 = n10756 ^ n10755 ;
  assign n10759 = n10758 ^ n10757 ;
  assign n10765 = n10764 ^ n10759 ;
  assign n10751 = n10077 ^ n9589 ;
  assign n10766 = n10765 ^ n10751 ;
  assign n10750 = ~n10701 & ~n10749 ;
  assign n10767 = n10766 ^ n10750 ;
  assign n10769 = n10768 ^ n10767 ;
  assign n10770 = ~n10700 & ~n10769 ;
  assign n10782 = x2 & ~n445 ;
  assign n10783 = n10782 ^ n485 ;
  assign n10784 = ~x1 & ~n10783 ;
  assign n10778 = n485 ^ x2 ;
  assign n10772 = n3943 ^ x1 ;
  assign n10773 = n10772 ^ n10703 ;
  assign n10774 = n3924 & n10773 ;
  assign n10775 = n10774 ^ n10772 ;
  assign n10779 = n10778 ^ n10775 ;
  assign n10785 = n10784 ^ n10779 ;
  assign n10786 = ~x0 & n10785 ;
  assign n10787 = n10786 ^ n10775 ;
  assign n10771 = n10697 ^ n10145 ;
  assign n10788 = n10787 ^ n10771 ;
  assign n10803 = x2 & ~n649 ;
  assign n10804 = n10803 ^ n317 ;
  assign n10805 = ~x1 & ~n10804 ;
  assign n10799 = n317 ^ x2 ;
  assign n10791 = n445 ^ x1 ;
  assign n10790 = n445 ^ x2 ;
  assign n10792 = n10791 ^ n10790 ;
  assign n10793 = n4072 & n10792 ;
  assign n10794 = n10793 ^ n10791 ;
  assign n10800 = n10799 ^ n10794 ;
  assign n10806 = n10805 ^ n10800 ;
  assign n10807 = ~x0 & n10806 ;
  assign n10795 = n10681 ^ n10160 ;
  assign n10796 = n10795 ^ n10794 ;
  assign n10808 = n10807 ^ n10796 ;
  assign n10821 = x2 & ~n3473 ;
  assign n10822 = n10821 ^ n649 ;
  assign n10823 = ~x1 & ~n10822 ;
  assign n10817 = n649 ^ x2 ;
  assign n10809 = n317 ^ x1 ;
  assign n10810 = n10809 ^ n10799 ;
  assign n10811 = n3955 & n10810 ;
  assign n10812 = n10811 ^ n10809 ;
  assign n10818 = n10817 ^ n10812 ;
  assign n10824 = n10823 ^ n10818 ;
  assign n10825 = ~x0 & n10824 ;
  assign n10813 = n10678 ^ n10173 ;
  assign n10814 = n10813 ^ n10812 ;
  assign n10826 = n10825 ^ n10814 ;
  assign n10840 = n10676 ^ n10665 ;
  assign n10828 = x2 ^ x1 ;
  assign n10829 = n3475 & n10828 ;
  assign n10830 = n10829 ^ n10817 ;
  assign n10841 = n10840 ^ n10830 ;
  assign n10832 = n3473 ^ x2 ;
  assign n10833 = n10832 ^ n10830 ;
  assign n10827 = x2 & n824 ;
  assign n10831 = n10830 ^ n10827 ;
  assign n10834 = n10833 ^ n10831 ;
  assign n10835 = n10831 ^ x1 ;
  assign n10836 = n10835 ^ n10831 ;
  assign n10837 = ~n10834 & n10836 ;
  assign n10838 = n10837 ^ n10831 ;
  assign n10839 = ~x0 & ~n10838 ;
  assign n10842 = n10841 ^ n10839 ;
  assign n11408 = n10631 & n10648 ;
  assign n10881 = x2 & ~n1433 ;
  assign n10882 = n10881 ^ n1540 ;
  assign n10883 = ~x1 & ~n10882 ;
  assign n10877 = n1540 ^ x2 ;
  assign n10873 = n3376 & n10828 ;
  assign n10866 = n1214 ^ x2 ;
  assign n10874 = n10873 ^ n10866 ;
  assign n10878 = n10877 ^ n10874 ;
  assign n10884 = n10883 ^ n10878 ;
  assign n10885 = ~x0 & n10884 ;
  assign n10871 = n10620 ^ n10206 ;
  assign n10875 = n10874 ^ n10871 ;
  assign n10886 = n10885 ^ n10875 ;
  assign n10899 = x2 & ~n1351 ;
  assign n10900 = n10899 ^ n1433 ;
  assign n10901 = ~x1 & ~n10900 ;
  assign n10895 = n1433 ^ x2 ;
  assign n10889 = n1540 ^ x1 ;
  assign n10890 = n10889 ^ n10877 ;
  assign n10891 = ~n3817 & n10890 ;
  assign n10892 = n10891 ^ n10889 ;
  assign n10896 = n10895 ^ n10892 ;
  assign n10902 = n10901 ^ n10896 ;
  assign n10903 = ~x0 & n10902 ;
  assign n10887 = n10617 ^ n10219 ;
  assign n10893 = n10892 ^ n10887 ;
  assign n10904 = n10903 ^ n10893 ;
  assign n11360 = x2 & n1703 ;
  assign n11353 = ~x2 & n3815 ;
  assign n11354 = n11353 ^ n3815 ;
  assign n11355 = n11354 ^ n1433 ;
  assign n11361 = n11360 ^ n11355 ;
  assign n11362 = ~x0 & ~n11361 ;
  assign n11363 = n11362 ^ n11355 ;
  assign n10906 = n1351 ^ x2 ;
  assign n11364 = n11363 ^ n10906 ;
  assign n11365 = n11364 ^ n1433 ;
  assign n11366 = n11365 ^ n11353 ;
  assign n11367 = n11366 ^ n11363 ;
  assign n11368 = x0 & ~n11367 ;
  assign n11369 = n11368 ^ n11364 ;
  assign n11370 = x1 & n11369 ;
  assign n11371 = n11370 ^ n11363 ;
  assign n11381 = n11371 ^ n10887 ;
  assign n10910 = n1703 ^ n1631 ;
  assign n10911 = n10910 ^ n1703 ;
  assign n10916 = x2 & ~n10911 ;
  assign n10917 = n10916 ^ n1703 ;
  assign n10918 = ~x1 & ~n10917 ;
  assign n10912 = n1703 ^ x2 ;
  assign n10907 = ~n4416 & n10828 ;
  assign n10908 = n10907 ^ n10906 ;
  assign n10913 = n10912 ^ n10908 ;
  assign n10919 = n10918 ^ n10913 ;
  assign n10920 = ~x0 & n10919 ;
  assign n10905 = n10611 ^ n10241 ;
  assign n10909 = n10908 ^ n10905 ;
  assign n10921 = n10920 ^ n10909 ;
  assign n11372 = n11371 ^ n10905 ;
  assign n11373 = n11372 ^ n11371 ;
  assign n10934 = x2 & ~n1871 ;
  assign n10935 = n10934 ^ n1631 ;
  assign n10936 = ~x1 & ~n10935 ;
  assign n10930 = n1631 ^ x2 ;
  assign n10922 = n1703 ^ x1 ;
  assign n10923 = n10922 ^ n10912 ;
  assign n10924 = ~n3808 & n10923 ;
  assign n10925 = n10924 ^ n10922 ;
  assign n10931 = n10930 ^ n10925 ;
  assign n10937 = n10936 ^ n10931 ;
  assign n10938 = ~x0 & n10937 ;
  assign n10926 = n10608 ^ n10251 ;
  assign n10927 = n10926 ^ n10925 ;
  assign n10939 = n10938 ^ n10927 ;
  assign n10944 = n10605 ^ n10261 ;
  assign n11349 = n10944 ^ n10926 ;
  assign n10950 = x2 & ~n1795 ;
  assign n10951 = n10950 ^ n1871 ;
  assign n10952 = ~x1 & ~n10951 ;
  assign n10946 = n1871 ^ x2 ;
  assign n10940 = n1631 ^ x1 ;
  assign n10941 = n10940 ^ n10930 ;
  assign n10942 = ~n4391 & n10941 ;
  assign n10943 = n10942 ^ n10940 ;
  assign n10947 = n10946 ^ n10943 ;
  assign n10953 = n10952 ^ n10947 ;
  assign n10954 = ~x0 & n10953 ;
  assign n10945 = n10944 ^ n10943 ;
  assign n10955 = n10954 ^ n10945 ;
  assign n10853 = ~x1 & x2 ;
  assign n10854 = ~x0 & n10853 ;
  assign n10966 = n1994 & n10854 ;
  assign n10964 = n1795 ^ x2 ;
  assign n10965 = n10850 & ~n10964 ;
  assign n10967 = n10966 ^ n10965 ;
  assign n10963 = n10603 ^ n10592 ;
  assign n10968 = n10967 ^ n10963 ;
  assign n10960 = n4858 & n10828 ;
  assign n10961 = n10960 ^ n10946 ;
  assign n10962 = x0 & ~n10961 ;
  assign n10969 = n10968 ^ n10962 ;
  assign n10972 = n10589 ^ n10271 ;
  assign n11343 = n10972 ^ n10963 ;
  assign n10980 = x2 & ~n2096 ;
  assign n10981 = n10980 ^ n1994 ;
  assign n10982 = ~x1 & ~n10981 ;
  assign n10976 = n1994 ^ x2 ;
  assign n10970 = ~n4384 & n10828 ;
  assign n10971 = n10970 ^ n10964 ;
  assign n10977 = n10976 ^ n10971 ;
  assign n10983 = n10982 ^ n10977 ;
  assign n10984 = ~x0 & n10983 ;
  assign n10973 = n10972 ^ n10971 ;
  assign n10985 = n10984 ^ n10973 ;
  assign n10997 = n10587 ^ n10576 ;
  assign n11340 = n10997 ^ n10972 ;
  assign n10995 = n2185 & n10854 ;
  assign n10993 = n2096 ^ x2 ;
  assign n10994 = n10850 & ~n10993 ;
  assign n10996 = n10995 ^ n10994 ;
  assign n10998 = n10997 ^ n10996 ;
  assign n10988 = n10976 ^ n10828 ;
  assign n10989 = n10988 ^ n10976 ;
  assign n10990 = ~n5408 & n10989 ;
  assign n10991 = n10990 ^ n10976 ;
  assign n10992 = x0 & ~n10991 ;
  assign n10999 = n10998 ^ n10992 ;
  assign n11004 = n10573 ^ n10281 ;
  assign n11337 = n11004 ^ n10997 ;
  assign n11012 = x2 & ~n2268 ;
  assign n11013 = n11012 ^ n2185 ;
  assign n11014 = ~x1 & ~n11013 ;
  assign n11008 = n2185 ^ x2 ;
  assign n11000 = n2096 ^ x1 ;
  assign n11001 = n11000 ^ n10993 ;
  assign n11002 = n5195 & n11001 ;
  assign n11003 = n11002 ^ n11000 ;
  assign n11009 = n11008 ^ n11003 ;
  assign n11015 = n11014 ^ n11009 ;
  assign n11016 = ~x0 & n11015 ;
  assign n11005 = n11004 ^ n11003 ;
  assign n11017 = n11016 ^ n11005 ;
  assign n11022 = n10571 ^ n10560 ;
  assign n11334 = n11022 ^ n11004 ;
  assign n11030 = x2 & ~n2364 ;
  assign n11031 = n11030 ^ n2268 ;
  assign n11032 = ~x1 & ~n11031 ;
  assign n11026 = n2268 ^ x2 ;
  assign n11018 = n2185 ^ x1 ;
  assign n11019 = n11018 ^ n11008 ;
  assign n11020 = n4930 & n11019 ;
  assign n11021 = n11020 ^ n11018 ;
  assign n11027 = n11026 ^ n11021 ;
  assign n11033 = n11032 ^ n11027 ;
  assign n11034 = ~x0 & n11033 ;
  assign n11023 = n11022 ^ n11021 ;
  assign n11035 = n11034 ^ n11023 ;
  assign n11043 = x2 & n2449 ;
  assign n11037 = n2268 ^ x1 ;
  assign n11038 = n11037 ^ n11026 ;
  assign n11039 = n5143 & n11038 ;
  assign n11040 = n11039 ^ n11037 ;
  assign n11044 = n11043 ^ n11040 ;
  assign n11041 = n2364 ^ x2 ;
  assign n11042 = n11041 ^ n11040 ;
  assign n11045 = n11044 ^ n11042 ;
  assign n11046 = n11044 ^ x1 ;
  assign n11047 = n11046 ^ n11044 ;
  assign n11048 = ~n11045 & n11047 ;
  assign n11049 = n11048 ^ n11044 ;
  assign n11050 = ~x0 & ~n11049 ;
  assign n11051 = n11050 ^ n11040 ;
  assign n11331 = n11051 ^ n11022 ;
  assign n11062 = x2 & ~n2486 ;
  assign n11063 = n11062 ^ n2449 ;
  assign n11064 = ~x1 & ~n11063 ;
  assign n11058 = n2449 ^ x2 ;
  assign n11053 = ~n5282 & n10828 ;
  assign n11054 = n11053 ^ n11041 ;
  assign n11059 = n11058 ^ n11054 ;
  assign n11065 = n11064 ^ n11059 ;
  assign n11066 = ~x0 & n11065 ;
  assign n11036 = n10555 ^ n10544 ;
  assign n11055 = n11054 ^ n11036 ;
  assign n11067 = n11066 ^ n11055 ;
  assign n11081 = x2 & ~n2554 ;
  assign n11082 = n11081 ^ n2486 ;
  assign n11083 = ~x1 & ~n11082 ;
  assign n11077 = n2486 ^ x2 ;
  assign n11070 = n2449 ^ x1 ;
  assign n11071 = n11070 ^ n11058 ;
  assign n11072 = n5519 & n11071 ;
  assign n11073 = n11072 ^ n11070 ;
  assign n11078 = n11077 ^ n11073 ;
  assign n11084 = n11083 ^ n11078 ;
  assign n11085 = ~x0 & n11084 ;
  assign n11068 = n10541 ^ n10301 ;
  assign n11074 = n11073 ^ n11068 ;
  assign n11086 = n11085 ^ n11074 ;
  assign n11091 = n10538 ^ n10314 ;
  assign n11322 = n11091 ^ n11068 ;
  assign n11093 = n2609 ^ n2554 ;
  assign n11094 = n11093 ^ n2554 ;
  assign n11099 = x2 & ~n11094 ;
  assign n11100 = n11099 ^ n2554 ;
  assign n11101 = ~x1 & ~n11100 ;
  assign n11095 = n2554 ^ x2 ;
  assign n11087 = n2486 ^ x1 ;
  assign n11088 = n11087 ^ n11077 ;
  assign n11089 = n5380 & n11088 ;
  assign n11090 = n11089 ^ n11087 ;
  assign n11096 = n11095 ^ n11090 ;
  assign n11102 = n11101 ^ n11096 ;
  assign n11103 = ~x0 & n11102 ;
  assign n11092 = n11091 ^ n11090 ;
  assign n11104 = n11103 ^ n11092 ;
  assign n11109 = n10536 ^ n10525 ;
  assign n11319 = n11109 ^ n11091 ;
  assign n11117 = x2 & ~n3227 ;
  assign n11118 = n11117 ^ n2609 ;
  assign n11119 = ~x1 & ~n11118 ;
  assign n11113 = n2609 ^ x2 ;
  assign n11105 = n2554 ^ x1 ;
  assign n11106 = n11105 ^ n11095 ;
  assign n11107 = n5540 & n11106 ;
  assign n11108 = n11107 ^ n11105 ;
  assign n11114 = n11113 ^ n11108 ;
  assign n11120 = n11119 ^ n11114 ;
  assign n11121 = ~x0 & n11120 ;
  assign n11110 = n11109 ^ n11108 ;
  assign n11122 = n11121 ^ n11110 ;
  assign n11292 = n2609 ^ x1 ;
  assign n11293 = n11292 ^ n11113 ;
  assign n11294 = n6171 & n11293 ;
  assign n11295 = n11294 ^ n11292 ;
  assign n11270 = n3227 ^ x2 ;
  assign n11298 = n11295 ^ n11270 ;
  assign n11299 = n11298 ^ n11295 ;
  assign n11300 = n11299 ^ n3227 ;
  assign n11301 = ~n2646 & n11300 ;
  assign n11302 = n11301 ^ n3227 ;
  assign n11303 = ~x1 & ~n11302 ;
  assign n11304 = n11303 ^ n11298 ;
  assign n11305 = ~x0 & n11304 ;
  assign n11306 = n11305 ^ n11295 ;
  assign n11316 = n11306 ^ n11109 ;
  assign n11154 = n2836 ^ x2 ;
  assign n11148 = x2 & n3151 ;
  assign n11142 = x2 & ~n3347 ;
  assign n11143 = n11142 ^ n2738 ;
  assign n11149 = n11148 ^ n11143 ;
  assign n11150 = ~x0 & ~n11149 ;
  assign n11151 = n11150 ^ n11143 ;
  assign n11157 = n11154 ^ n11151 ;
  assign n11153 = n11142 ^ n6907 ;
  assign n11155 = n11154 ^ n11153 ;
  assign n11156 = x0 & n11155 ;
  assign n11158 = n11157 ^ n11156 ;
  assign n11159 = x1 & n11158 ;
  assign n11140 = n10501 ^ n10489 ;
  assign n11152 = n11151 ^ n11140 ;
  assign n11160 = n11159 ^ n11152 ;
  assign n11176 = ~x1 & ~n3345 ;
  assign n11177 = n11176 ^ n2836 ;
  assign n11161 = n10359 ^ x5 ;
  assign n11162 = n11161 ^ n10352 ;
  assign n11163 = n11162 ^ x6 ;
  assign n11164 = n11163 ^ n10359 ;
  assign n11165 = n11164 ^ n10352 ;
  assign n11166 = ~n3337 & n11165 ;
  assign n11167 = n11166 ^ n11162 ;
  assign n11186 = n11177 ^ n11167 ;
  assign n11179 = n11177 ^ n2924 ;
  assign n11178 = n11177 ^ n3151 ;
  assign n11180 = n11179 ^ n11178 ;
  assign n11183 = x1 & n11180 ;
  assign n11184 = n11183 ^ n11179 ;
  assign n11185 = ~x0 & n11184 ;
  assign n11187 = n11186 ^ n11185 ;
  assign n11169 = n3345 ^ x0 ;
  assign n11170 = n11169 ^ n3345 ;
  assign n11171 = ~x1 & ~n2924 ;
  assign n11172 = n11171 ^ n3345 ;
  assign n11173 = ~n11170 & ~n11172 ;
  assign n11174 = n11173 ^ n3345 ;
  assign n11175 = ~x2 & n11174 ;
  assign n11188 = n11187 ^ n11175 ;
  assign n11219 = x2 & ~n3099 ;
  assign n11220 = n11219 ^ n2958 ;
  assign n11221 = ~x1 & ~n11220 ;
  assign n11215 = n2958 ^ x2 ;
  assign n11210 = n2924 ^ x1 ;
  assign n11196 = n2924 ^ x2 ;
  assign n11211 = n11210 ^ n11196 ;
  assign n11212 = n6343 & n11211 ;
  assign n11213 = n11212 ^ n11210 ;
  assign n11216 = n11215 ^ n11213 ;
  assign n11222 = n11221 ^ n11216 ;
  assign n11223 = ~x0 & n11222 ;
  assign n11206 = n9084 ^ x4 ;
  assign n11207 = ~n3337 & n11206 ;
  assign n11208 = n11207 ^ n10335 ;
  assign n11214 = n11213 ^ n11208 ;
  assign n11224 = n11223 ^ n11214 ;
  assign n11239 = x2 & n3027 ;
  assign n11240 = ~x0 & ~x1 ;
  assign n11241 = n11240 ^ n3337 ;
  assign n11229 = n3099 ^ x3 ;
  assign n11244 = n11229 & n11240 ;
  assign n11245 = n11244 ^ n3099 ;
  assign n11246 = n11241 & ~n11245 ;
  assign n11247 = n11246 ^ n3337 ;
  assign n11248 = n11239 & n11247 ;
  assign n11225 = ~x0 & n9077 ;
  assign n11234 = n11225 & n11229 ;
  assign n11235 = x1 & n11234 ;
  assign n11236 = n11235 ^ x1 ;
  assign n11226 = n11225 ^ n9077 ;
  assign n11227 = n11226 ^ x1 ;
  assign n11237 = n11236 ^ n11227 ;
  assign n11238 = ~n3337 & n11237 ;
  assign n11249 = n11248 ^ n11238 ;
  assign n11256 = n11249 ^ n11208 ;
  assign n11250 = x0 & n11249 ;
  assign n11251 = n2958 ^ x1 ;
  assign n11252 = n11251 ^ n11215 ;
  assign n11253 = n6439 & n11252 ;
  assign n11254 = n11253 ^ n11251 ;
  assign n11255 = n11250 & n11254 ;
  assign n11257 = n11256 ^ n11255 ;
  assign n11258 = ~n11224 & n11257 ;
  assign n11200 = x2 & ~n2958 ;
  assign n11201 = n11200 ^ n2924 ;
  assign n11202 = ~x1 & ~n11201 ;
  assign n11190 = n3151 ^ x1 ;
  assign n11189 = n3151 ^ x2 ;
  assign n11191 = n11190 ^ n11189 ;
  assign n11192 = n6282 & n11191 ;
  assign n11193 = n11192 ^ n11190 ;
  assign n11197 = n11196 ^ n11193 ;
  assign n11203 = n11202 ^ n11197 ;
  assign n11204 = ~x0 & n11203 ;
  assign n11205 = n11204 ^ n11193 ;
  assign n11209 = n11208 ^ n11205 ;
  assign n11259 = n11258 ^ n11209 ;
  assign n11260 = n11205 ^ n11167 ;
  assign n11261 = n11260 ^ n10351 ;
  assign n11262 = n11261 ^ n10339 ;
  assign n11263 = n11262 ^ n11167 ;
  assign n11264 = ~n11259 & ~n11263 ;
  assign n11265 = n11264 ^ n11260 ;
  assign n11266 = n11188 & ~n11265 ;
  assign n11168 = n11167 ^ n11140 ;
  assign n11267 = n11266 ^ n11168 ;
  assign n11268 = ~n11160 & n11267 ;
  assign n11134 = x2 & ~n2836 ;
  assign n11135 = n11134 ^ n2738 ;
  assign n11136 = ~x1 & ~n11135 ;
  assign n11130 = n2738 ^ x2 ;
  assign n11124 = n2646 ^ x2 ;
  assign n11123 = n2646 ^ x1 ;
  assign n11125 = n11124 ^ n11123 ;
  assign n11126 = ~n5650 & n11125 ;
  assign n11127 = n11126 ^ n11123 ;
  assign n11131 = n11130 ^ n11127 ;
  assign n11137 = n11136 ^ n11131 ;
  assign n11138 = ~x0 & n11137 ;
  assign n11139 = n11138 ^ n11127 ;
  assign n11141 = n11140 ^ n11139 ;
  assign n11269 = n11268 ^ n11141 ;
  assign n11271 = n3227 ^ x1 ;
  assign n11272 = n11271 ^ n11270 ;
  assign n11273 = n6176 & n11272 ;
  assign n11274 = n11273 ^ n11271 ;
  assign n11277 = n11274 ^ n11124 ;
  assign n11278 = n11277 ^ n11274 ;
  assign n11279 = n11278 ^ n2646 ;
  assign n11280 = ~n2738 & n11279 ;
  assign n11281 = n11280 ^ n2646 ;
  assign n11282 = ~x1 & ~n11281 ;
  assign n11283 = n11282 ^ n11277 ;
  assign n11284 = ~x0 & n11283 ;
  assign n11285 = n11284 ^ n11274 ;
  assign n11286 = n11285 ^ n11139 ;
  assign n11287 = n11286 ^ n10334 ;
  assign n11288 = n11287 ^ n11285 ;
  assign n11289 = n11288 ^ n10503 ;
  assign n11290 = ~n11269 & ~n11289 ;
  assign n11291 = n11290 ^ n11286 ;
  assign n11307 = n11306 ^ n11285 ;
  assign n11308 = n11307 ^ n10520 ;
  assign n11309 = n11308 ^ n11306 ;
  assign n11310 = n11309 ^ n10506 ;
  assign n11311 = n11291 & ~n11310 ;
  assign n11312 = n11311 ^ n11307 ;
  assign n11313 = n11306 ^ n10522 ;
  assign n11314 = n11313 ^ n10324 ;
  assign n11315 = n11312 & ~n11314 ;
  assign n11317 = n11316 ^ n11315 ;
  assign n11318 = ~n11122 & ~n11317 ;
  assign n11320 = n11319 ^ n11318 ;
  assign n11321 = ~n11104 & n11320 ;
  assign n11323 = n11322 ^ n11321 ;
  assign n11324 = ~n11086 & n11323 ;
  assign n11069 = n11068 ^ n11036 ;
  assign n11325 = n11324 ^ n11069 ;
  assign n11326 = ~n11067 & n11325 ;
  assign n11052 = n11051 ^ n11036 ;
  assign n11327 = n11326 ^ n11052 ;
  assign n11328 = n11051 ^ n10291 ;
  assign n11329 = n11328 ^ n10557 ;
  assign n11330 = ~n11327 & n11329 ;
  assign n11332 = n11331 ^ n11330 ;
  assign n11333 = ~n11035 & ~n11332 ;
  assign n11335 = n11334 ^ n11333 ;
  assign n11336 = n11017 & ~n11335 ;
  assign n11338 = n11337 ^ n11336 ;
  assign n11339 = n10999 & ~n11338 ;
  assign n11341 = n11340 ^ n11339 ;
  assign n11342 = ~n10985 & n11341 ;
  assign n11344 = n11343 ^ n11342 ;
  assign n11345 = n10969 & n11344 ;
  assign n11346 = n11345 ^ n10963 ;
  assign n11347 = n11346 ^ n10944 ;
  assign n11348 = n10955 & ~n11347 ;
  assign n11350 = n11349 ^ n11348 ;
  assign n11351 = n10939 & n11350 ;
  assign n11352 = n11351 ^ n10926 ;
  assign n11374 = n11373 ^ n11352 ;
  assign n11375 = n10921 & n11374 ;
  assign n11376 = n11375 ^ n11372 ;
  assign n11377 = n11371 ^ n10230 ;
  assign n11378 = n11377 ^ n10229 ;
  assign n11379 = n11378 ^ n10614 ;
  assign n11380 = n11376 & n11379 ;
  assign n11382 = n11381 ^ n11380 ;
  assign n11383 = n10904 & n11382 ;
  assign n10888 = n10887 ^ n10871 ;
  assign n11384 = n11383 ^ n10888 ;
  assign n11385 = n10886 & n11384 ;
  assign n10868 = n1540 & n10854 ;
  assign n10867 = n10850 & ~n10866 ;
  assign n10869 = n10868 ^ n10867 ;
  assign n10863 = ~n3381 & n10828 ;
  assign n10858 = n968 ^ x2 ;
  assign n10864 = n10863 ^ n10858 ;
  assign n10865 = x0 & ~n10864 ;
  assign n10870 = n10869 ^ n10865 ;
  assign n10872 = n10871 ^ n10870 ;
  assign n11386 = n11385 ^ n10872 ;
  assign n11387 = n10870 ^ n10623 ;
  assign n11388 = n11387 ^ n10196 ;
  assign n11389 = ~n11386 & ~n11388 ;
  assign n11390 = n11389 ^ n10870 ;
  assign n11392 = n1109 ^ x1 ;
  assign n11391 = n1109 ^ x2 ;
  assign n11393 = n11392 ^ n11391 ;
  assign n11394 = n3904 & n11393 ;
  assign n11395 = n11394 ^ n11392 ;
  assign n11398 = n11395 ^ n10858 ;
  assign n11399 = n11398 ^ n11395 ;
  assign n11400 = n11399 ^ n968 ;
  assign n11401 = ~n1214 & n11400 ;
  assign n11402 = n11401 ^ n968 ;
  assign n11403 = ~x1 & ~n11402 ;
  assign n11404 = n11403 ^ n11398 ;
  assign n11405 = ~x0 & n11404 ;
  assign n11406 = n11405 ^ n11395 ;
  assign n11407 = n11390 & ~n11406 ;
  assign n11409 = n11408 ^ n11407 ;
  assign n11410 = n824 ^ x1 ;
  assign n10851 = n824 ^ x2 ;
  assign n11411 = n11410 ^ n10851 ;
  assign n11412 = ~n4044 & n11411 ;
  assign n11413 = n11412 ^ n11410 ;
  assign n11416 = n11413 ^ n11391 ;
  assign n11417 = n11416 ^ n11413 ;
  assign n11418 = n11417 ^ n1109 ;
  assign n11419 = ~n968 & n11418 ;
  assign n11420 = n11419 ^ n1109 ;
  assign n11421 = ~x1 & ~n11420 ;
  assign n11422 = n11421 ^ n11416 ;
  assign n11423 = ~x0 & n11422 ;
  assign n11424 = n11423 ^ n11413 ;
  assign n11425 = n11424 ^ n10632 ;
  assign n11426 = n11425 ^ n10648 ;
  assign n11427 = n11424 ^ n11407 ;
  assign n11428 = n11427 ^ n10630 ;
  assign n11429 = n11427 ^ n11424 ;
  assign n11430 = n11428 & ~n11429 ;
  assign n11431 = ~n11426 & n11430 ;
  assign n11432 = n11431 ^ n11427 ;
  assign n11433 = ~n11409 & n11432 ;
  assign n11434 = n11433 ^ n11408 ;
  assign n11435 = n11406 ^ n11390 ;
  assign n11436 = n11435 ^ n11407 ;
  assign n11437 = n11436 ^ n11424 ;
  assign n11438 = n11408 ^ n10635 ;
  assign n11439 = n11438 ^ n11436 ;
  assign n11440 = n11439 ^ n10648 ;
  assign n11441 = n11437 & n11440 ;
  assign n11442 = n11441 ^ n11424 ;
  assign n11443 = ~n11434 & ~n11442 ;
  assign n11448 = n11443 ^ n10840 ;
  assign n10855 = n1109 & n10854 ;
  assign n10852 = n10850 & ~n10851 ;
  assign n10856 = n10855 ^ n10852 ;
  assign n10847 = n3388 & n10828 ;
  assign n10848 = n10847 ^ n10832 ;
  assign n10849 = x0 & ~n10848 ;
  assign n10857 = n10856 ^ n10849 ;
  assign n11444 = n11443 ^ n10857 ;
  assign n11445 = n10857 ^ n10663 ;
  assign n11446 = n11445 ^ n10650 ;
  assign n11447 = n11444 & ~n11446 ;
  assign n11449 = n11448 ^ n11447 ;
  assign n11450 = ~n10842 & n11449 ;
  assign n11451 = n11450 ^ n10840 ;
  assign n11452 = n11451 ^ n10813 ;
  assign n11453 = ~n10826 & n11452 ;
  assign n11454 = n11453 ^ n10813 ;
  assign n11455 = n11454 ^ n10795 ;
  assign n11456 = ~n10808 & n11455 ;
  assign n11457 = n11456 ^ n10795 ;
  assign n11476 = n11457 ^ n10787 ;
  assign n10789 = n10694 ^ n10684 ;
  assign n11458 = n11457 ^ n10789 ;
  assign n11459 = n485 ^ x1 ;
  assign n11460 = n11459 ^ n10778 ;
  assign n11461 = n3499 & n11460 ;
  assign n11462 = n11461 ^ n11459 ;
  assign n11466 = n11462 ^ n10790 ;
  assign n11467 = n11466 ^ n11462 ;
  assign n11468 = n11467 ^ n445 ;
  assign n11469 = ~n317 & n11468 ;
  assign n11470 = n11469 ^ n445 ;
  assign n11471 = ~x1 & ~n11470 ;
  assign n11472 = n11471 ^ n11466 ;
  assign n11473 = ~x0 & n11472 ;
  assign n11463 = n11462 ^ n10789 ;
  assign n11474 = n11473 ^ n11463 ;
  assign n11475 = ~n11458 & ~n11474 ;
  assign n11477 = n11476 ^ n11475 ;
  assign n11478 = n10788 & ~n11477 ;
  assign n11479 = n11478 ^ n10787 ;
  assign n11480 = n10767 ^ n10766 ;
  assign n11481 = n10699 ^ n10136 ;
  assign n11482 = n11481 ^ n10700 ;
  assign n11485 = n11480 & n11482 ;
  assign n11486 = n11485 ^ n10767 ;
  assign n11487 = ~n11479 & ~n11486 ;
  assign n11488 = n10770 & ~n11487 ;
  assign n11489 = n11479 ^ n10749 ;
  assign n11490 = n10768 & ~n11489 ;
  assign n11491 = n11490 ^ n10701 ;
  assign n11492 = ~n10766 & ~n11482 ;
  assign n11493 = n11491 & n11492 ;
  assign n11494 = n11493 ^ n11491 ;
  assign n11495 = ~n11488 & ~n11494 ;
  assign n11497 = n11496 ^ n11495 ;
  assign n11500 = n11496 ^ n10759 ;
  assign n11498 = n10759 ^ n10751 ;
  assign n11499 = ~n10765 & n11498 ;
  assign n11501 = n11500 ^ n11499 ;
  assign n11502 = ~n11497 & ~n11501 ;
  assign n11503 = n11502 ^ n11496 ;
  assign n11504 = ~n10120 & n11503 ;
  assign n11505 = n11504 ^ n11503 ;
  assign n11506 = n11505 ^ n11503 ;
  assign n11507 = n11505 ^ n10109 ;
  assign n11508 = n11507 ^ n11505 ;
  assign n11509 = n11505 ^ n10116 ;
  assign n11510 = n11509 ^ n11505 ;
  assign n11511 = n11508 & ~n11510 ;
  assign n11512 = n11506 & n11511 ;
  assign n11513 = n11512 ^ n11506 ;
  assign n11514 = n11513 ^ n11503 ;
  assign n11515 = ~n10127 & ~n11514 ;
  assign n11532 = n11518 ^ n11515 ;
  assign n11533 = ~n11520 & ~n11532 ;
  assign n11535 = n11534 ^ n11533 ;
  assign n8395 = n8394 ^ n8051 ;
  assign n8396 = n8061 & n8395 ;
  assign n8397 = n8396 ^ n8394 ;
  assign n11536 = n11522 ^ n8397 ;
  assign n11537 = n11536 ^ n11522 ;
  assign n8404 = ~n485 & n7141 ;
  assign n8402 = n3944 & n7135 ;
  assign n8399 = ~n3943 & n8054 ;
  assign n8398 = ~n445 & n7146 ;
  assign n8400 = n8399 ^ n8398 ;
  assign n8401 = n8400 ^ x8 ;
  assign n8403 = n8402 ^ n8401 ;
  assign n8405 = n8404 ^ n8403 ;
  assign n11538 = n11522 ^ n8405 ;
  assign n11539 = n11538 ^ n11522 ;
  assign n11540 = ~n11537 & n11539 ;
  assign n11541 = n11540 ^ n11522 ;
  assign n11542 = ~n11535 & ~n11541 ;
  assign n11543 = n11542 ^ n8405 ;
  assign n8406 = n8405 ^ n8397 ;
  assign n11521 = n11520 ^ n11515 ;
  assign n11523 = n11522 ^ n11515 ;
  assign n11524 = n11523 ^ n11522 ;
  assign n11525 = n11522 ^ n11518 ;
  assign n11526 = n11525 ^ n11522 ;
  assign n11527 = n11524 & n11526 ;
  assign n11528 = n11527 ^ n11522 ;
  assign n11529 = ~n11521 & ~n11528 ;
  assign n11530 = n11529 ^ n8397 ;
  assign n11531 = ~n8406 & n11530 ;
  assign n11544 = n11543 ^ n11531 ;
  assign n11545 = n11544 ^ n8021 ;
  assign n11546 = n8049 & ~n11545 ;
  assign n11547 = n11546 ^ n8021 ;
  assign n7127 = n7124 ^ n7113 ;
  assign n11548 = n11547 ^ n7127 ;
  assign n11549 = ~n7126 & n11548 ;
  assign n11550 = n8047 ^ n8037 ;
  assign n11551 = n8039 & n11550 ;
  assign n11552 = n11551 ^ n8047 ;
  assign n11553 = n8030 ^ n8026 ;
  assign n11554 = ~n8036 & n11553 ;
  assign n11555 = n11554 ^ n8030 ;
  assign n11557 = n11552 & ~n11555 ;
  assign n11556 = n11555 ^ n11552 ;
  assign n11558 = n11557 ^ n11556 ;
  assign n11559 = n11557 ^ n7112 ;
  assign n11561 = n11557 ^ n7124 ;
  assign n11560 = n11557 ^ n11547 ;
  assign n11562 = n11561 ^ n11560 ;
  assign n11563 = n11561 ^ n11547 ;
  assign n11564 = n11563 ^ n7113 ;
  assign n11565 = n11564 ^ n11561 ;
  assign n11566 = ~n11562 & ~n11565 ;
  assign n11567 = n11566 ^ n11561 ;
  assign n11568 = ~n11559 & ~n11567 ;
  assign n11569 = n11568 ^ n7112 ;
  assign n11570 = ~n11558 & n11569 ;
  assign n11571 = n11549 & n11570 ;
  assign n11572 = n11571 ^ n11569 ;
  assign n11573 = n11572 ^ n7109 ;
  assign n11574 = ~n7111 & n11573 ;
  assign n11575 = n11574 ^ n7109 ;
  assign n11577 = n6838 & ~n11575 ;
  assign n11576 = n11575 ^ n6838 ;
  assign n11578 = n11577 ^ n11576 ;
  assign n11592 = n5882 ^ n5863 ;
  assign n11580 = ~n3943 & ~n6074 ;
  assign n11579 = ~n485 & ~n6072 ;
  assign n11581 = n11580 ^ n11579 ;
  assign n11582 = n11581 ^ x14 ;
  assign n11583 = n11582 ^ x13 ;
  assign n11584 = n4515 & n4897 ;
  assign n11585 = n11583 & n11584 ;
  assign n11586 = n11585 ^ n11582 ;
  assign n11587 = n11586 ^ n6814 ;
  assign n11588 = n11587 ^ n6805 ;
  assign n11589 = n11588 ^ n11586 ;
  assign n11590 = ~n6811 & ~n11589 ;
  assign n11591 = n11590 ^ n11587 ;
  assign n11593 = n11592 ^ n11591 ;
  assign n11594 = n11593 ^ n6817 ;
  assign n11595 = n11593 ^ n11577 ;
  assign n11597 = n11593 ^ n6815 ;
  assign n11596 = n11593 ^ n6800 ;
  assign n11598 = n11597 ^ n11596 ;
  assign n11599 = n11593 ^ n6797 ;
  assign n11600 = n11599 ^ n11597 ;
  assign n11601 = n11598 & ~n11600 ;
  assign n11602 = n11601 ^ n11597 ;
  assign n11603 = ~n11595 & ~n11602 ;
  assign n11604 = n11603 ^ n11577 ;
  assign n11605 = ~n11594 & ~n11604 ;
  assign n11606 = ~n11578 & n11605 ;
  assign n11609 = n6818 & n11606 ;
  assign n11607 = n11606 ^ n11604 ;
  assign n11610 = n11609 ^ n11607 ;
  assign n11612 = n11611 ^ n11610 ;
  assign n11613 = n11592 ^ n11586 ;
  assign n11614 = ~n11591 & n11613 ;
  assign n11615 = n11614 ^ n11586 ;
  assign n11616 = n11615 ^ n11610 ;
  assign n11617 = n11612 & n11616 ;
  assign n11618 = n11617 ^ n11615 ;
  assign n11619 = n11618 ^ n6052 ;
  assign n11620 = ~n6054 & ~n11619 ;
  assign n11621 = n11620 ^ n6053 ;
  assign n11622 = n6049 & n11621 ;
  assign n11623 = ~n5899 & n11622 ;
  assign n11624 = n11623 ^ n11621 ;
  assign n11625 = n6053 & n6054 ;
  assign n11626 = n11625 ^ n6049 ;
  assign n11627 = ~n5898 & ~n11626 ;
  assign n11628 = ~n11624 & n11627 ;
  assign n11631 = n11626 ^ n6054 ;
  assign n11632 = n11631 ^ n6049 ;
  assign n11633 = n6049 ^ n5899 ;
  assign n11634 = n11633 ^ n6049 ;
  assign n11635 = n11632 & ~n11634 ;
  assign n11636 = n11635 ^ n6049 ;
  assign n11637 = n11618 & n11636 ;
  assign n11638 = n11628 & n11637 ;
  assign n11629 = n11628 ^ n11624 ;
  assign n11639 = n11638 ^ n11629 ;
  assign n11643 = n11642 ^ n11639 ;
  assign n11696 = ~n485 & n4916 ;
  assign n11689 = ~n3473 & n4504 ;
  assign n11685 = n4881 ^ n4723 ;
  assign n11686 = n11685 ^ x23 ;
  assign n11684 = n3956 & n4492 ;
  assign n11687 = n11686 ^ n11684 ;
  assign n11683 = ~n649 & ~n4496 ;
  assign n11688 = n11687 ^ n11683 ;
  assign n11690 = n11689 ^ n11688 ;
  assign n11682 = ~n317 & n4491 ;
  assign n11691 = n11690 ^ n11682 ;
  assign n11659 = ~n3473 & ~n4496 ;
  assign n11658 = ~n649 & n4491 ;
  assign n11660 = n11659 ^ n11658 ;
  assign n11655 = ~n824 & n4504 ;
  assign n11654 = ~n3476 & n4492 ;
  assign n11656 = n11655 ^ n11654 ;
  assign n11657 = n11656 ^ x23 ;
  assign n11661 = n11660 ^ n11657 ;
  assign n11653 = n4879 ^ n4732 ;
  assign n11662 = n11661 ^ n11653 ;
  assign n11650 = n5991 ^ n5982 ;
  assign n11651 = ~n5988 & n11650 ;
  assign n11652 = n11651 ^ n5991 ;
  assign n11679 = n11661 ^ n11652 ;
  assign n11680 = ~n11662 & n11679 ;
  assign n11681 = n11680 ^ n11661 ;
  assign n11692 = n11691 ^ n11681 ;
  assign n11693 = n11692 ^ x20 ;
  assign n11678 = ~n445 & n14027 ;
  assign n11694 = n11693 ^ n11678 ;
  assign n11677 = ~n3943 & n4683 ;
  assign n11695 = n11694 ^ n11677 ;
  assign n11697 = n11696 ^ n11695 ;
  assign n11676 = n3944 & n4684 ;
  assign n11698 = n11697 ^ n11676 ;
  assign n11667 = ~n317 & n14027 ;
  assign n11663 = n11662 ^ n11652 ;
  assign n11664 = n11663 ^ x20 ;
  assign n11649 = ~n445 & n4916 ;
  assign n11665 = n11664 ^ n11649 ;
  assign n11648 = ~n485 & n4683 ;
  assign n11666 = n11665 ^ n11648 ;
  assign n11668 = n11667 ^ n11666 ;
  assign n11647 = n3500 & n4684 ;
  assign n11669 = n11668 ^ n11647 ;
  assign n11670 = n5992 ^ n5975 ;
  assign n11671 = n5998 & n11670 ;
  assign n11672 = n11671 ^ n5992 ;
  assign n11673 = n11672 ^ n11663 ;
  assign n11674 = n11669 & ~n11673 ;
  assign n11675 = n11674 ^ n11672 ;
  assign n11699 = n11698 ^ n11675 ;
  assign n11644 = n6042 ^ n6025 ;
  assign n11645 = n6048 & n11644 ;
  assign n11646 = n11645 ^ n6042 ;
  assign n11700 = n11699 ^ n11646 ;
  assign n11706 = ~n3920 & n5703 ;
  assign n11707 = n20731 ^ n11706 ;
  assign n11708 = ~n3943 & n11707 ;
  assign n11709 = n11708 ^ x17 ;
  assign n11701 = n11672 ^ n11669 ;
  assign n11710 = n11709 ^ n11701 ;
  assign n11712 = n11701 ^ n11646 ;
  assign n11713 = ~n11710 & n11712 ;
  assign n11714 = n11713 ^ n11709 ;
  assign n11711 = n11710 ^ n11646 ;
  assign n11715 = n11714 ^ n11711 ;
  assign n11716 = n11700 & n11715 ;
  assign n11717 = n11716 ^ n11699 ;
  assign n11718 = n11717 ^ n11642 ;
  assign n11719 = n11714 ^ n11699 ;
  assign n11720 = n11718 & n11719 ;
  assign n11721 = n11643 & n11720 ;
  assign n11722 = n11721 ^ n11717 ;
  assign n11727 = ~n3943 & n4916 ;
  assign n11724 = ~n485 & n14027 ;
  assign n11723 = n4515 & n4684 ;
  assign n11725 = n11724 ^ n11723 ;
  assign n11726 = n11725 ^ x20 ;
  assign n11728 = n11727 ^ n11726 ;
  assign n11730 = n11722 & n11728 ;
  assign n11729 = n11728 ^ n11722 ;
  assign n11731 = n11730 ^ n11729 ;
  assign n11733 = n4890 ^ n4889 ;
  assign n11732 = n4884 ^ n4713 ;
  assign n11734 = n11733 ^ n11732 ;
  assign n11735 = n11734 ^ n11733 ;
  assign n11736 = n11733 ^ n11730 ;
  assign n11737 = n11736 ^ n11733 ;
  assign n11738 = ~n11735 & ~n11737 ;
  assign n11739 = n11738 ^ n11733 ;
  assign n11754 = n11737 ^ n11735 ;
  assign n11755 = n11754 ^ n11733 ;
  assign n11745 = n11685 ^ n11681 ;
  assign n11746 = n11691 & n11745 ;
  assign n11747 = n11746 ^ n11685 ;
  assign n11748 = n11747 ^ n11733 ;
  assign n11740 = n11692 ^ n11675 ;
  assign n11741 = n11698 & n11740 ;
  assign n11742 = n11741 ^ n11692 ;
  assign n11743 = n11742 ^ n11732 ;
  assign n11744 = n11743 ^ n11734 ;
  assign n11749 = n11748 ^ n11744 ;
  assign n11751 = n11743 ^ n11736 ;
  assign n11752 = n11751 ^ n11733 ;
  assign n11753 = ~n11749 & ~n11752 ;
  assign n11756 = n11755 ^ n11753 ;
  assign n11757 = n11739 & n11756 ;
  assign n11758 = n11757 ^ n11733 ;
  assign n11761 = n11747 ^ n11734 ;
  assign n11762 = n11761 ^ n11742 ;
  assign n11763 = n11762 ^ n11734 ;
  assign n11764 = n11743 & ~n11763 ;
  assign n11765 = n11764 ^ n11734 ;
  assign n11766 = ~n11758 & ~n11765 ;
  assign n11767 = ~n11731 & n11766 ;
  assign n11768 = n11767 ^ n11758 ;
  assign n11784 = n11768 ^ n4893 ;
  assign n11785 = ~n11783 & ~n11784 ;
  assign n4669 = n4667 ^ n4654 ;
  assign n4670 = ~n4668 & n4669 ;
  assign n4672 = n4671 ^ n4670 ;
  assign n4673 = n4672 ^ n4654 ;
  assign n11771 = n4893 & ~n11768 ;
  assign n4674 = n4670 ^ n4654 ;
  assign n11772 = n11771 ^ n4674 ;
  assign n11773 = n4673 & n11772 ;
  assign n11774 = n11773 ^ n11768 ;
  assign n11786 = n11785 ^ n11774 ;
  assign n11791 = n11790 ^ n11786 ;
  assign n11792 = ~n4487 & ~n4512 ;
  assign n11793 = n4569 & n11792 ;
  assign n11795 = n11793 ^ n4513 ;
  assign n11796 = n11795 ^ n4571 ;
  assign n11797 = n11796 ^ n11793 ;
  assign n11794 = n11793 ^ n11786 ;
  assign n11800 = n11794 ^ n4071 ;
  assign n11801 = n11800 ^ n11794 ;
  assign n11802 = n11797 & n11801 ;
  assign n11803 = n11802 ^ n11794 ;
  assign n11804 = n11791 & ~n11803 ;
  assign n11805 = n11804 ^ n11790 ;
  assign n11806 = ~n4573 & ~n11805 ;
  assign n12094 = n12093 ^ n11806 ;
  assign n12095 = n12091 & n12094 ;
  assign n12096 = n12089 ^ n11968 ;
  assign n12098 = n12089 ^ n11859 ;
  assign n12097 = n12089 ^ n11806 ;
  assign n12099 = n12098 ^ n12097 ;
  assign n12100 = n12098 ^ n11806 ;
  assign n12101 = n12100 ^ n11865 ;
  assign n12102 = n12101 ^ n12098 ;
  assign n12103 = n12099 & ~n12102 ;
  assign n12104 = n12103 ^ n12098 ;
  assign n12105 = n12096 & n12104 ;
  assign n12106 = n12105 ^ n11968 ;
  assign n12107 = ~n12095 & ~n12106 ;
  assign n11975 = n11850 & n11853 ;
  assign n11986 = n11975 ^ n11854 ;
  assign n11976 = n11975 ^ n11948 ;
  assign n11978 = n11975 ^ n11815 ;
  assign n11977 = n11975 ^ n11837 ;
  assign n11979 = n11978 ^ n11977 ;
  assign n11980 = n11978 ^ n11873 ;
  assign n11981 = n11980 ^ n11978 ;
  assign n11982 = ~n11979 & ~n11981 ;
  assign n11983 = n11982 ^ n11978 ;
  assign n11984 = ~n11976 & ~n11983 ;
  assign n11985 = n11984 ^ n11948 ;
  assign n11988 = n11987 ^ n11837 ;
  assign n11991 = n11988 ^ n11815 ;
  assign n11989 = n11988 ^ n11846 ;
  assign n11996 = n11987 & n11989 ;
  assign n11997 = ~n11991 & n11996 ;
  assign n11998 = n11997 ^ n11991 ;
  assign n11999 = n11998 ^ n11815 ;
  assign n12000 = n11985 & ~n11999 ;
  assign n12001 = n11986 & n12000 ;
  assign n12002 = n12001 ^ n11985 ;
  assign n12062 = n12061 ^ n12020 ;
  assign n12003 = ~n11928 & ~n11987 ;
  assign n12063 = n12062 ^ n12003 ;
  assign n12593 = ~n12002 & ~n12063 ;
  assign n12282 = n12063 ^ n12002 ;
  assign n12594 = n12593 ^ n12282 ;
  assign n12595 = ~n12278 & ~n12364 ;
  assign n12596 = n12594 & n12595 ;
  assign n12597 = n12596 ^ n12278 ;
  assign n12598 = ~n12107 & ~n12597 ;
  assign n12600 = n12592 ^ n12364 ;
  assign n12603 = ~n12593 & ~n12600 ;
  assign n12604 = n12603 ^ n12592 ;
  assign n12605 = n12598 & n12604 ;
  assign n12606 = n12605 ^ n12597 ;
  assign n12607 = n12592 & n12606 ;
  assign n12608 = n12107 ^ n12063 ;
  assign n12609 = n12282 & n12608 ;
  assign n12610 = n12609 ^ n12063 ;
  assign n12611 = n12607 & n12610 ;
  assign n12612 = n12611 ^ n12606 ;
  assign n12653 = n12612 ^ n12586 ;
  assign n12654 = n12591 & n12653 ;
  assign n12655 = n12654 ^ n12586 ;
  assign n12677 = n12666 ^ n12655 ;
  assign n12648 = n12647 ^ x29 ;
  assign n12649 = n12648 ^ n12572 ;
  assign n12622 = n3944 ^ n485 ;
  assign n12621 = n3944 ^ n445 ;
  assign n12623 = n12622 ^ n12621 ;
  assign n12626 = x30 & n12623 ;
  assign n12627 = n12626 ^ n12622 ;
  assign n12628 = ~n3520 & ~n12627 ;
  assign n12629 = n12628 ^ n3944 ;
  assign n12630 = x31 & n12629 ;
  assign n12650 = n12649 ^ n12630 ;
  assign n12726 = n12677 ^ n12650 ;
  assign n12727 = n12726 ^ n12677 ;
  assign n12728 = n12666 ^ n12649 ;
  assign n12729 = n12728 ^ n12677 ;
  assign n12730 = n12727 & n12729 ;
  assign n12731 = n12730 ^ n12677 ;
  assign n12732 = ~n12725 & n12731 ;
  assign n12733 = n12732 ^ n12701 ;
  assign n12734 = n12630 & ~n12655 ;
  assign n12735 = n12734 ^ n12701 ;
  assign n12736 = n12733 & ~n12735 ;
  assign n12665 = n12620 ^ n12617 ;
  assign n12667 = n12666 ^ n12665 ;
  assign n12738 = n12701 ^ n12649 ;
  assign n12739 = n12738 ^ n12734 ;
  assign n12737 = n12655 ^ n12630 ;
  assign n12740 = n12739 ^ n12737 ;
  assign n12741 = n12667 & n12740 ;
  assign n12742 = n12736 & n12741 ;
  assign n12743 = n12742 ^ n12733 ;
  assign n12854 = n508 & n12743 ;
  assign n12855 = ~n12746 & n12854 ;
  assign n12651 = n12650 ^ n12620 ;
  assign n12652 = n12651 ^ n12617 ;
  assign n12656 = n12655 ^ n12652 ;
  assign n12613 = n12612 ^ n12591 ;
  assign n12080 = n12079 ^ n12063 ;
  assign n12081 = n12080 ^ n12002 ;
  assign n12085 = n12084 ^ n12081 ;
  assign n12108 = n12107 ^ n12085 ;
  assign n11970 = n11869 ^ n11859 ;
  assign n11971 = ~n11866 & n11970 ;
  assign n11856 = n11855 ^ n11806 ;
  assign n11870 = n11869 ^ n11866 ;
  assign n11871 = n11870 ^ n11806 ;
  assign n11872 = n11856 & ~n11871 ;
  assign n11969 = n11968 ^ n11872 ;
  assign n11972 = n11971 ^ n11969 ;
  assign n12257 = n11865 ^ n11855 ;
  assign n12258 = n12257 ^ n11859 ;
  assign n12259 = n12258 ^ n11869 ;
  assign n12260 = n12259 ^ n11806 ;
  assign n12109 = n11775 ^ n4893 ;
  assign n12219 = n11784 & n12109 ;
  assign n12217 = n4671 ^ n4668 ;
  assign n12218 = n12217 ^ n4670 ;
  assign n12220 = n12219 ^ n12218 ;
  assign n12110 = n12109 ^ n11768 ;
  assign n12111 = n11742 ^ n11729 ;
  assign n12114 = n11747 ^ n11729 ;
  assign n12115 = ~n12111 & ~n12114 ;
  assign n12112 = n12111 ^ n11747 ;
  assign n12113 = ~n11732 & n12112 ;
  assign n12116 = n12115 ^ n12113 ;
  assign n12117 = n12116 ^ n11736 ;
  assign n12118 = n11747 ^ n11728 ;
  assign n12119 = n12118 ^ n11732 ;
  assign n12120 = n12119 ^ n11742 ;
  assign n12121 = n12120 ^ n11722 ;
  assign n12126 = n11701 ^ n11642 ;
  assign n12127 = n11710 & n12126 ;
  assign n12128 = n12127 ^ n11699 ;
  assign n12122 = n11710 ^ n11642 ;
  assign n12123 = n12122 ^ n11646 ;
  assign n12124 = n11646 ^ n11639 ;
  assign n12125 = ~n12123 & n12124 ;
  assign n12129 = n12128 ^ n12125 ;
  assign n12130 = n12123 ^ n11639 ;
  assign n12134 = n11625 ^ n5898 ;
  assign n12135 = n12134 ^ n6049 ;
  assign n12131 = n6054 ^ n5897 ;
  assign n12132 = n11618 ^ n5897 ;
  assign n12133 = n12131 & n12132 ;
  assign n12136 = n12135 ^ n12133 ;
  assign n12137 = n12131 ^ n11618 ;
  assign n12138 = n11615 ^ n11612 ;
  assign n12139 = n6838 ^ n6815 ;
  assign n12203 = n11576 ^ n6800 ;
  assign n12204 = n12203 ^ n6797 ;
  assign n12205 = n12139 & n12204 ;
  assign n12206 = n12205 ^ n11593 ;
  assign n12201 = n11575 ^ n6800 ;
  assign n12202 = n6801 & ~n12201 ;
  assign n12207 = n12206 ^ n12202 ;
  assign n12140 = n12139 ^ n6800 ;
  assign n12141 = n12140 ^ n6797 ;
  assign n12142 = n12141 ^ n11575 ;
  assign n12143 = n11572 ^ n7111 ;
  assign n12146 = n11552 ^ n7127 ;
  assign n12147 = ~n11548 & n12146 ;
  assign n12144 = n11552 ^ n11548 ;
  assign n12145 = n11555 & n12144 ;
  assign n12148 = n12147 ^ n12145 ;
  assign n12149 = n12148 ^ n7126 ;
  assign n12150 = n12146 ^ n11555 ;
  assign n12151 = n12150 ^ n11547 ;
  assign n12152 = n11544 ^ n8049 ;
  assign n12154 = n11518 ^ n8405 ;
  assign n12159 = ~n11532 & ~n12154 ;
  assign n12153 = n11519 ^ n8397 ;
  assign n12155 = n12154 ^ n11515 ;
  assign n12156 = n12155 ^ n8397 ;
  assign n12157 = ~n12153 & ~n12156 ;
  assign n12158 = n12157 ^ n11522 ;
  assign n12160 = n12159 ^ n12158 ;
  assign n12161 = n11519 ^ n8406 ;
  assign n12162 = n12161 ^ n11518 ;
  assign n12163 = n12162 ^ n11515 ;
  assign n12165 = n10120 ^ n10109 ;
  assign n12166 = n12165 ^ n10116 ;
  assign n12164 = ~n10123 & ~n11503 ;
  assign n12167 = n12166 ^ n12164 ;
  assign n12168 = n11503 ^ n10123 ;
  assign n12169 = n11501 ^ n11495 ;
  assign n12171 = n10768 ^ n10699 ;
  assign n12172 = n12171 ^ n11479 ;
  assign n12173 = n11481 & n12172 ;
  assign n12174 = n12173 ^ n10766 ;
  assign n12170 = ~n10768 & ~n11489 ;
  assign n12175 = n12174 ^ n12170 ;
  assign n12176 = n10749 ^ n10136 ;
  assign n12177 = n12176 ^ n10701 ;
  assign n12178 = n12177 ^ n10699 ;
  assign n12179 = n12178 ^ n11479 ;
  assign n12180 = n11477 ^ n10771 ;
  assign n12183 = n11451 ^ n10826 ;
  assign n12181 = n11474 ^ n11457 ;
  assign n12182 = n11454 ^ n10808 ;
  assign n12222 = n12182 ^ n12181 ;
  assign n12223 = ~n12181 & ~n12222 ;
  assign n12224 = n12183 & n12223 ;
  assign n12225 = n12224 ^ n12222 ;
  assign n12184 = n12182 & n12183 ;
  assign n12185 = n12184 ^ n12183 ;
  assign n12186 = n12185 ^ n12182 ;
  assign n12187 = ~n12181 & n12186 ;
  assign n12226 = n12225 ^ n12187 ;
  assign n12227 = ~n12180 & ~n12226 ;
  assign n12228 = n12179 & ~n12227 ;
  assign n12229 = ~n12175 & ~n12228 ;
  assign n12230 = ~n12169 & ~n12229 ;
  assign n12231 = ~n12168 & ~n12230 ;
  assign n12232 = n12167 & ~n12231 ;
  assign n12233 = ~n12163 & ~n12232 ;
  assign n12234 = n12160 & ~n12233 ;
  assign n12235 = ~n12152 & ~n12234 ;
  assign n12236 = ~n12151 & ~n12235 ;
  assign n12237 = ~n12149 & ~n12236 ;
  assign n12238 = n12143 & ~n12237 ;
  assign n12239 = n12142 & ~n12238 ;
  assign n12240 = n12207 & ~n12239 ;
  assign n12241 = n12138 & ~n12240 ;
  assign n12242 = n12137 & ~n12241 ;
  assign n12243 = n12136 & ~n12242 ;
  assign n12244 = n12130 & ~n12243 ;
  assign n12245 = n12129 & ~n12244 ;
  assign n12246 = n12121 & ~n12245 ;
  assign n12247 = ~n12117 & ~n12246 ;
  assign n12248 = ~n12110 & ~n12247 ;
  assign n12249 = n12220 & ~n12248 ;
  assign n12188 = n12180 & ~n12187 ;
  assign n12189 = ~n12179 & ~n12188 ;
  assign n12190 = n12175 & ~n12189 ;
  assign n12191 = n12169 & ~n12190 ;
  assign n12192 = n12168 & ~n12191 ;
  assign n12193 = ~n12167 & ~n12192 ;
  assign n12194 = n12163 & ~n12193 ;
  assign n12195 = ~n12160 & ~n12194 ;
  assign n12196 = n12152 & ~n12195 ;
  assign n12197 = n12151 & ~n12196 ;
  assign n12198 = n12149 & ~n12197 ;
  assign n12199 = ~n12143 & ~n12198 ;
  assign n12200 = ~n12142 & ~n12199 ;
  assign n12208 = ~n12200 & ~n12207 ;
  assign n12209 = ~n12138 & ~n12208 ;
  assign n12210 = ~n12137 & ~n12209 ;
  assign n12211 = ~n12136 & ~n12210 ;
  assign n12212 = ~n12130 & ~n12211 ;
  assign n12213 = ~n12129 & ~n12212 ;
  assign n12214 = ~n12121 & ~n12213 ;
  assign n12215 = n12117 & ~n12214 ;
  assign n12216 = n12110 & ~n12215 ;
  assign n12221 = ~n12216 & ~n12220 ;
  assign n12250 = n12249 ^ n12221 ;
  assign n12255 = n11797 ^ n4071 ;
  assign n12251 = n11787 ^ n4569 ;
  assign n12252 = n12251 ^ n4513 ;
  assign n12253 = n11787 ^ n11786 ;
  assign n12254 = n12252 & ~n12253 ;
  assign n12256 = n12255 ^ n12254 ;
  assign n12261 = n12260 ^ n12256 ;
  assign n12262 = n12252 ^ n11786 ;
  assign n12263 = n12262 ^ n12260 ;
  assign n12264 = ~n12261 & n12263 ;
  assign n12265 = n12250 & n12264 ;
  assign n12266 = n12264 ^ n12256 ;
  assign n12267 = n12266 ^ n12220 ;
  assign n12268 = n12265 & n12267 ;
  assign n12269 = n12268 ^ n12266 ;
  assign n12271 = ~n12260 & n12269 ;
  assign n12275 = n11972 & ~n12271 ;
  assign n12276 = n12108 & ~n12275 ;
  assign n12285 = n12084 ^ n12080 ;
  assign n12286 = n12285 ^ n12002 ;
  assign n12287 = n12107 & ~n12286 ;
  assign n12365 = n12364 ^ n12287 ;
  assign n12284 = ~n12081 & n12278 ;
  assign n12366 = n12365 ^ n12284 ;
  assign n12281 = n12280 ^ n12063 ;
  assign n12283 = ~n12281 & ~n12282 ;
  assign n12367 = n12366 ^ n12283 ;
  assign n12660 = ~n12276 & ~n12367 ;
  assign n12661 = n12613 & ~n12660 ;
  assign n12662 = n12656 & ~n12661 ;
  assign n12702 = n12701 ^ n12677 ;
  assign n12678 = n12677 ^ n12667 ;
  assign n12703 = n12702 ^ n12678 ;
  assign n12671 = n12630 & ~n12649 ;
  assign n12704 = n12703 ^ n12671 ;
  assign n12664 = n12655 ^ n12650 ;
  assign n12668 = n12667 ^ n12666 ;
  assign n12669 = n12668 ^ n12650 ;
  assign n12670 = n12669 ^ n12667 ;
  assign n12674 = ~n12670 & ~n12671 ;
  assign n12675 = n12674 ^ n12667 ;
  assign n12676 = ~n12664 & n12675 ;
  assign n12705 = n12704 ^ n12676 ;
  assign n12723 = ~n12662 & n12705 ;
  assign n12750 = ~n262 & ~n3935 ;
  assign n12747 = n12636 ^ n1408 ;
  assign n12748 = n12747 ^ n298 ;
  assign n12749 = n12748 ^ n256 ;
  assign n12751 = n12750 ^ n12749 ;
  assign n12752 = n476 & n12751 ;
  assign n12753 = n12752 ^ n12699 ;
  assign n12754 = n12753 ^ n12746 ;
  assign n12755 = n12754 ^ n12743 ;
  assign n12917 = ~n12723 & n12755 ;
  assign n12849 = n626 ^ n448 ;
  assign n12847 = n3592 ^ n433 ;
  assign n12846 = n298 ^ n119 ;
  assign n12848 = n12847 ^ n12846 ;
  assign n12850 = n12849 ^ n12848 ;
  assign n12851 = n12850 ^ n718 ;
  assign n12852 = ~n390 & ~n12851 ;
  assign n12932 = n12752 ^ n12689 ;
  assign n12933 = n12752 ^ n12685 ;
  assign n12934 = n12933 ^ n12743 ;
  assign n12935 = n12932 & ~n12934 ;
  assign n12926 = n12852 ^ n12752 ;
  assign n12936 = n12935 ^ n12926 ;
  assign n12937 = n12753 & n12936 ;
  assign n12919 = n254 & n12689 ;
  assign n12920 = ~n12699 & ~n12852 ;
  assign n12921 = ~n12685 & n12920 ;
  assign n12922 = n12921 ^ n12685 ;
  assign n12923 = n12919 & ~n12922 ;
  assign n12924 = n12923 ^ n12921 ;
  assign n12925 = n12924 ^ n12752 ;
  assign n12927 = n12926 ^ n12925 ;
  assign n12931 = n12927 ^ n12753 ;
  assign n12938 = n12937 ^ n12931 ;
  assign n12939 = n12938 ^ n12924 ;
  assign n12951 = n12752 & n12939 ;
  assign n12952 = ~n12937 & n12951 ;
  assign n12953 = n12952 ^ n12937 ;
  assign n12945 = n12938 ^ n12937 ;
  assign n12954 = n12953 ^ n12945 ;
  assign n12955 = ~n12743 & n12954 ;
  assign n12956 = n12955 ^ n12924 ;
  assign n12957 = ~n12852 & ~n12956 ;
  assign n12958 = n12752 ^ n12743 ;
  assign n12961 = n12700 & n12744 ;
  assign n12962 = n12961 ^ n12699 ;
  assign n12966 = ~n12743 & n12962 ;
  assign n12967 = n12966 ^ n12744 ;
  assign n12968 = ~n12958 & n12967 ;
  assign n12969 = n12968 ^ n12752 ;
  assign n12970 = n12957 & n12969 ;
  assign n12971 = n12970 ^ n12956 ;
  assign n12987 = ~n12917 & ~n12971 ;
  assign n14221 = ~n12855 & ~n12987 ;
  assign n24690 = n650 & ~n14221 ;
  assign n24689 = n12971 & ~n24688 ;
  assign n24691 = n24690 ^ n24689 ;
  assign n24692 = n24691 ^ n829 ;
  assign n24693 = x29 & ~n24692 ;
  assign n24695 = n24694 ^ n24693 ;
  assign n24686 = ~n47 & n650 ;
  assign n24687 = ~n14221 & n24686 ;
  assign n24696 = n24695 ^ n24687 ;
  assign n12270 = n12269 ^ n12260 ;
  assign n12272 = n12271 ^ n12270 ;
  assign n12273 = ~n11972 & ~n12272 ;
  assign n12274 = ~n12108 & ~n12273 ;
  assign n12657 = ~n12274 & n12367 ;
  assign n12658 = ~n12613 & ~n12657 ;
  assign n12659 = ~n12656 & ~n12658 ;
  assign n12663 = n12662 ^ n12659 ;
  assign n12706 = n12705 ^ n12663 ;
  assign n24055 = n12706 ^ n12656 ;
  assign n24056 = n23912 & n24055 ;
  assign n24053 = ~n35 & n12656 ;
  assign n24051 = n12656 ^ n3726 ;
  assign n12879 = ~n35 & ~n12613 ;
  assign n24052 = n24051 ^ n12879 ;
  assign n24054 = n24053 ^ n24052 ;
  assign n24057 = n24056 ^ n24054 ;
  assign n24043 = n12879 ^ n12656 ;
  assign n24044 = n24043 ^ n3726 ;
  assign n24045 = n24044 ^ n24043 ;
  assign n24046 = n24043 ^ n12705 ;
  assign n24047 = n24046 ^ n24043 ;
  assign n24048 = n24045 & n24047 ;
  assign n24049 = n24048 ^ n24043 ;
  assign n24050 = ~x31 & n24049 ;
  assign n24058 = n24057 ^ n24050 ;
  assign n24036 = n2663 ^ n1074 ;
  assign n24037 = n24036 ^ n667 ;
  assign n24034 = n2627 ^ n210 ;
  assign n14544 = n305 ^ n226 ;
  assign n24033 = n14544 ^ n478 ;
  assign n24035 = n24034 ^ n24033 ;
  assign n24038 = n24037 ^ n24035 ;
  assign n24039 = n24038 ^ n187 ;
  assign n24040 = n24039 ^ n437 ;
  assign n24041 = ~n648 & n12633 ;
  assign n24042 = ~n24040 & n24041 ;
  assign n24059 = n24058 ^ n24042 ;
  assign n12900 = n1987 ^ n228 ;
  assign n12901 = n12900 ^ n973 ;
  assign n12899 = n2694 ^ n994 ;
  assign n12902 = n12901 ^ n12899 ;
  assign n12903 = n12902 ^ n530 ;
  assign n12906 = n426 ^ n273 ;
  assign n12905 = n702 ^ n223 ;
  assign n12907 = n12906 ^ n12905 ;
  assign n12904 = n4263 ^ n193 ;
  assign n12908 = n12907 ^ n12904 ;
  assign n12909 = n12908 ^ n6399 ;
  assign n12910 = n12632 & ~n12909 ;
  assign n12911 = ~n12903 & n12910 ;
  assign n12912 = ~n3472 & n12911 ;
  assign n24683 = n24058 ^ n12912 ;
  assign n24684 = n24059 & n24683 ;
  assign n24675 = n3941 ^ n449 ;
  assign n24676 = n24675 ^ n483 ;
  assign n24677 = n24676 ^ n1074 ;
  assign n24678 = n24677 ^ n286 ;
  assign n24679 = n24678 ^ n389 ;
  assign n24680 = n24679 ^ n424 ;
  assign n24681 = n24680 ^ n12859 ;
  assign n24672 = n5208 ^ n35 ;
  assign n24673 = ~n12705 & ~n24672 ;
  assign n12722 = ~n12659 & ~n12705 ;
  assign n12724 = n12723 ^ n12722 ;
  assign n24670 = n3726 & ~n12724 ;
  assign n12756 = n12755 ^ n12724 ;
  assign n24669 = n3520 & ~n12756 ;
  assign n24671 = n24670 ^ n24669 ;
  assign n24674 = n24673 ^ n24671 ;
  assign n24682 = n24681 ^ n24674 ;
  assign n24685 = n24684 ^ n24682 ;
  assign n24697 = n24696 ^ n24685 ;
  assign n12837 = n4503 ^ x23 ;
  assign n12838 = n12837 ^ n4499 ;
  assign n12810 = n222 ^ n106 ;
  assign n12811 = n12810 ^ n5101 ;
  assign n12812 = n12811 ^ n2824 ;
  assign n12806 = n1059 ^ n814 ;
  assign n12807 = n12806 ^ n841 ;
  assign n12804 = n3973 ^ n88 ;
  assign n12805 = n12804 ^ n1215 ;
  assign n12808 = n12807 ^ n12805 ;
  assign n12803 = n3756 ^ n574 ;
  assign n12809 = n12808 ^ n12803 ;
  assign n12813 = n12812 ^ n12809 ;
  assign n12797 = n499 ^ n394 ;
  assign n12798 = n12797 ^ n1534 ;
  assign n12799 = n12798 ^ n3664 ;
  assign n12794 = n362 ^ n104 ;
  assign n12795 = n12794 ^ n2035 ;
  assign n12792 = n737 ^ n425 ;
  assign n12791 = n981 ^ n845 ;
  assign n12793 = n12792 ^ n12791 ;
  assign n12796 = n12795 ^ n12793 ;
  assign n12800 = n12799 ^ n12796 ;
  assign n12788 = n641 ^ n489 ;
  assign n12786 = n364 ^ n125 ;
  assign n12787 = n12786 ^ n742 ;
  assign n12789 = n12788 ^ n12787 ;
  assign n12790 = n12789 ^ n5624 ;
  assign n12801 = n12800 ^ n12790 ;
  assign n12802 = n12801 ^ n4314 ;
  assign n12814 = n12813 ^ n12802 ;
  assign n12832 = n1875 ^ n1123 ;
  assign n12831 = n4282 ^ n2213 ;
  assign n12833 = n12832 ^ n12831 ;
  assign n12828 = n964 ^ n882 ;
  assign n12829 = n12828 ^ n409 ;
  assign n12826 = n457 ^ n130 ;
  assign n12827 = n12826 ^ n2005 ;
  assign n12830 = n12829 ^ n12827 ;
  assign n12834 = n12833 ^ n12830 ;
  assign n12821 = n1640 ^ n496 ;
  assign n12819 = n1819 ^ n180 ;
  assign n12820 = n12819 ^ n550 ;
  assign n12822 = n12821 ^ n12820 ;
  assign n12823 = n12822 ^ n1292 ;
  assign n12815 = n1355 ^ n804 ;
  assign n12816 = n12815 ^ n2365 ;
  assign n12438 = n914 ^ n153 ;
  assign n12817 = n12816 ^ n12438 ;
  assign n12818 = n12817 ^ n2218 ;
  assign n12824 = n12823 ^ n12818 ;
  assign n12825 = n12824 ^ n4762 ;
  assign n12835 = n12834 ^ n12825 ;
  assign n12836 = ~n12814 & ~n12835 ;
  assign n12839 = n12838 ^ n12836 ;
  assign n12525 = n938 ^ n195 ;
  assign n12526 = n12525 ^ n3428 ;
  assign n12519 = n1020 ^ n689 ;
  assign n12518 = n6225 ^ n815 ;
  assign n12520 = n12519 ^ n12518 ;
  assign n12516 = n12308 ^ n1683 ;
  assign n12517 = n12516 ^ n872 ;
  assign n12521 = n12520 ^ n12517 ;
  assign n12522 = n12521 ^ n5310 ;
  assign n12513 = n1555 ^ n501 ;
  assign n12514 = n12513 ^ n1185 ;
  assign n12509 = n426 ^ n221 ;
  assign n12510 = n12509 ^ n4796 ;
  assign n12511 = n12510 ^ n4356 ;
  assign n12507 = n2374 ^ n490 ;
  assign n12505 = n791 ^ n172 ;
  assign n12506 = n12505 ^ n765 ;
  assign n12508 = n12507 ^ n12506 ;
  assign n12512 = n12511 ^ n12508 ;
  assign n12515 = n12514 ^ n12512 ;
  assign n12523 = n12522 ^ n12515 ;
  assign n12439 = n12438 ^ n2397 ;
  assign n12440 = n12439 ^ n2662 ;
  assign n12436 = n4092 ^ n280 ;
  assign n12435 = n6207 ^ n547 ;
  assign n12437 = n12436 ^ n12435 ;
  assign n12441 = n12440 ^ n12437 ;
  assign n12432 = n11890 ^ n351 ;
  assign n12430 = n2509 ^ n236 ;
  assign n12431 = n12430 ^ n298 ;
  assign n12433 = n12432 ^ n12431 ;
  assign n12426 = n954 ^ n117 ;
  assign n12427 = n12426 ^ n104 ;
  assign n12425 = n1510 ^ n161 ;
  assign n12428 = n12427 ^ n12425 ;
  assign n12424 = n5128 ^ n3128 ;
  assign n12429 = n12428 ^ n12424 ;
  assign n12434 = n12433 ^ n12429 ;
  assign n12442 = n12441 ^ n12434 ;
  assign n12524 = n12523 ^ n12442 ;
  assign n12527 = n12526 ^ n12524 ;
  assign n12528 = ~n4335 & ~n12527 ;
  assign n12885 = n12839 ^ n12528 ;
  assign n12783 = ~n35 & ~n12367 ;
  assign n12780 = ~n3520 & n12613 ;
  assign n12781 = n12780 ^ n3520 ;
  assign n12777 = n12660 ^ n12657 ;
  assign n12778 = ~n12777 & n23912 ;
  assign n12779 = n12778 ^ n12613 ;
  assign n12782 = n12781 ^ n12779 ;
  assign n12784 = n12783 ^ n12782 ;
  assign n12530 = ~n35 & ~n12108 ;
  assign n12772 = n12530 ^ n12367 ;
  assign n12773 = n12772 ^ n12530 ;
  assign n12774 = ~n3520 & ~n12773 ;
  assign n12775 = n12774 ^ n12530 ;
  assign n12776 = x31 & n12775 ;
  assign n12785 = n12784 ^ n12776 ;
  assign n12886 = n12885 ^ n12785 ;
  assign n12386 = ~n3520 & n12108 ;
  assign n12385 = n12108 ^ n3520 ;
  assign n12387 = n12386 ^ n12385 ;
  assign n11973 = ~n35 & n11972 ;
  assign n12388 = n12387 ^ n11973 ;
  assign n12375 = n12275 ^ n12273 ;
  assign n12376 = n12375 ^ n12108 ;
  assign n12389 = n12388 ^ n12376 ;
  assign n12378 = n12376 ^ n11972 ;
  assign n12377 = n12376 ^ n12260 ;
  assign n12379 = n12378 ^ n12377 ;
  assign n12380 = n12378 ^ x30 ;
  assign n12381 = n12380 ^ n12378 ;
  assign n12382 = n12379 & n12381 ;
  assign n12383 = n12382 ^ n12378 ;
  assign n12384 = ~n3520 & n12383 ;
  assign n12390 = n12389 ^ n12384 ;
  assign n12391 = x31 & n12390 ;
  assign n12392 = n12391 ^ n12388 ;
  assign n12417 = n2469 ^ n899 ;
  assign n12418 = n12417 ^ n3055 ;
  assign n12414 = n2574 ^ n1982 ;
  assign n12415 = n12414 ^ n1125 ;
  assign n12413 = n5115 ^ n1172 ;
  assign n12416 = n12415 ^ n12413 ;
  assign n12419 = n12418 ^ n12416 ;
  assign n12410 = n3390 ^ n1190 ;
  assign n12408 = n1029 ^ n797 ;
  assign n12406 = n1197 ^ n537 ;
  assign n12407 = n12406 ^ n737 ;
  assign n12409 = n12408 ^ n12407 ;
  assign n12411 = n12410 ^ n12409 ;
  assign n12412 = n12411 ^ n1895 ;
  assign n12420 = n12419 ^ n12412 ;
  assign n12401 = n455 ^ n296 ;
  assign n12402 = n12401 ^ n1428 ;
  assign n12400 = n1389 ^ n1202 ;
  assign n12403 = n12402 ^ n12400 ;
  assign n12397 = n3651 ^ n148 ;
  assign n12398 = n12397 ^ n673 ;
  assign n12394 = n1208 ^ n703 ;
  assign n12395 = n12394 ^ n137 ;
  assign n12396 = n12395 ^ n1298 ;
  assign n12399 = n12398 ^ n12396 ;
  assign n12404 = n12403 ^ n12399 ;
  assign n12393 = n3315 ^ n1567 ;
  assign n12405 = n12404 ^ n12393 ;
  assign n12421 = n12420 ^ n12405 ;
  assign n12422 = ~n2353 & ~n12421 ;
  assign n12423 = n12422 ^ n8212 ;
  assign n12471 = n920 ^ n760 ;
  assign n12469 = n3975 ^ n245 ;
  assign n12470 = n12469 ^ n1906 ;
  assign n12472 = n12471 ^ n12470 ;
  assign n12465 = n1088 ^ n359 ;
  assign n12464 = n1961 ^ n597 ;
  assign n12466 = n12465 ^ n12464 ;
  assign n12462 = n2213 ^ n1732 ;
  assign n12460 = n764 ^ n308 ;
  assign n12461 = n12460 ^ n844 ;
  assign n12463 = n12462 ^ n12461 ;
  assign n12467 = n12466 ^ n12463 ;
  assign n12456 = n642 ^ n378 ;
  assign n12457 = n12456 ^ n407 ;
  assign n12454 = n733 ^ n362 ;
  assign n12453 = n762 ^ n197 ;
  assign n12455 = n12454 ^ n12453 ;
  assign n12458 = n12457 ^ n12455 ;
  assign n12452 = n4352 ^ n845 ;
  assign n12459 = n12458 ^ n12452 ;
  assign n12468 = n12467 ^ n12459 ;
  assign n12473 = n12472 ^ n12468 ;
  assign n12449 = n4358 ^ n1171 ;
  assign n12450 = n12449 ^ n2262 ;
  assign n12446 = n3433 ^ n497 ;
  assign n12447 = n12446 ^ n550 ;
  assign n12443 = n1198 ^ n614 ;
  assign n12444 = n12443 ^ n403 ;
  assign n12445 = n12444 ^ n622 ;
  assign n12448 = n12447 ^ n12445 ;
  assign n12451 = n12450 ^ n12448 ;
  assign n12474 = n12473 ^ n12451 ;
  assign n12475 = ~n3062 & ~n12474 ;
  assign n12476 = ~n12442 & n12475 ;
  assign n12477 = n12476 ^ n8212 ;
  assign n12478 = n12423 & n12477 ;
  assign n12479 = n12478 ^ n8212 ;
  assign n12491 = n1014 ^ n391 ;
  assign n12492 = n12491 ^ n194 ;
  assign n12493 = n12492 ^ n116 ;
  assign n12490 = n2377 ^ n571 ;
  assign n12494 = n12493 ^ n12490 ;
  assign n12488 = n4747 ^ n203 ;
  assign n12487 = n2883 ^ n375 ;
  assign n12489 = n12488 ^ n12487 ;
  assign n12495 = n12494 ^ n12489 ;
  assign n12483 = n3442 ^ n849 ;
  assign n12484 = n12483 ^ n2325 ;
  assign n12485 = n12484 ^ n3294 ;
  assign n12481 = n1205 ^ n506 ;
  assign n12480 = n768 ^ n360 ;
  assign n12482 = n12481 ^ n12480 ;
  assign n12486 = n12485 ^ n12482 ;
  assign n12496 = n12495 ^ n12486 ;
  assign n12497 = n12496 ^ n11887 ;
  assign n12498 = ~n2154 & ~n12497 ;
  assign n12500 = n12479 & n12498 ;
  assign n12503 = ~n12392 & n12500 ;
  assign n12887 = n12785 ^ n12503 ;
  assign n12888 = n12887 ^ n12785 ;
  assign n12499 = n12498 ^ n12479 ;
  assign n12501 = n12500 ^ n12499 ;
  assign n12502 = n12392 & ~n12501 ;
  assign n12889 = n12887 ^ n12502 ;
  assign n12890 = n12889 ^ n12887 ;
  assign n12891 = n12887 ^ n12528 ;
  assign n12892 = n12891 ^ n12887 ;
  assign n12893 = ~n12890 & ~n12892 ;
  assign n12894 = ~n12888 & n12893 ;
  assign n12895 = n12894 ^ n12888 ;
  assign n12896 = n12895 ^ n12785 ;
  assign n12897 = n12886 & ~n12896 ;
  assign n12898 = n12897 ^ n12785 ;
  assign n12533 = n3726 ^ x31 ;
  assign n12881 = n12533 & ~n12780 ;
  assign n12871 = n12661 ^ n12658 ;
  assign n12876 = x31 & ~n12871 ;
  assign n12877 = n12876 ^ n12656 ;
  assign n12878 = n3520 & ~n12877 ;
  assign n12880 = n12879 ^ n12878 ;
  assign n12882 = n12881 ^ n12880 ;
  assign n12870 = x31 & n12783 ;
  assign n12883 = n12882 ^ n12870 ;
  assign n24612 = n12898 ^ n12883 ;
  assign n12981 = n831 & ~n12705 ;
  assign n12916 = ~n12722 & ~n12755 ;
  assign n12918 = n12917 ^ n12916 ;
  assign n12972 = n12971 ^ n12918 ;
  assign n12973 = n12972 ^ n12971 ;
  assign n12974 = n12971 ^ x29 ;
  assign n12975 = n12974 ^ x28 ;
  assign n12976 = n12975 ^ n12971 ;
  assign n12977 = ~n12973 & n12976 ;
  assign n12978 = n12977 ^ n12971 ;
  assign n12979 = n650 & n12978 ;
  assign n12980 = n12979 ^ x29 ;
  assign n12982 = n12981 ^ n12980 ;
  assign n12915 = n3484 & n12755 ;
  assign n12983 = n12982 ^ n12915 ;
  assign n24632 = ~n12983 & ~n24059 ;
  assign n24028 = n12983 ^ n12883 ;
  assign n12867 = n12838 ^ n12528 ;
  assign n12868 = ~n12839 & ~n12867 ;
  assign n12869 = n12868 ^ n12838 ;
  assign n24617 = n24028 ^ n12869 ;
  assign n24614 = n24612 ^ n12869 ;
  assign n24613 = n24059 ^ n12898 ;
  assign n24615 = n24614 ^ n24613 ;
  assign n24616 = n24615 ^ n24614 ;
  assign n24618 = n24617 ^ n24616 ;
  assign n24629 = n24618 ^ n24612 ;
  assign n24630 = n24629 ^ n24059 ;
  assign n24619 = n24618 ^ n24614 ;
  assign n24622 = n24619 ^ n12883 ;
  assign n24631 = n24630 ^ n24622 ;
  assign n24633 = n24632 ^ n24631 ;
  assign n24634 = ~n24612 & n24633 ;
  assign n24635 = n24634 ^ n24630 ;
  assign n24636 = n24635 ^ n24632 ;
  assign n24639 = n24635 ^ n24629 ;
  assign n24640 = n24639 ^ n24635 ;
  assign n24641 = ~n24634 & ~n24640 ;
  assign n24642 = n24636 & n24641 ;
  assign n24643 = n24642 ^ n24636 ;
  assign n24644 = n24643 ^ n24632 ;
  assign n24645 = ~n12912 & ~n24059 ;
  assign n24646 = n24645 ^ n12883 ;
  assign n24647 = n24646 ^ n24645 ;
  assign n24648 = n24645 ^ n12983 ;
  assign n24649 = n24648 ^ n24645 ;
  assign n24650 = n24647 & n24649 ;
  assign n24651 = n24650 ^ n24645 ;
  assign n24659 = n24649 ^ n24647 ;
  assign n24660 = n24659 ^ n24645 ;
  assign n24653 = n24645 ^ n12898 ;
  assign n24652 = n24645 ^ n12869 ;
  assign n24654 = n24653 ^ n24652 ;
  assign n24655 = n24653 ^ n24646 ;
  assign n24656 = n24655 ^ n24648 ;
  assign n24657 = n24656 ^ n24645 ;
  assign n24658 = ~n24654 & n24657 ;
  assign n24661 = n24660 ^ n24658 ;
  assign n24662 = n24651 & n24661 ;
  assign n24663 = n24662 ^ n24645 ;
  assign n24666 = n12912 & ~n24663 ;
  assign n24667 = ~n24644 & n24666 ;
  assign n24668 = n24667 ^ n24663 ;
  assign n24698 = n24697 ^ n24668 ;
  assign n24065 = n650 & ~n12855 ;
  assign n24066 = n24065 ^ x29 ;
  assign n24067 = n24066 ^ x28 ;
  assign n13005 = n12916 & n12971 ;
  assign n13006 = n13005 ^ n12971 ;
  assign n13007 = n13006 ^ n12987 ;
  assign n24068 = ~n13007 & n24065 ;
  assign n24069 = ~n24067 & n24068 ;
  assign n24070 = n24069 ^ n24066 ;
  assign n24064 = n3484 & n12971 ;
  assign n24071 = n24070 ^ n24064 ;
  assign n24063 = n831 & n12755 ;
  assign n24072 = n24071 ^ n24063 ;
  assign n24073 = n24072 ^ n12859 ;
  assign n24060 = n24059 ^ n12983 ;
  assign n12913 = n12912 ^ n12898 ;
  assign n24030 = n24028 ^ n12912 ;
  assign n24031 = n24030 ^ n12869 ;
  assign n24032 = n12913 & n24031 ;
  assign n24061 = n24060 ^ n24032 ;
  assign n12884 = n12883 ^ n12869 ;
  assign n24029 = ~n12884 & n24028 ;
  assign n24062 = n24061 ^ n24029 ;
  assign n24609 = n24062 ^ n12859 ;
  assign n24610 = n24073 & n24609 ;
  assign n24611 = n24610 ^ n24072 ;
  assign n24699 = n24698 ^ n24611 ;
  assign n12914 = n12913 ^ n12884 ;
  assign n12984 = n12983 ^ n12914 ;
  assign n12840 = n12839 ^ n12785 ;
  assign n12841 = n12840 ^ n12503 ;
  assign n12504 = n12503 ^ n12502 ;
  assign n12769 = n12504 & ~n12528 ;
  assign n12842 = n12841 ^ n12769 ;
  assign n12765 = n3484 & ~n12705 ;
  assign n12757 = n12756 ^ n12755 ;
  assign n12758 = n12755 ^ x29 ;
  assign n12759 = n12758 ^ x28 ;
  assign n12760 = n12759 ^ n12755 ;
  assign n12761 = ~n12757 & n12760 ;
  assign n12762 = n12761 ^ n12755 ;
  assign n12763 = n650 & n12762 ;
  assign n12764 = n12763 ^ x29 ;
  assign n12766 = n12765 ^ n12764 ;
  assign n12721 = n831 & n12656 ;
  assign n12767 = n12766 ^ n12721 ;
  assign n12996 = n12842 ^ n12767 ;
  assign n12534 = ~n12386 & n12533 ;
  assign n12529 = n12528 ^ n12504 ;
  assign n12531 = n12530 ^ n12529 ;
  assign n12277 = n12276 ^ n12274 ;
  assign n12368 = n12367 ^ n12277 ;
  assign n12369 = n12368 ^ n12367 ;
  assign n12370 = n12367 ^ x31 ;
  assign n12371 = n12370 ^ n12367 ;
  assign n12372 = ~n12369 & n12371 ;
  assign n12373 = n12372 ^ n12367 ;
  assign n12374 = n3520 & n12373 ;
  assign n12532 = n12531 ^ n12374 ;
  assign n12535 = n12534 ^ n12532 ;
  assign n11974 = x31 & n11973 ;
  assign n12536 = n12535 ^ n11974 ;
  assign n12715 = n3484 & n12656 ;
  assign n12707 = n12706 ^ n12705 ;
  assign n12708 = n12705 ^ x29 ;
  assign n12709 = n12708 ^ x28 ;
  assign n12710 = n12709 ^ n12705 ;
  assign n12711 = ~n12707 & n12710 ;
  assign n12712 = n12711 ^ n12705 ;
  assign n12713 = n650 & ~n12712 ;
  assign n12714 = n12713 ^ x29 ;
  assign n12716 = n12715 ^ n12714 ;
  assign n12614 = n831 & ~n12613 ;
  assign n12717 = n12716 ^ n12614 ;
  assign n12718 = n12717 ^ n12529 ;
  assign n12719 = ~n12536 & ~n12718 ;
  assign n12720 = n12719 ^ n12529 ;
  assign n12997 = n12996 ^ n12720 ;
  assign n12993 = n487 ^ x26 ;
  assign n12990 = ~n3501 & ~n12987 ;
  assign n12991 = n12990 ^ n446 ;
  assign n12992 = ~n12855 & n12991 ;
  assign n12994 = n12993 ^ n12992 ;
  assign n12986 = n12861 & n12971 ;
  assign n12995 = n12994 ^ n12986 ;
  assign n12998 = n12997 ^ n12995 ;
  assign n13002 = n64 & ~n12855 ;
  assign n13003 = n13002 ^ x26 ;
  assign n13004 = n13003 ^ x25 ;
  assign n13008 = n13002 & ~n13007 ;
  assign n13009 = ~n13004 & n13008 ;
  assign n13010 = n13009 ^ n13003 ;
  assign n13001 = n446 & n12971 ;
  assign n13011 = n13010 ^ n13001 ;
  assign n13000 = n12755 & n12861 ;
  assign n13012 = n13011 ^ n13000 ;
  assign n12999 = n12717 ^ n12536 ;
  assign n13013 = n13012 ^ n12999 ;
  assign n13082 = n12499 ^ n12392 ;
  assign n13098 = n13082 ^ n12999 ;
  assign n13078 = ~n3720 & n12260 ;
  assign n13073 = n12269 ^ n11972 ;
  assign n13074 = n13073 ^ n12256 ;
  assign n13075 = n13074 & n23912 ;
  assign n13072 = n4851 & ~n12256 ;
  assign n13076 = n13075 ^ n13072 ;
  assign n13071 = n3726 & n11972 ;
  assign n13077 = n13076 ^ n13071 ;
  assign n13079 = n13078 ^ n13077 ;
  assign n13083 = n13082 ^ n13079 ;
  assign n13038 = n838 ^ n592 ;
  assign n13037 = n1675 ^ n583 ;
  assign n13039 = n13038 ^ n13037 ;
  assign n13034 = n779 ^ n635 ;
  assign n13035 = n13034 ^ n1982 ;
  assign n13033 = n1482 ^ n218 ;
  assign n13036 = n13035 ^ n13033 ;
  assign n13040 = n13039 ^ n13036 ;
  assign n13041 = n13040 ^ n1755 ;
  assign n13031 = n6391 ^ n2387 ;
  assign n13029 = n2282 ^ n259 ;
  assign n13027 = n2269 ^ n280 ;
  assign n13028 = n13027 ^ n702 ;
  assign n13030 = n13029 ^ n13028 ;
  assign n13032 = n13031 ^ n13030 ;
  assign n13042 = n13041 ^ n13032 ;
  assign n13043 = n13042 ^ n2498 ;
  assign n13023 = n3401 ^ n1024 ;
  assign n13022 = n12490 ^ n2474 ;
  assign n13024 = n13023 ^ n13022 ;
  assign n13019 = n1321 ^ n239 ;
  assign n13017 = n1041 ^ n359 ;
  assign n13018 = n13017 ^ n149 ;
  assign n13020 = n13019 ^ n13018 ;
  assign n13014 = n426 ^ n194 ;
  assign n13015 = n13014 ^ n1798 ;
  assign n13016 = n13015 ^ n2969 ;
  assign n13021 = n13020 ^ n13016 ;
  assign n13025 = n13024 ^ n13021 ;
  assign n13026 = n13025 ^ n2505 ;
  assign n13044 = n13043 ^ n13026 ;
  assign n13045 = ~n4986 & ~n13044 ;
  assign n13046 = n13045 ^ n12476 ;
  assign n13048 = n12256 ^ n33 ;
  assign n13047 = ~n33 & ~n12256 ;
  assign n13049 = n13048 ^ n13047 ;
  assign n13050 = n12262 ^ n12256 ;
  assign n13062 = ~n13050 & n24214 ;
  assign n13061 = ~n35 & ~n12256 ;
  assign n13063 = n13062 ^ n13061 ;
  assign n13064 = n13063 ^ x31 ;
  assign n13051 = n12250 & n12262 ;
  assign n13052 = n13051 ^ n12249 ;
  assign n13053 = n13050 & ~n13052 ;
  assign n13056 = n12260 ^ x31 ;
  assign n13057 = n13056 ^ n12260 ;
  assign n13058 = ~n13053 & n13057 ;
  assign n13059 = n13058 ^ n12260 ;
  assign n13060 = n3520 & n13059 ;
  assign n13065 = n13064 ^ n13060 ;
  assign n13066 = n13049 & n13065 ;
  assign n13067 = n13066 ^ n13045 ;
  assign n13068 = ~n13046 & n13067 ;
  assign n13069 = n13068 ^ n12423 ;
  assign n13070 = n13068 ^ n12476 ;
  assign n13080 = n13079 ^ n13070 ;
  assign n13081 = n13069 & n13080 ;
  assign n13084 = n13083 ^ n13081 ;
  assign n13093 = n831 & ~n12367 ;
  assign n13086 = n12656 ^ x29 ;
  assign n13087 = n13086 ^ x28 ;
  assign n13088 = n13087 ^ n12656 ;
  assign n13089 = ~n12871 & n13088 ;
  assign n13090 = n13089 ^ n12656 ;
  assign n13091 = n650 & n13090 ;
  assign n13092 = n13091 ^ x29 ;
  assign n13094 = n13093 ^ n13092 ;
  assign n13085 = n3484 & ~n12613 ;
  assign n13095 = n13094 ^ n13085 ;
  assign n13096 = n13095 ^ n13082 ;
  assign n13097 = ~n13084 & ~n13096 ;
  assign n13099 = n13098 ^ n13097 ;
  assign n13100 = ~n13013 & ~n13099 ;
  assign n13101 = n13100 ^ n13012 ;
  assign n13102 = n13101 ^ n12995 ;
  assign n13103 = n12998 & ~n13102 ;
  assign n13104 = n13103 ^ n12995 ;
  assign n24006 = n12984 & ~n13104 ;
  assign n13353 = n13101 ^ n12998 ;
  assign n13106 = n13099 ^ n13012 ;
  assign n13107 = n13106 ^ n12838 ;
  assign n13119 = n3484 & ~n12367 ;
  assign n13110 = n12777 ^ n12613 ;
  assign n13111 = n13110 ^ n12613 ;
  assign n13112 = n12613 ^ x29 ;
  assign n13113 = n13112 ^ x28 ;
  assign n13114 = n13113 ^ n12613 ;
  assign n13115 = ~n13111 & n13114 ;
  assign n13116 = n13115 ^ n12613 ;
  assign n13117 = n650 & ~n13116 ;
  assign n13118 = n13117 ^ x29 ;
  assign n13120 = n13119 ^ n13118 ;
  assign n13109 = n831 & ~n12108 ;
  assign n13121 = n13120 ^ n13109 ;
  assign n13108 = n13079 ^ n12423 ;
  assign n13122 = n13121 ^ n13108 ;
  assign n13123 = n13122 ^ n13068 ;
  assign n13141 = n3775 ^ n3600 ;
  assign n13158 = n5081 ^ n1089 ;
  assign n13155 = n5565 ^ n413 ;
  assign n13154 = n768 ^ n141 ;
  assign n13156 = n13155 ^ n13154 ;
  assign n13151 = n2002 ^ n745 ;
  assign n13150 = n3331 ^ n906 ;
  assign n13152 = n13151 ^ n13150 ;
  assign n13147 = n4341 ^ n223 ;
  assign n13146 = n3390 ^ n451 ;
  assign n13148 = n13147 ^ n13146 ;
  assign n13143 = n1249 ^ n570 ;
  assign n13144 = n13143 ^ n260 ;
  assign n13142 = n1128 ^ n837 ;
  assign n13145 = n13144 ^ n13142 ;
  assign n13149 = n13148 ^ n13145 ;
  assign n13153 = n13152 ^ n13149 ;
  assign n13157 = n13156 ^ n13153 ;
  assign n13159 = n13158 ^ n13157 ;
  assign n13160 = n13159 ^ n2808 ;
  assign n13161 = ~n13141 & ~n13160 ;
  assign n13134 = n5299 ^ n3104 ;
  assign n13135 = n13134 ^ n2848 ;
  assign n13129 = n3119 ^ n175 ;
  assign n13130 = n13129 ^ n673 ;
  assign n13131 = n13130 ^ n283 ;
  assign n13132 = n13131 ^ n2240 ;
  assign n13127 = n842 ^ n818 ;
  assign n13126 = n12426 ^ n1113 ;
  assign n13128 = n13127 ^ n13126 ;
  assign n13133 = n13132 ^ n13128 ;
  assign n13136 = n13135 ^ n13133 ;
  assign n13137 = n13136 ^ n12451 ;
  assign n13125 = n12549 ^ n3061 ;
  assign n13138 = n13137 ^ n13125 ;
  assign n13139 = ~n4811 & ~n13138 ;
  assign n5708 = x17 & n5707 ;
  assign n5709 = n5705 & n5708 ;
  assign n5710 = n5709 ^ n5707 ;
  assign n13140 = n13139 ^ n5710 ;
  assign n13189 = n13161 ^ n13140 ;
  assign n13183 = n3520 & ~n12110 ;
  assign n13184 = n13183 ^ n12220 ;
  assign n13185 = x31 & n13184 ;
  assign n13181 = n3720 ^ n33 ;
  assign n13165 = n12220 ^ n12110 ;
  assign n13172 = n12248 ^ n12216 ;
  assign n13173 = x31 & ~n13172 ;
  assign n13174 = n13173 ^ n12262 ;
  assign n13175 = n13174 ^ n12262 ;
  assign n13178 = n13165 & n13175 ;
  assign n13179 = n13178 ^ n12262 ;
  assign n13180 = n3520 & n13179 ;
  assign n13182 = n13181 ^ n13180 ;
  assign n13186 = n13185 ^ n13182 ;
  assign n13187 = n24214 ^ n13186 ;
  assign n13166 = n13165 ^ n12220 ;
  assign n13169 = n13166 & ~n24214 ;
  assign n13170 = n13169 ^ n13165 ;
  assign n13171 = ~n35 & ~n13170 ;
  assign n13188 = n13187 ^ n13171 ;
  assign n13190 = n13189 ^ n13188 ;
  assign n13221 = n4228 ^ n759 ;
  assign n13222 = n13221 ^ n1415 ;
  assign n13219 = n2937 ^ n1920 ;
  assign n13218 = n1986 ^ n844 ;
  assign n13220 = n13219 ^ n13218 ;
  assign n13223 = n13222 ^ n13220 ;
  assign n13214 = n4004 ^ n397 ;
  assign n13213 = n6208 ^ n1798 ;
  assign n13215 = n13214 ^ n13213 ;
  assign n13211 = n2890 ^ n2208 ;
  assign n13212 = n13211 ^ n2541 ;
  assign n13216 = n13215 ^ n13212 ;
  assign n13208 = n5006 ^ n4223 ;
  assign n13209 = n13208 ^ n1336 ;
  assign n13210 = n13209 ^ n5351 ;
  assign n13217 = n13216 ^ n13210 ;
  assign n13224 = n13223 ^ n13217 ;
  assign n13225 = n13224 ^ n3306 ;
  assign n13226 = n2969 ^ n625 ;
  assign n13227 = n13226 ^ n12802 ;
  assign n13228 = ~n13225 & ~n13227 ;
  assign n13204 = ~n35 & n12117 ;
  assign n13203 = n13183 ^ n12117 ;
  assign n13205 = n13204 ^ n13203 ;
  assign n13206 = ~x31 & n13205 ;
  assign n13195 = n12247 ^ n12215 ;
  assign n13196 = n13195 ^ n12110 ;
  assign n13197 = n13196 ^ n12117 ;
  assign n13192 = n12121 ^ n12117 ;
  assign n13198 = n13197 ^ n13192 ;
  assign n13199 = n35 & n13198 ;
  assign n13200 = n13199 ^ n13192 ;
  assign n13201 = n4851 & n13200 ;
  assign n13202 = n13201 ^ n12117 ;
  assign n13207 = n13206 ^ n13202 ;
  assign n13229 = n13228 ^ n13207 ;
  assign n13259 = n4944 ^ n204 ;
  assign n13256 = n3444 ^ n1375 ;
  assign n13257 = n13256 ^ n1725 ;
  assign n13253 = n641 ^ n221 ;
  assign n13254 = n13253 ^ n3171 ;
  assign n13255 = n13254 ^ n4244 ;
  assign n13258 = n13257 ^ n13255 ;
  assign n13260 = n13259 ^ n13258 ;
  assign n13261 = n13260 ^ n1846 ;
  assign n13262 = n13261 ^ n3005 ;
  assign n13251 = n955 ^ n635 ;
  assign n13252 = n13251 ^ n5261 ;
  assign n13263 = n13262 ^ n13252 ;
  assign n13264 = ~n1011 & ~n13263 ;
  assign n13267 = n13264 ^ n13228 ;
  assign n13242 = n1222 ^ n1015 ;
  assign n13243 = n13242 ^ n1896 ;
  assign n13244 = n13243 ^ n4304 ;
  assign n13240 = n1450 ^ n797 ;
  assign n13238 = n5332 ^ n285 ;
  assign n13239 = n13238 ^ n2035 ;
  assign n13241 = n13240 ^ n13239 ;
  assign n13245 = n13244 ^ n13241 ;
  assign n13236 = n4343 ^ n1468 ;
  assign n13233 = n737 ^ n218 ;
  assign n13231 = n359 ^ n106 ;
  assign n13232 = n13231 ^ n190 ;
  assign n13234 = n13233 ^ n13232 ;
  assign n13230 = n4021 ^ n3540 ;
  assign n13235 = n13234 ^ n13230 ;
  assign n13237 = n13236 ^ n13235 ;
  assign n13246 = n13245 ^ n13237 ;
  assign n13247 = n13246 ^ n2382 ;
  assign n13248 = n6233 ^ n2447 ;
  assign n13249 = ~n13247 & ~n13248 ;
  assign n13250 = n13249 ^ n6070 ;
  assign n13265 = n13264 ^ n6070 ;
  assign n13266 = ~n13250 & n13265 ;
  assign n13268 = n13267 ^ n13266 ;
  assign n13269 = n13229 & ~n13268 ;
  assign n13270 = n13269 ^ n13228 ;
  assign n13271 = n13270 ^ n13188 ;
  assign n13191 = n13188 ^ n13161 ;
  assign n13272 = n13271 ^ n13191 ;
  assign n13276 = n13269 & n13272 ;
  assign n13277 = n13276 ^ n13191 ;
  assign n13278 = ~n13190 & n13277 ;
  assign n13279 = n13278 ^ n13188 ;
  assign n13162 = n13161 ^ n5710 ;
  assign n13163 = ~n13140 & n13162 ;
  assign n13164 = n13163 ^ n13161 ;
  assign n13319 = n13279 ^ n13164 ;
  assign n13280 = ~n13164 & n13279 ;
  assign n13320 = n13319 ^ n13280 ;
  assign n13124 = n13066 ^ n13046 ;
  assign n13281 = n13280 ^ n13124 ;
  assign n13291 = ~n3732 & n12262 ;
  assign n13294 = n3725 & ~n13047 ;
  assign n13295 = ~n13291 & n13294 ;
  assign n13283 = n13052 ^ n12256 ;
  assign n13284 = n13283 ^ n3520 ;
  assign n13285 = n13284 ^ n13283 ;
  assign n13286 = x30 & n12220 ;
  assign n13287 = n13286 ^ n13283 ;
  assign n13288 = ~n13285 & n13287 ;
  assign n13289 = n13288 ^ n13283 ;
  assign n13290 = x31 & n13289 ;
  assign n13292 = n13291 ^ n13290 ;
  assign n13296 = n13295 ^ n13292 ;
  assign n13297 = n13296 ^ n13124 ;
  assign n13282 = n13124 ^ n12476 ;
  assign n13298 = n13297 ^ n13282 ;
  assign n13310 = n3484 & n11972 ;
  assign n13308 = n13296 ^ x29 ;
  assign n13300 = n12376 ^ n12108 ;
  assign n13303 = n12108 ^ n4536 ;
  assign n13304 = n13303 ^ n12108 ;
  assign n13305 = ~n13300 & n13304 ;
  assign n13306 = n13305 ^ n12108 ;
  assign n13307 = n650 & ~n13306 ;
  assign n13309 = n13308 ^ n13307 ;
  assign n13311 = n13310 ^ n13309 ;
  assign n13299 = n831 & n12260 ;
  assign n13312 = n13311 ^ n13299 ;
  assign n13315 = ~n13298 & ~n13312 ;
  assign n13316 = n13315 ^ n13297 ;
  assign n13317 = ~n13281 & ~n13316 ;
  assign n13318 = n13317 ^ n13280 ;
  assign n13327 = ~n13282 & n13312 ;
  assign n13328 = n13297 & n13327 ;
  assign n13329 = n13328 ^ n13297 ;
  assign n13330 = n13329 ^ n13296 ;
  assign n13331 = ~n13318 & ~n13330 ;
  assign n13332 = ~n13320 & n13331 ;
  assign n13333 = n13332 ^ n13318 ;
  assign n13334 = n13333 ^ n13121 ;
  assign n13335 = ~n13123 & n13334 ;
  assign n13336 = n13335 ^ n13121 ;
  assign n13349 = n13336 ^ n13106 ;
  assign n13337 = n13095 ^ n13084 ;
  assign n13338 = n13337 ^ n13336 ;
  assign n13342 = n446 & n12755 ;
  assign n13341 = ~n12705 & n12861 ;
  assign n13343 = n13342 ^ n13341 ;
  assign n13344 = n13343 ^ x26 ;
  assign n13340 = ~n487 & n12971 ;
  assign n13345 = n13344 ^ n13340 ;
  assign n13339 = ~n3501 & ~n12972 ;
  assign n13346 = n13345 ^ n13339 ;
  assign n13347 = n13346 ^ n13336 ;
  assign n13348 = ~n13338 & n13347 ;
  assign n13350 = n13349 ^ n13348 ;
  assign n13351 = ~n13107 & ~n13350 ;
  assign n13352 = n13351 ^ n12838 ;
  assign n13354 = n13353 ^ n13352 ;
  assign n20822 = n13350 ^ n12838 ;
  assign n20808 = n4504 & ~n12855 ;
  assign n13355 = n13346 ^ n13338 ;
  assign n20807 = n13355 ^ n4502 ;
  assign n20809 = n20808 ^ n20807 ;
  assign n13430 = n4488 & ~n12855 ;
  assign n13431 = n13430 ^ x23 ;
  assign n13432 = n13431 ^ x22 ;
  assign n13433 = ~n13007 & n13430 ;
  assign n13434 = ~n13432 & n13433 ;
  assign n13435 = n13434 ^ n13431 ;
  assign n13429 = ~n4496 & n12971 ;
  assign n13436 = n13435 ^ n13429 ;
  assign n13428 = n4504 & n12755 ;
  assign n13437 = n13436 ^ n13428 ;
  assign n13383 = ~n12613 & n12861 ;
  assign n13382 = n446 & n12656 ;
  assign n13384 = n13383 ^ n13382 ;
  assign n13385 = n13384 ^ n65 ;
  assign n13386 = n13384 ^ x26 ;
  assign n13387 = n13386 ^ n67 ;
  assign n13388 = n13387 ^ x25 ;
  assign n13389 = n13388 ^ n12705 ;
  assign n13390 = n13389 ^ n13386 ;
  assign n13391 = n13390 ^ n12663 ;
  assign n13392 = n13391 ^ n13390 ;
  assign n13393 = n13386 & ~n13392 ;
  assign n13394 = n13393 ^ n13387 ;
  assign n13395 = n13390 ^ n12705 ;
  assign n13396 = ~n13392 & ~n13395 ;
  assign n13397 = n13396 ^ n12705 ;
  assign n13398 = ~n13387 & n13397 ;
  assign n13399 = ~n13394 & n13398 ;
  assign n13400 = n13399 ^ n13396 ;
  assign n13401 = n13400 ^ n67 ;
  assign n13402 = n13401 ^ n12705 ;
  assign n13403 = ~n13385 & ~n13402 ;
  assign n13373 = n13296 ^ n12476 ;
  assign n13374 = n13373 ^ n13319 ;
  assign n13375 = n13312 & n13374 ;
  assign n13376 = n13375 ^ n13124 ;
  assign n13371 = n13164 ^ n12476 ;
  assign n13372 = n13319 & n13371 ;
  assign n13377 = n13376 ^ n13372 ;
  assign n13378 = n13377 ^ x29 ;
  assign n13366 = n12367 ^ n4536 ;
  assign n13367 = n13366 ^ n12367 ;
  assign n13368 = ~n12369 & n13367 ;
  assign n13369 = n13368 ^ n12367 ;
  assign n13370 = n650 & ~n13369 ;
  assign n13379 = n13378 ^ n13370 ;
  assign n13363 = n3484 & ~n12108 ;
  assign n13380 = n13379 ^ n13363 ;
  assign n13362 = n831 & n11972 ;
  assign n13381 = n13380 ^ n13362 ;
  assign n13427 = n13403 ^ n13381 ;
  assign n13438 = n13437 ^ n13427 ;
  assign n13484 = n13319 ^ n12476 ;
  assign n13485 = n13484 ^ n13312 ;
  assign n13525 = n13485 ^ n13427 ;
  assign n13490 = n831 & ~n12256 ;
  assign n13489 = n3484 & n12260 ;
  assign n13491 = n13490 ^ n13489 ;
  assign n13492 = n13491 ^ x29 ;
  assign n13493 = n13492 ^ n653 ;
  assign n13502 = ~n11972 & n13493 ;
  assign n13498 = ~x28 & n13493 ;
  assign n13499 = n13498 ^ n653 ;
  assign n13500 = ~n12270 & n13499 ;
  assign n13501 = n13500 ^ n653 ;
  assign n13503 = n13502 ^ n13501 ;
  assign n13504 = n13491 ^ n651 ;
  assign n13505 = ~n13503 & ~n13504 ;
  assign n13508 = n13228 ^ n13161 ;
  assign n13456 = ~n3733 & ~n12110 ;
  assign n13453 = n13173 ^ n12220 ;
  assign n13454 = n3520 & ~n13453 ;
  assign n13452 = x31 & n13204 ;
  assign n13455 = n13454 ^ n13452 ;
  assign n13457 = n13456 ^ n13455 ;
  assign n13449 = n3484 & ~n12256 ;
  assign n13442 = n12260 ^ x29 ;
  assign n13443 = n13442 ^ x28 ;
  assign n13444 = n13443 ^ n12260 ;
  assign n13445 = n13053 & n13444 ;
  assign n13446 = n13445 ^ n12260 ;
  assign n13447 = n650 & n13446 ;
  assign n13448 = n13447 ^ x29 ;
  assign n13450 = n13449 ^ n13448 ;
  assign n13441 = n831 & ~n12262 ;
  assign n13451 = n13450 ^ n13441 ;
  assign n13462 = n13457 ^ n13451 ;
  assign n13509 = n13462 ^ n13269 ;
  assign n13510 = n13508 & ~n13509 ;
  assign n13511 = n13510 ^ n13190 ;
  assign n13506 = n13457 ^ n13270 ;
  assign n13507 = ~n13462 & ~n13506 ;
  assign n13512 = n13511 ^ n13507 ;
  assign n13513 = ~n13505 & n13512 ;
  assign n13439 = n13228 & ~n13270 ;
  assign n13440 = n13439 ^ n13269 ;
  assign n13458 = n13451 & n13457 ;
  assign n13459 = n13439 & n13458 ;
  assign n13460 = n13459 ^ n13190 ;
  assign n13461 = ~n13440 & ~n13460 ;
  assign n13463 = n13462 ^ n13458 ;
  assign n13464 = n13439 ^ n13161 ;
  assign n13465 = n13463 & ~n13464 ;
  assign n13466 = n13461 & n13465 ;
  assign n13467 = n13466 ^ n13460 ;
  assign n13486 = n13485 ^ n13467 ;
  assign n13468 = n13439 ^ n13190 ;
  assign n13469 = n13468 ^ n13190 ;
  assign n13474 = n13161 & n13458 ;
  assign n13475 = ~n13469 & n13474 ;
  assign n13476 = n13475 ^ n13469 ;
  assign n13477 = n13476 ^ n13468 ;
  assign n13478 = n13467 & n13477 ;
  assign n13487 = n13486 ^ n13478 ;
  assign n13479 = n13451 ^ n13161 ;
  assign n13480 = ~n13462 & n13479 ;
  assign n13481 = n13480 ^ n13161 ;
  assign n13482 = n13440 & n13481 ;
  assign n13483 = n13478 & n13482 ;
  assign n13488 = n13487 ^ n13483 ;
  assign n13514 = n13513 ^ n13488 ;
  assign n13518 = n446 & ~n12613 ;
  assign n13517 = ~n12367 & n12861 ;
  assign n13519 = n13518 ^ n13517 ;
  assign n13520 = n13519 ^ x26 ;
  assign n13516 = ~n487 & n12656 ;
  assign n13521 = n13520 ^ n13516 ;
  assign n12872 = n12871 ^ n12656 ;
  assign n13515 = ~n3501 & ~n12872 ;
  assign n13522 = n13521 ^ n13515 ;
  assign n13523 = n13522 ^ n13485 ;
  assign n13524 = n13514 & n13523 ;
  assign n13526 = n13525 ^ n13524 ;
  assign n13527 = ~n13438 & n13526 ;
  assign n13528 = n13527 ^ n13437 ;
  assign n13425 = n4504 & n12971 ;
  assign n13420 = n13333 ^ n13123 ;
  assign n13408 = n12656 & n12861 ;
  assign n13407 = n446 & ~n12705 ;
  assign n13409 = n13408 ^ n13407 ;
  assign n13410 = n13409 ^ n65 ;
  assign n13411 = n13409 ^ x26 ;
  assign n13415 = n13411 ^ n67 ;
  assign n13416 = ~x25 & ~n12724 ;
  assign n13417 = n13415 & n13416 ;
  assign n13413 = n67 & ~n12756 ;
  assign n13412 = ~n12755 & n13411 ;
  assign n13414 = n13413 ^ n13412 ;
  assign n13418 = n13417 ^ n13414 ;
  assign n13419 = ~n13410 & ~n13418 ;
  assign n13421 = n13420 ^ n13419 ;
  assign n13404 = n13403 ^ n13377 ;
  assign n13405 = n13381 & ~n13404 ;
  assign n13406 = n13405 ^ n13377 ;
  assign n13422 = n13421 ^ n13406 ;
  assign n13361 = n4491 ^ x23 ;
  assign n13423 = n13422 ^ n13361 ;
  assign n13358 = n4492 & ~n12987 ;
  assign n13359 = n13358 ^ n4496 ;
  assign n13360 = ~n12855 & ~n13359 ;
  assign n13424 = n13423 ^ n13360 ;
  assign n13426 = n13425 ^ n13424 ;
  assign n13533 = n13528 ^ n13426 ;
  assign n13534 = n13526 ^ n13437 ;
  assign n13680 = n13522 ^ n13514 ;
  assign n13542 = ~n487 & ~n12613 ;
  assign n13538 = n13512 ^ n13505 ;
  assign n13539 = n13538 ^ x26 ;
  assign n13537 = n446 & ~n12367 ;
  assign n13540 = n13539 ^ n13537 ;
  assign n13536 = ~n12108 & n12861 ;
  assign n13541 = n13540 ^ n13536 ;
  assign n13543 = n13542 ^ n13541 ;
  assign n13535 = ~n3501 & n13110 ;
  assign n13544 = n13543 ^ n13535 ;
  assign n13567 = n13508 ^ n13457 ;
  assign n13568 = n13567 ^ n13270 ;
  assign n13569 = n13568 ^ n13451 ;
  assign n13546 = n11972 & n12861 ;
  assign n13545 = n446 & ~n12108 ;
  assign n13547 = n13546 ^ n13545 ;
  assign n13548 = n13547 ^ n65 ;
  assign n13549 = n13547 ^ x26 ;
  assign n13550 = n13549 ^ n67 ;
  assign n13551 = n13550 ^ x25 ;
  assign n13552 = n13551 ^ n12367 ;
  assign n13553 = n13552 ^ n13549 ;
  assign n13554 = n13553 ^ n12277 ;
  assign n13555 = n13554 ^ n13553 ;
  assign n13556 = n13549 & ~n13555 ;
  assign n13557 = n13556 ^ n13550 ;
  assign n13558 = n13553 ^ n12367 ;
  assign n13559 = ~n13555 & ~n13558 ;
  assign n13560 = n13559 ^ n12367 ;
  assign n13561 = ~n13550 & n13560 ;
  assign n13562 = ~n13557 & n13561 ;
  assign n13563 = n13562 ^ n13559 ;
  assign n13564 = n13563 ^ n67 ;
  assign n13565 = n13564 ^ n12367 ;
  assign n13566 = ~n13548 & ~n13565 ;
  assign n13570 = n13569 ^ n13566 ;
  assign n13581 = n3484 & ~n12262 ;
  assign n13577 = n4536 & n13052 ;
  assign n13578 = n13577 ^ n12256 ;
  assign n13579 = n650 & ~n13578 ;
  assign n13580 = n13579 ^ x29 ;
  assign n13582 = n13581 ^ n13580 ;
  assign n13572 = n831 & ~n12220 ;
  assign n13583 = n13582 ^ n13572 ;
  assign n13673 = n13583 ^ n13569 ;
  assign n13571 = n13268 ^ n13207 ;
  assign n13584 = n13583 ^ n13571 ;
  assign n13637 = n1104 ^ n1029 ;
  assign n13635 = n693 ^ n674 ;
  assign n13634 = n1215 ^ n1017 ;
  assign n13636 = n13635 ^ n13634 ;
  assign n13638 = n13637 ^ n13636 ;
  assign n13630 = n394 ^ n300 ;
  assign n13629 = n5223 ^ n143 ;
  assign n13631 = n13630 ^ n13629 ;
  assign n13628 = n1318 ^ n1159 ;
  assign n13632 = n13631 ^ n13628 ;
  assign n13625 = n3603 ^ n1835 ;
  assign n13626 = n13625 ^ n2129 ;
  assign n13627 = n13626 ^ n1635 ;
  assign n13633 = n13632 ^ n13627 ;
  assign n13639 = n13638 ^ n13633 ;
  assign n13640 = n13639 ^ n3190 ;
  assign n13658 = n245 ^ n201 ;
  assign n13659 = n13658 ^ n211 ;
  assign n13660 = n13659 ^ n2397 ;
  assign n13655 = n602 ^ n407 ;
  assign n13653 = n2539 ^ n194 ;
  assign n13654 = n13653 ^ n409 ;
  assign n13656 = n13655 ^ n13654 ;
  assign n13657 = n13656 ^ n3674 ;
  assign n13661 = n13660 ^ n13657 ;
  assign n13649 = n4132 ^ n558 ;
  assign n13647 = n660 ^ n507 ;
  assign n13648 = n13647 ^ n2830 ;
  assign n13650 = n13649 ^ n13648 ;
  assign n13644 = n1366 ^ n1093 ;
  assign n13642 = n12810 ^ n180 ;
  assign n13643 = n13642 ^ n1925 ;
  assign n13645 = n13644 ^ n13643 ;
  assign n13641 = n2594 ^ n1429 ;
  assign n13646 = n13645 ^ n13641 ;
  assign n13651 = n13650 ^ n13646 ;
  assign n13652 = n13651 ^ n3847 ;
  assign n13662 = n13661 ^ n13652 ;
  assign n13663 = ~n13640 & ~n13662 ;
  assign n13605 = n12245 ^ n12213 ;
  assign n13587 = ~n35 & ~n12129 ;
  assign n13617 = n13605 ^ n13587 ;
  assign n13606 = n13605 ^ n12121 ;
  assign n13608 = n13606 ^ n12129 ;
  assign n13607 = n13606 ^ n12130 ;
  assign n13609 = n13608 ^ n13607 ;
  assign n13610 = n13608 ^ x30 ;
  assign n13611 = n13610 ^ n13608 ;
  assign n13612 = ~n13609 & n13611 ;
  assign n13613 = n13612 ^ n13608 ;
  assign n13614 = ~n3520 & n13613 ;
  assign n13615 = n13614 ^ n13606 ;
  assign n13616 = n13615 ^ n13587 ;
  assign n13618 = n13617 ^ n13616 ;
  assign n13619 = n13617 ^ n3520 ;
  assign n13620 = n13619 ^ n13617 ;
  assign n13621 = n13618 & ~n13620 ;
  assign n13622 = n13621 ^ n13617 ;
  assign n13623 = ~x31 & ~n13622 ;
  assign n13624 = n13623 ^ n13615 ;
  assign n13664 = n13663 ^ n13624 ;
  assign n13665 = n13624 ^ n13264 ;
  assign n13666 = ~n13664 & ~n13665 ;
  assign n13667 = n13666 ^ n13250 ;
  assign n13668 = n13666 ^ n13264 ;
  assign n13599 = n12121 ^ n3726 ;
  assign n13600 = n13599 ^ n13587 ;
  assign n13586 = n12246 ^ n12214 ;
  assign n13596 = n13586 ^ n12117 ;
  assign n13597 = n13596 ^ n12121 ;
  assign n13598 = ~n12015 & ~n13597 ;
  assign n13601 = n13600 ^ n13598 ;
  assign n13588 = n13587 ^ n13586 ;
  assign n13589 = n13588 ^ n3726 ;
  assign n13590 = n13589 ^ n13588 ;
  assign n13591 = n13588 ^ n12117 ;
  assign n13592 = n13591 ^ n13588 ;
  assign n13593 = ~n13590 & ~n13592 ;
  assign n13594 = n13593 ^ n13588 ;
  assign n13595 = ~x31 & n13594 ;
  assign n13602 = n13601 ^ n13595 ;
  assign n13585 = ~n35 & n12121 ;
  assign n13603 = n13602 ^ n13585 ;
  assign n13669 = n13668 ^ n13603 ;
  assign n13670 = n13667 & n13669 ;
  assign n13604 = n13603 ^ n13583 ;
  assign n13671 = n13670 ^ n13604 ;
  assign n13672 = ~n13584 & n13671 ;
  assign n13674 = n13673 ^ n13672 ;
  assign n13675 = n13570 & ~n13674 ;
  assign n13676 = n13675 ^ n13569 ;
  assign n13677 = n13676 ^ n13538 ;
  assign n13678 = ~n13544 & n13677 ;
  assign n13679 = n13678 ^ n13538 ;
  assign n13681 = n13680 ^ n13679 ;
  assign n13690 = ~n4496 & n12755 ;
  assign n13683 = n12971 ^ x23 ;
  assign n13684 = n13683 ^ x22 ;
  assign n13685 = n13684 ^ n12971 ;
  assign n13686 = ~n12973 & n13685 ;
  assign n13687 = n13686 ^ n12971 ;
  assign n13688 = n4488 & n13687 ;
  assign n13689 = n13688 ^ x23 ;
  assign n13691 = n13690 ^ n13689 ;
  assign n13682 = n4504 & ~n12705 ;
  assign n13692 = n13691 ^ n13682 ;
  assign n13693 = n13692 ^ n13679 ;
  assign n13694 = ~n13681 & ~n13693 ;
  assign n13695 = n13694 ^ n13679 ;
  assign n13697 = n13534 & n13695 ;
  assign n13696 = n13695 ^ n13534 ;
  assign n13698 = n13697 ^ n13696 ;
  assign n13699 = n13533 & ~n13698 ;
  assign n14000 = n13676 ^ n13544 ;
  assign n13709 = n13674 ^ n13566 ;
  assign n13704 = n4504 & ~n12613 ;
  assign n13703 = n4491 & ~n12705 ;
  assign n13705 = n13704 ^ n13703 ;
  assign n13706 = n13705 ^ x23 ;
  assign n13702 = n4492 & n12706 ;
  assign n13707 = n13706 ^ n13702 ;
  assign n13701 = ~n4496 & n12656 ;
  assign n13708 = n13707 ^ n13701 ;
  assign n13710 = n13709 ^ n13708 ;
  assign n13989 = n12260 & n12861 ;
  assign n13988 = n446 & n11972 ;
  assign n13990 = n13989 ^ n13988 ;
  assign n13991 = n13990 ^ x26 ;
  assign n13987 = ~n487 & ~n12108 ;
  assign n13992 = n13991 ^ n13987 ;
  assign n13986 = ~n3501 & n12376 ;
  assign n13993 = n13992 ^ n13986 ;
  assign n13996 = n13993 ^ n13709 ;
  assign n13984 = n13671 ^ n13571 ;
  assign n13967 = n13664 ^ n13264 ;
  assign n13762 = n12452 ^ n3267 ;
  assign n13761 = n1009 ^ n581 ;
  assign n13763 = n13762 ^ n13761 ;
  assign n13758 = n1739 ^ n663 ;
  assign n13757 = n12509 ^ n1482 ;
  assign n13759 = n13758 ^ n13757 ;
  assign n13754 = n673 ^ n282 ;
  assign n13755 = n13754 ^ n176 ;
  assign n13752 = n1650 ^ n109 ;
  assign n13753 = n13752 ^ n625 ;
  assign n13756 = n13755 ^ n13753 ;
  assign n13760 = n13759 ^ n13756 ;
  assign n13764 = n13763 ^ n13760 ;
  assign n13765 = n13764 ^ n3447 ;
  assign n13766 = n5312 ^ n1831 ;
  assign n13767 = n13766 ^ n1211 ;
  assign n13768 = ~n13765 & ~n13767 ;
  assign n13769 = n13768 ^ n6653 ;
  assign n13778 = n2228 ^ n217 ;
  assign n13775 = n1116 ^ n141 ;
  assign n13773 = n607 ^ n560 ;
  assign n13774 = n13773 ^ n3215 ;
  assign n13776 = n13775 ^ n13774 ;
  assign n13770 = n773 ^ n255 ;
  assign n13771 = n13770 ^ n1473 ;
  assign n13772 = n13771 ^ n1059 ;
  assign n13777 = n13776 ^ n13772 ;
  assign n13779 = n13778 ^ n13777 ;
  assign n13795 = n5257 ^ n848 ;
  assign n13794 = n1383 ^ n774 ;
  assign n13796 = n13795 ^ n13794 ;
  assign n13791 = n1078 ^ n260 ;
  assign n13790 = n5129 ^ n1476 ;
  assign n13792 = n13791 ^ n13790 ;
  assign n13789 = n3630 ^ n2200 ;
  assign n13793 = n13792 ^ n13789 ;
  assign n13797 = n13796 ^ n13793 ;
  assign n13786 = n2586 ^ n1305 ;
  assign n13785 = n1739 ^ n228 ;
  assign n13787 = n13786 ^ n13785 ;
  assign n13783 = n1494 ^ n129 ;
  assign n13780 = n1104 ^ n933 ;
  assign n13781 = n13780 ^ n356 ;
  assign n13782 = n13781 ^ n838 ;
  assign n13784 = n13783 ^ n13782 ;
  assign n13788 = n13787 ^ n13784 ;
  assign n13798 = n13797 ^ n13788 ;
  assign n13799 = n13798 ^ n5588 ;
  assign n13800 = ~n3282 & ~n13799 ;
  assign n13801 = ~n13779 & n13800 ;
  assign n13802 = n13801 ^ n6653 ;
  assign n13803 = n13769 & n13802 ;
  assign n13804 = n13803 ^ n6653 ;
  assign n13805 = n13804 ^ n13264 ;
  assign n13749 = ~n3724 & n12130 ;
  assign n13748 = n3726 & ~n12129 ;
  assign n13750 = n13749 ^ n13748 ;
  assign n13736 = n12244 ^ n12212 ;
  assign n13737 = n13736 ^ n12129 ;
  assign n13739 = n13737 ^ n12130 ;
  assign n13738 = n13737 ^ n12136 ;
  assign n13740 = n13739 ^ n13738 ;
  assign n13743 = x30 & ~n13740 ;
  assign n13744 = n13743 ^ n13739 ;
  assign n13745 = ~n3520 & n13744 ;
  assign n13746 = n13745 ^ n13737 ;
  assign n13747 = x31 & n13746 ;
  assign n13751 = n13750 ^ n13747 ;
  assign n13806 = n13805 ^ n13751 ;
  assign n13733 = n3484 & n12117 ;
  assign n13726 = n12110 ^ x29 ;
  assign n13727 = n13726 ^ x28 ;
  assign n13728 = n13727 ^ n12110 ;
  assign n13729 = ~n13195 & n13728 ;
  assign n13730 = n13729 ^ n12110 ;
  assign n13731 = n650 & ~n13730 ;
  assign n13732 = n13731 ^ x29 ;
  assign n13734 = n13733 ^ n13732 ;
  assign n13724 = n831 & n12121 ;
  assign n13735 = n13734 ^ n13724 ;
  assign n13807 = n13806 ^ n13735 ;
  assign n13817 = n12243 ^ n12211 ;
  assign n13818 = n13817 ^ n12130 ;
  assign n13820 = n13818 ^ n12137 ;
  assign n13819 = n13818 ^ n12136 ;
  assign n13821 = n13820 ^ n13819 ;
  assign n13824 = ~x30 & ~n13821 ;
  assign n13825 = n13824 ^ n13820 ;
  assign n13826 = ~n3520 & ~n13825 ;
  assign n13827 = n13826 ^ n13818 ;
  assign n13828 = x31 & ~n13827 ;
  assign n13809 = n12136 ^ n12130 ;
  assign n13814 = ~n35 & ~n13809 ;
  assign n13815 = n13814 ^ n12130 ;
  assign n13816 = ~n3514 & n13815 ;
  assign n13829 = n13828 ^ n13816 ;
  assign n13963 = n13829 ^ n13806 ;
  assign n13808 = n13801 ^ n13769 ;
  assign n13830 = n13829 ^ n13808 ;
  assign n13847 = n1494 ^ n1059 ;
  assign n13846 = n1036 ^ n751 ;
  assign n13848 = n13847 ^ n13846 ;
  assign n13844 = n1176 ^ n99 ;
  assign n13842 = n1758 ^ n841 ;
  assign n13843 = n13842 ^ n732 ;
  assign n13845 = n13844 ^ n13843 ;
  assign n13849 = n13848 ^ n13845 ;
  assign n13838 = n867 ^ n745 ;
  assign n13837 = n1516 ^ n513 ;
  assign n13839 = n13838 ^ n13837 ;
  assign n13840 = n13839 ^ n686 ;
  assign n13834 = n12539 ^ n1898 ;
  assign n13835 = n13834 ^ n2069 ;
  assign n13832 = n5359 ^ n848 ;
  assign n13831 = n12509 ^ n1956 ;
  assign n13833 = n13832 ^ n13831 ;
  assign n13836 = n13835 ^ n13833 ;
  assign n13841 = n13840 ^ n13836 ;
  assign n13850 = n13849 ^ n13841 ;
  assign n13851 = n13850 ^ n2535 ;
  assign n13863 = n1372 ^ n811 ;
  assign n13864 = n13863 ^ n1041 ;
  assign n13860 = n13034 ^ n2114 ;
  assign n13859 = n1405 ^ n1250 ;
  assign n13861 = n13860 ^ n13859 ;
  assign n13858 = n13628 ^ n1453 ;
  assign n13862 = n13861 ^ n13858 ;
  assign n13865 = n13864 ^ n13862 ;
  assign n13853 = n2037 ^ n360 ;
  assign n13854 = n13853 ^ n1408 ;
  assign n13852 = n3259 ^ n362 ;
  assign n13855 = n13854 ^ n13852 ;
  assign n13856 = n13855 ^ n2909 ;
  assign n13857 = n13856 ^ n2820 ;
  assign n13866 = n13865 ^ n13857 ;
  assign n13867 = n13866 ^ n4227 ;
  assign n13868 = ~n13851 & ~n13867 ;
  assign n13899 = ~n18156 ^ n7144 ;
  assign n13900 = n13899 ^ n7138 ;
  assign n13869 = n12058 ^ n1867 ;
  assign n13892 = n2325 ^ n225 ;
  assign n13893 = n13892 ^ n1311 ;
  assign n13894 = n13893 ^ n2191 ;
  assign n13890 = n2228 ^ n130 ;
  assign n13891 = n13890 ^ n1534 ;
  assign n13895 = n13894 ^ n13891 ;
  assign n13896 = n13895 ^ n2566 ;
  assign n13885 = n1494 ^ n229 ;
  assign n13886 = n13885 ^ n2677 ;
  assign n13883 = n567 ^ n109 ;
  assign n13884 = n13883 ^ n1343 ;
  assign n13887 = n13886 ^ n13884 ;
  assign n13880 = n526 ^ n409 ;
  assign n13881 = n13880 ^ n1809 ;
  assign n13879 = n1956 ^ n835 ;
  assign n13882 = n13881 ^ n13879 ;
  assign n13888 = n13887 ^ n13882 ;
  assign n13874 = n773 ^ n391 ;
  assign n13875 = n13874 ^ n1157 ;
  assign n13876 = n13875 ^ n2334 ;
  assign n13872 = n1058 ^ n265 ;
  assign n13870 = n362 ^ n270 ;
  assign n13871 = n13870 ^ n547 ;
  assign n13873 = n13872 ^ n13871 ;
  assign n13877 = n13876 ^ n13873 ;
  assign n13878 = n13877 ^ n5637 ;
  assign n13889 = n13888 ^ n13878 ;
  assign n13897 = n13896 ^ n13889 ;
  assign n13898 = ~n13869 & ~n13897 ;
  assign n13901 = n13900 ^ n13898 ;
  assign n13930 = n12834 ^ n621 ;
  assign n13927 = n3128 ^ n1260 ;
  assign n13925 = n810 ^ n183 ;
  assign n13924 = n931 ^ n221 ;
  assign n13926 = n13925 ^ n13924 ;
  assign n13928 = n13927 ^ n13926 ;
  assign n13919 = n2511 ^ n720 ;
  assign n13920 = n13919 ^ n987 ;
  assign n13917 = n2544 ^ n579 ;
  assign n13916 = n12035 ^ n940 ;
  assign n13918 = n13917 ^ n13916 ;
  assign n13921 = n13920 ^ n13918 ;
  assign n13913 = n4217 ^ n899 ;
  assign n13912 = n1159 ^ n1100 ;
  assign n13914 = n13913 ^ n13912 ;
  assign n13915 = n13914 ^ n3627 ;
  assign n13922 = n13921 ^ n13915 ;
  assign n13909 = n1428 ^ n1206 ;
  assign n13908 = n2713 ^ n1500 ;
  assign n13910 = n13909 ^ n13908 ;
  assign n13905 = n11828 ^ n932 ;
  assign n13902 = n981 ^ n88 ;
  assign n13903 = n13902 ^ n702 ;
  assign n13904 = n13903 ^ n1931 ;
  assign n13906 = n13905 ^ n13904 ;
  assign n13907 = n13906 ^ n4102 ;
  assign n13911 = n13910 ^ n13907 ;
  assign n13923 = n13922 ^ n13911 ;
  assign n13929 = n13928 ^ n13923 ;
  assign n13931 = n13930 ^ n13929 ;
  assign n13932 = ~n3533 & ~n13931 ;
  assign n13933 = n13932 ^ n13900 ;
  assign n13934 = n13901 & n13933 ;
  assign n13935 = n13934 ^ n13900 ;
  assign n13951 = ~n12207 & n24214 ;
  assign n13949 = ~n35 & n12138 ;
  assign n13936 = n12241 ^ n12209 ;
  assign n13939 = n13936 ^ n12137 ;
  assign n13946 = n13939 ^ n12138 ;
  assign n13947 = ~n12015 & n13946 ;
  assign n13944 = n12138 ^ n3724 ;
  assign n13937 = n13936 ^ n3726 ;
  assign n13938 = n13937 ^ n13936 ;
  assign n13940 = n13939 ^ n13936 ;
  assign n13941 = ~n13938 & n13940 ;
  assign n13942 = n13941 ^ n13936 ;
  assign n13943 = ~x31 & ~n13942 ;
  assign n13945 = n13944 ^ n13943 ;
  assign n13948 = n13947 ^ n13945 ;
  assign n13950 = n13949 ^ n13948 ;
  assign n13952 = n13951 ^ n13950 ;
  assign n13953 = ~n13935 & n13952 ;
  assign n13954 = ~n13801 & ~n13953 ;
  assign n13955 = ~n13868 & ~n13954 ;
  assign n13956 = n13952 ^ n13935 ;
  assign n13957 = n13956 ^ n13953 ;
  assign n13958 = n13801 & ~n13957 ;
  assign n13959 = n13955 & ~n13958 ;
  assign n13960 = n13959 ^ n13958 ;
  assign n13961 = n13960 ^ n13829 ;
  assign n13962 = ~n13830 & n13961 ;
  assign n13964 = n13963 ^ n13962 ;
  assign n13965 = ~n13807 & ~n13964 ;
  assign n13966 = n13965 ^ n13806 ;
  assign n13968 = n13967 ^ n13966 ;
  assign n13969 = n13966 ^ n13751 ;
  assign n13970 = n13969 ^ n13664 ;
  assign n13971 = n13804 ^ n13751 ;
  assign n13974 = n13970 & n13971 ;
  assign n13975 = n13974 ^ n13664 ;
  assign n13976 = ~n13968 & n13975 ;
  assign n13977 = n13976 ^ n13967 ;
  assign n13721 = n3484 & ~n12220 ;
  assign n13712 = n12262 ^ n12250 ;
  assign n13713 = n13712 ^ n12262 ;
  assign n13714 = n12262 ^ x29 ;
  assign n13715 = n13714 ^ x28 ;
  assign n13716 = n13715 ^ n12262 ;
  assign n13717 = ~n13713 & n13716 ;
  assign n13718 = n13717 ^ n12262 ;
  assign n13719 = n650 & ~n13718 ;
  assign n13720 = n13719 ^ x29 ;
  assign n13722 = n13721 ^ n13720 ;
  assign n13711 = n831 & ~n12110 ;
  assign n13723 = n13722 ^ n13711 ;
  assign n13978 = n13977 ^ n13723 ;
  assign n13979 = n13603 ^ n13250 ;
  assign n13980 = n13979 ^ n13723 ;
  assign n13981 = n13980 ^ n13666 ;
  assign n13982 = n13978 & n13981 ;
  assign n13983 = n13982 ^ n13977 ;
  assign n13985 = n13984 ^ n13983 ;
  assign n13994 = n13993 ^ n13983 ;
  assign n13995 = n13985 & n13994 ;
  assign n13997 = n13996 ^ n13995 ;
  assign n13998 = n13710 & n13997 ;
  assign n13999 = n13998 ^ n13709 ;
  assign n14001 = n14000 ^ n13999 ;
  assign n14003 = n4504 & n12656 ;
  assign n14002 = ~n4496 & ~n12705 ;
  assign n14004 = n14003 ^ n14002 ;
  assign n14006 = n14005 ^ n14004 ;
  assign n14018 = n12724 & n14008 ;
  assign n14009 = n14004 ^ x23 ;
  assign n14010 = n14009 ^ n14008 ;
  assign n14011 = n12755 ^ x22 ;
  assign n14012 = n14011 ^ n12755 ;
  assign n14015 = ~n12757 & ~n14012 ;
  assign n14016 = n14015 ^ n12755 ;
  assign n14017 = n14010 & ~n14016 ;
  assign n14019 = n14018 ^ n14017 ;
  assign n14020 = ~n14006 & ~n14019 ;
  assign n14021 = n14020 ^ n13999 ;
  assign n14022 = ~n14001 & ~n14021 ;
  assign n14023 = n14022 ^ n14020 ;
  assign n13700 = n13692 ^ n13681 ;
  assign n14024 = n14023 ^ n13700 ;
  assign n14029 = n14023 ^ n8212 ;
  assign n14028 = n12855 & n14027 ;
  assign n14030 = n14029 ^ n14028 ;
  assign n14031 = n14024 & ~n14030 ;
  assign n14032 = n14031 ^ n14023 ;
  assign n14034 = n14032 ^ n8212 ;
  assign n14033 = ~n8212 & n14032 ;
  assign n14035 = n14034 ^ n14033 ;
  assign n14205 = n12755 & n14027 ;
  assign n14204 = n4916 & n12971 ;
  assign n14206 = n14205 ^ n14204 ;
  assign n14207 = n14206 ^ x20 ;
  assign n14203 = n4678 & ~n12855 ;
  assign n14208 = n14207 ^ n14203 ;
  assign n14209 = n14208 ^ n14207 ;
  assign n14210 = n4685 & ~n13007 ;
  assign n14211 = n14209 & n14210 ;
  assign n14212 = n14211 ^ n14208 ;
  assign n14087 = n13981 ^ n13977 ;
  assign n14082 = ~n12256 & n12861 ;
  assign n14081 = n446 & n12260 ;
  assign n14083 = n14082 ^ n14081 ;
  assign n14084 = n14083 ^ x26 ;
  assign n14080 = ~n487 & n11972 ;
  assign n14085 = n14084 ^ n14080 ;
  assign n14078 = n13073 ^ n12260 ;
  assign n14079 = ~n3501 & ~n14078 ;
  assign n14086 = n14085 ^ n14079 ;
  assign n14088 = n14087 ^ n14086 ;
  assign n14167 = n13993 ^ n13985 ;
  assign n14168 = n14167 ^ n14086 ;
  assign n14169 = n14168 ^ n14167 ;
  assign n14059 = n3484 & ~n12110 ;
  assign n14055 = ~n13805 & n13971 ;
  assign n14054 = n13966 ^ n13664 ;
  assign n14056 = n14055 ^ n14054 ;
  assign n14057 = n14056 ^ x29 ;
  assign n14047 = n13172 ^ n12220 ;
  assign n14049 = n14047 ^ n4536 ;
  assign n14050 = n14049 ^ n14047 ;
  assign n14051 = ~n13172 & ~n14050 ;
  assign n14052 = n14051 ^ n14047 ;
  assign n14053 = n650 & n14052 ;
  assign n14058 = n14057 ^ n14053 ;
  assign n14060 = n14059 ^ n14058 ;
  assign n14046 = n831 & n12117 ;
  assign n14061 = n14060 ^ n14046 ;
  assign n14063 = ~n12262 & n12861 ;
  assign n14062 = n446 & ~n12256 ;
  assign n14064 = n14063 ^ n14062 ;
  assign n14065 = n14064 ^ n65 ;
  assign n14066 = n14064 ^ x26 ;
  assign n14070 = n14066 ^ n67 ;
  assign n14071 = ~x25 & n13053 ;
  assign n14072 = n14070 & n14071 ;
  assign n13054 = n13053 ^ n12260 ;
  assign n14068 = n67 & n13054 ;
  assign n14067 = ~n12260 & n14066 ;
  assign n14069 = n14068 ^ n14067 ;
  assign n14073 = n14072 ^ n14069 ;
  assign n14074 = ~n14065 & ~n14073 ;
  assign n14075 = n14074 ^ n14056 ;
  assign n14076 = n14061 & n14075 ;
  assign n14077 = n14076 ^ n14074 ;
  assign n14170 = n14169 ^ n14077 ;
  assign n14171 = ~n14088 & ~n14170 ;
  assign n14172 = n14171 ^ n14168 ;
  assign n14197 = n13997 ^ n13708 ;
  assign n14199 = n14197 ^ n14167 ;
  assign n14179 = ~n4496 & ~n12613 ;
  assign n14177 = n4492 & ~n12872 ;
  assign n14174 = n4504 & ~n12367 ;
  assign n14173 = n4491 & n12656 ;
  assign n14175 = n14174 ^ n14173 ;
  assign n14176 = n14175 ^ x23 ;
  assign n14178 = n14177 ^ n14176 ;
  assign n14180 = n14179 ^ n14178 ;
  assign n14198 = n14197 ^ n14180 ;
  assign n14200 = n14199 ^ n14198 ;
  assign n14201 = ~n14172 & ~n14200 ;
  assign n14202 = n14201 ^ n14199 ;
  assign n14213 = n14212 ^ n14202 ;
  assign n14181 = n14180 ^ n14172 ;
  assign n14089 = n14088 ^ n14077 ;
  assign n14044 = ~n4496 & ~n12367 ;
  assign n14042 = n4492 & n13110 ;
  assign n14039 = n4504 & ~n12108 ;
  assign n14038 = n4491 & ~n12613 ;
  assign n14040 = n14039 ^ n14038 ;
  assign n14041 = n14040 ^ x23 ;
  assign n14043 = n14042 ^ n14041 ;
  assign n14045 = n14044 ^ n14043 ;
  assign n14090 = n14089 ^ n14045 ;
  assign n14099 = n14074 ^ n14061 ;
  assign n14094 = n4504 & n11972 ;
  assign n14093 = n4491 & ~n12367 ;
  assign n14095 = n14094 ^ n14093 ;
  assign n14096 = n14095 ^ x23 ;
  assign n14092 = n4492 & n12368 ;
  assign n14097 = n14096 ^ n14092 ;
  assign n14091 = ~n4496 & ~n12108 ;
  assign n14098 = n14097 ^ n14091 ;
  assign n14100 = n14099 ^ n14098 ;
  assign n14109 = n13964 ^ n13735 ;
  assign n14160 = n14109 ^ n14099 ;
  assign n14104 = ~n12220 & n12861 ;
  assign n14103 = n446 & ~n12262 ;
  assign n14105 = n14104 ^ n14103 ;
  assign n14106 = n14105 ^ x26 ;
  assign n14102 = ~n487 & ~n12256 ;
  assign n14107 = n14106 ^ n14102 ;
  assign n14101 = ~n3501 & ~n13283 ;
  assign n14108 = n14107 ^ n14101 ;
  assign n14110 = n14109 ^ n14108 ;
  assign n14124 = n13960 ^ n13830 ;
  assign n14120 = n3484 & n12121 ;
  assign n14113 = n12117 ^ x29 ;
  assign n14114 = n14113 ^ x28 ;
  assign n14115 = n14114 ^ n12117 ;
  assign n14116 = ~n13586 & n14115 ;
  assign n14117 = n14116 ^ n12117 ;
  assign n14118 = n650 & n14117 ;
  assign n14119 = n14118 ^ x29 ;
  assign n14121 = n14120 ^ n14119 ;
  assign n14111 = n831 & ~n12129 ;
  assign n14122 = n14121 ^ n14111 ;
  assign n14125 = n14124 ^ n14122 ;
  assign n14137 = ~n3733 & n12137 ;
  assign n14128 = n12242 ^ n12210 ;
  assign n14129 = n14128 ^ n12136 ;
  assign n14134 = n14129 ^ n12138 ;
  assign n14135 = ~n14134 & n24214 ;
  assign n14132 = n4851 & n14129 ;
  assign n14130 = n14129 ^ n14128 ;
  assign n14131 = n3726 & ~n14130 ;
  assign n14133 = n14132 ^ n14131 ;
  assign n14136 = n14135 ^ n14133 ;
  assign n14138 = n14137 ^ n14136 ;
  assign n14126 = n13958 ^ n13954 ;
  assign n14127 = n14126 ^ n13868 ;
  assign n14139 = n14138 ^ n14127 ;
  assign n14141 = n831 & n12130 ;
  assign n14140 = n3484 & ~n12129 ;
  assign n14142 = n14141 ^ n14140 ;
  assign n14143 = n14142 ^ n651 ;
  assign n14145 = n14142 ^ x29 ;
  assign n14148 = n14145 ^ n653 ;
  assign n14149 = ~x28 & ~n13605 ;
  assign n14150 = n14148 & n14149 ;
  assign n14146 = ~n12121 & n14145 ;
  assign n14144 = n653 & ~n13606 ;
  assign n14147 = n14146 ^ n14144 ;
  assign n14151 = n14150 ^ n14147 ;
  assign n14152 = ~n14143 & ~n14151 ;
  assign n14153 = n14152 ^ n14138 ;
  assign n14154 = n14139 & ~n14153 ;
  assign n14155 = n14154 ^ n14138 ;
  assign n14156 = n14155 ^ n14122 ;
  assign n14157 = ~n14125 & n14156 ;
  assign n14123 = n14122 ^ n14108 ;
  assign n14158 = n14157 ^ n14123 ;
  assign n14159 = ~n14110 & ~n14158 ;
  assign n14161 = n14160 ^ n14159 ;
  assign n14162 = n14100 & ~n14161 ;
  assign n14163 = n14162 ^ n14099 ;
  assign n14164 = n14163 ^ n14045 ;
  assign n14165 = n14090 & n14164 ;
  assign n14166 = n14165 ^ n14045 ;
  assign n14182 = n14181 ^ n14166 ;
  assign n14191 = ~n12705 & n14027 ;
  assign n14184 = n12971 ^ x20 ;
  assign n14185 = n14184 ^ x19 ;
  assign n14186 = n14185 ^ n12971 ;
  assign n14187 = ~n12973 & n14186 ;
  assign n14188 = n14187 ^ n12971 ;
  assign n14189 = n4678 & n14188 ;
  assign n14190 = n14189 ^ x20 ;
  assign n14192 = n14191 ^ n14190 ;
  assign n14183 = n4916 & n12755 ;
  assign n14193 = n14192 ^ n14183 ;
  assign n14194 = n14193 ^ n14166 ;
  assign n14195 = ~n14182 & n14194 ;
  assign n14196 = n14195 ^ n14166 ;
  assign n14214 = n14213 ^ n14196 ;
  assign n14215 = n14196 ^ n5710 ;
  assign n14216 = ~n14214 & ~n14215 ;
  assign n14217 = n14216 ^ n14213 ;
  assign n14037 = n14020 ^ n14001 ;
  assign n20778 = n14217 ^ n14037 ;
  assign n14218 = n14037 & n14217 ;
  assign n20779 = n20778 ^ n14218 ;
  assign n14036 = n14030 ^ n13700 ;
  assign n14219 = n14218 ^ n14036 ;
  assign n20740 = n14215 ^ n14213 ;
  assign n14405 = n14161 ^ n14098 ;
  assign n14246 = n14158 ^ n14109 ;
  assign n14244 = ~n4496 & n11972 ;
  assign n14242 = n4492 & n12376 ;
  assign n14239 = n4504 & n12260 ;
  assign n14238 = n4491 & ~n12108 ;
  assign n14240 = n14239 ^ n14238 ;
  assign n14241 = n14240 ^ x23 ;
  assign n14243 = n14242 ^ n14241 ;
  assign n14245 = n14244 ^ n14243 ;
  assign n14247 = n14246 ^ n14245 ;
  assign n14249 = n14155 ^ n14125 ;
  assign n14401 = n14249 ^ n14246 ;
  assign n14256 = ~n3501 & n13712 ;
  assign n14253 = ~n487 & ~n12262 ;
  assign n14251 = n446 & ~n12220 ;
  assign n14250 = n14249 ^ x26 ;
  assign n14252 = n14251 ^ n14250 ;
  assign n14254 = n14253 ^ n14252 ;
  assign n14248 = ~n12110 & n12861 ;
  assign n14255 = n14254 ^ n14248 ;
  assign n14257 = n14256 ^ n14255 ;
  assign n14266 = n14153 ^ n14127 ;
  assign n14261 = n12117 & n12861 ;
  assign n14260 = n446 & ~n12110 ;
  assign n14262 = n14261 ^ n14260 ;
  assign n14263 = n14262 ^ x26 ;
  assign n14259 = ~n487 & ~n12220 ;
  assign n14264 = n14263 ^ n14259 ;
  assign n14258 = ~n3501 & n14047 ;
  assign n14265 = n14264 ^ n14258 ;
  assign n14267 = n14266 ^ n14265 ;
  assign n14279 = n3484 & n12130 ;
  assign n14271 = n13737 ^ n12129 ;
  assign n14272 = n12129 ^ x29 ;
  assign n14273 = n14272 ^ x28 ;
  assign n14274 = n14273 ^ n12129 ;
  assign n14275 = ~n14271 & n14274 ;
  assign n14276 = n14275 ^ n12129 ;
  assign n14277 = n650 & ~n14276 ;
  assign n14278 = n14277 ^ x29 ;
  assign n14280 = n14279 ^ n14278 ;
  assign n14270 = n831 & ~n12136 ;
  assign n14281 = n14280 ^ n14270 ;
  assign n14395 = n14281 ^ n14266 ;
  assign n14268 = n13935 ^ n13801 ;
  assign n14269 = n14268 ^ n13952 ;
  assign n14282 = n14281 ^ n14269 ;
  assign n14365 = n13932 ^ n13901 ;
  assign n14291 = n3542 ^ n1202 ;
  assign n14290 = n12794 ^ n1835 ;
  assign n14292 = n14291 ^ n14290 ;
  assign n14288 = n13773 ^ n309 ;
  assign n14289 = n14288 ^ n2114 ;
  assign n14293 = n14292 ^ n14289 ;
  assign n14294 = n14293 ^ n750 ;
  assign n14284 = n1739 ^ n1050 ;
  assign n14285 = n14284 ^ n2215 ;
  assign n14283 = n3755 ^ n2627 ;
  assign n14286 = n14285 ^ n14283 ;
  assign n14287 = n14286 ^ n700 ;
  assign n14295 = n14294 ^ n14287 ;
  assign n14296 = n14295 ^ n2395 ;
  assign n14297 = ~n2552 & ~n14296 ;
  assign n14311 = ~n3724 & n12143 ;
  assign n14310 = n3726 & ~n12142 ;
  assign n14312 = n14311 ^ n14310 ;
  assign n14298 = n12238 ^ n12199 ;
  assign n14299 = n14298 ^ n12142 ;
  assign n14301 = n14299 ^ n12143 ;
  assign n14300 = n14299 ^ n12149 ;
  assign n14302 = n14301 ^ n14300 ;
  assign n14305 = x30 & n14302 ;
  assign n14306 = n14305 ^ n14301 ;
  assign n14307 = ~n3520 & n14306 ;
  assign n14308 = n14307 ^ n14299 ;
  assign n14309 = x31 & n14308 ;
  assign n14313 = n14312 ^ n14309 ;
  assign n14315 = ~x2 & ~n11240 ;
  assign n14314 = n9091 ^ x5 ;
  assign n14316 = n14315 ^ n14314 ;
  assign n14335 = n12460 ^ n1172 ;
  assign n14336 = n14335 ^ n12308 ;
  assign n14333 = n3655 ^ n1130 ;
  assign n14334 = n14333 ^ n2667 ;
  assign n14337 = n14336 ^ n14334 ;
  assign n14330 = n1197 ^ n1036 ;
  assign n14331 = n14330 ^ n782 ;
  assign n14332 = n14331 ^ n13843 ;
  assign n14338 = n14337 ^ n14332 ;
  assign n14326 = n5369 ^ n231 ;
  assign n14324 = n2303 ^ n937 ;
  assign n14323 = n1457 ^ n244 ;
  assign n14325 = n14324 ^ n14323 ;
  assign n14327 = n14326 ^ n14325 ;
  assign n14320 = n12401 ^ n2037 ;
  assign n14321 = n14320 ^ n4371 ;
  assign n14322 = n14321 ^ n807 ;
  assign n14328 = n14327 ^ n14322 ;
  assign n14317 = n13242 ^ n4209 ;
  assign n14318 = n14317 ^ n11896 ;
  assign n14319 = n14318 ^ n3044 ;
  assign n14329 = n14328 ^ n14319 ;
  assign n14339 = n14338 ^ n14329 ;
  assign n14347 = n2111 ^ n527 ;
  assign n14344 = n952 ^ n122 ;
  assign n14345 = n14344 ^ n363 ;
  assign n14346 = n14345 ^ n1142 ;
  assign n14348 = n14347 ^ n14346 ;
  assign n14349 = n14348 ^ n5559 ;
  assign n14340 = n3651 ^ n1188 ;
  assign n14341 = n14340 ^ n3799 ;
  assign n14342 = n14341 ^ n6369 ;
  assign n14343 = n14342 ^ n3970 ;
  assign n14350 = n14349 ^ n14343 ;
  assign n14351 = n14350 ^ n13779 ;
  assign n14352 = ~n14339 & ~n14351 ;
  assign n14353 = n14352 ^ n14314 ;
  assign n14354 = ~n14316 & n14353 ;
  assign n14355 = n14354 ^ n14315 ;
  assign n14356 = n14313 & ~n14355 ;
  assign n14357 = ~n13932 & ~n14356 ;
  assign n14358 = ~n14297 & ~n14357 ;
  assign n14359 = n14355 ^ n14313 ;
  assign n14360 = n14359 ^ n14356 ;
  assign n14361 = n13932 & ~n14360 ;
  assign n14362 = n14358 & ~n14361 ;
  assign n14363 = n14362 ^ n14361 ;
  assign n14366 = n14365 ^ n14363 ;
  assign n14388 = ~n3724 & n12207 ;
  assign n14387 = n3726 & ~n12138 ;
  assign n14389 = n14388 ^ n14387 ;
  assign n14379 = n12240 ^ n12138 ;
  assign n14382 = n33 & ~n14379 ;
  assign n14383 = n14382 ^ n12138 ;
  assign n14384 = n3722 & n14383 ;
  assign n14367 = x31 & ~n12142 ;
  assign n14385 = n14384 ^ n14367 ;
  assign n14368 = n12239 ^ n12208 ;
  assign n14369 = n14368 ^ n12240 ;
  assign n14370 = n14369 ^ n12239 ;
  assign n14371 = n14370 ^ n14367 ;
  assign n14376 = n33 & n14367 ;
  assign n14377 = n14376 ^ n3722 ;
  assign n14378 = n14371 & n14377 ;
  assign n14386 = n14385 ^ n14378 ;
  assign n14390 = n14389 ^ n14386 ;
  assign n14391 = n14390 ^ n14363 ;
  assign n14392 = ~n14366 & n14391 ;
  assign n14364 = n14363 ^ n14269 ;
  assign n14393 = n14392 ^ n14364 ;
  assign n14394 = ~n14282 & n14393 ;
  assign n14396 = n14395 ^ n14394 ;
  assign n14397 = ~n14267 & ~n14396 ;
  assign n14398 = n14397 ^ n14266 ;
  assign n14399 = n14398 ^ n14249 ;
  assign n14400 = ~n14257 & n14399 ;
  assign n14402 = n14401 ^ n14400 ;
  assign n14403 = ~n14247 & n14402 ;
  assign n14404 = n14403 ^ n14246 ;
  assign n14406 = n14405 ^ n14404 ;
  assign n14415 = n4916 & n12656 ;
  assign n14408 = n12705 ^ x20 ;
  assign n14409 = n14408 ^ x19 ;
  assign n14410 = n14409 ^ n12705 ;
  assign n14411 = ~n12707 & n14410 ;
  assign n14412 = n14411 ^ n12705 ;
  assign n14413 = n4678 & ~n14412 ;
  assign n14414 = n14413 ^ x20 ;
  assign n14416 = n14415 ^ n14414 ;
  assign n14407 = ~n12613 & n14027 ;
  assign n14417 = n14416 ^ n14407 ;
  assign n14418 = n14417 ^ n14404 ;
  assign n14419 = ~n14406 & ~n14418 ;
  assign n14420 = n14419 ^ n14417 ;
  assign n14236 = n4916 & ~n12705 ;
  assign n14233 = n4684 & ~n12756 ;
  assign n14231 = n12656 & n14027 ;
  assign n14229 = n14163 ^ n14090 ;
  assign n14230 = n14229 ^ x20 ;
  assign n14232 = n14231 ^ n14230 ;
  assign n14234 = n14233 ^ n14232 ;
  assign n14228 = n4683 & n12755 ;
  assign n14235 = n14234 ^ n14228 ;
  assign n14237 = n14236 ^ n14235 ;
  assign n14684 = n14420 ^ n14237 ;
  assign n14680 = n5693 ^ x17 ;
  assign n14679 = n5703 & ~n14221 ;
  assign n14681 = n14680 ^ n14679 ;
  assign n14678 = n12971 & n20731 ;
  assign n14682 = n14681 ^ n14678 ;
  assign n14677 = n5700 & ~n12855 ;
  assign n14683 = n14682 ^ n14677 ;
  assign n14685 = n14684 ^ n14683 ;
  assign n14434 = n14417 ^ n14406 ;
  assign n14426 = n5693 & ~n12855 ;
  assign n14427 = n14426 ^ x17 ;
  assign n14428 = n14427 ^ x16 ;
  assign n14429 = ~n13007 & n14426 ;
  assign n14430 = ~n14428 & n14429 ;
  assign n14431 = n14430 ^ n14427 ;
  assign n14425 = n12755 & n20731 ;
  assign n14432 = n14431 ^ n14425 ;
  assign n14424 = n5700 & n12971 ;
  assign n14433 = n14432 ^ n14424 ;
  assign n14435 = n14434 ^ n14433 ;
  assign n14446 = ~n12367 & n14027 ;
  assign n14439 = n12656 ^ x20 ;
  assign n14440 = n14439 ^ x19 ;
  assign n14441 = n14440 ^ n12656 ;
  assign n14442 = ~n12871 & n14441 ;
  assign n14443 = n14442 ^ n12656 ;
  assign n14444 = n4678 & n14443 ;
  assign n14445 = n14444 ^ x20 ;
  assign n14447 = n14446 ^ n14445 ;
  assign n14438 = n4916 & ~n12613 ;
  assign n14448 = n14447 ^ n14438 ;
  assign n14436 = n14402 ^ n14245 ;
  assign n14449 = n14448 ^ n14436 ;
  assign n14462 = n14390 ^ n14366 ;
  assign n14459 = n3484 & ~n12136 ;
  assign n14452 = n12130 ^ x29 ;
  assign n14453 = n14452 ^ x28 ;
  assign n14454 = n14453 ^ n12130 ;
  assign n14455 = ~n13817 & n14454 ;
  assign n14456 = n14455 ^ n12130 ;
  assign n14457 = n650 & n14456 ;
  assign n14458 = n14457 ^ x29 ;
  assign n14460 = n14459 ^ n14458 ;
  assign n14450 = n831 & n12137 ;
  assign n14461 = n14460 ^ n14450 ;
  assign n14463 = n14462 ^ n14461 ;
  assign n14476 = n12239 ^ n12200 ;
  assign n14478 = n14476 ^ n14367 ;
  assign n14479 = n14478 ^ n12207 ;
  assign n14480 = n3520 & ~n14479 ;
  assign n14477 = n3726 & ~n14476 ;
  assign n14481 = n14480 ^ n14477 ;
  assign n14482 = n14481 ^ n14367 ;
  assign n14471 = n12142 ^ n4851 ;
  assign n14472 = n14471 ^ n12142 ;
  assign n14473 = n12143 & n14472 ;
  assign n14474 = n14473 ^ n12142 ;
  assign n14475 = ~n35 & ~n14474 ;
  assign n14483 = n14482 ^ n14475 ;
  assign n14467 = n14361 ^ n14357 ;
  assign n14468 = n14467 ^ n14297 ;
  assign n14484 = n14483 ^ n14468 ;
  assign n14609 = n14355 ^ n13932 ;
  assign n14610 = n14609 ^ n14313 ;
  assign n14505 = n14352 ^ n14316 ;
  assign n14503 = ~n35 & n12149 ;
  assign n14497 = n12237 ^ n12198 ;
  assign n14498 = n14497 ^ n12143 ;
  assign n14499 = n14498 ^ n12149 ;
  assign n14500 = ~n14499 & n23912 ;
  assign n14494 = n12149 ^ n3726 ;
  assign n14485 = ~n35 & ~n12151 ;
  assign n14495 = n14494 ^ n14485 ;
  assign n14501 = n14500 ^ n14495 ;
  assign n14486 = n14485 ^ n12149 ;
  assign n14487 = n14486 ^ n3726 ;
  assign n14488 = n14487 ^ n14486 ;
  assign n14489 = n14486 ^ n12143 ;
  assign n14490 = n14489 ^ n14486 ;
  assign n14491 = n14488 & ~n14490 ;
  assign n14492 = n14491 ^ n14486 ;
  assign n14493 = ~x31 & n14492 ;
  assign n14502 = n14501 ^ n14493 ;
  assign n14504 = n14503 ^ n14502 ;
  assign n14506 = n14505 ^ n14504 ;
  assign n14515 = n12417 ^ n819 ;
  assign n14514 = n456 ^ n396 ;
  assign n14516 = n14515 ^ n14514 ;
  assign n14511 = n1205 ^ n291 ;
  assign n14512 = n14511 ^ n403 ;
  assign n14510 = n13770 ^ n2771 ;
  assign n14513 = n14512 ^ n14510 ;
  assign n14517 = n14516 ^ n14513 ;
  assign n14507 = n4304 ^ n507 ;
  assign n14508 = n14507 ^ n3323 ;
  assign n14509 = n14508 ^ n3288 ;
  assign n14518 = n14517 ^ n14509 ;
  assign n14519 = n14518 ^ n5372 ;
  assign n14520 = n14519 ^ n595 ;
  assign n14521 = ~n3897 & ~n14520 ;
  assign n14522 = n14521 ^ n14315 ;
  assign n14535 = n4132 ^ n2912 ;
  assign n14534 = n3433 ^ n1004 ;
  assign n14536 = n14535 ^ n14534 ;
  assign n14531 = n378 ^ n104 ;
  assign n14532 = n14531 ^ n1184 ;
  assign n14530 = n4356 ^ n682 ;
  assign n14533 = n14532 ^ n14530 ;
  assign n14537 = n14536 ^ n14533 ;
  assign n14538 = n14537 ^ n12482 ;
  assign n14526 = n12797 ^ n961 ;
  assign n14527 = n14526 ^ n11919 ;
  assign n14528 = n14527 ^ n1507 ;
  assign n14523 = n1783 ^ n379 ;
  assign n14524 = n14523 ^ n6215 ;
  assign n14525 = n14524 ^ n1275 ;
  assign n14529 = n14528 ^ n14525 ;
  assign n14539 = n14538 ^ n14529 ;
  assign n14540 = ~n14339 & ~n14539 ;
  assign n14552 = n2481 ^ n1435 ;
  assign n14551 = n3212 ^ n1564 ;
  assign n14553 = n14552 ^ n14551 ;
  assign n14549 = n945 ^ n153 ;
  assign n14550 = n14549 ^ n2098 ;
  assign n14554 = n14553 ^ n14550 ;
  assign n14547 = n6491 ^ n2167 ;
  assign n14545 = n14544 ^ n3444 ;
  assign n14546 = n14545 ^ n6333 ;
  assign n14548 = n14547 ^ n14546 ;
  assign n14555 = n14554 ^ n14548 ;
  assign n14542 = n13843 ^ n1906 ;
  assign n14541 = n2292 ^ n1088 ;
  assign n14543 = n14542 ^ n14541 ;
  assign n14556 = n14555 ^ n14543 ;
  assign n14557 = n14556 ^ n13026 ;
  assign n14576 = n4089 ^ n625 ;
  assign n14575 = n2067 ^ n122 ;
  assign n14577 = n14576 ^ n14575 ;
  assign n14570 = n641 ^ n417 ;
  assign n14571 = n14570 ^ n668 ;
  assign n14572 = n14571 ^ n2082 ;
  assign n14567 = n2764 ^ n550 ;
  assign n14568 = n14567 ^ n5226 ;
  assign n14565 = n2171 ^ n1148 ;
  assign n14563 = n4336 ^ n505 ;
  assign n14564 = n14563 ^ n3442 ;
  assign n14566 = n14565 ^ n14564 ;
  assign n14569 = n14568 ^ n14566 ;
  assign n14573 = n14572 ^ n14569 ;
  assign n14559 = n4121 ^ n137 ;
  assign n14560 = n14559 ^ n2724 ;
  assign n14558 = n2177 ^ n600 ;
  assign n14561 = n14560 ^ n14558 ;
  assign n14562 = n14561 ^ n2275 ;
  assign n14574 = n14573 ^ n14562 ;
  assign n14578 = n14577 ^ n14574 ;
  assign n14579 = ~n14557 & ~n14578 ;
  assign n14591 = n3726 & n12152 ;
  assign n14590 = ~n3733 & n12160 ;
  assign n14592 = n14591 ^ n14590 ;
  assign n14582 = ~n35 & n12163 ;
  assign n14580 = n12234 ^ n12195 ;
  assign n14581 = n14580 ^ n12152 ;
  assign n14583 = n14582 ^ n14581 ;
  assign n14584 = n14583 ^ n14582 ;
  assign n14585 = n14582 ^ n3520 ;
  assign n14586 = n14585 ^ n14582 ;
  assign n14587 = ~n14584 & n14586 ;
  assign n14588 = n14587 ^ n14582 ;
  assign n14589 = x31 & n14588 ;
  assign n14593 = n14592 ^ n14589 ;
  assign n14594 = ~n14579 & n14593 ;
  assign n14595 = ~n14315 & ~n14594 ;
  assign n14596 = ~n14540 & ~n14595 ;
  assign n14597 = n14593 ^ n14579 ;
  assign n14598 = n14597 ^ n14594 ;
  assign n14599 = n14315 & ~n14598 ;
  assign n14600 = n14596 & ~n14599 ;
  assign n14601 = n14600 ^ n14599 ;
  assign n14602 = n14601 ^ n14521 ;
  assign n14603 = ~n14522 & n14602 ;
  assign n14604 = n14603 ^ n14315 ;
  assign n14605 = n14604 ^ n14504 ;
  assign n14606 = n14506 & n14605 ;
  assign n14607 = n14606 ^ n14504 ;
  assign n14611 = n14610 ^ n14607 ;
  assign n14621 = n3484 & ~n12138 ;
  assign n14614 = n12137 ^ x29 ;
  assign n14615 = n14614 ^ x28 ;
  assign n14616 = n14615 ^ n12137 ;
  assign n14617 = ~n13936 & n14616 ;
  assign n14618 = n14617 ^ n12137 ;
  assign n14619 = n650 & n14618 ;
  assign n14620 = n14619 ^ x29 ;
  assign n14622 = n14621 ^ n14620 ;
  assign n14612 = n831 & n12207 ;
  assign n14623 = n14622 ^ n14612 ;
  assign n14624 = n14623 ^ n14607 ;
  assign n14625 = ~n14611 & n14624 ;
  assign n14608 = n14607 ^ n14483 ;
  assign n14626 = n14625 ^ n14608 ;
  assign n14627 = n14484 & n14626 ;
  assign n14628 = n14627 ^ n14483 ;
  assign n14464 = n14393 ^ n14281 ;
  assign n14465 = n14464 ^ n14461 ;
  assign n14466 = n14465 ^ n14464 ;
  assign n14629 = n14628 ^ n14466 ;
  assign n14630 = ~n14463 & n14629 ;
  assign n14631 = n14630 ^ n14465 ;
  assign n14632 = n14396 ^ n14265 ;
  assign n14642 = n14632 ^ n14464 ;
  assign n14636 = n12121 & n12861 ;
  assign n14635 = n446 & n12117 ;
  assign n14637 = n14636 ^ n14635 ;
  assign n14638 = n14637 ^ x26 ;
  assign n14634 = ~n487 & ~n12110 ;
  assign n14639 = n14638 ^ n14634 ;
  assign n14633 = ~n3501 & n13196 ;
  assign n14640 = n14639 ^ n14633 ;
  assign n14641 = n14640 ^ n14632 ;
  assign n14643 = n14642 ^ n14641 ;
  assign n14644 = ~n14631 & ~n14643 ;
  assign n14645 = n14644 ^ n14642 ;
  assign n14651 = n4491 & n11972 ;
  assign n14648 = n4492 & ~n14078 ;
  assign n14647 = ~n4496 & n12260 ;
  assign n14649 = n14648 ^ n14647 ;
  assign n14650 = n14649 ^ x23 ;
  assign n14652 = n14651 ^ n14650 ;
  assign n14646 = n4504 & ~n12256 ;
  assign n14653 = n14652 ^ n14646 ;
  assign n14663 = n14653 ^ n14632 ;
  assign n14660 = ~n4496 & ~n12256 ;
  assign n14658 = n4492 & n13054 ;
  assign n14655 = n4504 & ~n12262 ;
  assign n14654 = n4491 & n12260 ;
  assign n14656 = n14655 ^ n14654 ;
  assign n14657 = n14656 ^ x23 ;
  assign n14659 = n14658 ^ n14657 ;
  assign n14661 = n14660 ^ n14659 ;
  assign n14662 = n14661 ^ n14653 ;
  assign n14664 = n14663 ^ n14662 ;
  assign n14665 = n14645 & ~n14664 ;
  assign n14666 = n14665 ^ n14663 ;
  assign n14669 = n14653 ^ n14436 ;
  assign n14667 = n14398 ^ n14257 ;
  assign n14668 = n14667 ^ n14436 ;
  assign n14670 = n14669 ^ n14668 ;
  assign n14671 = ~n14666 & n14670 ;
  assign n14672 = n14671 ^ n14669 ;
  assign n14673 = n14449 & n14672 ;
  assign n14437 = n14436 ^ n14434 ;
  assign n14674 = n14673 ^ n14437 ;
  assign n14675 = n14435 & n14674 ;
  assign n14676 = n14675 ^ n14434 ;
  assign n20735 = n14683 ^ n14676 ;
  assign n20736 = n14685 & n20735 ;
  assign n20737 = n20736 ^ n14683 ;
  assign n20752 = n20740 ^ n20737 ;
  assign n20734 = n14193 ^ n14182 ;
  assign n20738 = n20737 ^ n20734 ;
  assign n20732 = ~n12855 & n20731 ;
  assign n20733 = n20732 ^ n20727 ;
  assign n20750 = n20734 ^ n20733 ;
  assign n20751 = ~n20738 & n20750 ;
  assign n20753 = n20752 ^ n20751 ;
  assign n20754 = n20751 ^ n20737 ;
  assign n14421 = n14420 ^ n14229 ;
  assign n14422 = ~n14237 & n14421 ;
  assign n14423 = n14422 ^ n14420 ;
  assign n20755 = n20754 ^ n14423 ;
  assign n20756 = n20755 ^ n20754 ;
  assign n14687 = n14674 ^ n14433 ;
  assign n14723 = n14661 ^ n14645 ;
  assign n14720 = n4916 & ~n12108 ;
  assign n14713 = n12367 ^ x20 ;
  assign n14714 = n14713 ^ x19 ;
  assign n14715 = n14714 ^ n12367 ;
  assign n14716 = ~n12369 & n14715 ;
  assign n14717 = n14716 ^ n12367 ;
  assign n14718 = n4678 & ~n14717 ;
  assign n14719 = n14718 ^ x20 ;
  assign n14721 = n14720 ^ n14719 ;
  assign n14712 = n11972 & n14027 ;
  assign n14722 = n14721 ^ n14712 ;
  assign n14724 = n14723 ^ n14722 ;
  assign n14734 = n14628 ^ n14463 ;
  assign n14729 = ~n12129 & n12861 ;
  assign n14728 = n446 & n12121 ;
  assign n14730 = n14729 ^ n14728 ;
  assign n14731 = n14730 ^ x26 ;
  assign n14727 = ~n487 & n12117 ;
  assign n14732 = n14731 ^ n14727 ;
  assign n14726 = ~n3501 & ~n13596 ;
  assign n14733 = n14732 ^ n14726 ;
  assign n14735 = n14734 ^ n14733 ;
  assign n14749 = n14626 ^ n14468 ;
  assign n14737 = n12130 & n12861 ;
  assign n14736 = n446 & ~n12129 ;
  assign n14738 = n14737 ^ n14736 ;
  assign n14739 = n14738 ^ n65 ;
  assign n14741 = n14738 ^ x26 ;
  assign n14744 = n14741 ^ n67 ;
  assign n14745 = ~x25 & ~n13605 ;
  assign n14746 = n14744 & n14745 ;
  assign n14742 = ~n12121 & n14741 ;
  assign n14740 = n67 & ~n13606 ;
  assign n14743 = n14742 ^ n14740 ;
  assign n14747 = n14746 ^ n14743 ;
  assign n14748 = ~n14739 & ~n14747 ;
  assign n14750 = n14749 ^ n14748 ;
  assign n14761 = n14749 ^ x29 ;
  assign n14753 = n14129 ^ n12136 ;
  assign n14756 = n12136 ^ n4536 ;
  assign n14757 = n14756 ^ n12136 ;
  assign n14758 = ~n14753 & n14757 ;
  assign n14759 = n14758 ^ n12136 ;
  assign n14760 = n650 & ~n14759 ;
  assign n14762 = n14761 ^ n14760 ;
  assign n14752 = n3484 & n12137 ;
  assign n14763 = n14762 ^ n14752 ;
  assign n14751 = n831 & ~n12138 ;
  assign n14764 = n14763 ^ n14751 ;
  assign n14765 = ~n14750 & n14764 ;
  assign n14766 = n14765 ^ n14749 ;
  assign n14767 = n14766 ^ n14733 ;
  assign n14768 = ~n14735 & n14767 ;
  assign n14769 = n14768 ^ n14733 ;
  assign n14725 = n14640 ^ n14631 ;
  assign n14770 = n14769 ^ n14725 ;
  assign n14775 = n4504 & ~n12220 ;
  assign n14774 = n4491 & ~n12256 ;
  assign n14776 = n14775 ^ n14774 ;
  assign n14777 = n14776 ^ x23 ;
  assign n14773 = n4492 & ~n13283 ;
  assign n14778 = n14777 ^ n14773 ;
  assign n14772 = ~n4496 & ~n12262 ;
  assign n14779 = n14778 ^ n14772 ;
  assign n14771 = n14769 ^ n14723 ;
  assign n14780 = n14779 ^ n14771 ;
  assign n14781 = n14780 ^ n14723 ;
  assign n14782 = ~n14770 & n14781 ;
  assign n14783 = n14782 ^ n14771 ;
  assign n14784 = n14724 & n14783 ;
  assign n14785 = n14784 ^ n14723 ;
  assign n14710 = n14667 ^ n14666 ;
  assign n14707 = n4916 & ~n12367 ;
  assign n14700 = n12613 ^ x20 ;
  assign n14701 = n14700 ^ x19 ;
  assign n14702 = n14701 ^ n12613 ;
  assign n14703 = ~n13111 & n14702 ;
  assign n14704 = n14703 ^ n12613 ;
  assign n14705 = n4678 & ~n14704 ;
  assign n14706 = n14705 ^ x20 ;
  assign n14708 = n14707 ^ n14706 ;
  assign n14699 = ~n12108 & n14027 ;
  assign n14709 = n14708 ^ n14699 ;
  assign n14711 = n14710 ^ n14709 ;
  assign n15363 = n14785 ^ n14711 ;
  assign n14800 = n14783 ^ n14722 ;
  assign n14795 = n5700 & n12656 ;
  assign n14794 = n5702 & ~n12705 ;
  assign n14796 = n14795 ^ n14794 ;
  assign n14797 = n14796 ^ x17 ;
  assign n14793 = n5703 & n12706 ;
  assign n14798 = n14797 ^ n14793 ;
  assign n14792 = ~n12613 & n20731 ;
  assign n14799 = n14798 ^ n14792 ;
  assign n14801 = n14800 ^ n14799 ;
  assign n15356 = n14779 ^ n14770 ;
  assign n14819 = n14766 ^ n14735 ;
  assign n14817 = ~n4496 & ~n12220 ;
  assign n14815 = n4492 & n13712 ;
  assign n14812 = n4504 & ~n12110 ;
  assign n14811 = n4491 & ~n12262 ;
  assign n14813 = n14812 ^ n14811 ;
  assign n14814 = n14813 ^ x23 ;
  assign n14816 = n14815 ^ n14814 ;
  assign n14818 = n14817 ^ n14816 ;
  assign n14820 = n14819 ^ n14818 ;
  assign n14829 = n14764 ^ n14748 ;
  assign n14824 = n4504 & n12117 ;
  assign n14823 = n4491 & ~n12220 ;
  assign n14825 = n14824 ^ n14823 ;
  assign n14826 = n14825 ^ x23 ;
  assign n14822 = n4492 & n14047 ;
  assign n14827 = n14826 ^ n14822 ;
  assign n14821 = ~n4496 & ~n12110 ;
  assign n14828 = n14827 ^ n14821 ;
  assign n14830 = n14829 ^ n14828 ;
  assign n15338 = n14623 ^ n14611 ;
  assign n14844 = n14604 ^ n14506 ;
  assign n14841 = n3484 & n12207 ;
  assign n14837 = n4536 & ~n14370 ;
  assign n14838 = n14837 ^ n12138 ;
  assign n14839 = n650 & ~n14838 ;
  assign n14840 = n14839 ^ x29 ;
  assign n14842 = n14841 ^ n14840 ;
  assign n14831 = n831 & ~n12142 ;
  assign n14843 = n14842 ^ n14831 ;
  assign n14845 = n14844 ^ n14843 ;
  assign n15309 = n14601 ^ n14522 ;
  assign n15294 = n14599 ^ n14595 ;
  assign n15295 = n15294 ^ n14540 ;
  assign n15276 = n14579 ^ n14315 ;
  assign n15277 = n15276 ^ n14593 ;
  assign n14864 = ~n35 & n12167 ;
  assign n14876 = n14864 ^ n14585 ;
  assign n14863 = n3726 & ~n12160 ;
  assign n14865 = n14864 ^ n14863 ;
  assign n14877 = n14876 ^ n14865 ;
  assign n14869 = n14865 ^ n12163 ;
  assign n14866 = n12233 ^ n12194 ;
  assign n14867 = n14866 ^ n12160 ;
  assign n14868 = n14867 ^ n14865 ;
  assign n14870 = n14869 ^ n14868 ;
  assign n14871 = n14869 ^ n3520 ;
  assign n14872 = n14871 ^ n14869 ;
  assign n14873 = n14870 & n14872 ;
  assign n14874 = n14873 ^ n14869 ;
  assign n14875 = x31 & n14874 ;
  assign n14878 = n14877 ^ n14875 ;
  assign n14856 = n11911 ^ n1247 ;
  assign n14855 = n13902 ^ n2133 ;
  assign n14857 = n14856 ^ n14855 ;
  assign n14858 = n14857 ^ n13796 ;
  assign n14859 = n14858 ^ n2700 ;
  assign n14851 = n2814 ^ n565 ;
  assign n14852 = n14851 ^ n3303 ;
  assign n14853 = n14852 ^ n11816 ;
  assign n14848 = n1492 ^ n407 ;
  assign n14849 = n14848 ^ n888 ;
  assign n14846 = n3675 ^ n304 ;
  assign n14847 = n14846 ^ n857 ;
  assign n14850 = n14849 ^ n14847 ;
  assign n14854 = n14853 ^ n14850 ;
  assign n14860 = n14859 ^ n14854 ;
  assign n14861 = n14860 ^ n1431 ;
  assign n14862 = ~n4812 & ~n14861 ;
  assign n14879 = n14878 ^ n14862 ;
  assign n14906 = n3973 ^ n3002 ;
  assign n14907 = n14906 ^ n3323 ;
  assign n14908 = n14907 ^ n2871 ;
  assign n14904 = n12443 ^ n2345 ;
  assign n14902 = n940 ^ n577 ;
  assign n14900 = n2432 ^ n161 ;
  assign n14901 = n14900 ^ n1050 ;
  assign n14903 = n14902 ^ n14901 ;
  assign n14905 = n14904 ^ n14903 ;
  assign n14909 = n14908 ^ n14905 ;
  assign n14899 = n12312 ^ n5636 ;
  assign n14910 = n14909 ^ n14899 ;
  assign n14911 = ~n1538 & ~n1596 ;
  assign n14912 = ~n14910 & n14911 ;
  assign n14893 = n12163 ^ n3726 ;
  assign n14894 = n14893 ^ n14864 ;
  assign n14880 = n12232 ^ n12193 ;
  assign n14895 = n14894 ^ n14880 ;
  assign n14881 = ~n35 & n12168 ;
  assign n14896 = n14895 ^ n14881 ;
  assign n14890 = n14880 ^ n12163 ;
  assign n14891 = n14890 ^ n12167 ;
  assign n14892 = n12015 & ~n14891 ;
  assign n14897 = n14896 ^ n14892 ;
  assign n14882 = n14881 ^ n14880 ;
  assign n14883 = n14882 ^ n3726 ;
  assign n14884 = n14883 ^ n14882 ;
  assign n14885 = n14882 ^ n12163 ;
  assign n14886 = n14885 ^ n14882 ;
  assign n14887 = ~n14884 & ~n14886 ;
  assign n14888 = n14887 ^ n14882 ;
  assign n14889 = ~x31 & n14888 ;
  assign n14898 = n14897 ^ n14889 ;
  assign n14913 = n14912 ^ n14898 ;
  assign n14941 = n4352 ^ n2180 ;
  assign n14942 = n14941 ^ n2533 ;
  assign n14938 = n13034 ^ n1608 ;
  assign n14937 = n2720 ^ n2243 ;
  assign n14939 = n14938 ^ n14937 ;
  assign n14935 = n11830 ^ n797 ;
  assign n14934 = n4318 ^ n297 ;
  assign n14936 = n14935 ^ n14934 ;
  assign n14940 = n14939 ^ n14936 ;
  assign n14943 = n14942 ^ n14940 ;
  assign n14944 = n14943 ^ n2934 ;
  assign n14945 = n14944 ^ n2318 ;
  assign n14946 = ~n14578 & ~n14945 ;
  assign n14914 = n12231 ^ n12192 ;
  assign n14915 = n14914 ^ n12167 ;
  assign n14917 = n14915 ^ n12168 ;
  assign n14916 = n14915 ^ n12169 ;
  assign n14918 = n14917 ^ n14916 ;
  assign n14921 = x30 & ~n14918 ;
  assign n14922 = n14921 ^ n14917 ;
  assign n14923 = ~n3520 & ~n14922 ;
  assign n14924 = n14923 ^ n14915 ;
  assign n14925 = n14924 ^ n14881 ;
  assign n14928 = n14925 ^ n12167 ;
  assign n14929 = n14928 ^ n14925 ;
  assign n14930 = n3520 & n14929 ;
  assign n14931 = n14930 ^ n14925 ;
  assign n14932 = ~x31 & ~n14931 ;
  assign n14933 = n14932 ^ n14924 ;
  assign n14947 = n14946 ^ n14933 ;
  assign n14972 = n2180 ^ n1425 ;
  assign n14970 = n769 ^ n192 ;
  assign n14971 = n14970 ^ n1050 ;
  assign n14973 = n14972 ^ n14971 ;
  assign n14968 = n1004 ^ n953 ;
  assign n14967 = n12320 ^ n1023 ;
  assign n14969 = n14968 ^ n14967 ;
  assign n14974 = n14973 ^ n14969 ;
  assign n14963 = n5069 ^ n772 ;
  assign n14964 = n14963 ^ n1122 ;
  assign n14965 = n14964 ^ n2507 ;
  assign n14966 = n14965 ^ n3695 ;
  assign n14975 = n14974 ^ n14966 ;
  assign n14976 = n14975 ^ n3454 ;
  assign n14977 = ~n4037 & ~n14976 ;
  assign n14960 = ~n3733 & ~n12169 ;
  assign n14958 = ~n35 & n12175 ;
  assign n14959 = x31 & n14958 ;
  assign n14961 = n14960 ^ n14959 ;
  assign n14948 = n12230 ^ n12191 ;
  assign n14953 = n12168 ^ x31 ;
  assign n14954 = n14953 ^ n12168 ;
  assign n14955 = ~n14948 & n14954 ;
  assign n14956 = n14955 ^ n12168 ;
  assign n14957 = n3520 & n14956 ;
  assign n14962 = n14961 ^ n14957 ;
  assign n14978 = n14977 ^ n14962 ;
  assign n15032 = n12229 ^ n12190 ;
  assign n15035 = n15032 ^ n12169 ;
  assign n15043 = n15035 ^ n12175 ;
  assign n15044 = ~n12015 & n15043 ;
  assign n15040 = n12175 ^ n3726 ;
  assign n15041 = n15040 ^ n14958 ;
  assign n15033 = n15032 ^ n3726 ;
  assign n15034 = n15033 ^ n15032 ;
  assign n15036 = n15035 ^ n15032 ;
  assign n15037 = ~n15034 & n15036 ;
  assign n15038 = n15037 ^ n15032 ;
  assign n15039 = ~x31 & n15038 ;
  assign n15042 = n15041 ^ n15039 ;
  assign n15045 = n15044 ^ n15042 ;
  assign n15031 = n12179 & n24214 ;
  assign n15046 = n15045 ^ n15031 ;
  assign n15011 = n2912 ^ n285 ;
  assign n15012 = n15011 ^ n425 ;
  assign n15008 = n2269 ^ n704 ;
  assign n15006 = n12690 ^ n124 ;
  assign n15007 = n15006 ^ n403 ;
  assign n15009 = n15008 ^ n15007 ;
  assign n15010 = n15009 ^ n6213 ;
  assign n15013 = n15012 ^ n15010 ;
  assign n15000 = n11823 ^ n212 ;
  assign n15001 = n15000 ^ n627 ;
  assign n15002 = n15001 ^ n1969 ;
  assign n15003 = n15002 ^ n3534 ;
  assign n15004 = n15003 ^ n3009 ;
  assign n15005 = n15004 ^ n13661 ;
  assign n15014 = n15013 ^ n15005 ;
  assign n14994 = n1822 ^ n507 ;
  assign n14993 = n698 ^ n371 ;
  assign n14995 = n14994 ^ n14993 ;
  assign n14991 = n4973 ^ n2744 ;
  assign n14992 = n14991 ^ n5605 ;
  assign n14996 = n14995 ^ n14992 ;
  assign n14988 = n11921 ^ n683 ;
  assign n14989 = n14988 ^ n3086 ;
  assign n14986 = n6419 ^ n632 ;
  assign n14987 = n14986 ^ n940 ;
  assign n14990 = n14989 ^ n14987 ;
  assign n14997 = n14996 ^ n14990 ;
  assign n14982 = n73 ^ n70 ;
  assign n14983 = ~n338 & ~n14982 ;
  assign n14998 = n14997 ^ n14983 ;
  assign n14980 = n138 & n358 ;
  assign n14979 = n72 & ~n338 ;
  assign n14981 = n14980 ^ n14979 ;
  assign n14984 = x26 & ~n14983 ;
  assign n14985 = n14981 & n14984 ;
  assign n14999 = n14998 ^ n14985 ;
  assign n15015 = n15014 ^ n14999 ;
  assign n15025 = n13649 ^ n2090 ;
  assign n15022 = n14570 ^ n541 ;
  assign n15023 = n15022 ^ n893 ;
  assign n15020 = n3689 ^ n1129 ;
  assign n15021 = n15020 ^ n151 ;
  assign n15024 = n15023 ^ n15021 ;
  assign n15026 = n15025 ^ n15024 ;
  assign n15017 = n3602 ^ n2888 ;
  assign n15016 = n3671 ^ n1476 ;
  assign n15018 = n15017 ^ n15016 ;
  assign n15019 = n15018 ^ n6323 ;
  assign n15027 = n15026 ^ n15019 ;
  assign n15028 = n15027 ^ n1732 ;
  assign n15029 = ~n15015 & ~n15028 ;
  assign n15047 = n15046 ^ n15029 ;
  assign n15074 = n2423 ^ n805 ;
  assign n15073 = n1933 ^ n1188 ;
  assign n15075 = n15074 ^ n15073 ;
  assign n15070 = n512 ^ n190 ;
  assign n15068 = n1392 ^ n774 ;
  assign n15069 = n15068 ^ n760 ;
  assign n15071 = n15070 ^ n15069 ;
  assign n15066 = n11890 ^ n2849 ;
  assign n15065 = n1847 ^ n1783 ;
  assign n15067 = n15066 ^ n15065 ;
  assign n15072 = n15071 ^ n15067 ;
  assign n15076 = n15075 ^ n15072 ;
  assign n15064 = n13896 ^ n1992 ;
  assign n15077 = n15076 ^ n15064 ;
  assign n15090 = n697 ^ n542 ;
  assign n15091 = n15090 ^ n12055 ;
  assign n15092 = n15091 ^ n13637 ;
  assign n15093 = n15092 ^ n2431 ;
  assign n15086 = n3973 ^ n3601 ;
  assign n15087 = n15086 ^ n3995 ;
  assign n15084 = n1305 ^ n1021 ;
  assign n15083 = n1254 ^ n118 ;
  assign n15085 = n15084 ^ n15083 ;
  assign n15088 = n15087 ^ n15085 ;
  assign n15080 = n835 ^ n376 ;
  assign n15081 = n15080 ^ n229 ;
  assign n15078 = n4118 ^ n496 ;
  assign n15079 = n15078 ^ n798 ;
  assign n15082 = n15081 ^ n15079 ;
  assign n15089 = n15088 ^ n15082 ;
  assign n15094 = n15093 ^ n15089 ;
  assign n15095 = n15094 ^ n11908 ;
  assign n15096 = ~n15077 & ~n15095 ;
  assign n15057 = ~x31 & ~n12180 ;
  assign n15056 = n12180 ^ x31 ;
  assign n15058 = n15057 ^ n15056 ;
  assign n15059 = n15058 ^ n12179 ;
  assign n15060 = ~n35 & ~n15059 ;
  assign n15053 = x31 & n12179 ;
  assign n15061 = n15060 ^ n15053 ;
  assign n15062 = n15061 ^ n3726 ;
  assign n15051 = n12175 & ~n23912 ;
  assign n15048 = n12228 ^ n12189 ;
  assign n15049 = n15048 ^ n12175 ;
  assign n15050 = x31 & n15049 ;
  assign n15052 = n15051 ^ n15050 ;
  assign n15054 = n15053 ^ n15052 ;
  assign n15055 = n3520 & ~n15054 ;
  assign n15063 = n15062 ^ n15055 ;
  assign n15097 = n15096 ^ n15063 ;
  assign n15144 = x30 & n12180 ;
  assign n15127 = n12227 ^ n12188 ;
  assign n15128 = n15127 ^ n12179 ;
  assign n15130 = n15128 ^ n12180 ;
  assign n15129 = n15128 ^ n12181 ;
  assign n15131 = n15130 ^ n15129 ;
  assign n15134 = x30 & n15131 ;
  assign n15135 = n15134 ^ n15130 ;
  assign n15136 = ~n3520 & ~n15135 ;
  assign n15137 = n15136 ^ n15128 ;
  assign n15138 = n15137 ^ n12179 ;
  assign n15139 = n15138 ^ n15137 ;
  assign n15145 = n15144 ^ n15139 ;
  assign n15146 = ~n3520 & n15145 ;
  assign n15147 = n15146 ^ n15138 ;
  assign n15148 = ~x31 & ~n15147 ;
  assign n15149 = n15148 ^ n15137 ;
  assign n15103 = n1986 ^ n725 ;
  assign n15104 = n15103 ^ n1746 ;
  assign n15105 = n15104 ^ n13892 ;
  assign n15101 = n4754 ^ n4140 ;
  assign n15098 = n5605 ^ n602 ;
  assign n15099 = n15098 ^ n410 ;
  assign n15100 = n15099 ^ n1448 ;
  assign n15102 = n15101 ^ n15100 ;
  assign n15106 = n15105 ^ n15102 ;
  assign n15107 = n15106 ^ n2778 ;
  assign n15120 = n308 ^ n210 ;
  assign n15121 = n15120 ^ n952 ;
  assign n15122 = n15121 ^ n1278 ;
  assign n15117 = n13231 ^ n1379 ;
  assign n15118 = n15117 ^ n878 ;
  assign n15115 = n13658 ^ n2336 ;
  assign n15114 = n3664 ^ n3432 ;
  assign n15116 = n15115 ^ n15114 ;
  assign n15119 = n15118 ^ n15116 ;
  assign n15123 = n15122 ^ n15119 ;
  assign n15110 = n453 ^ n226 ;
  assign n15111 = n15110 ^ n455 ;
  assign n15108 = n3128 ^ n355 ;
  assign n15109 = n15108 ^ n1148 ;
  assign n15112 = n15111 ^ n15109 ;
  assign n15113 = n15112 ^ n13856 ;
  assign n15124 = n15123 ^ n15113 ;
  assign n15125 = ~n2122 & ~n15124 ;
  assign n15126 = ~n15107 & n15125 ;
  assign n15150 = n15149 ^ n15126 ;
  assign n15175 = n3985 ^ n2618 ;
  assign n15172 = n835 ^ n405 ;
  assign n15173 = n15172 ^ n1236 ;
  assign n15171 = n2937 ^ n589 ;
  assign n15174 = n15173 ^ n15171 ;
  assign n15176 = n15175 ^ n15174 ;
  assign n15177 = n15176 ^ n5044 ;
  assign n15169 = n6272 ^ n168 ;
  assign n15170 = n15169 ^ n3073 ;
  assign n15178 = n15177 ^ n15170 ;
  assign n15179 = n12546 ^ n12339 ;
  assign n15180 = ~n15178 & ~n15179 ;
  assign n15181 = ~n3659 & n15180 ;
  assign n15160 = n12222 ^ n12182 ;
  assign n15163 = ~n35 & n15160 ;
  assign n15164 = n15163 ^ n12182 ;
  assign n15165 = n15164 & ~n24214 ;
  assign n15166 = n15165 ^ n12182 ;
  assign n15159 = n12533 & ~n15057 ;
  assign n15167 = n15166 ^ n15159 ;
  assign n15151 = n12225 ^ n12180 ;
  assign n15152 = n15151 ^ n3520 ;
  assign n15153 = n15152 ^ n15151 ;
  assign n15154 = ~x30 & ~n12181 ;
  assign n15155 = n15154 ^ n15151 ;
  assign n15156 = ~n15153 & n15155 ;
  assign n15157 = n15156 ^ n15151 ;
  assign n15158 = x31 & n15157 ;
  assign n15168 = n15167 ^ n15158 ;
  assign n15182 = n15181 ^ n15168 ;
  assign n15226 = n11900 ^ n2506 ;
  assign n15225 = n2051 ^ n964 ;
  assign n15227 = n15226 ^ n15225 ;
  assign n15221 = n5226 ^ n871 ;
  assign n15222 = n15221 ^ n613 ;
  assign n15220 = n773 ^ n273 ;
  assign n15223 = n15222 ^ n15220 ;
  assign n15184 = n597 ^ n203 ;
  assign n15218 = n15184 ^ n883 ;
  assign n15217 = n4356 ^ n2135 ;
  assign n15219 = n15218 ^ n15217 ;
  assign n15224 = n15223 ^ n15219 ;
  assign n15228 = n15227 ^ n15224 ;
  assign n15229 = n15228 ^ n14548 ;
  assign n15230 = n15229 ^ n12824 ;
  assign n15231 = ~n13851 & ~n15230 ;
  assign n15185 = n15184 ^ n2190 ;
  assign n15183 = n4980 ^ n610 ;
  assign n15186 = n15185 ^ n15183 ;
  assign n15199 = n3606 ^ n158 ;
  assign n15198 = n13844 ^ n12041 ;
  assign n15200 = n15199 ^ n15198 ;
  assign n15195 = n4342 ^ n2510 ;
  assign n15192 = n678 ^ n144 ;
  assign n15193 = n15192 ^ n364 ;
  assign n15194 = n15193 ^ n1169 ;
  assign n15196 = n15195 ^ n15194 ;
  assign n15189 = n2059 ^ n627 ;
  assign n15190 = n15189 ^ n797 ;
  assign n15187 = n14965 ^ n592 ;
  assign n15188 = n15187 ^ n775 ;
  assign n15191 = n15190 ^ n15188 ;
  assign n15197 = n15196 ^ n15191 ;
  assign n15201 = n15200 ^ n15197 ;
  assign n15207 = n3209 ^ n3184 ;
  assign n15205 = n12336 ^ n5245 ;
  assign n15203 = n2627 ^ n226 ;
  assign n15202 = n14567 ^ n577 ;
  assign n15204 = n15203 ^ n15202 ;
  assign n15206 = n15205 ^ n15204 ;
  assign n15208 = n15207 ^ n15206 ;
  assign n15209 = n15208 ^ n6394 ;
  assign n15210 = n15209 ^ n2881 ;
  assign n15211 = ~n15201 & ~n15210 ;
  assign n15212 = ~n15186 & n15211 ;
  assign n15214 = ~n3720 & ~n12183 ;
  assign n15213 = n3520 & ~n12182 ;
  assign n15215 = n15214 ^ n15213 ;
  assign n15216 = ~n15212 & n15215 ;
  assign n15232 = n15231 ^ n15216 ;
  assign n15244 = n12182 & n23912 ;
  assign n15245 = n15244 ^ n4851 ;
  assign n15246 = n12183 & n15245 ;
  assign n15239 = n24214 ^ n12181 ;
  assign n15247 = n15246 ^ n15239 ;
  assign n15234 = n12181 ^ n3720 ;
  assign n15235 = n15234 ^ n12181 ;
  assign n15236 = ~n12182 & ~n15235 ;
  assign n15237 = n15236 ^ n12181 ;
  assign n15238 = ~n3520 & n15237 ;
  assign n15248 = n15247 ^ n15238 ;
  assign n15249 = n15248 ^ n15216 ;
  assign n15250 = ~n15232 & n15249 ;
  assign n15251 = n15250 ^ n15216 ;
  assign n15252 = n15251 ^ n15168 ;
  assign n15253 = ~n15182 & ~n15252 ;
  assign n15254 = n15253 ^ n15181 ;
  assign n15255 = n15254 ^ n15149 ;
  assign n15256 = n15150 & n15255 ;
  assign n15257 = n15256 ^ n15149 ;
  assign n15258 = n15257 ^ n15063 ;
  assign n15259 = ~n15097 & ~n15258 ;
  assign n15260 = n15259 ^ n15063 ;
  assign n15261 = n15260 ^ n15046 ;
  assign n15262 = ~n15047 & n15261 ;
  assign n15263 = n15262 ^ n15046 ;
  assign n15264 = n15263 ^ n14962 ;
  assign n15265 = ~n14978 & n15264 ;
  assign n15266 = n15265 ^ n14962 ;
  assign n15267 = n15266 ^ n14933 ;
  assign n15268 = n14947 & ~n15267 ;
  assign n15269 = n15268 ^ n14933 ;
  assign n15270 = n15269 ^ n14898 ;
  assign n15271 = n14913 & n15270 ;
  assign n15272 = n15271 ^ n14898 ;
  assign n15273 = n15272 ^ n14878 ;
  assign n15274 = ~n14879 & ~n15273 ;
  assign n15275 = n15274 ^ n14878 ;
  assign n15278 = n15277 ^ n15275 ;
  assign n15288 = n3484 & n12149 ;
  assign n15280 = n14498 ^ n12143 ;
  assign n15281 = n12143 ^ x29 ;
  assign n15282 = n15281 ^ x28 ;
  assign n15283 = n15282 ^ n12143 ;
  assign n15284 = ~n15280 & n15283 ;
  assign n15285 = n15284 ^ n12143 ;
  assign n15286 = n650 & n15285 ;
  assign n15287 = n15286 ^ x29 ;
  assign n15289 = n15288 ^ n15287 ;
  assign n15279 = n831 & ~n12151 ;
  assign n15290 = n15289 ^ n15279 ;
  assign n15291 = n15290 ^ n15275 ;
  assign n15292 = ~n15278 & n15291 ;
  assign n15293 = n15292 ^ n15275 ;
  assign n15296 = n15295 ^ n15293 ;
  assign n15299 = n12235 ^ n12196 ;
  assign n15302 = n3726 & ~n15299 ;
  assign n15300 = n15299 ^ n12151 ;
  assign n15301 = n3520 & n15300 ;
  assign n15303 = n15302 ^ n15301 ;
  assign n15304 = n15303 ^ n15295 ;
  assign n15298 = n12160 & n24214 ;
  assign n15305 = n15304 ^ n15298 ;
  assign n15297 = ~n3733 & n12152 ;
  assign n15306 = n15305 ^ n15297 ;
  assign n15307 = n15296 & n15306 ;
  assign n15308 = n15307 ^ n15295 ;
  assign n15310 = n15309 ^ n15308 ;
  assign n15311 = n12236 ^ n12197 ;
  assign n15312 = n15311 ^ n12149 ;
  assign n15314 = n15312 ^ n12151 ;
  assign n15313 = n15312 ^ n12152 ;
  assign n15315 = n15314 ^ n15313 ;
  assign n15316 = n15314 ^ x30 ;
  assign n15317 = n15316 ^ n15314 ;
  assign n15318 = ~n15315 & n15317 ;
  assign n15319 = n15318 ^ n15314 ;
  assign n15320 = ~n3520 & n15319 ;
  assign n15321 = n15320 ^ n15312 ;
  assign n15330 = n15321 ^ n15309 ;
  assign n15322 = n15321 ^ n14485 ;
  assign n15325 = n15322 ^ n12149 ;
  assign n15326 = n15325 ^ n15322 ;
  assign n15327 = n3520 & n15326 ;
  assign n15328 = n15327 ^ n15322 ;
  assign n15329 = ~x31 & ~n15328 ;
  assign n15331 = n15330 ^ n15329 ;
  assign n15332 = ~n15310 & n15331 ;
  assign n15333 = n15332 ^ n15309 ;
  assign n15334 = n15333 ^ n14843 ;
  assign n15335 = n14845 & ~n15334 ;
  assign n15336 = n15335 ^ n14843 ;
  assign n15339 = n15338 ^ n15336 ;
  assign n15343 = ~n12136 & n12861 ;
  assign n15342 = n446 & n12130 ;
  assign n15344 = n15343 ^ n15342 ;
  assign n15345 = n15344 ^ x26 ;
  assign n15341 = ~n487 & ~n12129 ;
  assign n15346 = n15345 ^ n15341 ;
  assign n15340 = ~n3501 & n13737 ;
  assign n15347 = n15346 ^ n15340 ;
  assign n15348 = n15347 ^ n15336 ;
  assign n15349 = ~n15339 & n15348 ;
  assign n15337 = n15336 ^ n14829 ;
  assign n15350 = n15349 ^ n15337 ;
  assign n15351 = ~n14830 & ~n15350 ;
  assign n15352 = n15351 ^ n14829 ;
  assign n15353 = n15352 ^ n14818 ;
  assign n15354 = ~n14820 & n15353 ;
  assign n15355 = n15354 ^ n14819 ;
  assign n15357 = n15356 ^ n15355 ;
  assign n14805 = n12260 & n14027 ;
  assign n14804 = n4684 & n12376 ;
  assign n14806 = n14805 ^ n14804 ;
  assign n14807 = n14806 ^ x20 ;
  assign n14803 = n4683 & ~n12108 ;
  assign n14808 = n14807 ^ n14803 ;
  assign n14802 = n4916 & n11972 ;
  assign n14809 = n14808 ^ n14802 ;
  assign n15358 = n15355 ^ n14809 ;
  assign n15359 = ~n15357 & ~n15358 ;
  assign n14810 = n14809 ^ n14800 ;
  assign n15360 = n15359 ^ n14810 ;
  assign n15361 = n14801 & n15360 ;
  assign n15362 = n15361 ^ n14800 ;
  assign n15364 = n15363 ^ n15362 ;
  assign n15366 = n12656 & n20731 ;
  assign n15365 = n5700 & ~n12705 ;
  assign n15367 = n15366 ^ n15365 ;
  assign n15368 = n15367 ^ n5694 ;
  assign n15369 = n15367 ^ x17 ;
  assign n15373 = n15369 ^ n5696 ;
  assign n15374 = ~x16 & ~n12724 ;
  assign n15375 = n15373 & n15374 ;
  assign n15371 = n5696 & ~n12756 ;
  assign n15370 = ~n12755 & n15369 ;
  assign n15372 = n15371 ^ n15370 ;
  assign n15376 = n15375 ^ n15372 ;
  assign n15377 = ~n15368 & ~n15376 ;
  assign n15378 = n15377 ^ n15362 ;
  assign n15379 = n15364 & ~n15378 ;
  assign n15380 = n15379 ^ n15377 ;
  assign n14789 = n14672 ^ n14448 ;
  assign n14786 = n14785 ^ n14709 ;
  assign n14787 = ~n14711 & n14786 ;
  assign n14788 = n14787 ^ n14709 ;
  assign n14790 = n14789 ^ n14788 ;
  assign n14696 = n5700 & n12755 ;
  assign n14689 = n12971 ^ x17 ;
  assign n14690 = n14689 ^ x16 ;
  assign n14691 = n14690 ^ n12971 ;
  assign n14692 = ~n12973 & n14691 ;
  assign n14693 = n14692 ^ n12971 ;
  assign n14694 = n5693 & n14693 ;
  assign n14695 = n14694 ^ x17 ;
  assign n14697 = n14696 ^ n14695 ;
  assign n14688 = ~n12705 & n20731 ;
  assign n14698 = n14697 ^ n14688 ;
  assign n14791 = n14790 ^ n14698 ;
  assign n15381 = n15380 ^ n14791 ;
  assign n15383 = ~n12855 & n15382 ;
  assign n15386 = n15385 ^ n15380 ;
  assign n15384 = n15380 ^ x13 ;
  assign n15387 = n15386 ^ n15384 ;
  assign n15388 = n15383 & ~n15387 ;
  assign n15389 = n15388 ^ n15386 ;
  assign n15390 = ~n15381 & n15389 ;
  assign n15391 = n15390 ^ n15380 ;
  assign n15392 = n14687 & ~n15391 ;
  assign n14686 = n14685 ^ n14676 ;
  assign n15393 = n15392 ^ n14686 ;
  assign n15394 = n15391 ^ n14687 ;
  assign n15395 = n15394 ^ n15392 ;
  assign n15396 = n6070 & ~n15395 ;
  assign n15397 = n15396 ^ n14686 ;
  assign n15398 = n15397 ^ n15396 ;
  assign n15405 = n15377 ^ n15364 ;
  assign n15403 = n8435 & ~n14221 ;
  assign n15400 = ~n6074 & ~n12855 ;
  assign n15399 = ~n6072 & n12971 ;
  assign n15401 = n15400 ^ n15399 ;
  assign n15402 = n15401 ^ n6061 ;
  assign n15404 = n15403 ^ n15402 ;
  assign n20688 = n15405 ^ n15404 ;
  assign n15406 = ~n15404 & ~n15405 ;
  assign n20689 = n20688 ^ n15406 ;
  assign n16323 = ~n12367 & n20731 ;
  assign n16321 = n5703 & ~n12872 ;
  assign n16318 = n5700 & ~n12613 ;
  assign n16317 = n5702 & n12656 ;
  assign n16319 = n16318 ^ n16317 ;
  assign n16320 = n16319 ^ x17 ;
  assign n16322 = n16321 ^ n16320 ;
  assign n16324 = n16323 ^ n16322 ;
  assign n15603 = n15350 ^ n14828 ;
  assign n15515 = n12137 & n12861 ;
  assign n15514 = n446 & ~n12136 ;
  assign n15516 = n15515 ^ n15514 ;
  assign n15517 = n15516 ^ n65 ;
  assign n15518 = n15516 ^ x26 ;
  assign n15522 = n15518 ^ n67 ;
  assign n15523 = ~x25 & ~n13817 ;
  assign n15524 = n15522 & n15523 ;
  assign n15520 = n67 & ~n13818 ;
  assign n15519 = ~n12130 & n15518 ;
  assign n15521 = n15520 ^ n15519 ;
  assign n15525 = n15524 ^ n15521 ;
  assign n15526 = ~n15517 & ~n15525 ;
  assign n15497 = n15331 ^ n15308 ;
  assign n15476 = ~n12138 & n12861 ;
  assign n15475 = n446 & n12137 ;
  assign n15477 = n15476 ^ n15475 ;
  assign n15478 = n15477 ^ n65 ;
  assign n15479 = n15477 ^ x26 ;
  assign n15480 = n15479 ^ n67 ;
  assign n15481 = n15480 ^ x25 ;
  assign n15482 = n15481 ^ n12136 ;
  assign n15483 = n15482 ^ n15479 ;
  assign n15484 = n15483 ^ n14128 ;
  assign n15485 = n15484 ^ n15483 ;
  assign n15486 = n15479 & ~n15485 ;
  assign n15487 = n15486 ^ n15480 ;
  assign n15488 = n15483 ^ n12136 ;
  assign n15489 = ~n15485 & ~n15488 ;
  assign n15490 = n15489 ^ n12136 ;
  assign n15491 = ~n15480 & n15490 ;
  assign n15492 = ~n15487 & n15491 ;
  assign n15493 = n15492 ^ n15489 ;
  assign n15494 = n15493 ^ n67 ;
  assign n15495 = n15494 ^ n12136 ;
  assign n15496 = ~n15478 & ~n15495 ;
  assign n15498 = n15497 ^ n15496 ;
  assign n15509 = n3484 & ~n12142 ;
  assign n15507 = n15497 ^ x29 ;
  assign n15500 = n14476 ^ n12207 ;
  assign n15502 = n15500 ^ n4536 ;
  assign n15503 = n15502 ^ n15500 ;
  assign n15504 = ~n14476 & ~n15503 ;
  assign n15505 = n15504 ^ n15500 ;
  assign n15506 = n650 & ~n15505 ;
  assign n15508 = n15507 ^ n15506 ;
  assign n15510 = n15509 ^ n15508 ;
  assign n15499 = n831 & n12143 ;
  assign n15511 = n15510 ^ n15499 ;
  assign n15512 = ~n15498 & n15511 ;
  assign n15513 = n15512 ^ n15497 ;
  assign n15527 = n15526 ^ n15513 ;
  assign n15528 = n15333 ^ n14845 ;
  assign n15529 = n15528 ^ n15513 ;
  assign n15530 = n15527 & ~n15529 ;
  assign n15531 = n15530 ^ n15528 ;
  assign n15604 = n15603 ^ n15531 ;
  assign n15474 = n15347 ^ n15339 ;
  assign n15532 = n15531 ^ n15474 ;
  assign n15472 = ~n4496 & n12117 ;
  assign n15470 = n4492 & n13196 ;
  assign n15467 = n4504 & n12121 ;
  assign n15466 = n4491 & ~n12110 ;
  assign n15468 = n15467 ^ n15466 ;
  assign n15469 = n15468 ^ x23 ;
  assign n15471 = n15470 ^ n15469 ;
  assign n15473 = n15472 ^ n15471 ;
  assign n15601 = n15531 ^ n15473 ;
  assign n15602 = n15532 & ~n15601 ;
  assign n15605 = n15604 ^ n15602 ;
  assign n15614 = n4916 & ~n12256 ;
  assign n15607 = n12260 ^ x20 ;
  assign n15608 = n15607 ^ x19 ;
  assign n15609 = n15608 ^ n12260 ;
  assign n15610 = n13053 & n15609 ;
  assign n15611 = n15610 ^ n12260 ;
  assign n15612 = n4678 & n15611 ;
  assign n15613 = n15612 ^ x20 ;
  assign n15615 = n15614 ^ n15613 ;
  assign n15606 = ~n12262 & n14027 ;
  assign n15616 = n15615 ^ n15606 ;
  assign n16264 = n15616 ^ n15603 ;
  assign n16265 = n15605 & ~n16264 ;
  assign n16266 = n16265 ^ n15603 ;
  assign n16267 = n16266 ^ x20 ;
  assign n16259 = n11972 ^ n4685 ;
  assign n16260 = n16259 ^ n11972 ;
  assign n16261 = ~n12270 & n16260 ;
  assign n16262 = n16261 ^ n11972 ;
  assign n16263 = n4678 & n16262 ;
  assign n16268 = n16267 ^ n16263 ;
  assign n16256 = n4916 & n12260 ;
  assign n16269 = n16268 ^ n16256 ;
  assign n16255 = ~n12256 & n14027 ;
  assign n16270 = n16269 ^ n16255 ;
  assign n16311 = n15357 ^ n14809 ;
  assign n16254 = n15352 ^ n14820 ;
  assign n16312 = n16311 ^ n16254 ;
  assign n16313 = n16312 ^ n16311 ;
  assign n16314 = n16313 ^ n16266 ;
  assign n16315 = n16270 & ~n16314 ;
  assign n16316 = n16315 ^ n16312 ;
  assign n16325 = n16324 ^ n16316 ;
  assign n16280 = n5700 & ~n12367 ;
  assign n16273 = n12613 ^ x17 ;
  assign n16274 = n16273 ^ x16 ;
  assign n16275 = n16274 ^ n12613 ;
  assign n16276 = ~n13111 & n16275 ;
  assign n16277 = n16276 ^ n12613 ;
  assign n16278 = n5693 & ~n16277 ;
  assign n16279 = n16278 ^ x17 ;
  assign n16281 = n16280 ^ n16279 ;
  assign n16272 = ~n12108 & n20731 ;
  assign n16282 = n16281 ^ n16272 ;
  assign n16271 = n16270 ^ n16254 ;
  assign n16283 = n16282 ^ n16271 ;
  assign n15617 = n15616 ^ n15605 ;
  assign n15571 = n15528 ^ n15527 ;
  assign n15542 = n15511 ^ n15496 ;
  assign n15537 = n4504 & n12130 ;
  assign n15536 = n4491 & n12121 ;
  assign n15538 = n15537 ^ n15536 ;
  assign n15539 = n15538 ^ x23 ;
  assign n15535 = n4492 & ~n13606 ;
  assign n15540 = n15539 ^ n15535 ;
  assign n15534 = ~n4496 & ~n12129 ;
  assign n15541 = n15540 ^ n15534 ;
  assign n15543 = n15542 ^ n15541 ;
  assign n15555 = n3484 & n12143 ;
  assign n15544 = n15306 ^ n15293 ;
  assign n15553 = n15544 ^ x29 ;
  assign n15548 = n12142 ^ n4536 ;
  assign n15549 = n15548 ^ n12142 ;
  assign n15550 = ~n14298 & n15549 ;
  assign n15551 = n15550 ^ n12142 ;
  assign n15552 = n650 & ~n15551 ;
  assign n15554 = n15553 ^ n15552 ;
  assign n15556 = n15555 ^ n15554 ;
  assign n15546 = n831 & n12149 ;
  assign n15557 = n15556 ^ n15546 ;
  assign n15561 = n12207 & n12861 ;
  assign n15560 = n446 & ~n12138 ;
  assign n15562 = n15561 ^ n15560 ;
  assign n15563 = n15562 ^ x26 ;
  assign n15559 = ~n487 & n12137 ;
  assign n15564 = n15563 ^ n15559 ;
  assign n15558 = ~n3501 & ~n13939 ;
  assign n15565 = n15564 ^ n15558 ;
  assign n15566 = n15565 ^ n15544 ;
  assign n15567 = n15557 & n15566 ;
  assign n15545 = n15544 ^ n15542 ;
  assign n15568 = n15567 ^ n15545 ;
  assign n15569 = ~n15543 & ~n15568 ;
  assign n15570 = n15569 ^ n15542 ;
  assign n15572 = n15571 ^ n15570 ;
  assign n15581 = ~n4496 & n12121 ;
  assign n15574 = n12117 ^ x23 ;
  assign n15575 = n15574 ^ x22 ;
  assign n15576 = n15575 ^ n12117 ;
  assign n15577 = ~n13586 & n15576 ;
  assign n15578 = n15577 ^ n12117 ;
  assign n15579 = n4488 & n15578 ;
  assign n15580 = n15579 ^ x23 ;
  assign n15582 = n15581 ^ n15580 ;
  assign n15573 = n4504 & ~n12129 ;
  assign n15583 = n15582 ^ n15573 ;
  assign n15584 = n15583 ^ n15570 ;
  assign n15585 = n15572 & ~n15584 ;
  assign n15586 = n15585 ^ n15583 ;
  assign n15618 = n15617 ^ n15586 ;
  assign n15533 = n15532 ^ n15473 ;
  assign n15587 = n15586 ^ n15533 ;
  assign n15596 = n4916 & ~n12262 ;
  assign n15589 = n12256 ^ x20 ;
  assign n15590 = n15589 ^ x19 ;
  assign n15591 = n15590 ^ n12256 ;
  assign n15592 = n13052 & n15591 ;
  assign n15593 = n15592 ^ n12256 ;
  assign n15594 = n4678 & ~n15593 ;
  assign n15595 = n15594 ^ x20 ;
  assign n15597 = n15596 ^ n15595 ;
  assign n15588 = ~n12220 & n14027 ;
  assign n15598 = n15597 ^ n15588 ;
  assign n15599 = n15598 ^ n15586 ;
  assign n15600 = n15587 & n15599 ;
  assign n15619 = n15618 ^ n15600 ;
  assign n15623 = n5700 & ~n12108 ;
  assign n15622 = n5702 & ~n12367 ;
  assign n15624 = n15623 ^ n15622 ;
  assign n15625 = n15624 ^ x17 ;
  assign n15621 = n5703 & n12368 ;
  assign n15626 = n15625 ^ n15621 ;
  assign n15620 = n11972 & n20731 ;
  assign n15627 = n15626 ^ n15620 ;
  assign n16251 = n15627 ^ n15617 ;
  assign n16252 = n15619 & n16251 ;
  assign n16253 = n16252 ^ n15617 ;
  assign n16308 = n16271 ^ n16253 ;
  assign n16309 = ~n16283 & n16308 ;
  assign n16310 = n16309 ^ n16282 ;
  assign n16326 = n16325 ^ n16310 ;
  assign n16303 = n12755 ^ x14 ;
  assign n16292 = n12971 ^ x13 ;
  assign n16291 = n12971 ^ x14 ;
  assign n16293 = n16292 ^ n16291 ;
  assign n16294 = n12918 & n16293 ;
  assign n16295 = n16294 ^ n16292 ;
  assign n16304 = n16303 ^ n16295 ;
  assign n16296 = n12755 ^ n12705 ;
  assign n16297 = n16296 ^ n12755 ;
  assign n16298 = n12755 ^ n4899 ;
  assign n16299 = n16298 ^ n12755 ;
  assign n16300 = ~n16297 & n16299 ;
  assign n16301 = n16300 ^ n12755 ;
  assign n16302 = ~n6066 & n16301 ;
  assign n16305 = n16304 ^ n16302 ;
  assign n16306 = ~n4897 & n16305 ;
  assign n16307 = n16306 ^ n16295 ;
  assign n20661 = n16310 ^ n16307 ;
  assign n20662 = ~n16326 & n20661 ;
  assign n20663 = n20662 ^ n16307 ;
  assign n20664 = n20663 ^ n6653 ;
  assign n20647 = n4897 & ~n12855 ;
  assign n20643 = ~n6072 & n12755 ;
  assign n20642 = ~n6074 & n12971 ;
  assign n20644 = n20643 ^ n20642 ;
  assign n20648 = n20647 ^ n20644 ;
  assign n20658 = n20648 ^ x14 ;
  assign n20645 = ~n12855 & n13007 ;
  assign n20646 = n20645 ^ n20644 ;
  assign n20649 = n20648 ^ n20646 ;
  assign n20650 = n20644 ^ n6060 ;
  assign n20651 = n20650 ^ n20648 ;
  assign n20652 = n20651 ^ n6060 ;
  assign n20655 = x13 & n20652 ;
  assign n20656 = n20655 ^ n6060 ;
  assign n20657 = n20649 & n20656 ;
  assign n20659 = n20658 ^ n20657 ;
  assign n20636 = n15360 ^ n14799 ;
  assign n20638 = n20636 ^ n16324 ;
  assign n20637 = n20636 ^ n16311 ;
  assign n20639 = n20638 ^ n20637 ;
  assign n20640 = n16316 & n20639 ;
  assign n20641 = n20640 ^ n20637 ;
  assign n20660 = n20659 ^ n20641 ;
  assign n20679 = n20663 ^ n20660 ;
  assign n20680 = n20664 & ~n20679 ;
  assign n20681 = n20680 ^ n6653 ;
  assign n20674 = n20659 ^ n20636 ;
  assign n20675 = n20641 & n20674 ;
  assign n20676 = n20675 ^ n20636 ;
  assign n20691 = n20681 ^ n20676 ;
  assign n20690 = ~n20676 & ~n20681 ;
  assign n20692 = n20691 ^ n20690 ;
  assign n15407 = n15389 ^ n14791 ;
  assign n20693 = n20692 ^ n15407 ;
  assign n20665 = n20664 ^ n20660 ;
  assign n16327 = n16326 ^ n16307 ;
  assign n16329 = n16327 ^ x10 ;
  assign n16328 = n16327 ^ n16290 ;
  assign n16330 = n16329 ^ n16328 ;
  assign n16331 = ~n12855 & n16289 ;
  assign n16332 = ~n16330 & n16331 ;
  assign n16333 = n16332 ^ n16328 ;
  assign n16234 = ~x13 & ~n12724 ;
  assign n16246 = n16234 ^ n12755 ;
  assign n16248 = n6060 & ~n16246 ;
  assign n16242 = n6060 ^ x14 ;
  assign n15890 = n15598 ^ n15587 ;
  assign n15640 = n15583 ^ n15572 ;
  assign n15637 = n4916 & ~n12220 ;
  assign n15630 = n12262 ^ x20 ;
  assign n15631 = n15630 ^ x19 ;
  assign n15632 = n15631 ^ n12262 ;
  assign n15633 = ~n13713 & n15632 ;
  assign n15634 = n15633 ^ n12262 ;
  assign n15635 = n4678 & ~n15634 ;
  assign n15636 = n15635 ^ x20 ;
  assign n15638 = n15637 ^ n15636 ;
  assign n15629 = ~n12110 & n14027 ;
  assign n15639 = n15638 ^ n15629 ;
  assign n15641 = n15640 ^ n15639 ;
  assign n15653 = n15568 ^ n15541 ;
  assign n15650 = n4916 & ~n12110 ;
  assign n15643 = n14047 ^ x20 ;
  assign n15644 = n15643 ^ x19 ;
  assign n15645 = n15644 ^ n14047 ;
  assign n15646 = ~n13172 & ~n15645 ;
  assign n15647 = n15646 ^ n14047 ;
  assign n15648 = n4678 & n15647 ;
  assign n15649 = n15648 ^ x20 ;
  assign n15651 = n15650 ^ n15649 ;
  assign n15642 = n12117 & n14027 ;
  assign n15652 = n15651 ^ n15642 ;
  assign n15654 = n15653 ^ n15652 ;
  assign n15662 = ~n4496 & n12130 ;
  assign n15660 = n4492 & n13737 ;
  assign n15657 = n4504 & ~n12136 ;
  assign n15656 = n4491 & ~n12129 ;
  assign n15658 = n15657 ^ n15656 ;
  assign n15659 = n15658 ^ x23 ;
  assign n15661 = n15660 ^ n15659 ;
  assign n15663 = n15662 ^ n15661 ;
  assign n15883 = n15663 ^ n15653 ;
  assign n15655 = n15565 ^ n15557 ;
  assign n15664 = n15663 ^ n15655 ;
  assign n14832 = n14370 ^ n12138 ;
  assign n15876 = ~n3501 & n14832 ;
  assign n15669 = n3481 & ~n15312 ;
  assign n15668 = n656 & n12149 ;
  assign n15670 = n15669 ^ n15668 ;
  assign n15666 = n831 & n12152 ;
  assign n15665 = n3484 & ~n12151 ;
  assign n15667 = n15666 ^ n15665 ;
  assign n15671 = n15670 ^ n15667 ;
  assign n15672 = n15272 ^ n14879 ;
  assign n15673 = n15671 & n15672 ;
  assign n15863 = ~x29 & ~n15673 ;
  assign n15676 = n15269 ^ n14913 ;
  assign n15681 = n3481 & n15300 ;
  assign n15680 = n656 & ~n12151 ;
  assign n15682 = n15681 ^ n15680 ;
  assign n15678 = n3484 & n12152 ;
  assign n15677 = n831 & n12160 ;
  assign n15679 = n15678 ^ n15677 ;
  assign n15683 = n15682 ^ n15679 ;
  assign n15684 = n15683 ^ x29 ;
  assign n15685 = ~n15676 & n15684 ;
  assign n15698 = n15266 ^ n14947 ;
  assign n15695 = n3484 & n12160 ;
  assign n15691 = n4536 & ~n14580 ;
  assign n15692 = n15691 ^ n12152 ;
  assign n15693 = n650 & n15692 ;
  assign n15694 = n15693 ^ x29 ;
  assign n15696 = n15695 ^ n15694 ;
  assign n15686 = n831 & n12163 ;
  assign n15697 = n15696 ^ n15686 ;
  assign n15699 = n15698 ^ n15697 ;
  assign n15712 = n15263 ^ n14978 ;
  assign n15709 = n3484 & n12163 ;
  assign n15702 = n12160 ^ x29 ;
  assign n15703 = n15702 ^ x28 ;
  assign n15704 = n15703 ^ n12160 ;
  assign n15705 = ~n14866 & n15704 ;
  assign n15706 = n15705 ^ n12160 ;
  assign n15707 = n650 & n15706 ;
  assign n15708 = n15707 ^ x29 ;
  assign n15710 = n15709 ^ n15708 ;
  assign n15700 = n831 & n12167 ;
  assign n15711 = n15710 ^ n15700 ;
  assign n15713 = n15712 ^ n15711 ;
  assign n15832 = n15260 ^ n15047 ;
  assign n15726 = n15257 ^ n15097 ;
  assign n15723 = n3484 & n12168 ;
  assign n15716 = n12167 ^ x29 ;
  assign n15717 = n15716 ^ x28 ;
  assign n15718 = n15717 ^ n12167 ;
  assign n15719 = ~n14914 & n15718 ;
  assign n15720 = n15719 ^ n12167 ;
  assign n15721 = n650 & n15720 ;
  assign n15722 = n15721 ^ x29 ;
  assign n15724 = n15723 ^ n15722 ;
  assign n15714 = n831 & ~n12169 ;
  assign n15725 = n15724 ^ n15714 ;
  assign n15727 = n15726 ^ n15725 ;
  assign n15739 = n15254 ^ n15150 ;
  assign n15736 = n831 & n12175 ;
  assign n15729 = n12168 ^ x29 ;
  assign n15730 = n15729 ^ x28 ;
  assign n15731 = n15730 ^ n12168 ;
  assign n15732 = ~n14948 & n15731 ;
  assign n15733 = n15732 ^ n12168 ;
  assign n15734 = n650 & n15733 ;
  assign n15735 = n15734 ^ x29 ;
  assign n15737 = n15736 ^ n15735 ;
  assign n15728 = n3484 & ~n12169 ;
  assign n15738 = n15737 ^ n15728 ;
  assign n15740 = n15739 ^ n15738 ;
  assign n15753 = n15251 ^ n15182 ;
  assign n15750 = n3484 & n12175 ;
  assign n15743 = n12169 ^ x29 ;
  assign n15744 = n15743 ^ x28 ;
  assign n15745 = n15744 ^ n12169 ;
  assign n15746 = ~n15032 & n15745 ;
  assign n15747 = n15746 ^ n12169 ;
  assign n15748 = n650 & ~n15747 ;
  assign n15749 = n15748 ^ x29 ;
  assign n15751 = n15750 ^ n15749 ;
  assign n15741 = n831 & n12179 ;
  assign n15752 = n15751 ^ n15741 ;
  assign n15754 = n15753 ^ n15752 ;
  assign n15806 = n15248 ^ n15232 ;
  assign n15789 = n15215 ^ n15212 ;
  assign n15755 = n3520 & ~n12183 ;
  assign n15761 = n831 & ~n12183 ;
  assign n15760 = n656 & n12181 ;
  assign n15762 = n15761 ^ n15760 ;
  assign n15758 = n3484 & ~n12182 ;
  assign n15756 = n12185 ^ n12181 ;
  assign n15757 = n3481 & n15756 ;
  assign n15759 = n15758 ^ n15757 ;
  assign n15763 = n15762 ^ n15759 ;
  assign n15764 = n12182 ^ n826 ;
  assign n15765 = n650 & n15764 ;
  assign n15766 = n15765 ^ n826 ;
  assign n15767 = n12183 ^ n650 ;
  assign n15768 = n15767 ^ x29 ;
  assign n15769 = n15766 & n15768 ;
  assign n15770 = n15769 ^ n650 ;
  assign n15771 = x29 & n15770 ;
  assign n15772 = n15771 ^ x29 ;
  assign n15773 = ~n15763 & n15772 ;
  assign n15774 = ~n15755 & ~n15773 ;
  assign n15784 = n3484 & n12181 ;
  assign n15777 = n12180 ^ x29 ;
  assign n15778 = n15777 ^ x28 ;
  assign n15779 = n15778 ^ n12180 ;
  assign n15780 = ~n12225 & n15779 ;
  assign n15781 = n15780 ^ n12180 ;
  assign n15782 = n650 & n15781 ;
  assign n15783 = n15782 ^ x29 ;
  assign n15785 = n15784 ^ n15783 ;
  assign n15775 = n831 & ~n12182 ;
  assign n15786 = n15785 ^ n15775 ;
  assign n15787 = n15774 & n15786 ;
  assign n15788 = n15787 ^ n15786 ;
  assign n15790 = n15789 ^ n15788 ;
  assign n15800 = n3484 & n12180 ;
  assign n15793 = n12179 ^ x29 ;
  assign n15794 = n15793 ^ x28 ;
  assign n15795 = n15794 ^ n12179 ;
  assign n15796 = ~n15127 & n15795 ;
  assign n15797 = n15796 ^ n12179 ;
  assign n15798 = n650 & n15797 ;
  assign n15799 = n15798 ^ x29 ;
  assign n15801 = n15800 ^ n15799 ;
  assign n15791 = n831 & n12181 ;
  assign n15802 = n15801 ^ n15791 ;
  assign n15803 = n15802 ^ n15788 ;
  assign n15804 = ~n15790 & n15803 ;
  assign n15805 = n15804 ^ n15788 ;
  assign n15807 = n15806 ^ n15805 ;
  assign n15817 = n3484 & n12179 ;
  assign n15810 = n12175 ^ x29 ;
  assign n15811 = n15810 ^ x28 ;
  assign n15812 = n15811 ^ n12175 ;
  assign n15813 = ~n15048 & n15812 ;
  assign n15814 = n15813 ^ n12175 ;
  assign n15815 = n650 & n15814 ;
  assign n15816 = n15815 ^ x29 ;
  assign n15818 = n15817 ^ n15816 ;
  assign n15808 = n831 & n12180 ;
  assign n15819 = n15818 ^ n15808 ;
  assign n15820 = n15819 ^ n15805 ;
  assign n15821 = ~n15807 & ~n15820 ;
  assign n15822 = n15821 ^ n15806 ;
  assign n15823 = n15822 ^ n15752 ;
  assign n15824 = ~n15754 & ~n15823 ;
  assign n15825 = n15824 ^ n15752 ;
  assign n15826 = n15825 ^ n15738 ;
  assign n15827 = ~n15740 & n15826 ;
  assign n15828 = n15827 ^ n15738 ;
  assign n15829 = n15828 ^ n15725 ;
  assign n15830 = n15727 & n15829 ;
  assign n15831 = n15830 ^ n15725 ;
  assign n15833 = n15832 ^ n15831 ;
  assign n15843 = n3484 & n12167 ;
  assign n15841 = n15832 ^ x29 ;
  assign n15836 = n12163 ^ n4536 ;
  assign n15837 = n15836 ^ n12163 ;
  assign n15838 = ~n14880 & n15837 ;
  assign n15839 = n15838 ^ n12163 ;
  assign n15840 = n650 & n15839 ;
  assign n15842 = n15841 ^ n15840 ;
  assign n15844 = n15843 ^ n15842 ;
  assign n15834 = n831 & n12168 ;
  assign n15845 = n15844 ^ n15834 ;
  assign n15846 = ~n15833 & ~n15845 ;
  assign n15847 = n15846 ^ n15832 ;
  assign n15848 = n15847 ^ n15711 ;
  assign n15849 = ~n15713 & ~n15848 ;
  assign n15850 = n15849 ^ n15711 ;
  assign n15851 = n15850 ^ n15697 ;
  assign n15852 = n15699 & n15851 ;
  assign n15853 = n15852 ^ n15697 ;
  assign n15854 = n15685 & ~n15853 ;
  assign n15855 = n15854 ^ n15853 ;
  assign n15856 = n15676 & ~n15683 ;
  assign n15674 = n15673 ^ n15672 ;
  assign n15858 = n15674 ^ n15671 ;
  assign n15864 = ~n15856 & n15858 ;
  assign n15865 = n15855 & n15864 ;
  assign n15866 = n15863 & ~n15865 ;
  assign n15675 = x29 & ~n15674 ;
  assign n15857 = n15856 ^ n15676 ;
  assign n15859 = n15858 ^ n15672 ;
  assign n15860 = ~n15857 & ~n15859 ;
  assign n15861 = n15855 & n15860 ;
  assign n15862 = n15675 & ~n15861 ;
  assign n15867 = n15866 ^ n15862 ;
  assign n15872 = n15867 ^ x26 ;
  assign n15871 = ~n12142 & n12861 ;
  assign n15873 = n15872 ^ n15871 ;
  assign n15870 = n446 & n12207 ;
  assign n15874 = n15873 ^ n15870 ;
  assign n15869 = ~n487 & ~n12138 ;
  assign n15875 = n15874 ^ n15869 ;
  assign n15877 = n15876 ^ n15875 ;
  assign n15878 = n15290 ^ n15278 ;
  assign n15879 = n15878 ^ n15867 ;
  assign n15880 = ~n15877 & n15879 ;
  assign n15868 = n15867 ^ n15655 ;
  assign n15881 = n15880 ^ n15868 ;
  assign n15882 = n15664 & n15881 ;
  assign n15884 = n15883 ^ n15882 ;
  assign n15885 = ~n15654 & ~n15884 ;
  assign n15886 = n15885 ^ n15653 ;
  assign n15887 = n15886 ^ n15639 ;
  assign n15888 = ~n15641 & n15887 ;
  assign n15889 = n15888 ^ n15640 ;
  assign n15891 = n15890 ^ n15889 ;
  assign n15898 = n12260 & n20731 ;
  assign n15896 = n5703 & n12376 ;
  assign n15893 = n5700 & n11972 ;
  assign n15892 = n5702 & ~n12108 ;
  assign n15894 = n15893 ^ n15892 ;
  assign n15895 = n15894 ^ x17 ;
  assign n15897 = n15896 ^ n15895 ;
  assign n15899 = n15898 ^ n15897 ;
  assign n15900 = n15899 ^ n15889 ;
  assign n15901 = n15891 & ~n15900 ;
  assign n15902 = n15901 ^ n15899 ;
  assign n15628 = n15627 ^ n15619 ;
  assign n15903 = n15902 ^ n15628 ;
  assign n15431 = n12656 ^ x12 ;
  assign n15432 = n15431 ^ n12656 ;
  assign n15433 = ~x13 & x14 ;
  assign n15434 = ~n12613 & n15433 ;
  assign n15435 = n15434 ^ n12656 ;
  assign n15436 = ~n15432 & n15435 ;
  assign n15437 = n15436 ^ n12656 ;
  assign n15438 = ~n4897 & n15437 ;
  assign n15439 = n15438 ^ n4897 ;
  assign n15442 = n12656 ^ x14 ;
  assign n15443 = n15442 ^ n12656 ;
  assign n19710 = n12656 ^ n12613 ;
  assign n19711 = n19710 ^ n12656 ;
  assign n15446 = ~n15443 & ~n19711 ;
  assign n15447 = n15446 ^ n12656 ;
  assign n15448 = x11 & n15447 ;
  assign n15440 = n15439 ^ n12656 ;
  assign n15449 = n15448 ^ n15440 ;
  assign n15450 = x13 & n15449 ;
  assign n15453 = n4898 & n15450 ;
  assign n15454 = n15439 & n15453 ;
  assign n15451 = n15450 ^ x14 ;
  assign n15452 = n15451 ^ n15439 ;
  assign n15455 = n15454 ^ n15452 ;
  assign n15430 = n12705 ^ x13 ;
  assign n15456 = n15455 ^ n15430 ;
  assign n15457 = n15456 ^ n12663 ;
  assign n15458 = n15457 ^ n15456 ;
  assign n15459 = n15456 ^ n4899 ;
  assign n15460 = n12705 & ~n15459 ;
  assign n15461 = n15460 ^ n15456 ;
  assign n15462 = n15458 & ~n15461 ;
  assign n15463 = n15462 ^ n15456 ;
  assign n15464 = n4897 & ~n15463 ;
  assign n15465 = n15464 ^ n15455 ;
  assign n16239 = n15902 ^ n15465 ;
  assign n16240 = n15903 & n16239 ;
  assign n16241 = n16240 ^ n15902 ;
  assign n16243 = n16242 ^ n16241 ;
  assign n16238 = ~n6074 & ~n12705 ;
  assign n16244 = n16243 ^ n16238 ;
  assign n16237 = ~n6072 & n12656 ;
  assign n16245 = n16244 ^ n16237 ;
  assign n16249 = n16248 ^ n16245 ;
  assign n16235 = n16234 ^ n12756 ;
  assign n16236 = n6063 & ~n16235 ;
  assign n16250 = n16249 ^ n16236 ;
  assign n16284 = n16283 ^ n16253 ;
  assign n16285 = n16284 ^ n16241 ;
  assign n16286 = ~n16250 & ~n16285 ;
  assign n16287 = n16286 ^ n16284 ;
  assign n16334 = n16333 ^ n16287 ;
  assign n15417 = n6658 ^ x11 ;
  assign n15410 = n12987 ^ n6650 ;
  assign n15411 = n15410 ^ n6650 ;
  assign n15414 = ~n15411 & n15413 ;
  assign n15415 = n15414 ^ n6650 ;
  assign n15416 = ~n12855 & n15415 ;
  assign n15418 = n15417 ^ n15416 ;
  assign n15409 = n6655 & n12971 ;
  assign n15419 = n15418 ^ n15409 ;
  assign n15904 = n15903 ^ n15465 ;
  assign n15422 = n6648 & ~n12855 ;
  assign n15423 = n15422 ^ x11 ;
  assign n15424 = n15423 ^ x10 ;
  assign n15425 = ~n13007 & n15422 ;
  assign n15426 = ~n15424 & n15425 ;
  assign n15427 = n15426 ^ n15423 ;
  assign n15421 = n6650 & n12971 ;
  assign n15428 = n15427 ^ n15421 ;
  assign n15420 = n6655 & n12755 ;
  assign n15429 = n15428 ^ n15420 ;
  assign n15905 = n15904 ^ n15429 ;
  assign n16184 = n15886 ^ n15641 ;
  assign n15915 = n15884 ^ n15652 ;
  assign n15913 = ~n12262 & n20731 ;
  assign n15911 = n5703 & n13054 ;
  assign n15908 = n5700 & ~n12256 ;
  assign n15907 = n5702 & n12260 ;
  assign n15909 = n15908 ^ n15907 ;
  assign n15910 = n15909 ^ x17 ;
  assign n15912 = n15911 ^ n15910 ;
  assign n15914 = n15913 ^ n15912 ;
  assign n15916 = n15915 ^ n15914 ;
  assign n15921 = n12121 & n14027 ;
  assign n15920 = n4684 & n13196 ;
  assign n15922 = n15921 ^ n15920 ;
  assign n15923 = n15922 ^ x20 ;
  assign n15919 = n4683 & ~n12110 ;
  assign n15924 = n15923 ^ n15919 ;
  assign n15918 = n4916 & n12117 ;
  assign n15925 = n15924 ^ n15918 ;
  assign n16180 = n15925 ^ n15915 ;
  assign n15917 = n15881 ^ n15663 ;
  assign n15926 = n15925 ^ n15917 ;
  assign n15928 = n15878 ^ n15877 ;
  assign n16177 = n15928 ^ n15917 ;
  assign n15935 = ~n4496 & ~n12136 ;
  assign n15932 = n4491 & n12130 ;
  assign n15930 = n4504 & n12137 ;
  assign n15929 = n15928 ^ x23 ;
  assign n15931 = n15930 ^ n15929 ;
  assign n15933 = n15932 ^ n15931 ;
  assign n15927 = n4492 & ~n13818 ;
  assign n15934 = n15933 ^ n15927 ;
  assign n15936 = n15935 ^ n15934 ;
  assign n16159 = n15853 ^ n15684 ;
  assign n16160 = n15684 ^ n15676 ;
  assign n16161 = n16159 & ~n16160 ;
  assign n16157 = n15683 ^ n15671 ;
  assign n16158 = n16157 ^ n15672 ;
  assign n16162 = n16161 ^ n16158 ;
  assign n15945 = ~n487 & ~n12142 ;
  assign n15940 = n15853 ^ n15676 ;
  assign n15941 = n15940 ^ n15684 ;
  assign n15942 = n15941 ^ x26 ;
  assign n15939 = n446 & n12143 ;
  assign n15943 = n15942 ^ n15939 ;
  assign n15938 = n12149 & n12861 ;
  assign n15944 = n15943 ^ n15938 ;
  assign n15946 = n15945 ^ n15944 ;
  assign n15937 = ~n3501 & n14299 ;
  assign n15947 = n15946 ^ n15937 ;
  assign n15955 = n446 & n12149 ;
  assign n15951 = n15850 ^ n15699 ;
  assign n15952 = n15951 ^ x26 ;
  assign n15950 = ~n487 & n12143 ;
  assign n15953 = n15952 ^ n15950 ;
  assign n15949 = ~n12151 & n12861 ;
  assign n15954 = n15953 ^ n15949 ;
  assign n15956 = n15955 ^ n15954 ;
  assign n15948 = ~n3501 & ~n14498 ;
  assign n15957 = n15956 ^ n15948 ;
  assign n15966 = n15847 ^ n15713 ;
  assign n15961 = n12152 & n12861 ;
  assign n15960 = n446 & ~n12151 ;
  assign n15962 = n15961 ^ n15960 ;
  assign n15963 = n15962 ^ x26 ;
  assign n15959 = ~n487 & n12149 ;
  assign n15964 = n15963 ^ n15959 ;
  assign n15958 = ~n3501 & ~n15312 ;
  assign n15965 = n15964 ^ n15958 ;
  assign n15967 = n15966 ^ n15965 ;
  assign n15976 = n15845 ^ n15831 ;
  assign n15971 = n446 & n12152 ;
  assign n15970 = n12160 & n12861 ;
  assign n15972 = n15971 ^ n15970 ;
  assign n15973 = n15972 ^ x26 ;
  assign n15969 = ~n487 & ~n12151 ;
  assign n15974 = n15973 ^ n15969 ;
  assign n15968 = ~n3501 & n15300 ;
  assign n15975 = n15974 ^ n15968 ;
  assign n15977 = n15976 ^ n15975 ;
  assign n15986 = n15828 ^ n15727 ;
  assign n15981 = n12163 & n12861 ;
  assign n15980 = ~n487 & n12152 ;
  assign n15982 = n15981 ^ n15980 ;
  assign n15983 = n15982 ^ x26 ;
  assign n15979 = n446 & n12160 ;
  assign n15984 = n15983 ^ n15979 ;
  assign n15978 = ~n3501 & ~n14581 ;
  assign n15985 = n15984 ^ n15978 ;
  assign n15987 = n15986 ^ n15985 ;
  assign n16115 = n15825 ^ n15740 ;
  assign n16001 = n15822 ^ n15754 ;
  assign n15989 = n12168 & n12861 ;
  assign n15988 = n446 & n12167 ;
  assign n15990 = n15989 ^ n15988 ;
  assign n15991 = n15990 ^ n65 ;
  assign n15992 = n15990 ^ x26 ;
  assign n15996 = n15992 ^ n67 ;
  assign n15997 = ~x25 & ~n14880 ;
  assign n15998 = n15996 & n15997 ;
  assign n15994 = n67 & ~n14890 ;
  assign n15993 = ~n12163 & n15992 ;
  assign n15995 = n15994 ^ n15993 ;
  assign n15999 = n15998 ^ n15995 ;
  assign n16000 = ~n15991 & ~n15999 ;
  assign n16002 = n16001 ^ n16000 ;
  assign n16011 = n15819 ^ n15807 ;
  assign n16006 = ~n12169 & n12861 ;
  assign n16005 = n446 & n12168 ;
  assign n16007 = n16006 ^ n16005 ;
  assign n16008 = n16007 ^ x26 ;
  assign n16004 = ~n487 & n12167 ;
  assign n16009 = n16008 ^ n16004 ;
  assign n16003 = ~n3501 & ~n14915 ;
  assign n16010 = n16009 ^ n16003 ;
  assign n16012 = n16011 ^ n16010 ;
  assign n16035 = n15802 ^ n15790 ;
  assign n16014 = n446 & ~n12169 ;
  assign n16013 = n12175 & n12861 ;
  assign n16015 = n16014 ^ n16013 ;
  assign n16016 = n16015 ^ n65 ;
  assign n16017 = n16015 ^ x26 ;
  assign n16018 = n16017 ^ n67 ;
  assign n16019 = n16018 ^ x25 ;
  assign n16020 = n16019 ^ n12168 ;
  assign n16021 = n16020 ^ n16017 ;
  assign n16022 = n16021 ^ n14948 ;
  assign n16023 = n16022 ^ n16021 ;
  assign n16024 = n16017 & ~n16023 ;
  assign n16025 = n16024 ^ n16018 ;
  assign n16026 = n16021 ^ n12168 ;
  assign n16027 = ~n16023 & ~n16026 ;
  assign n16028 = n16027 ^ n12168 ;
  assign n16029 = ~n16018 & ~n16028 ;
  assign n16030 = ~n16025 & n16029 ;
  assign n16031 = n16030 ^ n16027 ;
  assign n16032 = n16031 ^ n67 ;
  assign n16033 = n16032 ^ n12168 ;
  assign n16034 = ~n16016 & n16033 ;
  assign n16036 = n16035 ^ n16034 ;
  assign n16042 = n12179 & n12861 ;
  assign n16041 = ~n487 & ~n12169 ;
  assign n16043 = n16042 ^ n16041 ;
  assign n16044 = n16043 ^ x26 ;
  assign n16040 = n446 & n12175 ;
  assign n16045 = n16044 ^ n16040 ;
  assign n16039 = ~n3501 & n15035 ;
  assign n16046 = n16045 ^ n16039 ;
  assign n16105 = n16046 ^ n16034 ;
  assign n16037 = n15786 ^ n15773 ;
  assign n16038 = n16037 ^ n15755 ;
  assign n16047 = n16046 ^ n16038 ;
  assign n16052 = n12180 & n12861 ;
  assign n16051 = n446 & n12179 ;
  assign n16053 = n16052 ^ n16051 ;
  assign n16054 = n16053 ^ x26 ;
  assign n16050 = ~n487 & n12175 ;
  assign n16055 = n16054 ^ n16050 ;
  assign n16049 = ~n3501 & ~n15049 ;
  assign n16056 = n16055 ^ n16049 ;
  assign n16048 = n15771 ^ n15763 ;
  assign n16057 = n16056 ^ n16048 ;
  assign n16069 = ~n3501 & ~n15128 ;
  assign n16066 = n446 & n12180 ;
  assign n16064 = n12181 & n12861 ;
  assign n16059 = n826 & ~n12183 ;
  assign n16058 = n650 & ~n12182 ;
  assign n16060 = n16059 ^ n16058 ;
  assign n16063 = n16060 ^ x26 ;
  assign n16065 = n16064 ^ n16063 ;
  assign n16067 = n16066 ^ n16065 ;
  assign n16062 = ~n487 & n12179 ;
  assign n16068 = n16067 ^ n16062 ;
  assign n16070 = n16069 ^ n16068 ;
  assign n16071 = n650 & ~n12183 ;
  assign n16072 = n64 & ~n12182 ;
  assign n16073 = x26 & ~n16072 ;
  assign n16074 = ~n12183 & n16073 ;
  assign n16075 = n7214 & n16074 ;
  assign n16076 = n16075 ^ n16073 ;
  assign n16084 = ~n3501 & n15756 ;
  assign n16081 = ~n12183 & n12861 ;
  assign n16080 = n446 & ~n12182 ;
  assign n16082 = n16081 ^ n16080 ;
  assign n16079 = ~n487 & n12181 ;
  assign n16083 = n16082 ^ n16079 ;
  assign n16085 = n16084 ^ n16083 ;
  assign n16086 = n16076 & ~n16085 ;
  assign n16087 = ~n16071 & ~n16086 ;
  assign n16091 = ~n12182 & n12861 ;
  assign n16090 = n446 & n12181 ;
  assign n16092 = n16091 ^ n16090 ;
  assign n16093 = n16092 ^ x26 ;
  assign n16089 = ~n487 & n12180 ;
  assign n16094 = n16093 ^ n16089 ;
  assign n16088 = ~n3501 & ~n15151 ;
  assign n16095 = n16094 ^ n16088 ;
  assign n16096 = n16087 & n16095 ;
  assign n16097 = n16096 ^ n16095 ;
  assign n16098 = n16097 ^ n16060 ;
  assign n16099 = n16070 & n16098 ;
  assign n16061 = n16060 ^ n16048 ;
  assign n16100 = n16099 ^ n16061 ;
  assign n16101 = n16057 & ~n16100 ;
  assign n16102 = n16101 ^ n16056 ;
  assign n16103 = n16102 ^ n16046 ;
  assign n16104 = n16047 & n16103 ;
  assign n16106 = n16105 ^ n16104 ;
  assign n16107 = n16036 & n16106 ;
  assign n16108 = n16107 ^ n16035 ;
  assign n16109 = n16108 ^ n16010 ;
  assign n16110 = ~n16012 & ~n16109 ;
  assign n16111 = n16110 ^ n16010 ;
  assign n16112 = n16111 ^ n16000 ;
  assign n16113 = ~n16002 & ~n16112 ;
  assign n16114 = n16113 ^ n16000 ;
  assign n16116 = n16115 ^ n16114 ;
  assign n16118 = n12167 & n12861 ;
  assign n16117 = n446 & n12163 ;
  assign n16119 = n16118 ^ n16117 ;
  assign n16120 = n16119 ^ n65 ;
  assign n16121 = n16119 ^ x26 ;
  assign n16122 = n16121 ^ n67 ;
  assign n16123 = n16122 ^ x25 ;
  assign n16124 = n16123 ^ n12160 ;
  assign n16125 = n16124 ^ n16121 ;
  assign n16126 = n16125 ^ n14866 ;
  assign n16127 = n16126 ^ n16125 ;
  assign n16128 = n16121 & ~n16127 ;
  assign n16129 = n16128 ^ n16122 ;
  assign n16130 = n16125 ^ n12160 ;
  assign n16131 = ~n16127 & ~n16130 ;
  assign n16132 = n16131 ^ n12160 ;
  assign n16133 = ~n16122 & ~n16132 ;
  assign n16134 = ~n16129 & n16133 ;
  assign n16135 = n16134 ^ n16131 ;
  assign n16136 = n16135 ^ n67 ;
  assign n16137 = n16136 ^ n12160 ;
  assign n16138 = ~n16120 & n16137 ;
  assign n16139 = n16138 ^ n16114 ;
  assign n16140 = n16116 & ~n16139 ;
  assign n16141 = n16140 ^ n16115 ;
  assign n16142 = n16141 ^ n15985 ;
  assign n16143 = n15987 & ~n16142 ;
  assign n16144 = n16143 ^ n15985 ;
  assign n16145 = n16144 ^ n15975 ;
  assign n16146 = ~n15977 & n16145 ;
  assign n16147 = n16146 ^ n15975 ;
  assign n16148 = n16147 ^ n15965 ;
  assign n16149 = n15967 & n16148 ;
  assign n16150 = n16149 ^ n15965 ;
  assign n16151 = n16150 ^ n15951 ;
  assign n16152 = n15957 & n16151 ;
  assign n16153 = n16152 ^ n15951 ;
  assign n16154 = n16153 ^ n15941 ;
  assign n16155 = ~n15947 & ~n16154 ;
  assign n16156 = n16155 ^ n15941 ;
  assign n16163 = n16162 ^ n16156 ;
  assign n16170 = ~n487 & n12207 ;
  assign n16168 = n12143 & n12861 ;
  assign n16166 = n446 & ~n12142 ;
  assign n16165 = n16162 ^ x26 ;
  assign n16167 = n16166 ^ n16165 ;
  assign n16169 = n16168 ^ n16167 ;
  assign n16171 = n16170 ^ n16169 ;
  assign n16164 = ~n3501 & ~n15500 ;
  assign n16172 = n16171 ^ n16164 ;
  assign n16173 = ~n16163 & n16172 ;
  assign n16174 = n16173 ^ n16162 ;
  assign n16175 = n16174 ^ n15928 ;
  assign n16176 = n15936 & n16175 ;
  assign n16178 = n16177 ^ n16176 ;
  assign n16179 = ~n15926 & n16178 ;
  assign n16181 = n16180 ^ n16179 ;
  assign n16182 = ~n15916 & ~n16181 ;
  assign n16183 = n16182 ^ n15915 ;
  assign n16185 = n16184 ^ n16183 ;
  assign n16187 = ~n12256 & n20731 ;
  assign n16186 = n5700 & n12260 ;
  assign n16188 = n16187 ^ n16186 ;
  assign n16189 = n16188 ^ n5694 ;
  assign n16190 = n16188 ^ x17 ;
  assign n16191 = n16190 ^ n5696 ;
  assign n16192 = n14078 & n16191 ;
  assign n16193 = n16192 ^ n5696 ;
  assign n16194 = n16193 ^ x16 ;
  assign n16195 = n16194 ^ n11972 ;
  assign n16196 = n16195 ^ n16193 ;
  assign n16197 = n16193 ^ n16191 ;
  assign n16198 = n16197 ^ n16193 ;
  assign n16199 = n16196 & n16198 ;
  assign n16200 = n16199 ^ n16193 ;
  assign n16201 = ~n12270 & n16200 ;
  assign n16202 = n16201 ^ n16193 ;
  assign n16203 = ~n16189 & ~n16202 ;
  assign n16204 = n16203 ^ n16183 ;
  assign n16205 = n16185 & n16204 ;
  assign n16206 = n16205 ^ n16203 ;
  assign n16229 = n16206 ^ n15904 ;
  assign n15906 = n15899 ^ n15891 ;
  assign n16207 = n16206 ^ n15906 ;
  assign n16209 = ~n6074 & ~n12613 ;
  assign n16208 = ~n6072 & ~n12367 ;
  assign n16210 = n16209 ^ n16208 ;
  assign n16211 = n16210 ^ n6060 ;
  assign n16212 = n16211 ^ x14 ;
  assign n16222 = n8465 & n12656 ;
  assign n16221 = x13 & n12872 ;
  assign n16223 = n16222 ^ n16221 ;
  assign n16224 = ~n6063 & n16223 ;
  assign n16219 = n12871 ^ n8465 ;
  assign n16213 = n16210 ^ x14 ;
  assign n16214 = n12656 ^ x13 ;
  assign n16215 = n16214 ^ n12656 ;
  assign n16216 = ~n12871 & ~n16215 ;
  assign n16217 = n16216 ^ n12656 ;
  assign n16218 = ~n16213 & ~n16217 ;
  assign n16220 = n16219 ^ n16218 ;
  assign n16225 = n16224 ^ n16220 ;
  assign n16226 = ~n16212 & n16225 ;
  assign n16227 = n16226 ^ n16206 ;
  assign n16228 = n16207 & n16227 ;
  assign n16230 = n16229 ^ n16228 ;
  assign n16231 = n15905 & ~n16230 ;
  assign n16232 = n16231 ^ n15904 ;
  assign n16233 = n15419 & n16232 ;
  assign n16335 = n16334 ^ n16233 ;
  assign n16338 = n16230 ^ n15429 ;
  assign n16339 = n16338 ^ n13900 ;
  assign n16691 = n16226 ^ n16207 ;
  assign n16351 = n12367 ^ n12108 ;
  assign n16352 = x14 & ~n16351 ;
  assign n16353 = n16352 ^ n12108 ;
  assign n16354 = ~n4898 & n4899 ;
  assign n16355 = n16353 & n16354 ;
  assign n16356 = n16355 ^ n6068 ;
  assign n16349 = ~n6065 & n6068 ;
  assign n16350 = ~n12367 & n16349 ;
  assign n16357 = n16356 ^ n16350 ;
  assign n16358 = n4896 & ~n16357 ;
  assign n16360 = n12108 ^ x14 ;
  assign n16361 = n16360 ^ n12108 ;
  assign n16362 = ~n12367 & n16361 ;
  assign n16363 = n16362 ^ n12108 ;
  assign n16364 = x13 & ~n16363 ;
  assign n16365 = n16364 ^ n12108 ;
  assign n16366 = n16358 & ~n16365 ;
  assign n16367 = n16366 ^ n16357 ;
  assign n16342 = n12613 ^ x14 ;
  assign n16341 = n12613 ^ x13 ;
  assign n16343 = n16342 ^ n16341 ;
  assign n16344 = n16342 ^ n12777 ;
  assign n16345 = n16344 ^ n16342 ;
  assign n16346 = n16343 & ~n16345 ;
  assign n16347 = n16346 ^ n16342 ;
  assign n16348 = n4897 & n16347 ;
  assign n16368 = n16367 ^ n16348 ;
  assign n16340 = n16203 ^ n16185 ;
  assign n16369 = n16368 ^ n16340 ;
  assign n16372 = x13 ^ x11 ;
  assign n16384 = n16372 ^ x14 ;
  assign n16374 = n12367 ^ x13 ;
  assign n16373 = n12367 ^ x14 ;
  assign n16375 = n16374 ^ n16373 ;
  assign n16376 = n12277 & n16375 ;
  assign n16377 = n16376 ^ n16374 ;
  assign n16378 = n16377 ^ n12108 ;
  assign n16379 = n16378 ^ x13 ;
  assign n16380 = n16379 ^ n11972 ;
  assign n16381 = n16380 ^ n16377 ;
  assign n16382 = ~n16372 & ~n16381 ;
  assign n16383 = n16382 ^ n16378 ;
  assign n16385 = n16383 ^ n16377 ;
  assign n16386 = ~n16384 & ~n16385 ;
  assign n16387 = n16386 ^ n16377 ;
  assign n16388 = n16387 ^ n16383 ;
  assign n16389 = n16388 ^ n16383 ;
  assign n16391 = n16389 ^ n11972 ;
  assign n16392 = n16391 ^ n16389 ;
  assign n16395 = ~n16372 & n16392 ;
  assign n16396 = ~n16388 & n16395 ;
  assign n16397 = n16396 ^ n16388 ;
  assign n16398 = n16397 ^ n16383 ;
  assign n16399 = ~n4897 & n16398 ;
  assign n16400 = n16399 ^ n16377 ;
  assign n16405 = ~n12108 & n16349 ;
  assign n16406 = n16405 ^ n6068 ;
  assign n16407 = ~n16400 & ~n16406 ;
  assign n16370 = n16181 ^ n15914 ;
  assign n16408 = n16407 ^ n16370 ;
  assign n16674 = n16178 ^ n15925 ;
  assign n16420 = n16174 ^ n15936 ;
  assign n16417 = n4916 & n12121 ;
  assign n16410 = n12117 ^ x20 ;
  assign n16411 = n16410 ^ x19 ;
  assign n16412 = n16411 ^ n12117 ;
  assign n16413 = ~n13586 & n16412 ;
  assign n16414 = n16413 ^ n12117 ;
  assign n16415 = n4678 & n16414 ;
  assign n16416 = n16415 ^ x20 ;
  assign n16418 = n16417 ^ n16416 ;
  assign n16409 = ~n12129 & n14027 ;
  assign n16419 = n16418 ^ n16409 ;
  assign n16421 = n16420 ^ n16419 ;
  assign n16430 = n16172 ^ n16156 ;
  assign n16425 = n4504 & ~n12138 ;
  assign n16424 = n4491 & ~n12136 ;
  assign n16426 = n16425 ^ n16424 ;
  assign n16427 = n16426 ^ x23 ;
  assign n16423 = n4492 & n14129 ;
  assign n16428 = n16427 ^ n16423 ;
  assign n16422 = ~n4496 & n12137 ;
  assign n16429 = n16428 ^ n16422 ;
  assign n16431 = n16430 ^ n16429 ;
  assign n16440 = n16153 ^ n15947 ;
  assign n16438 = ~n4496 & ~n12138 ;
  assign n16436 = n4492 & ~n13939 ;
  assign n16433 = n4504 & n12207 ;
  assign n16432 = n4491 & n12137 ;
  assign n16434 = n16433 ^ n16432 ;
  assign n16435 = n16434 ^ x23 ;
  assign n16437 = n16436 ^ n16435 ;
  assign n16439 = n16438 ^ n16437 ;
  assign n16441 = n16440 ^ n16439 ;
  assign n16450 = n16150 ^ n15957 ;
  assign n16448 = ~n4496 & n12207 ;
  assign n16446 = n4492 & n14832 ;
  assign n16443 = n4504 & ~n12142 ;
  assign n16442 = n4491 & ~n12138 ;
  assign n16444 = n16443 ^ n16442 ;
  assign n16445 = n16444 ^ x23 ;
  assign n16447 = n16446 ^ n16445 ;
  assign n16449 = n16448 ^ n16447 ;
  assign n16451 = n16450 ^ n16449 ;
  assign n16460 = n16147 ^ n15967 ;
  assign n16455 = n4504 & n12143 ;
  assign n16454 = n4491 & n12207 ;
  assign n16456 = n16455 ^ n16454 ;
  assign n16457 = n16456 ^ x23 ;
  assign n16453 = n4492 & ~n15500 ;
  assign n16458 = n16457 ^ n16453 ;
  assign n16452 = ~n4496 & ~n12142 ;
  assign n16459 = n16458 ^ n16452 ;
  assign n16461 = n16460 ^ n16459 ;
  assign n16470 = n16144 ^ n15977 ;
  assign n16465 = n4504 & n12149 ;
  assign n16464 = n4491 & ~n12142 ;
  assign n16466 = n16465 ^ n16464 ;
  assign n16467 = n16466 ^ x23 ;
  assign n16463 = n4492 & n14299 ;
  assign n16468 = n16467 ^ n16463 ;
  assign n16462 = ~n4496 & n12143 ;
  assign n16469 = n16468 ^ n16462 ;
  assign n16471 = n16470 ^ n16469 ;
  assign n16480 = n16141 ^ n15987 ;
  assign n16475 = n4504 & ~n12151 ;
  assign n16474 = n4491 & n12143 ;
  assign n16476 = n16475 ^ n16474 ;
  assign n16477 = n16476 ^ x23 ;
  assign n16473 = n4492 & ~n14498 ;
  assign n16478 = n16477 ^ n16473 ;
  assign n16472 = ~n4496 & n12149 ;
  assign n16479 = n16478 ^ n16472 ;
  assign n16481 = n16480 ^ n16479 ;
  assign n16490 = n16139 ^ n16115 ;
  assign n16485 = n4504 & n12152 ;
  assign n16484 = n4491 & n12149 ;
  assign n16486 = n16485 ^ n16484 ;
  assign n16487 = n16486 ^ x23 ;
  assign n16483 = n4492 & ~n15312 ;
  assign n16488 = n16487 ^ n16483 ;
  assign n16482 = ~n4496 & ~n12151 ;
  assign n16489 = n16488 ^ n16482 ;
  assign n16491 = n16490 ^ n16489 ;
  assign n16500 = n16111 ^ n16002 ;
  assign n16498 = ~n4496 & n12152 ;
  assign n16496 = n4492 & n15300 ;
  assign n16493 = n4504 & n12160 ;
  assign n16492 = n4491 & ~n12151 ;
  assign n16494 = n16493 ^ n16492 ;
  assign n16495 = n16494 ^ x23 ;
  assign n16497 = n16496 ^ n16495 ;
  assign n16499 = n16498 ^ n16497 ;
  assign n16501 = n16500 ^ n16499 ;
  assign n16506 = n4504 & n12167 ;
  assign n16505 = n4491 & n12160 ;
  assign n16507 = n16506 ^ n16505 ;
  assign n16503 = ~n4496 & n12163 ;
  assign n16502 = n4492 & ~n14867 ;
  assign n16504 = n16503 ^ n16502 ;
  assign n16508 = n16507 ^ n16504 ;
  assign n16509 = n16508 ^ x23 ;
  assign n16516 = n4504 & n12163 ;
  assign n16515 = n4491 & n12152 ;
  assign n16517 = n16516 ^ n16515 ;
  assign n16513 = ~n4496 & n12160 ;
  assign n16512 = n4492 & ~n14581 ;
  assign n16514 = n16513 ^ n16512 ;
  assign n16518 = n16517 ^ n16514 ;
  assign n16510 = n16108 ^ n16012 ;
  assign n16511 = n16510 ^ n16508 ;
  assign n16519 = n16518 ^ n16511 ;
  assign n16520 = n16509 & ~n16519 ;
  assign n16532 = n16102 ^ n16047 ;
  assign n16530 = n4504 & n12168 ;
  assign n16528 = ~n4496 & n12167 ;
  assign n16521 = n12163 ^ x23 ;
  assign n16522 = n16521 ^ x22 ;
  assign n16523 = n16522 ^ n12163 ;
  assign n16524 = ~n14880 & n16523 ;
  assign n16525 = n16524 ^ n12163 ;
  assign n16526 = n4488 & n16525 ;
  assign n16527 = n16526 ^ x23 ;
  assign n16529 = n16528 ^ n16527 ;
  assign n16531 = n16530 ^ n16529 ;
  assign n16533 = n16532 ^ n16531 ;
  assign n16545 = n16100 ^ n16056 ;
  assign n16542 = ~n4496 & n12168 ;
  assign n16535 = n12167 ^ x23 ;
  assign n16536 = n16535 ^ x22 ;
  assign n16537 = n16536 ^ n12167 ;
  assign n16538 = ~n14914 & n16537 ;
  assign n16539 = n16538 ^ n12167 ;
  assign n16540 = n4488 & n16539 ;
  assign n16541 = n16540 ^ x23 ;
  assign n16543 = n16542 ^ n16541 ;
  assign n16534 = n4504 & ~n12169 ;
  assign n16544 = n16543 ^ n16534 ;
  assign n16546 = n16545 ^ n16544 ;
  assign n16554 = ~n4496 & ~n12169 ;
  assign n14949 = n14948 ^ n12168 ;
  assign n16552 = n4492 & ~n14949 ;
  assign n16549 = n4504 & n12175 ;
  assign n16548 = n4491 & n12168 ;
  assign n16550 = n16549 ^ n16548 ;
  assign n16551 = n16550 ^ x23 ;
  assign n16553 = n16552 ^ n16551 ;
  assign n16555 = n16554 ^ n16553 ;
  assign n16627 = n16555 ^ n16544 ;
  assign n16547 = n16097 ^ n16070 ;
  assign n16556 = n16555 ^ n16547 ;
  assign n16565 = n16086 ^ n16071 ;
  assign n16566 = n16565 ^ n16095 ;
  assign n16563 = ~n4496 & n12175 ;
  assign n16561 = n4492 & n15035 ;
  assign n16558 = n4504 & n12179 ;
  assign n16557 = n4491 & ~n12169 ;
  assign n16559 = n16558 ^ n16557 ;
  assign n16560 = n16559 ^ x23 ;
  assign n16562 = n16561 ^ n16560 ;
  assign n16564 = n16563 ^ n16562 ;
  assign n16567 = n16566 ^ n16564 ;
  assign n16077 = n16076 ^ x26 ;
  assign n16609 = n16085 ^ n16077 ;
  assign n16576 = n64 & ~n12183 ;
  assign n16577 = n4488 & ~n12182 ;
  assign n16578 = x23 & ~n16577 ;
  assign n16579 = ~n12183 & n16578 ;
  assign n16580 = ~n4500 & n16579 ;
  assign n16581 = n16580 ^ n16578 ;
  assign n16588 = ~n4496 & ~n12182 ;
  assign n16587 = n4491 & n12181 ;
  assign n16589 = n16588 ^ n16587 ;
  assign n16585 = n4504 & ~n12183 ;
  assign n16584 = n4492 & n15756 ;
  assign n16586 = n16585 ^ n16584 ;
  assign n16590 = n16589 ^ n16586 ;
  assign n16591 = n16581 & ~n16590 ;
  assign n16592 = ~n16576 & ~n16591 ;
  assign n16596 = n4504 & ~n12182 ;
  assign n16595 = n4491 & n12180 ;
  assign n16597 = n16596 ^ n16595 ;
  assign n16598 = n16597 ^ x23 ;
  assign n16594 = n4492 & ~n15151 ;
  assign n16599 = n16598 ^ n16594 ;
  assign n16593 = ~n4496 & n12181 ;
  assign n16600 = n16599 ^ n16593 ;
  assign n16601 = n16592 & n16600 ;
  assign n16602 = n16601 ^ n16600 ;
  assign n16574 = ~n4496 & n12180 ;
  assign n16572 = n4492 & ~n15128 ;
  assign n16569 = n4504 & n12181 ;
  assign n16568 = n4491 & n12179 ;
  assign n16570 = n16569 ^ n16568 ;
  assign n16571 = n16570 ^ x23 ;
  assign n16573 = n16572 ^ n16571 ;
  assign n16575 = n16574 ^ n16573 ;
  assign n16603 = n16602 ^ n16575 ;
  assign n16605 = ~n7434 & ~n12183 ;
  assign n16604 = n16602 ^ n16072 ;
  assign n16606 = n16605 ^ n16604 ;
  assign n16607 = n16603 & n16606 ;
  assign n16608 = n16607 ^ n16602 ;
  assign n16610 = n16609 ^ n16608 ;
  assign n16614 = n4504 & n12180 ;
  assign n16613 = n4491 & n12175 ;
  assign n16615 = n16614 ^ n16613 ;
  assign n16616 = n16615 ^ x23 ;
  assign n16612 = n4492 & ~n15049 ;
  assign n16617 = n16616 ^ n16612 ;
  assign n16611 = ~n4496 & n12179 ;
  assign n16618 = n16617 ^ n16611 ;
  assign n16619 = n16618 ^ n16608 ;
  assign n16620 = ~n16610 & n16619 ;
  assign n16621 = n16620 ^ n16618 ;
  assign n16622 = n16621 ^ n16564 ;
  assign n16623 = n16567 & ~n16622 ;
  assign n16624 = n16623 ^ n16566 ;
  assign n16625 = n16624 ^ n16555 ;
  assign n16626 = n16556 & n16625 ;
  assign n16628 = n16627 ^ n16626 ;
  assign n16629 = n16546 & ~n16628 ;
  assign n16630 = n16629 ^ n16545 ;
  assign n16631 = n16630 ^ n16531 ;
  assign n16632 = n16533 & n16631 ;
  assign n16633 = n16632 ^ n16531 ;
  assign n16634 = n16106 ^ n16035 ;
  assign n16636 = n16633 & n16634 ;
  assign n16635 = n16634 ^ n16633 ;
  assign n16637 = n16636 ^ n16635 ;
  assign n16638 = n16636 ^ n16510 ;
  assign n16639 = n16518 ^ x23 ;
  assign n16640 = n16639 ^ n16636 ;
  assign n16641 = n16638 & ~n16640 ;
  assign n16642 = n16641 ^ n16510 ;
  assign n16643 = n16637 & ~n16642 ;
  assign n16644 = n16520 & n16643 ;
  assign n16645 = n16644 ^ n16642 ;
  assign n16646 = n16645 ^ n16499 ;
  assign n16647 = ~n16501 & n16646 ;
  assign n16648 = n16647 ^ n16499 ;
  assign n16649 = n16648 ^ n16489 ;
  assign n16650 = ~n16491 & n16649 ;
  assign n16651 = n16650 ^ n16489 ;
  assign n16652 = n16651 ^ n16479 ;
  assign n16653 = ~n16481 & n16652 ;
  assign n16654 = n16653 ^ n16479 ;
  assign n16655 = n16654 ^ n16469 ;
  assign n16656 = ~n16471 & n16655 ;
  assign n16657 = n16656 ^ n16469 ;
  assign n16658 = n16657 ^ n16459 ;
  assign n16659 = n16461 & n16658 ;
  assign n16660 = n16659 ^ n16459 ;
  assign n16661 = n16660 ^ n16449 ;
  assign n16662 = n16451 & n16661 ;
  assign n16663 = n16662 ^ n16449 ;
  assign n16664 = n16663 ^ n16439 ;
  assign n16665 = ~n16441 & n16664 ;
  assign n16666 = n16665 ^ n16439 ;
  assign n16667 = n16666 ^ n16429 ;
  assign n16668 = ~n16431 & n16667 ;
  assign n16669 = n16668 ^ n16429 ;
  assign n16670 = n16669 ^ n16419 ;
  assign n16671 = n16421 & n16670 ;
  assign n16672 = n16671 ^ n16419 ;
  assign n16675 = n16674 ^ n16672 ;
  assign n16679 = n5700 & ~n12262 ;
  assign n16678 = n5702 & ~n12256 ;
  assign n16680 = n16679 ^ n16678 ;
  assign n16681 = n16680 ^ x17 ;
  assign n16677 = n5703 & ~n13283 ;
  assign n16682 = n16681 ^ n16677 ;
  assign n16676 = ~n12220 & n20731 ;
  assign n16683 = n16682 ^ n16676 ;
  assign n16684 = n16683 ^ n16672 ;
  assign n16685 = ~n16675 & n16684 ;
  assign n16673 = n16672 ^ n16370 ;
  assign n16686 = n16685 ^ n16673 ;
  assign n16687 = ~n16408 & ~n16686 ;
  assign n16371 = n16370 ^ n16368 ;
  assign n16688 = n16687 ^ n16371 ;
  assign n16689 = ~n16369 & n16688 ;
  assign n16690 = n16689 ^ n16368 ;
  assign n16692 = n16691 ^ n16690 ;
  assign n16701 = n6650 & n12755 ;
  assign n16694 = n12971 ^ x11 ;
  assign n16695 = n16694 ^ x10 ;
  assign n16696 = n16695 ^ n12971 ;
  assign n16697 = ~n12973 & n16696 ;
  assign n16698 = n16697 ^ n12971 ;
  assign n16699 = n6648 & n16698 ;
  assign n16700 = n16699 ^ x11 ;
  assign n16702 = n16701 ^ n16700 ;
  assign n16693 = n6655 & ~n12705 ;
  assign n16703 = n16702 ^ n16693 ;
  assign n16704 = n16703 ^ n16690 ;
  assign n16705 = ~n16692 & ~n16704 ;
  assign n16706 = n16705 ^ n16703 ;
  assign n20610 = n16706 ^ n16338 ;
  assign n20611 = ~n16339 & n20610 ;
  assign n20612 = n20611 ^ n13900 ;
  assign n18113 = n7128 & ~n12855 ;
  assign n18114 = n18113 ^ x8 ;
  assign n18115 = n18114 ^ x7 ;
  assign n18116 = ~n13007 & n18113 ;
  assign n18117 = ~n18115 & n18116 ;
  assign n18118 = n18117 ^ n18114 ;
  assign n18112 = n7141 & n12971 ;
  assign n18119 = n18118 ^ n18112 ;
  assign n18111 = n7146 & n12755 ;
  assign n18120 = n18119 ^ n18111 ;
  assign n17035 = n4916 & ~n12129 ;
  assign n17032 = n16666 ^ n16431 ;
  assign n17033 = n17032 ^ x20 ;
  assign n17027 = n12121 ^ n4685 ;
  assign n17028 = n17027 ^ n12121 ;
  assign n17029 = ~n13605 & n17028 ;
  assign n17030 = n17029 ^ n12121 ;
  assign n17031 = n4678 & n17030 ;
  assign n17034 = n17033 ^ n17031 ;
  assign n17036 = n17035 ^ n17034 ;
  assign n17025 = n12130 & n14027 ;
  assign n17037 = n17036 ^ n17025 ;
  assign n16717 = n16663 ^ n16441 ;
  assign n16712 = ~n12136 & n14027 ;
  assign n16711 = n4684 & n13737 ;
  assign n16713 = n16712 ^ n16711 ;
  assign n16714 = n16713 ^ x20 ;
  assign n16710 = n4683 & ~n12129 ;
  assign n16715 = n16714 ^ n16710 ;
  assign n16709 = n4916 & n12130 ;
  assign n16716 = n16715 ^ n16709 ;
  assign n16718 = n16717 ^ n16716 ;
  assign n16730 = n16660 ^ n16451 ;
  assign n16727 = n4916 & ~n12136 ;
  assign n16720 = n12130 ^ x20 ;
  assign n16721 = n16720 ^ x19 ;
  assign n16722 = n16721 ^ n12130 ;
  assign n16723 = ~n13817 & n16722 ;
  assign n16724 = n16723 ^ n12130 ;
  assign n16725 = n4678 & n16724 ;
  assign n16726 = n16725 ^ x20 ;
  assign n16728 = n16727 ^ n16726 ;
  assign n16719 = n12137 & n14027 ;
  assign n16729 = n16728 ^ n16719 ;
  assign n16731 = n16730 ^ n16729 ;
  assign n16744 = n16654 ^ n16471 ;
  assign n16741 = n4916 & ~n12138 ;
  assign n16734 = n12137 ^ x20 ;
  assign n16735 = n16734 ^ x19 ;
  assign n16736 = n16735 ^ n12137 ;
  assign n16737 = ~n13936 & n16736 ;
  assign n16738 = n16737 ^ n12137 ;
  assign n16739 = n4678 & n16738 ;
  assign n16740 = n16739 ^ x20 ;
  assign n16742 = n16741 ^ n16740 ;
  assign n16733 = n12207 & n14027 ;
  assign n16743 = n16742 ^ n16733 ;
  assign n16745 = n16744 ^ n16743 ;
  assign n16987 = n16651 ^ n16481 ;
  assign n16980 = ~n12142 & n14027 ;
  assign n16979 = n4916 & n12207 ;
  assign n16981 = n16980 ^ n16979 ;
  assign n16977 = n4683 & ~n14370 ;
  assign n16976 = n4678 & n14832 ;
  assign n16978 = n16977 ^ n16976 ;
  assign n16982 = n16981 ^ n16978 ;
  assign n16988 = n16987 ^ n16982 ;
  assign n16973 = n12143 & n14027 ;
  assign n16972 = n4916 & ~n12142 ;
  assign n16974 = n16973 ^ n16972 ;
  assign n16970 = n4683 & ~n14476 ;
  assign n16969 = n4678 & ~n15500 ;
  assign n16971 = n16970 ^ n16969 ;
  assign n16975 = n16974 ^ n16971 ;
  assign n16983 = n16982 ^ n16975 ;
  assign n16967 = n16648 ^ n16491 ;
  assign n16757 = n16645 ^ n16501 ;
  assign n16754 = n4916 & n12143 ;
  assign n16747 = n12142 ^ x20 ;
  assign n16748 = n16747 ^ x19 ;
  assign n16749 = n16748 ^ n12142 ;
  assign n16750 = ~n14298 & n16749 ;
  assign n16751 = n16750 ^ n12142 ;
  assign n16752 = n4678 & ~n16751 ;
  assign n16753 = n16752 ^ x20 ;
  assign n16755 = n16754 ^ n16753 ;
  assign n16746 = n12149 & n14027 ;
  assign n16756 = n16755 ^ n16746 ;
  assign n16758 = n16757 ^ n16756 ;
  assign n16778 = n16635 ^ n16509 ;
  assign n16773 = n12152 & n14027 ;
  assign n16772 = n4684 & ~n15312 ;
  assign n16774 = n16773 ^ n16772 ;
  assign n16775 = n16774 ^ x20 ;
  assign n16771 = n4683 & n12149 ;
  assign n16776 = n16775 ^ n16771 ;
  assign n16770 = n4916 & ~n12151 ;
  assign n16777 = n16776 ^ n16770 ;
  assign n16779 = n16778 ^ n16777 ;
  assign n16792 = n16630 ^ n16533 ;
  assign n16789 = n12160 & n14027 ;
  assign n16782 = n12151 ^ x20 ;
  assign n16783 = n16782 ^ x19 ;
  assign n16784 = n16783 ^ n12151 ;
  assign n16785 = ~n15299 & n16784 ;
  assign n16786 = n16785 ^ n12151 ;
  assign n16787 = n4678 & ~n16786 ;
  assign n16788 = n16787 ^ x20 ;
  assign n16790 = n16789 ^ n16788 ;
  assign n16780 = n4916 & n12152 ;
  assign n16791 = n16790 ^ n16780 ;
  assign n16793 = n16792 ^ n16791 ;
  assign n16805 = n16628 ^ n16545 ;
  assign n16802 = n4916 & n12160 ;
  assign n16798 = n4685 & ~n14580 ;
  assign n16799 = n16798 ^ n12152 ;
  assign n16800 = n4678 & n16799 ;
  assign n16801 = n16800 ^ x20 ;
  assign n16803 = n16802 ^ n16801 ;
  assign n16794 = n12163 & n14027 ;
  assign n16804 = n16803 ^ n16794 ;
  assign n16806 = n16805 ^ n16804 ;
  assign n16818 = n16624 ^ n16556 ;
  assign n16815 = n4916 & n12163 ;
  assign n16808 = n12160 ^ x20 ;
  assign n16809 = n16808 ^ x19 ;
  assign n16810 = n16809 ^ n12160 ;
  assign n16811 = ~n14866 & n16810 ;
  assign n16812 = n16811 ^ n12160 ;
  assign n16813 = n4678 & n16812 ;
  assign n16814 = n16813 ^ x20 ;
  assign n16816 = n16815 ^ n16814 ;
  assign n16807 = n12167 & n14027 ;
  assign n16817 = n16816 ^ n16807 ;
  assign n16819 = n16818 ^ n16817 ;
  assign n16831 = n16621 ^ n16567 ;
  assign n16828 = n4916 & n12167 ;
  assign n16821 = n12163 ^ x20 ;
  assign n16822 = n16821 ^ x19 ;
  assign n16823 = n16822 ^ n12163 ;
  assign n16824 = ~n14880 & n16823 ;
  assign n16825 = n16824 ^ n12163 ;
  assign n16826 = n4678 & n16825 ;
  assign n16827 = n16826 ^ x20 ;
  assign n16829 = n16828 ^ n16827 ;
  assign n16820 = n12168 & n14027 ;
  assign n16830 = n16829 ^ n16820 ;
  assign n16832 = n16831 ^ n16830 ;
  assign n16844 = n16618 ^ n16610 ;
  assign n16841 = n4916 & n12168 ;
  assign n16834 = n12167 ^ x20 ;
  assign n16835 = n16834 ^ x19 ;
  assign n16836 = n16835 ^ n12167 ;
  assign n16837 = ~n14914 & n16836 ;
  assign n16838 = n16837 ^ n12167 ;
  assign n16839 = n4678 & n16838 ;
  assign n16840 = n16839 ^ x20 ;
  assign n16842 = n16841 ^ n16840 ;
  assign n16833 = ~n12169 & n14027 ;
  assign n16843 = n16842 ^ n16833 ;
  assign n16845 = n16844 ^ n16843 ;
  assign n16857 = n16606 ^ n16575 ;
  assign n16854 = n12175 & n14027 ;
  assign n16847 = n12168 ^ x20 ;
  assign n16848 = n16847 ^ x19 ;
  assign n16849 = n16848 ^ n12168 ;
  assign n16850 = ~n14948 & n16849 ;
  assign n16851 = n16850 ^ n12168 ;
  assign n16852 = n4678 & n16851 ;
  assign n16853 = n16852 ^ x20 ;
  assign n16855 = n16854 ^ n16853 ;
  assign n16846 = n4916 & ~n12169 ;
  assign n16856 = n16855 ^ n16846 ;
  assign n16858 = n16857 ^ n16856 ;
  assign n16870 = n16591 ^ n16576 ;
  assign n16871 = n16870 ^ n16600 ;
  assign n16867 = n4916 & n12175 ;
  assign n16860 = n12169 ^ x20 ;
  assign n16861 = n16860 ^ x19 ;
  assign n16862 = n16861 ^ n12169 ;
  assign n16863 = ~n15032 & n16862 ;
  assign n16864 = n16863 ^ n12169 ;
  assign n16865 = n4678 & ~n16864 ;
  assign n16866 = n16865 ^ x20 ;
  assign n16868 = n16867 ^ n16866 ;
  assign n16859 = n12179 & n14027 ;
  assign n16869 = n16868 ^ n16859 ;
  assign n16872 = n16871 ^ n16869 ;
  assign n16582 = n16581 ^ x23 ;
  assign n16920 = n16590 ^ n16582 ;
  assign n16884 = n4488 & ~n12183 ;
  assign n16885 = n4678 & ~n12182 ;
  assign n16886 = x20 & ~n16885 ;
  assign n16887 = ~n12183 & n16886 ;
  assign n16888 = n7824 & n16887 ;
  assign n16889 = n16888 ^ n16886 ;
  assign n16896 = ~n12183 & n14027 ;
  assign n16895 = n4683 & n12181 ;
  assign n16897 = n16896 ^ n16895 ;
  assign n16893 = n4916 & ~n12182 ;
  assign n16892 = n4684 & n15756 ;
  assign n16894 = n16893 ^ n16892 ;
  assign n16898 = n16897 ^ n16894 ;
  assign n16899 = n16889 & ~n16898 ;
  assign n16900 = ~n16884 & ~n16899 ;
  assign n16909 = n4916 & n12181 ;
  assign n16902 = n12180 ^ x20 ;
  assign n16903 = n16902 ^ x19 ;
  assign n16904 = n16903 ^ n12180 ;
  assign n16905 = ~n12225 & n16904 ;
  assign n16906 = n16905 ^ n12180 ;
  assign n16907 = n4678 & n16906 ;
  assign n16908 = n16907 ^ x20 ;
  assign n16910 = n16909 ^ n16908 ;
  assign n16901 = ~n12182 & n14027 ;
  assign n16911 = n16910 ^ n16901 ;
  assign n16912 = n16900 & n16911 ;
  assign n16913 = n16912 ^ n16911 ;
  assign n16881 = n4916 & n12180 ;
  assign n16874 = n12179 ^ x20 ;
  assign n16875 = n16874 ^ x19 ;
  assign n16876 = n16875 ^ n12179 ;
  assign n16877 = ~n15127 & n16876 ;
  assign n16878 = n16877 ^ n12179 ;
  assign n16879 = n4678 & n16878 ;
  assign n16880 = n16879 ^ x20 ;
  assign n16882 = n16881 ^ n16880 ;
  assign n16873 = n12181 & n14027 ;
  assign n16883 = n16882 ^ n16873 ;
  assign n16914 = n16913 ^ n16883 ;
  assign n16916 = ~n7810 & ~n12183 ;
  assign n16915 = n16913 ^ n16577 ;
  assign n16917 = n16916 ^ n16915 ;
  assign n16918 = n16914 & n16917 ;
  assign n16919 = n16918 ^ n16913 ;
  assign n16921 = n16920 ^ n16919 ;
  assign n16926 = n4916 & n12179 ;
  assign n16925 = n4683 & n12175 ;
  assign n16927 = n16926 ^ n16925 ;
  assign n16923 = n12180 & n14027 ;
  assign n16922 = n4684 & ~n15049 ;
  assign n16924 = n16923 ^ n16922 ;
  assign n16928 = n16927 ^ n16924 ;
  assign n16929 = n16928 ^ x20 ;
  assign n16930 = n16929 ^ n16919 ;
  assign n16931 = n16921 & ~n16930 ;
  assign n16932 = n16931 ^ n16920 ;
  assign n16933 = n16932 ^ n16869 ;
  assign n16934 = n16872 & n16933 ;
  assign n16935 = n16934 ^ n16869 ;
  assign n16936 = n16935 ^ n16856 ;
  assign n16937 = n16858 & n16936 ;
  assign n16938 = n16937 ^ n16856 ;
  assign n16939 = n16938 ^ n16843 ;
  assign n16940 = n16845 & n16939 ;
  assign n16941 = n16940 ^ n16843 ;
  assign n16942 = n16941 ^ n16830 ;
  assign n16943 = n16832 & n16942 ;
  assign n16944 = n16943 ^ n16830 ;
  assign n16945 = n16944 ^ n16817 ;
  assign n16946 = n16819 & n16945 ;
  assign n16947 = n16946 ^ n16817 ;
  assign n16948 = n16947 ^ n16804 ;
  assign n16949 = n16806 & n16948 ;
  assign n16950 = n16949 ^ n16804 ;
  assign n16951 = n16950 ^ n16791 ;
  assign n16952 = n16793 & n16951 ;
  assign n16953 = n16952 ^ n16791 ;
  assign n16954 = n16953 ^ n16777 ;
  assign n16955 = n16779 & n16954 ;
  assign n16956 = n16955 ^ n16777 ;
  assign n16767 = n4916 & n12149 ;
  assign n16760 = n12143 ^ x20 ;
  assign n16761 = n16760 ^ x19 ;
  assign n16762 = n16761 ^ n12143 ;
  assign n16763 = ~n15280 & n16762 ;
  assign n16764 = n16763 ^ n12143 ;
  assign n16765 = n4678 & n16764 ;
  assign n16766 = n16765 ^ x20 ;
  assign n16768 = n16767 ^ n16766 ;
  assign n16759 = ~n12151 & n14027 ;
  assign n16769 = n16768 ^ n16759 ;
  assign n16957 = n16956 ^ n16769 ;
  assign n16959 = n16634 ^ n16509 ;
  assign n16960 = ~n16635 & n16959 ;
  assign n16958 = n16769 ^ n16519 ;
  assign n16961 = n16960 ^ n16958 ;
  assign n16962 = n16957 & ~n16961 ;
  assign n16963 = n16962 ^ n16956 ;
  assign n16964 = n16963 ^ n16756 ;
  assign n16965 = ~n16758 & n16964 ;
  assign n16966 = n16965 ^ n16756 ;
  assign n16968 = n16967 ^ n16966 ;
  assign n16984 = n16983 ^ n16968 ;
  assign n16985 = n16984 ^ n16983 ;
  assign n16995 = n16982 ^ n16967 ;
  assign n16996 = n16995 ^ n16983 ;
  assign n16997 = n16985 & ~n16996 ;
  assign n16998 = n16997 ^ n16983 ;
  assign n16999 = ~n16988 & n16998 ;
  assign n17000 = n16999 ^ n16982 ;
  assign n16989 = n16988 ^ n16975 ;
  assign n16986 = n16983 ^ n16966 ;
  assign n16990 = n16989 ^ n16986 ;
  assign n16991 = n16990 ^ n16983 ;
  assign n16992 = n16985 & n16991 ;
  assign n16993 = n16992 ^ n16983 ;
  assign n16994 = x20 & ~n16993 ;
  assign n17001 = n17000 ^ n16994 ;
  assign n17002 = n17001 ^ n16743 ;
  assign n17003 = ~n16745 & n17002 ;
  assign n17004 = n17003 ^ n16743 ;
  assign n16732 = n16657 ^ n16461 ;
  assign n17005 = n17004 ^ n16732 ;
  assign n17014 = n4916 & n12137 ;
  assign n17012 = n16732 ^ x20 ;
  assign n17007 = n12136 ^ n4685 ;
  assign n17008 = n17007 ^ n12136 ;
  assign n17009 = ~n14753 & n17008 ;
  assign n17010 = n17009 ^ n12136 ;
  assign n17011 = n4678 & ~n17010 ;
  assign n17013 = n17012 ^ n17011 ;
  assign n17015 = n17014 ^ n17013 ;
  assign n17006 = ~n12138 & n14027 ;
  assign n17016 = n17015 ^ n17006 ;
  assign n17017 = n17005 & ~n17016 ;
  assign n17018 = n17017 ^ n17004 ;
  assign n17019 = n17018 ^ n16729 ;
  assign n17020 = n16731 & n17019 ;
  assign n17021 = n17020 ^ n16729 ;
  assign n17022 = n17021 ^ n16716 ;
  assign n17023 = ~n16718 & n17022 ;
  assign n17024 = n17023 ^ n16716 ;
  assign n17384 = n17032 ^ n17024 ;
  assign n17385 = ~n17037 & ~n17384 ;
  assign n17386 = n17385 ^ n17032 ;
  assign n17382 = n16669 ^ n16421 ;
  assign n17380 = ~n12110 & n20731 ;
  assign n17378 = n5703 & n13712 ;
  assign n17375 = n5700 & ~n12220 ;
  assign n17374 = n5702 & ~n12262 ;
  assign n17376 = n17375 ^ n17374 ;
  assign n17377 = n17376 ^ x17 ;
  assign n17379 = n17378 ^ n17377 ;
  assign n17381 = n17380 ^ n17379 ;
  assign n17383 = n17382 ^ n17381 ;
  assign n17387 = n17386 ^ n17383 ;
  assign n17044 = n5703 & n14047 ;
  assign n17042 = n5700 & ~n12110 ;
  assign n17040 = n5702 & ~n12220 ;
  assign n17038 = n17037 ^ n17024 ;
  assign n17039 = n17038 ^ x17 ;
  assign n17041 = n17040 ^ n17039 ;
  assign n17043 = n17042 ^ n17041 ;
  assign n17045 = n17044 ^ n17043 ;
  assign n16708 = n12117 & n20731 ;
  assign n17046 = n17045 ^ n16708 ;
  assign n17054 = n5703 & n13196 ;
  assign n17052 = n5700 & n12117 ;
  assign n17050 = n5702 & ~n12110 ;
  assign n17048 = n17021 ^ n16718 ;
  assign n17049 = n17048 ^ x17 ;
  assign n17051 = n17050 ^ n17049 ;
  assign n17053 = n17052 ^ n17051 ;
  assign n17055 = n17054 ^ n17053 ;
  assign n17047 = n12121 & n20731 ;
  assign n17056 = n17055 ^ n17047 ;
  assign n17355 = n17018 ^ n16731 ;
  assign n17070 = n17016 ^ n17004 ;
  assign n17058 = n12130 & n20731 ;
  assign n17057 = n5700 & ~n12129 ;
  assign n17059 = n17058 ^ n17057 ;
  assign n17060 = n17059 ^ n5694 ;
  assign n17062 = n17059 ^ x17 ;
  assign n17065 = n17062 ^ n5696 ;
  assign n17066 = ~x16 & ~n13605 ;
  assign n17067 = n17065 & n17066 ;
  assign n17063 = ~n12121 & n17062 ;
  assign n17061 = n5696 & ~n13606 ;
  assign n17064 = n17063 ^ n17061 ;
  assign n17068 = n17067 ^ n17064 ;
  assign n17069 = ~n17060 & ~n17068 ;
  assign n17071 = n17070 ^ n17069 ;
  assign n17080 = n17001 ^ n16745 ;
  assign n17078 = ~n12136 & n20731 ;
  assign n17076 = n5703 & n13737 ;
  assign n17073 = n5700 & n12130 ;
  assign n17072 = n5702 & ~n12129 ;
  assign n17074 = n17073 ^ n17072 ;
  assign n17075 = n17074 ^ x17 ;
  assign n17077 = n17076 ^ n17075 ;
  assign n17079 = n17078 ^ n17077 ;
  assign n17081 = n17080 ^ n17079 ;
  assign n17091 = n12137 & n20731 ;
  assign n17089 = n5703 & ~n13818 ;
  assign n17086 = n5700 & ~n12136 ;
  assign n17085 = n5702 & n12130 ;
  assign n17087 = n17086 ^ n17085 ;
  assign n17088 = n17087 ^ x17 ;
  assign n17090 = n17089 ^ n17088 ;
  assign n17092 = n17091 ^ n17090 ;
  assign n17093 = n17092 ^ n16989 ;
  assign n17082 = n16975 ^ n16966 ;
  assign n17083 = n17082 ^ x20 ;
  assign n17084 = n16968 & n17083 ;
  assign n17094 = n17093 ^ n17084 ;
  assign n17103 = n16967 ^ x20 ;
  assign n17104 = n17103 ^ n16975 ;
  assign n17105 = n17104 ^ n16966 ;
  assign n17098 = n5700 & n12137 ;
  assign n17097 = n5702 & ~n12136 ;
  assign n17099 = n17098 ^ n17097 ;
  assign n17100 = n17099 ^ x17 ;
  assign n17096 = n5703 & n14129 ;
  assign n17101 = n17100 ^ n17096 ;
  assign n17095 = ~n12138 & n20731 ;
  assign n17102 = n17101 ^ n17095 ;
  assign n17106 = n17105 ^ n17102 ;
  assign n17115 = n16963 ^ n16758 ;
  assign n17113 = n12207 & n20731 ;
  assign n17111 = n5703 & ~n13939 ;
  assign n17108 = n5700 & ~n12138 ;
  assign n17107 = n5702 & n12137 ;
  assign n17109 = n17108 ^ n17107 ;
  assign n17110 = n17109 ^ x17 ;
  assign n17112 = n17111 ^ n17110 ;
  assign n17114 = n17113 ^ n17112 ;
  assign n17116 = n17115 ^ n17114 ;
  assign n17125 = n16961 ^ n16956 ;
  assign n17123 = ~n12142 & n20731 ;
  assign n17121 = n5703 & n14832 ;
  assign n17118 = n5700 & n12207 ;
  assign n17117 = n5702 & ~n12138 ;
  assign n17119 = n17118 ^ n17117 ;
  assign n17120 = n17119 ^ x17 ;
  assign n17122 = n17121 ^ n17120 ;
  assign n17124 = n17123 ^ n17122 ;
  assign n17126 = n17125 ^ n17124 ;
  assign n17135 = n16953 ^ n16779 ;
  assign n17130 = n5700 & ~n12142 ;
  assign n17129 = n5702 & n12207 ;
  assign n17131 = n17130 ^ n17129 ;
  assign n17132 = n17131 ^ x17 ;
  assign n17128 = n5703 & ~n15500 ;
  assign n17133 = n17132 ^ n17128 ;
  assign n17127 = n12143 & n20731 ;
  assign n17134 = n17133 ^ n17127 ;
  assign n17136 = n17135 ^ n17134 ;
  assign n17145 = n16950 ^ n16793 ;
  assign n17140 = n5700 & n12143 ;
  assign n17139 = n5702 & ~n12142 ;
  assign n17141 = n17140 ^ n17139 ;
  assign n17142 = n17141 ^ x17 ;
  assign n17138 = n5703 & n14299 ;
  assign n17143 = n17142 ^ n17138 ;
  assign n17137 = n12149 & n20731 ;
  assign n17144 = n17143 ^ n17137 ;
  assign n17146 = n17145 ^ n17144 ;
  assign n17155 = n16947 ^ n16806 ;
  assign n17150 = n5700 & n12149 ;
  assign n17149 = n5702 & n12143 ;
  assign n17151 = n17150 ^ n17149 ;
  assign n17152 = n17151 ^ x17 ;
  assign n17148 = n5703 & ~n14498 ;
  assign n17153 = n17152 ^ n17148 ;
  assign n17147 = ~n12151 & n20731 ;
  assign n17154 = n17153 ^ n17147 ;
  assign n17156 = n17155 ^ n17154 ;
  assign n17169 = n16944 ^ n16819 ;
  assign n17161 = ~x16 & ~n15311 ;
  assign n17166 = n17161 ^ n15312 ;
  assign n17167 = n5696 & ~n17166 ;
  assign n17162 = n17161 ^ n12149 ;
  assign n17164 = n17162 & n17163 ;
  assign n17158 = n12152 & n20731 ;
  assign n17157 = n5700 & ~n12151 ;
  assign n17159 = n17158 ^ n17157 ;
  assign n17160 = n17159 ^ x17 ;
  assign n17165 = n17164 ^ n17160 ;
  assign n17168 = n17167 ^ n17165 ;
  assign n17170 = n17169 ^ n17168 ;
  assign n17307 = n16941 ^ n16832 ;
  assign n17179 = n16938 ^ n16845 ;
  assign n17177 = n12163 & n20731 ;
  assign n17175 = n5703 & ~n14581 ;
  assign n17172 = n5702 & n12152 ;
  assign n17171 = n5700 & n12160 ;
  assign n17173 = n17172 ^ n17171 ;
  assign n17174 = n17173 ^ x17 ;
  assign n17176 = n17175 ^ n17174 ;
  assign n17178 = n17177 ^ n17176 ;
  assign n17180 = n17179 ^ n17178 ;
  assign n17189 = n16935 ^ n16858 ;
  assign n17184 = n5700 & n12163 ;
  assign n17183 = n5702 & n12160 ;
  assign n17185 = n17184 ^ n17183 ;
  assign n17186 = n17185 ^ x17 ;
  assign n17182 = n5703 & ~n14867 ;
  assign n17187 = n17186 ^ n17182 ;
  assign n17181 = n12167 & n20731 ;
  assign n17188 = n17187 ^ n17181 ;
  assign n17190 = n17189 ^ n17188 ;
  assign n17199 = n16932 ^ n16872 ;
  assign n17197 = n12168 & n20731 ;
  assign n17195 = n5703 & ~n14890 ;
  assign n17192 = n5700 & n12167 ;
  assign n17191 = n5702 & n12163 ;
  assign n17193 = n17192 ^ n17191 ;
  assign n17194 = n17193 ^ x17 ;
  assign n17196 = n17195 ^ n17194 ;
  assign n17198 = n17197 ^ n17196 ;
  assign n17200 = n17199 ^ n17198 ;
  assign n17212 = n16920 ^ x20 ;
  assign n17213 = n17212 ^ n16928 ;
  assign n17214 = n17213 ^ n16919 ;
  assign n17209 = n5700 & n12168 ;
  assign n17202 = n12167 ^ x17 ;
  assign n17203 = n17202 ^ x16 ;
  assign n17204 = n17203 ^ n12167 ;
  assign n17205 = ~n14914 & n17204 ;
  assign n17206 = n17205 ^ n12167 ;
  assign n17207 = n5693 & n17206 ;
  assign n17208 = n17207 ^ x17 ;
  assign n17210 = n17209 ^ n17208 ;
  assign n17201 = ~n12169 & n20731 ;
  assign n17211 = n17210 ^ n17201 ;
  assign n17215 = n17214 ^ n17211 ;
  assign n17224 = n16917 ^ n16883 ;
  assign n17222 = n12175 & n20731 ;
  assign n17220 = n5703 & ~n14949 ;
  assign n17217 = n5700 & ~n12169 ;
  assign n17216 = n5702 & n12168 ;
  assign n17218 = n17217 ^ n17216 ;
  assign n17219 = n17218 ^ x17 ;
  assign n17221 = n17220 ^ n17219 ;
  assign n17223 = n17222 ^ n17221 ;
  assign n17225 = n17224 ^ n17223 ;
  assign n17234 = n16899 ^ n16884 ;
  assign n17235 = n17234 ^ n16911 ;
  assign n17232 = n12179 & n20731 ;
  assign n17230 = n5703 & n15035 ;
  assign n17227 = n5702 & ~n12169 ;
  assign n17226 = n5700 & n12175 ;
  assign n17228 = n17227 ^ n17226 ;
  assign n17229 = n17228 ^ x17 ;
  assign n17231 = n17230 ^ n17229 ;
  assign n17233 = n17232 ^ n17231 ;
  assign n17236 = n17235 ^ n17233 ;
  assign n16890 = n16889 ^ x20 ;
  assign n17276 = n16898 ^ n16890 ;
  assign n17263 = n8156 & ~n12183 ;
  assign n17241 = n5700 & n12181 ;
  assign n17240 = n5702 & n12180 ;
  assign n17242 = n17241 ^ n17240 ;
  assign n17238 = ~n12182 & n20731 ;
  assign n17237 = n5703 & ~n15151 ;
  assign n17239 = n17238 ^ n17237 ;
  assign n17243 = n17242 ^ n17239 ;
  assign n17245 = n4675 & ~n12183 ;
  assign n17244 = n4678 & ~n12183 ;
  assign n17246 = n17245 ^ n17244 ;
  assign n17247 = n5705 & ~n12184 ;
  assign n17251 = n5702 & n12181 ;
  assign n17249 = ~n12183 & n20731 ;
  assign n17248 = n5703 & n15756 ;
  assign n17250 = n17249 ^ n17248 ;
  assign n17252 = n17251 ^ n17250 ;
  assign n17253 = x17 & ~n17252 ;
  assign n17254 = n17247 & n17253 ;
  assign n17255 = n17254 ^ n17253 ;
  assign n17258 = ~n17246 & ~n17255 ;
  assign n17259 = n17258 ^ n17245 ;
  assign n17260 = ~n17243 & ~n17259 ;
  assign n17261 = n17260 ^ n17245 ;
  assign n17262 = n17261 ^ n16885 ;
  assign n17264 = n17263 ^ n17262 ;
  assign n17271 = n12181 & n20731 ;
  assign n17269 = n5703 & ~n15128 ;
  assign n17266 = n5700 & n12180 ;
  assign n17265 = n5702 & n12179 ;
  assign n17267 = n17266 ^ n17265 ;
  assign n17268 = n17267 ^ x17 ;
  assign n17270 = n17269 ^ n17268 ;
  assign n17272 = n17271 ^ n17270 ;
  assign n17273 = n17272 ^ n17261 ;
  assign n17274 = n17264 & n17273 ;
  assign n17275 = n17274 ^ n17261 ;
  assign n17277 = n17276 ^ n17275 ;
  assign n17285 = n12180 & n20731 ;
  assign n17281 = n17276 ^ x17 ;
  assign n17280 = n5700 & n12179 ;
  assign n17282 = n17281 ^ n17280 ;
  assign n17279 = n5702 & n12175 ;
  assign n17283 = n17282 ^ n17279 ;
  assign n17278 = n5703 & ~n15049 ;
  assign n17284 = n17283 ^ n17278 ;
  assign n17286 = n17285 ^ n17284 ;
  assign n17287 = n17277 & n17286 ;
  assign n17288 = n17287 ^ n17276 ;
  assign n17289 = n17288 ^ n17233 ;
  assign n17290 = n17236 & n17289 ;
  assign n17291 = n17290 ^ n17233 ;
  assign n17292 = n17291 ^ n17223 ;
  assign n17293 = n17225 & n17292 ;
  assign n17294 = n17293 ^ n17223 ;
  assign n17295 = n17294 ^ n17211 ;
  assign n17296 = n17215 & n17295 ;
  assign n17297 = n17296 ^ n17211 ;
  assign n17298 = n17297 ^ n17198 ;
  assign n17299 = n17200 & n17298 ;
  assign n17300 = n17299 ^ n17198 ;
  assign n17301 = n17300 ^ n17188 ;
  assign n17302 = n17190 & n17301 ;
  assign n17303 = n17302 ^ n17188 ;
  assign n17304 = n17303 ^ n17178 ;
  assign n17305 = n17180 & n17304 ;
  assign n17306 = n17305 ^ n17178 ;
  assign n17308 = n17307 ^ n17306 ;
  assign n17318 = n5700 & n12152 ;
  assign n17317 = n12160 & n20731 ;
  assign n17319 = n17318 ^ n17317 ;
  assign n17320 = n17319 ^ x17 ;
  assign n17309 = n12151 ^ x17 ;
  assign n17310 = n17309 ^ x16 ;
  assign n17311 = n17310 ^ n12151 ;
  assign n17313 = n15300 ^ n12151 ;
  assign n17314 = n17311 & ~n17313 ;
  assign n17315 = n17314 ^ n12151 ;
  assign n17316 = n5693 & ~n17315 ;
  assign n17321 = n17320 ^ n17316 ;
  assign n17322 = n17321 ^ n17306 ;
  assign n17323 = n17308 & ~n17322 ;
  assign n17324 = n17323 ^ n17307 ;
  assign n17325 = n17324 ^ n17168 ;
  assign n17326 = n17170 & ~n17325 ;
  assign n17327 = n17326 ^ n17169 ;
  assign n17328 = n17327 ^ n17154 ;
  assign n17329 = n17156 & n17328 ;
  assign n17330 = n17329 ^ n17154 ;
  assign n17331 = n17330 ^ n17144 ;
  assign n17332 = n17146 & n17331 ;
  assign n17333 = n17332 ^ n17144 ;
  assign n17334 = n17333 ^ n17134 ;
  assign n17335 = n17136 & n17334 ;
  assign n17336 = n17335 ^ n17134 ;
  assign n17337 = n17336 ^ n17124 ;
  assign n17338 = n17126 & n17337 ;
  assign n17339 = n17338 ^ n17124 ;
  assign n17340 = n17339 ^ n17114 ;
  assign n17341 = ~n17116 & n17340 ;
  assign n17342 = n17341 ^ n17114 ;
  assign n17343 = n17342 ^ n17102 ;
  assign n17344 = ~n17106 & n17343 ;
  assign n17345 = n17344 ^ n17102 ;
  assign n17346 = n17345 ^ n17092 ;
  assign n17347 = ~n17094 & n17346 ;
  assign n17348 = n17347 ^ n17092 ;
  assign n17349 = n17348 ^ n17079 ;
  assign n17350 = ~n17081 & n17349 ;
  assign n17351 = n17350 ^ n17079 ;
  assign n17352 = n17351 ^ n17069 ;
  assign n17353 = ~n17071 & ~n17352 ;
  assign n17354 = n17353 ^ n17069 ;
  assign n17356 = n17355 ^ n17354 ;
  assign n17363 = n5703 & ~n13596 ;
  assign n17361 = n5700 & n12121 ;
  assign n17359 = n5702 & n12117 ;
  assign n17358 = n17355 ^ x17 ;
  assign n17360 = n17359 ^ n17358 ;
  assign n17362 = n17361 ^ n17360 ;
  assign n17364 = n17363 ^ n17362 ;
  assign n17357 = ~n12129 & n20731 ;
  assign n17365 = n17364 ^ n17357 ;
  assign n17366 = ~n17356 & n17365 ;
  assign n17367 = n17366 ^ n17355 ;
  assign n17368 = n17367 ^ n17048 ;
  assign n17369 = ~n17056 & ~n17368 ;
  assign n17370 = n17369 ^ n17048 ;
  assign n17371 = n17370 ^ n17038 ;
  assign n17372 = ~n17046 & n17371 ;
  assign n17373 = n17372 ^ n17038 ;
  assign n17388 = n17387 ^ n17373 ;
  assign n17413 = ~n6072 & ~n12256 ;
  assign n17412 = ~n6074 & n12260 ;
  assign n17414 = n17413 ^ n17412 ;
  assign n17415 = n17414 ^ x14 ;
  assign n17407 = ~x13 & ~n12270 ;
  assign n17408 = n17407 ^ n11972 ;
  assign n17411 = n6060 & n17408 ;
  assign n17416 = n17415 ^ n17411 ;
  assign n17409 = n17408 ^ n12270 ;
  assign n17410 = n6063 & ~n17409 ;
  assign n17417 = n17416 ^ n17410 ;
  assign n17401 = ~n6072 & n12260 ;
  assign n17395 = n16360 ^ x13 ;
  assign n17396 = n17395 ^ n12108 ;
  assign n17397 = ~n13300 & n17396 ;
  assign n17398 = n17397 ^ n12108 ;
  assign n17399 = n4897 & ~n17398 ;
  assign n17400 = n17399 ^ x14 ;
  assign n17402 = n17401 ^ n17400 ;
  assign n17394 = ~n6074 & n11972 ;
  assign n17403 = n17402 ^ n17394 ;
  assign n17392 = n16683 ^ n16675 ;
  assign n17389 = n17386 ^ n17381 ;
  assign n17390 = ~n17383 & ~n17389 ;
  assign n17391 = n17390 ^ n17386 ;
  assign n17393 = n17392 ^ n17391 ;
  assign n17404 = n17403 ^ n17393 ;
  assign n17405 = n17404 ^ n17373 ;
  assign n17406 = n17405 ^ n17404 ;
  assign n17418 = n17417 ^ n17406 ;
  assign n17419 = n17388 & ~n17418 ;
  assign n17420 = n17419 ^ n17405 ;
  assign n18100 = n6655 & ~n12613 ;
  assign n18099 = n6658 & ~n12705 ;
  assign n18101 = n18100 ^ n18099 ;
  assign n18102 = n18101 ^ x11 ;
  assign n18098 = n12706 & n15413 ;
  assign n18103 = n18102 ^ n18098 ;
  assign n18097 = n6650 & n12656 ;
  assign n18104 = n18103 ^ n18097 ;
  assign n18091 = n16686 ^ n16407 ;
  assign n18092 = n18091 ^ n17403 ;
  assign n18093 = n18092 ^ n18091 ;
  assign n18094 = n18093 ^ n17391 ;
  assign n18095 = ~n17393 & ~n18094 ;
  assign n18096 = n18095 ^ n18092 ;
  assign n18105 = n18104 ^ n18096 ;
  assign n18107 = n18105 ^ n17404 ;
  assign n17427 = n6650 & ~n12613 ;
  assign n17425 = ~n12872 & n15413 ;
  assign n17422 = n6655 & ~n12367 ;
  assign n17421 = n6658 & n12656 ;
  assign n17423 = n17422 ^ n17421 ;
  assign n17424 = n17423 ^ x11 ;
  assign n17426 = n17425 ^ n17424 ;
  assign n17428 = n17427 ^ n17426 ;
  assign n18106 = n18105 ^ n17428 ;
  assign n18108 = n18107 ^ n18106 ;
  assign n18109 = ~n17420 & n18108 ;
  assign n18110 = n18109 ^ n18107 ;
  assign n18121 = n18120 ^ n18110 ;
  assign n17441 = n17417 ^ n17388 ;
  assign n17438 = n6650 & ~n12367 ;
  assign n17431 = n12613 ^ x11 ;
  assign n17432 = n17431 ^ x10 ;
  assign n17433 = n17432 ^ n12613 ;
  assign n17434 = ~n13111 & n17433 ;
  assign n17435 = n17434 ^ n12613 ;
  assign n17436 = n6648 & ~n17435 ;
  assign n17437 = n17436 ^ x11 ;
  assign n17439 = n17438 ^ n17437 ;
  assign n17430 = n6655 & ~n12108 ;
  assign n17440 = n17439 ^ n17430 ;
  assign n17442 = n17441 ^ n17440 ;
  assign n17445 = ~n6072 & ~n12262 ;
  assign n17444 = ~n6074 & ~n12256 ;
  assign n17446 = n17445 ^ n17444 ;
  assign n17447 = n17446 ^ n6060 ;
  assign n17448 = n17447 ^ x14 ;
  assign n17457 = n6063 & ~n13053 ;
  assign n17449 = n17446 ^ n6062 ;
  assign n17452 = n12260 ^ x13 ;
  assign n17453 = n17452 ^ n12260 ;
  assign n17454 = n13053 & ~n17453 ;
  assign n17455 = n17454 ^ n12260 ;
  assign n17456 = n17449 & ~n17455 ;
  assign n17458 = n17457 ^ n17456 ;
  assign n17459 = ~n17448 & ~n17458 ;
  assign n17443 = n17370 ^ n17046 ;
  assign n17460 = n17459 ^ n17443 ;
  assign n17480 = n17367 ^ n17056 ;
  assign n17462 = ~n6072 & ~n12220 ;
  assign n17461 = ~n6074 & ~n12262 ;
  assign n17463 = n17462 ^ n17461 ;
  assign n17464 = n17463 ^ n6060 ;
  assign n17465 = n17464 ^ x14 ;
  assign n17475 = n8465 & ~n12256 ;
  assign n17474 = x13 & n13283 ;
  assign n17476 = n17475 ^ n17474 ;
  assign n17477 = ~n6063 & n17476 ;
  assign n17472 = n13052 ^ n8465 ;
  assign n17466 = n17463 ^ x14 ;
  assign n17467 = n12256 ^ x13 ;
  assign n17468 = n17467 ^ n12256 ;
  assign n17469 = n13052 & ~n17468 ;
  assign n17470 = n17469 ^ n12256 ;
  assign n17471 = ~n17466 & n17470 ;
  assign n17473 = n17472 ^ n17471 ;
  assign n17478 = n17477 ^ n17473 ;
  assign n17479 = ~n17465 & ~n17478 ;
  assign n17481 = n17480 ^ n17479 ;
  assign n17501 = n17365 ^ n17354 ;
  assign n17483 = ~n6072 & ~n12110 ;
  assign n17482 = ~n6074 & ~n12220 ;
  assign n17484 = n17483 ^ n17482 ;
  assign n17486 = n12262 ^ x13 ;
  assign n17485 = n12262 ^ n6063 ;
  assign n17487 = n17486 ^ n17485 ;
  assign n17488 = n17485 ^ n12250 ;
  assign n17489 = n17488 ^ n17485 ;
  assign n17490 = ~n17487 & ~n17489 ;
  assign n17491 = n17490 ^ n17485 ;
  assign n17492 = ~n17484 & n17491 ;
  assign n17495 = n17492 ^ x14 ;
  assign n17496 = n4897 & n17495 ;
  assign n17493 = n17484 ^ x14 ;
  assign n17500 = n17496 ^ n17493 ;
  assign n17502 = n17501 ^ n17500 ;
  assign n17513 = n17351 ^ n17071 ;
  assign n17509 = ~n6072 & n12117 ;
  assign n17508 = ~n6074 & ~n12110 ;
  assign n17510 = n17509 ^ n17508 ;
  assign n17511 = n17510 ^ x14 ;
  assign n17503 = n14047 ^ n4899 ;
  assign n17504 = n17503 ^ n14047 ;
  assign n17505 = ~n13172 & ~n17504 ;
  assign n17506 = n17505 ^ n14047 ;
  assign n17507 = n4897 & n17506 ;
  assign n17512 = n17511 ^ n17507 ;
  assign n17514 = n17513 ^ n17512 ;
  assign n17531 = n17348 ^ n17081 ;
  assign n17516 = ~n6072 & n12121 ;
  assign n17515 = ~n6074 & n12117 ;
  assign n17517 = n17516 ^ n17515 ;
  assign n17518 = n17517 ^ n6060 ;
  assign n17519 = n17518 ^ x14 ;
  assign n17528 = n6063 & n13195 ;
  assign n17520 = n17517 ^ n6062 ;
  assign n17522 = n13196 ^ n12110 ;
  assign n17523 = n12110 ^ x13 ;
  assign n17524 = n17523 ^ n12110 ;
  assign n17525 = ~n17522 & ~n17524 ;
  assign n17526 = n17525 ^ n12110 ;
  assign n17527 = n17520 & n17526 ;
  assign n17529 = n17528 ^ n17527 ;
  assign n17530 = ~n17519 & ~n17529 ;
  assign n17532 = n17531 ^ n17530 ;
  assign n17559 = n17345 ^ n17094 ;
  assign n17534 = ~n6072 & ~n12129 ;
  assign n17533 = ~n6074 & n12121 ;
  assign n17535 = n17534 ^ n17533 ;
  assign n17536 = n17535 ^ n6060 ;
  assign n17537 = n17536 ^ x14 ;
  assign n17555 = n12117 ^ n6063 ;
  assign n17541 = n17535 ^ n6062 ;
  assign n17554 = ~n13586 & ~n17542 ;
  assign n17548 = n17554 ^ n12117 ;
  assign n17549 = ~n17541 & ~n17548 ;
  assign n17556 = n17555 ^ n17549 ;
  assign n17557 = n17556 ^ n17554 ;
  assign n17558 = ~n17537 & n17557 ;
  assign n17560 = n17559 ^ n17558 ;
  assign n17563 = ~n6072 & n12130 ;
  assign n17562 = ~n6074 & ~n12129 ;
  assign n17564 = n17563 ^ n17562 ;
  assign n17565 = n17564 ^ n6060 ;
  assign n17566 = n17565 ^ x14 ;
  assign n17568 = n17564 ^ n6062 ;
  assign n17575 = ~n12121 & n17568 ;
  assign n17571 = ~x13 & n17568 ;
  assign n17572 = n17571 ^ n6063 ;
  assign n17573 = ~n13605 & n17572 ;
  assign n17574 = n17573 ^ n6063 ;
  assign n17576 = n17575 ^ n17574 ;
  assign n17577 = ~n17566 & ~n17576 ;
  assign n17561 = n17342 ^ n17106 ;
  assign n17578 = n17577 ^ n17561 ;
  assign n17598 = n17339 ^ n17116 ;
  assign n17580 = ~n6072 & ~n12136 ;
  assign n17579 = ~n6074 & n12130 ;
  assign n17581 = n17580 ^ n17579 ;
  assign n17582 = n17581 ^ n6060 ;
  assign n17583 = n17582 ^ x14 ;
  assign n17593 = n8465 & ~n12129 ;
  assign n17592 = x13 & ~n13737 ;
  assign n17594 = n17593 ^ n17592 ;
  assign n17595 = ~n6063 & n17594 ;
  assign n17590 = n13736 ^ n8465 ;
  assign n17584 = n17581 ^ x14 ;
  assign n17585 = n12129 ^ x13 ;
  assign n17586 = n17585 ^ n12129 ;
  assign n17587 = ~n14271 & ~n17586 ;
  assign n17588 = n17587 ^ n12129 ;
  assign n17589 = ~n17584 & n17588 ;
  assign n17591 = n17590 ^ n17589 ;
  assign n17596 = n17595 ^ n17591 ;
  assign n17597 = ~n17583 & n17596 ;
  assign n17599 = n17598 ^ n17597 ;
  assign n17616 = n17336 ^ n17126 ;
  assign n17601 = ~n6072 & n12137 ;
  assign n17600 = ~n6074 & ~n12136 ;
  assign n17602 = n17601 ^ n17600 ;
  assign n17603 = n17602 ^ n6060 ;
  assign n17604 = n17603 ^ x14 ;
  assign n17613 = n6063 & n13817 ;
  assign n17605 = n17602 ^ n6062 ;
  assign n17608 = n12130 ^ x13 ;
  assign n17609 = n17608 ^ n12130 ;
  assign n17610 = ~n13817 & ~n17609 ;
  assign n17611 = n17610 ^ n12130 ;
  assign n17612 = n17605 & ~n17611 ;
  assign n17614 = n17613 ^ n17612 ;
  assign n17615 = ~n17604 & ~n17614 ;
  assign n17617 = n17616 ^ n17615 ;
  assign n17641 = n17333 ^ n17136 ;
  assign n17619 = ~n6072 & ~n12138 ;
  assign n17618 = ~n6074 & n12137 ;
  assign n17620 = n17619 ^ n17618 ;
  assign n17621 = n17620 ^ n6060 ;
  assign n17622 = n17621 ^ x14 ;
  assign n17637 = n12136 ^ n6063 ;
  assign n17626 = n17620 ^ n6062 ;
  assign n17629 = ~n14753 & ~n17542 ;
  assign n17630 = n17629 ^ n12136 ;
  assign n17631 = ~n17626 & n17630 ;
  assign n17638 = n17637 ^ n17631 ;
  assign n17636 = ~n14128 & ~n17542 ;
  assign n17639 = n17638 ^ n17636 ;
  assign n17640 = ~n17622 & ~n17639 ;
  assign n17642 = n17641 ^ n17640 ;
  assign n17662 = n17330 ^ n17146 ;
  assign n17644 = ~n6072 & n12207 ;
  assign n17643 = ~n6074 & ~n12138 ;
  assign n17645 = n17644 ^ n17643 ;
  assign n17646 = n17645 ^ n6060 ;
  assign n17647 = n17646 ^ x14 ;
  assign n17657 = n8465 & n12137 ;
  assign n17656 = x13 & n13939 ;
  assign n17658 = n17657 ^ n17656 ;
  assign n17659 = ~n6063 & n17658 ;
  assign n17654 = n13936 ^ n8465 ;
  assign n17648 = n17645 ^ x14 ;
  assign n17649 = n12137 ^ x13 ;
  assign n17650 = n17649 ^ n12137 ;
  assign n17651 = ~n13936 & ~n17650 ;
  assign n17652 = n17651 ^ n12137 ;
  assign n17653 = ~n17648 & ~n17652 ;
  assign n17655 = n17654 ^ n17653 ;
  assign n17660 = n17659 ^ n17655 ;
  assign n17661 = ~n17647 & n17660 ;
  assign n17663 = n17662 ^ n17661 ;
  assign n17684 = n17327 ^ n17156 ;
  assign n17665 = ~n6072 & ~n12142 ;
  assign n17664 = ~n6074 & n12207 ;
  assign n17666 = n17665 ^ n17664 ;
  assign n17667 = n17666 ^ n6060 ;
  assign n17668 = n17667 ^ x14 ;
  assign n17670 = n12138 ^ n6063 ;
  assign n17671 = n17670 ^ x13 ;
  assign n17672 = n17671 ^ n12138 ;
  assign n17676 = ~n14370 & ~n17672 ;
  assign n17677 = ~x13 & n17676 ;
  assign n17680 = n17677 ^ n17676 ;
  assign n17669 = n17666 ^ n6062 ;
  assign n17673 = n17672 ^ n17669 ;
  assign n17675 = n17673 ^ n17672 ;
  assign n17678 = n17677 ^ n12138 ;
  assign n17679 = n17675 & n17678 ;
  assign n17681 = n17680 ^ n17679 ;
  assign n17682 = n17681 ^ n6063 ;
  assign n17683 = ~n17668 & ~n17682 ;
  assign n17685 = n17684 ^ n17683 ;
  assign n17709 = n17324 ^ n17170 ;
  assign n17687 = ~n6072 & n12143 ;
  assign n17686 = ~n6074 & ~n12142 ;
  assign n17688 = n17687 ^ n17686 ;
  assign n17689 = n17688 ^ n6060 ;
  assign n17690 = n17689 ^ x14 ;
  assign n17705 = n12207 ^ n6063 ;
  assign n17694 = n17688 ^ n6062 ;
  assign n17704 = ~n14476 & ~n17542 ;
  assign n17698 = n17704 ^ n12207 ;
  assign n17699 = ~n17694 & ~n17698 ;
  assign n17706 = n17705 ^ n17699 ;
  assign n17707 = n17706 ^ n17704 ;
  assign n17708 = ~n17690 & n17707 ;
  assign n17710 = n17709 ^ n17708 ;
  assign n17736 = n17321 ^ n17308 ;
  assign n17712 = ~n6072 & n12149 ;
  assign n17711 = ~n6074 & n12143 ;
  assign n17713 = n17712 ^ n17711 ;
  assign n17714 = n17713 ^ n6060 ;
  assign n17715 = n17714 ^ x14 ;
  assign n17732 = n12142 ^ n6063 ;
  assign n17719 = n17713 ^ n6062 ;
  assign n17731 = ~n14298 & ~n17542 ;
  assign n17725 = n17731 ^ n12142 ;
  assign n17726 = ~n17719 & n17725 ;
  assign n17733 = n17732 ^ n17726 ;
  assign n17734 = n17733 ^ n17731 ;
  assign n17735 = ~n17715 & ~n17734 ;
  assign n17737 = n17736 ^ n17735 ;
  assign n18019 = n17303 ^ n17180 ;
  assign n17755 = n17300 ^ n17190 ;
  assign n17745 = ~n6072 & n12152 ;
  assign n17744 = ~n6074 & ~n12151 ;
  assign n17746 = n17745 ^ n17744 ;
  assign n17738 = n12149 ^ x13 ;
  assign n17739 = n17738 ^ n12149 ;
  assign n17747 = ~n15311 & ~n17739 ;
  assign n17748 = n17747 ^ n12149 ;
  assign n17749 = n6060 & ~n17748 ;
  assign n17750 = n17749 ^ n16242 ;
  assign n17751 = n17750 ^ x14 ;
  assign n17752 = ~n17746 & ~n17751 ;
  assign n17753 = n17752 ^ x14 ;
  assign n17741 = ~n15311 & n17739 ;
  assign n17742 = n17741 ^ n12149 ;
  assign n17743 = n6063 & n17742 ;
  assign n17754 = n17753 ^ n17743 ;
  assign n17756 = n17755 ^ n17754 ;
  assign n17765 = n17297 ^ n17200 ;
  assign n17760 = ~n6074 & n12152 ;
  assign n17759 = ~n6072 & n12160 ;
  assign n17761 = n17760 ^ n17759 ;
  assign n17762 = n17761 ^ x14 ;
  assign n17758 = n8435 & ~n15299 ;
  assign n17763 = n17762 ^ n17758 ;
  assign n17757 = n4897 & ~n12151 ;
  assign n17764 = n17763 ^ n17757 ;
  assign n17766 = n17765 ^ n17764 ;
  assign n17783 = n17294 ^ n17215 ;
  assign n17768 = ~n6072 & n12163 ;
  assign n17767 = ~n6074 & n12160 ;
  assign n17769 = n17768 ^ n17767 ;
  assign n17770 = n17769 ^ n6060 ;
  assign n17771 = n17770 ^ x14 ;
  assign n17780 = n6063 & n14580 ;
  assign n17772 = n17769 ^ n6062 ;
  assign n17775 = n12152 ^ x13 ;
  assign n17776 = n17775 ^ n12152 ;
  assign n17777 = ~n14580 & ~n17776 ;
  assign n17778 = n17777 ^ n12152 ;
  assign n17779 = n17772 & ~n17778 ;
  assign n17781 = n17780 ^ n17779 ;
  assign n17782 = ~n17771 & ~n17781 ;
  assign n17784 = n17783 ^ n17782 ;
  assign n17804 = n17291 ^ n17225 ;
  assign n17786 = ~n6072 & n12167 ;
  assign n17785 = ~n6074 & n12163 ;
  assign n17787 = n17786 ^ n17785 ;
  assign n17788 = n17787 ^ n6060 ;
  assign n17789 = n17788 ^ x14 ;
  assign n17799 = n8465 & n12160 ;
  assign n17798 = x13 & n14867 ;
  assign n17800 = n17799 ^ n17798 ;
  assign n17801 = ~n6063 & n17800 ;
  assign n17796 = n14866 ^ n8465 ;
  assign n17790 = n17787 ^ x14 ;
  assign n17793 = ~x13 & ~n14866 ;
  assign n17794 = n17793 ^ n12160 ;
  assign n17795 = ~n17790 & ~n17794 ;
  assign n17797 = n17796 ^ n17795 ;
  assign n17802 = n17801 ^ n17797 ;
  assign n17803 = ~n17789 & n17802 ;
  assign n17805 = n17804 ^ n17803 ;
  assign n17808 = ~n6072 & n12168 ;
  assign n17807 = ~n6074 & n12167 ;
  assign n17809 = n17808 ^ n17807 ;
  assign n17810 = n17809 ^ n6060 ;
  assign n17811 = n17810 ^ x14 ;
  assign n17820 = n6063 & n14880 ;
  assign n17812 = n17809 ^ n6062 ;
  assign n17815 = n12163 ^ x13 ;
  assign n17816 = n17815 ^ n12163 ;
  assign n17817 = ~n14880 & ~n17816 ;
  assign n17818 = n17817 ^ n12163 ;
  assign n17819 = n17812 & ~n17818 ;
  assign n17821 = n17820 ^ n17819 ;
  assign n17822 = ~n17811 & ~n17821 ;
  assign n18006 = n17822 ^ n17803 ;
  assign n17806 = n17288 ^ n17236 ;
  assign n17823 = n17822 ^ n17806 ;
  assign n17843 = n17286 ^ n17275 ;
  assign n17825 = ~n6072 & ~n12169 ;
  assign n17824 = ~n6074 & n12168 ;
  assign n17826 = n17825 ^ n17824 ;
  assign n17827 = n17826 ^ n6060 ;
  assign n17828 = n17827 ^ x14 ;
  assign n17839 = n14914 ^ n8465 ;
  assign n17833 = n17826 ^ x14 ;
  assign n17834 = n12167 ^ x13 ;
  assign n17835 = n17834 ^ n12167 ;
  assign n17836 = ~n14914 & ~n17835 ;
  assign n17837 = n17836 ^ n12167 ;
  assign n17838 = ~n17833 & ~n17837 ;
  assign n17840 = n17839 ^ n17838 ;
  assign n17830 = n8465 & n12167 ;
  assign n17829 = x13 & n14915 ;
  assign n17831 = n17830 ^ n17829 ;
  assign n17832 = ~n6063 & n17831 ;
  assign n17841 = n17840 ^ n17832 ;
  assign n17842 = ~n17828 & n17841 ;
  assign n17844 = n17843 ^ n17842 ;
  assign n17864 = n17272 ^ n17264 ;
  assign n17846 = ~n6074 & ~n12169 ;
  assign n17845 = ~n6072 & n12175 ;
  assign n17847 = n17846 ^ n17845 ;
  assign n17848 = n17847 ^ n6060 ;
  assign n17849 = n17848 ^ x14 ;
  assign n17859 = n8465 & n12168 ;
  assign n17858 = x13 & n14949 ;
  assign n17860 = n17859 ^ n17858 ;
  assign n17861 = ~n6063 & n17860 ;
  assign n17856 = n14948 ^ n8465 ;
  assign n17850 = n17847 ^ x14 ;
  assign n17851 = n12168 ^ x13 ;
  assign n17852 = n17851 ^ n12168 ;
  assign n17853 = ~n14948 & ~n17852 ;
  assign n17854 = n17853 ^ n12168 ;
  assign n17855 = ~n17850 & ~n17854 ;
  assign n17857 = n17856 ^ n17855 ;
  assign n17862 = n17861 ^ n17857 ;
  assign n17863 = ~n17849 & n17862 ;
  assign n17865 = n17864 ^ n17863 ;
  assign n17882 = n17244 ^ x17 ;
  assign n17883 = n17882 ^ n17255 ;
  assign n17884 = n17883 ^ n17243 ;
  assign n17872 = n12169 ^ x13 ;
  assign n17871 = n12169 ^ n6063 ;
  assign n17873 = n17872 ^ n17871 ;
  assign n17874 = n15032 & ~n17873 ;
  assign n17875 = n17874 ^ n17872 ;
  assign n17876 = n4897 & ~n17875 ;
  assign n17867 = ~n6072 & n12179 ;
  assign n17866 = ~n6074 & n12175 ;
  assign n17868 = n17867 ^ n17866 ;
  assign n17869 = n17868 ^ n16242 ;
  assign n17877 = n17876 ^ n17869 ;
  assign n17885 = n17884 ^ n17877 ;
  assign n17907 = n5706 ^ n5696 ;
  assign n17908 = n17907 ^ n5710 ;
  assign n17909 = ~n12182 & n17908 ;
  assign n17905 = x17 & ~n12184 ;
  assign n17906 = n17252 & ~n17905 ;
  assign n17910 = n17909 ^ n17906 ;
  assign n17915 = n17252 ^ n5693 ;
  assign n17916 = n17906 ^ n17905 ;
  assign n17917 = n17915 & n17916 ;
  assign n17911 = n12183 ^ n12182 ;
  assign n17912 = n5700 & n17911 ;
  assign n17918 = n17917 ^ n17912 ;
  assign n17913 = ~n12183 & ~n17253 ;
  assign n17914 = n17912 & n17913 ;
  assign n17919 = n17918 ^ n17914 ;
  assign n17920 = ~n17910 & ~n17919 ;
  assign n17887 = ~n6072 & n12180 ;
  assign n17886 = ~n6074 & n12179 ;
  assign n17888 = n17887 ^ n17886 ;
  assign n17889 = n17888 ^ n6060 ;
  assign n17890 = n17889 ^ x14 ;
  assign n17900 = n8465 & n12175 ;
  assign n17899 = x13 & n15049 ;
  assign n17901 = n17900 ^ n17899 ;
  assign n17902 = ~n6063 & n17901 ;
  assign n17897 = n15048 ^ n8465 ;
  assign n17891 = n17888 ^ x14 ;
  assign n17894 = ~x13 & ~n15048 ;
  assign n17895 = n17894 ^ n12175 ;
  assign n17896 = ~n17891 & ~n17895 ;
  assign n17898 = n17897 ^ n17896 ;
  assign n17903 = n17902 ^ n17898 ;
  assign n17904 = ~n17890 & n17903 ;
  assign n17921 = n17920 ^ n17904 ;
  assign n17926 = ~n6072 & n12181 ;
  assign n17925 = ~n6074 & n12180 ;
  assign n17927 = n17926 ^ n17925 ;
  assign n17928 = n17927 ^ n6060 ;
  assign n17929 = n17928 ^ x14 ;
  assign n17938 = n6063 & n15127 ;
  assign n17930 = n17927 ^ n6062 ;
  assign n17933 = n12179 ^ x13 ;
  assign n17934 = n17933 ^ n12179 ;
  assign n17935 = ~n15127 & ~n17934 ;
  assign n17936 = n17935 ^ n12179 ;
  assign n17937 = n17930 & ~n17936 ;
  assign n17939 = n17938 ^ n17937 ;
  assign n17940 = ~n17929 & ~n17939 ;
  assign n17991 = n17940 ^ n17920 ;
  assign n17923 = n5698 & ~n12183 ;
  assign n17922 = n5693 & ~n12182 ;
  assign n17924 = n17923 ^ n17922 ;
  assign n17941 = n17940 ^ n17924 ;
  assign n17983 = ~n6072 & ~n12182 ;
  assign n17982 = ~n6074 & n12181 ;
  assign n17984 = n17983 ^ n17982 ;
  assign n17985 = n17984 ^ x14 ;
  assign n17977 = n12180 ^ n4899 ;
  assign n17978 = n17977 ^ n12180 ;
  assign n17979 = ~n12225 & n17978 ;
  assign n17980 = n17979 ^ n12180 ;
  assign n17981 = n4897 & n17980 ;
  assign n17986 = n17985 ^ n17981 ;
  assign n17988 = n17986 ^ n17940 ;
  assign n17942 = n5693 & ~n12183 ;
  assign n17944 = ~n6072 & ~n12183 ;
  assign n17943 = ~n6074 & ~n12182 ;
  assign n17945 = n17944 ^ n17943 ;
  assign n17946 = n17945 ^ n6060 ;
  assign n17947 = n17946 ^ x14 ;
  assign n17963 = n12181 ^ n6063 ;
  assign n17951 = n17945 ^ n6062 ;
  assign n17962 = n12185 & ~n17542 ;
  assign n17956 = n17962 ^ n12181 ;
  assign n17957 = ~n17951 & ~n17956 ;
  assign n17964 = n17963 ^ n17957 ;
  assign n17965 = n17964 ^ n17962 ;
  assign n17966 = ~n17947 & n17965 ;
  assign n17967 = n12182 ^ n4907 ;
  assign n17968 = ~n4897 & ~n17967 ;
  assign n17969 = n17968 ^ n12182 ;
  assign n17970 = n12183 ^ n4897 ;
  assign n17971 = n17970 ^ x14 ;
  assign n17972 = n17969 & n17971 ;
  assign n17973 = n17972 ^ n4897 ;
  assign n17974 = x14 & ~n17973 ;
  assign n17975 = ~n17966 & n17974 ;
  assign n17976 = ~n17942 & ~n17975 ;
  assign n17987 = n17976 & n17986 ;
  assign n17989 = n17988 ^ n17987 ;
  assign n17990 = ~n17941 & ~n17989 ;
  assign n17992 = n17991 ^ n17990 ;
  assign n17993 = n17921 & n17992 ;
  assign n17994 = n17993 ^ n17920 ;
  assign n17995 = n17994 ^ n17877 ;
  assign n17996 = n17885 & n17995 ;
  assign n17997 = n17996 ^ n17884 ;
  assign n17998 = n17997 ^ n17863 ;
  assign n17999 = ~n17865 & ~n17998 ;
  assign n18000 = n17999 ^ n17863 ;
  assign n18001 = n18000 ^ n17842 ;
  assign n18002 = ~n17844 & n18001 ;
  assign n18003 = n18002 ^ n17842 ;
  assign n18004 = n18003 ^ n17822 ;
  assign n18005 = ~n17823 & n18004 ;
  assign n18007 = n18006 ^ n18005 ;
  assign n18008 = ~n17805 & ~n18007 ;
  assign n18009 = n18008 ^ n17804 ;
  assign n18010 = n18009 ^ n17782 ;
  assign n18011 = ~n17784 & ~n18010 ;
  assign n18012 = n18011 ^ n17782 ;
  assign n18013 = n18012 ^ n17764 ;
  assign n18014 = n17766 & ~n18013 ;
  assign n18015 = n18014 ^ n17764 ;
  assign n18016 = n18015 ^ n17754 ;
  assign n18017 = n17756 & ~n18016 ;
  assign n18018 = n18017 ^ n18015 ;
  assign n18020 = n18019 ^ n18018 ;
  assign n18027 = ~n6072 & ~n12151 ;
  assign n18026 = ~n6074 & n12149 ;
  assign n18028 = n18027 ^ n18026 ;
  assign n18029 = n18028 ^ x14 ;
  assign n18021 = n12143 ^ n4899 ;
  assign n18022 = n18021 ^ n12143 ;
  assign n18023 = ~n15280 & n18022 ;
  assign n18024 = n18023 ^ n12143 ;
  assign n18025 = n4897 & n18024 ;
  assign n18030 = n18029 ^ n18025 ;
  assign n18031 = n18030 ^ n18019 ;
  assign n18032 = n18020 & n18031 ;
  assign n18033 = n18032 ^ n18019 ;
  assign n18034 = n18033 ^ n17735 ;
  assign n18035 = ~n17737 & ~n18034 ;
  assign n18036 = n18035 ^ n17735 ;
  assign n18037 = n18036 ^ n17708 ;
  assign n18038 = ~n17710 & n18037 ;
  assign n18039 = n18038 ^ n17708 ;
  assign n18040 = n18039 ^ n17683 ;
  assign n18041 = ~n17685 & n18040 ;
  assign n18042 = n18041 ^ n17683 ;
  assign n18043 = n18042 ^ n17661 ;
  assign n18044 = ~n17663 & n18043 ;
  assign n18045 = n18044 ^ n17661 ;
  assign n18046 = n18045 ^ n17640 ;
  assign n18047 = ~n17642 & n18046 ;
  assign n18048 = n18047 ^ n17640 ;
  assign n18049 = n18048 ^ n17615 ;
  assign n18050 = ~n17617 & n18049 ;
  assign n18051 = n18050 ^ n17615 ;
  assign n18052 = n18051 ^ n17597 ;
  assign n18053 = n17599 & n18052 ;
  assign n18054 = n18053 ^ n17597 ;
  assign n18055 = n18054 ^ n17577 ;
  assign n18056 = n17578 & n18055 ;
  assign n18057 = n18056 ^ n17577 ;
  assign n18058 = n18057 ^ n17558 ;
  assign n18059 = n17560 & n18058 ;
  assign n18060 = n18059 ^ n17558 ;
  assign n18061 = n18060 ^ n17530 ;
  assign n18062 = n17532 & n18061 ;
  assign n18063 = n18062 ^ n17530 ;
  assign n18064 = n18063 ^ n17512 ;
  assign n18065 = n17514 & ~n18064 ;
  assign n18066 = n18065 ^ n18063 ;
  assign n18067 = n18066 ^ n17500 ;
  assign n18068 = n17502 & ~n18067 ;
  assign n18069 = n18068 ^ n18066 ;
  assign n18070 = n18069 ^ n17479 ;
  assign n18071 = n17481 & n18070 ;
  assign n18072 = n18071 ^ n17479 ;
  assign n18073 = n18072 ^ n17459 ;
  assign n18074 = ~n17460 & n18073 ;
  assign n18075 = n18074 ^ n17459 ;
  assign n18076 = n18075 ^ n17440 ;
  assign n18077 = n17442 & ~n18076 ;
  assign n18078 = n18077 ^ n17440 ;
  assign n17429 = n17428 ^ n17420 ;
  assign n18079 = n18078 ^ n17429 ;
  assign n18083 = n7146 & ~n12705 ;
  assign n18082 = n8054 & n12971 ;
  assign n18084 = n18083 ^ n18082 ;
  assign n18085 = n18084 ^ x8 ;
  assign n18081 = n7135 & ~n12972 ;
  assign n18086 = n18085 ^ n18081 ;
  assign n18080 = n7141 & n12755 ;
  assign n18087 = n18086 ^ n18080 ;
  assign n18088 = n18087 ^ n18078 ;
  assign n18089 = ~n18079 & n18088 ;
  assign n18090 = n18089 ^ n18078 ;
  assign n18122 = n18121 ^ n18090 ;
  assign n18123 = n18121 ^ n14314 ;
  assign n18124 = n18122 & n18123 ;
  assign n18125 = n18124 ^ n14314 ;
  assign n18126 = n18120 ^ n18105 ;
  assign n18127 = ~n18110 & ~n18126 ;
  assign n18128 = n18127 ^ n18105 ;
  assign n18129 = n18125 & n18128 ;
  assign n18167 = n16703 ^ n16692 ;
  assign n18157 = ~n12855 & n18156 ;
  assign n18161 = n18156 ^ x8 ;
  assign n18145 = n6650 & ~n12705 ;
  assign n18143 = ~n12756 & n15413 ;
  assign n18140 = n6655 & n12656 ;
  assign n18139 = n6658 & n12755 ;
  assign n18141 = n18140 ^ n18139 ;
  assign n18142 = n18141 ^ x11 ;
  assign n18144 = n18143 ^ n18142 ;
  assign n18146 = n18145 ^ n18144 ;
  assign n18148 = n18146 ^ n18104 ;
  assign n18147 = n18146 ^ n18091 ;
  assign n18149 = n18148 ^ n18147 ;
  assign n18150 = ~n18096 & ~n18149 ;
  assign n18151 = n18150 ^ n18147 ;
  assign n18152 = n16688 ^ n16340 ;
  assign n18158 = n18152 ^ n18146 ;
  assign n18159 = n18151 & n18158 ;
  assign n18160 = n18159 ^ n18152 ;
  assign n18162 = n18161 ^ n18160 ;
  assign n18163 = n18162 ^ x7 ;
  assign n18164 = n18163 ^ n18160 ;
  assign n18165 = n18157 & ~n18164 ;
  assign n18166 = n18165 ^ n18162 ;
  assign n18168 = n18167 ^ n18166 ;
  assign n18136 = n8054 ^ x8 ;
  assign n18131 = n12987 ^ n7141 ;
  assign n18132 = n18131 ^ n7141 ;
  assign n18133 = n7135 & ~n18132 ;
  assign n18134 = n18133 ^ n7141 ;
  assign n18135 = ~n12855 & n18134 ;
  assign n18137 = n18136 ^ n18135 ;
  assign n18130 = n7146 & n12971 ;
  assign n18138 = n18137 ^ n18130 ;
  assign n18153 = n18152 ^ n18151 ;
  assign n18154 = ~n18138 & n18153 ;
  assign n18169 = n18168 ^ n18154 ;
  assign n18170 = n18128 ^ n18125 ;
  assign n18171 = n18170 ^ n18129 ;
  assign n18172 = n18171 ^ n18168 ;
  assign n18173 = n18169 & ~n18172 ;
  assign n18174 = n18173 ^ n18154 ;
  assign n18189 = n18075 ^ n17442 ;
  assign n18176 = n7146 & n12656 ;
  assign n18175 = n7141 & ~n12705 ;
  assign n18177 = n18176 ^ n18175 ;
  assign n18178 = n18177 ^ n7129 ;
  assign n18179 = n18178 ^ x8 ;
  assign n18180 = n18177 ^ x8 ;
  assign n18184 = n18180 ^ n7130 ;
  assign n18185 = ~x7 & ~n12724 ;
  assign n18186 = n18184 & n18185 ;
  assign n18182 = n7130 & ~n12756 ;
  assign n18181 = ~n12755 & n18180 ;
  assign n18183 = n18182 ^ n18181 ;
  assign n18187 = n18186 ^ n18183 ;
  assign n18188 = ~n18179 & ~n18187 ;
  assign n18190 = n18189 ^ n18188 ;
  assign n18198 = n12368 & n15413 ;
  assign n18196 = n6655 & n11972 ;
  assign n18194 = n6658 & ~n12367 ;
  assign n18192 = n18072 ^ n17460 ;
  assign n18193 = n18192 ^ x11 ;
  assign n18195 = n18194 ^ n18193 ;
  assign n18197 = n18196 ^ n18195 ;
  assign n18199 = n18198 ^ n18197 ;
  assign n18191 = n6650 & ~n12108 ;
  assign n18200 = n18199 ^ n18191 ;
  assign n18208 = n12376 & n15413 ;
  assign n18206 = n6655 & n12260 ;
  assign n18204 = n6658 & ~n12108 ;
  assign n18202 = n18069 ^ n17481 ;
  assign n18203 = n18202 ^ x11 ;
  assign n18205 = n18204 ^ n18203 ;
  assign n18207 = n18206 ^ n18205 ;
  assign n18209 = n18208 ^ n18207 ;
  assign n18201 = n6650 & n11972 ;
  assign n18210 = n18209 ^ n18201 ;
  assign n18215 = n18066 ^ n17502 ;
  assign n18216 = n18215 ^ x11 ;
  assign n18214 = n6650 & n12260 ;
  assign n18217 = n18216 ^ n18214 ;
  assign n18213 = ~n14078 & n15413 ;
  assign n18218 = n18217 ^ n18213 ;
  assign n18212 = n6658 & n11972 ;
  assign n18219 = n18218 ^ n18212 ;
  assign n18211 = n6655 & ~n12256 ;
  assign n18220 = n18219 ^ n18211 ;
  assign n18223 = n6655 & ~n12262 ;
  assign n18222 = n6650 & ~n12256 ;
  assign n18224 = n18223 ^ n18222 ;
  assign n18225 = n18224 ^ n6656 ;
  assign n18226 = n18225 ^ x11 ;
  assign n18227 = n18224 ^ x11 ;
  assign n18231 = n18227 ^ n6657 ;
  assign n18232 = ~x10 & n13053 ;
  assign n18233 = n18231 & n18232 ;
  assign n18229 = n6657 & n13054 ;
  assign n18228 = ~n12260 & n18227 ;
  assign n18230 = n18229 ^ n18228 ;
  assign n18234 = n18233 ^ n18230 ;
  assign n18235 = ~n18226 & ~n18234 ;
  assign n18221 = n18063 ^ n17514 ;
  assign n18236 = n18235 ^ n18221 ;
  assign n18598 = n18060 ^ n17532 ;
  assign n18244 = n13712 & n15413 ;
  assign n18242 = n6655 & ~n12110 ;
  assign n18240 = n6658 & ~n12262 ;
  assign n18238 = n18057 ^ n17560 ;
  assign n18239 = n18238 ^ x11 ;
  assign n18241 = n18240 ^ n18239 ;
  assign n18243 = n18242 ^ n18241 ;
  assign n18245 = n18244 ^ n18243 ;
  assign n18237 = n6650 & ~n12220 ;
  assign n18246 = n18245 ^ n18237 ;
  assign n18255 = n18054 ^ n17578 ;
  assign n18250 = n6655 & n12117 ;
  assign n18249 = n6658 & ~n12220 ;
  assign n18251 = n18250 ^ n18249 ;
  assign n18252 = n18251 ^ x11 ;
  assign n18248 = n14047 & n15413 ;
  assign n18253 = n18252 ^ n18248 ;
  assign n18247 = n6650 & ~n12110 ;
  assign n18254 = n18253 ^ n18247 ;
  assign n18256 = n18255 ^ n18254 ;
  assign n18264 = n13196 & n15413 ;
  assign n18262 = n6655 & n12121 ;
  assign n18260 = n6658 & ~n12110 ;
  assign n18258 = n18051 ^ n17599 ;
  assign n18259 = n18258 ^ x11 ;
  assign n18261 = n18260 ^ n18259 ;
  assign n18263 = n18262 ^ n18261 ;
  assign n18265 = n18264 ^ n18263 ;
  assign n18257 = n6650 & n12117 ;
  assign n18266 = n18265 ^ n18257 ;
  assign n18275 = n18048 ^ n17617 ;
  assign n18270 = n6655 & ~n12129 ;
  assign n18269 = n6658 & n12117 ;
  assign n18271 = n18270 ^ n18269 ;
  assign n18272 = n18271 ^ x11 ;
  assign n18268 = ~n13596 & n15413 ;
  assign n18273 = n18272 ^ n18268 ;
  assign n18267 = n6650 & n12121 ;
  assign n18274 = n18273 ^ n18267 ;
  assign n18276 = n18275 ^ n18274 ;
  assign n18285 = n18045 ^ n17642 ;
  assign n18280 = n6655 & n12130 ;
  assign n18279 = n6658 & n12121 ;
  assign n18281 = n18280 ^ n18279 ;
  assign n18282 = n18281 ^ x11 ;
  assign n18278 = ~n13606 & n15413 ;
  assign n18283 = n18282 ^ n18278 ;
  assign n18277 = n6650 & ~n12129 ;
  assign n18284 = n18283 ^ n18277 ;
  assign n18286 = n18285 ^ n18284 ;
  assign n18295 = n18042 ^ n17663 ;
  assign n18293 = n6650 & n12130 ;
  assign n18291 = n13737 & n15413 ;
  assign n18288 = n6655 & ~n12136 ;
  assign n18287 = n6658 & ~n12129 ;
  assign n18289 = n18288 ^ n18287 ;
  assign n18290 = n18289 ^ x11 ;
  assign n18292 = n18291 ^ n18290 ;
  assign n18294 = n18293 ^ n18292 ;
  assign n18296 = n18295 ^ n18294 ;
  assign n18304 = ~n13818 & n15413 ;
  assign n18302 = n6655 & n12137 ;
  assign n18300 = n6658 & n12130 ;
  assign n18298 = n18039 ^ n17685 ;
  assign n18299 = n18298 ^ x11 ;
  assign n18301 = n18300 ^ n18299 ;
  assign n18303 = n18302 ^ n18301 ;
  assign n18305 = n18304 ^ n18303 ;
  assign n18297 = n6650 & ~n12136 ;
  assign n18306 = n18305 ^ n18297 ;
  assign n18315 = n18036 ^ n17710 ;
  assign n18310 = n6655 & ~n12138 ;
  assign n18309 = n6658 & ~n12136 ;
  assign n18311 = n18310 ^ n18309 ;
  assign n18312 = n18311 ^ x11 ;
  assign n18308 = n14129 & n15413 ;
  assign n18313 = n18312 ^ n18308 ;
  assign n18307 = n6650 & n12137 ;
  assign n18314 = n18313 ^ n18307 ;
  assign n18316 = n18315 ^ n18314 ;
  assign n18325 = n18033 ^ n17737 ;
  assign n18323 = n6650 & ~n12138 ;
  assign n18321 = ~n13939 & n15413 ;
  assign n18318 = n6655 & n12207 ;
  assign n18317 = n6658 & n12137 ;
  assign n18319 = n18318 ^ n18317 ;
  assign n18320 = n18319 ^ x11 ;
  assign n18322 = n18321 ^ n18320 ;
  assign n18324 = n18323 ^ n18322 ;
  assign n18326 = n18325 ^ n18324 ;
  assign n18335 = n18031 ^ n18018 ;
  assign n18333 = n6650 & n12207 ;
  assign n18331 = n14832 & n15413 ;
  assign n18328 = n6655 & ~n12142 ;
  assign n18327 = n6658 & ~n12138 ;
  assign n18329 = n18328 ^ n18327 ;
  assign n18330 = n18329 ^ x11 ;
  assign n18332 = n18331 ^ n18330 ;
  assign n18334 = n18333 ^ n18332 ;
  assign n18336 = n18335 ^ n18334 ;
  assign n18345 = n18015 ^ n17756 ;
  assign n18340 = n6655 & n12143 ;
  assign n18339 = n6658 & n12207 ;
  assign n18341 = n18340 ^ n18339 ;
  assign n18342 = n18341 ^ x11 ;
  assign n18338 = n15413 & ~n15500 ;
  assign n18343 = n18342 ^ n18338 ;
  assign n18337 = n6650 & ~n12142 ;
  assign n18344 = n18343 ^ n18337 ;
  assign n18346 = n18345 ^ n18344 ;
  assign n18355 = n18012 ^ n17766 ;
  assign n18350 = n6655 & n12149 ;
  assign n18349 = n6658 & ~n12142 ;
  assign n18351 = n18350 ^ n18349 ;
  assign n18352 = n18351 ^ x11 ;
  assign n18348 = n14299 & n15413 ;
  assign n18353 = n18352 ^ n18348 ;
  assign n18347 = n6650 & n12143 ;
  assign n18354 = n18353 ^ n18347 ;
  assign n18356 = n18355 ^ n18354 ;
  assign n18365 = n18009 ^ n17784 ;
  assign n18360 = n6655 & ~n12151 ;
  assign n18359 = n6658 & n12143 ;
  assign n18361 = n18360 ^ n18359 ;
  assign n18362 = n18361 ^ x11 ;
  assign n18358 = ~n14498 & n15413 ;
  assign n18363 = n18362 ^ n18358 ;
  assign n18357 = n6650 & n12149 ;
  assign n18364 = n18363 ^ n18357 ;
  assign n18366 = n18365 ^ n18364 ;
  assign n18378 = n18007 ^ n17804 ;
  assign n18373 = n6655 & n12152 ;
  assign n18372 = n6650 & ~n12151 ;
  assign n18374 = n18373 ^ n18372 ;
  assign n18375 = n18374 ^ x11 ;
  assign n18367 = ~x10 & ~n15311 ;
  assign n18370 = n18367 ^ n12149 ;
  assign n18371 = n6656 & n18370 ;
  assign n18376 = n18375 ^ n18371 ;
  assign n18368 = n18367 ^ n15312 ;
  assign n18369 = n6657 & ~n18368 ;
  assign n18377 = n18376 ^ n18369 ;
  assign n18379 = n18378 ^ n18377 ;
  assign n18390 = n18003 ^ n17823 ;
  assign n18386 = n6650 & n12152 ;
  assign n18385 = n6655 & n12160 ;
  assign n18387 = n18386 ^ n18385 ;
  assign n18388 = n18387 ^ x11 ;
  assign n18380 = n12151 ^ n9154 ;
  assign n18381 = n18380 ^ n12151 ;
  assign n18382 = ~n15299 & n18381 ;
  assign n18383 = n18382 ^ n12151 ;
  assign n18384 = n6648 & ~n18383 ;
  assign n18389 = n18388 ^ n18384 ;
  assign n18391 = n18390 ^ n18389 ;
  assign n18406 = n18000 ^ n17844 ;
  assign n18393 = n6655 & n12163 ;
  assign n18392 = n6650 & n12160 ;
  assign n18394 = n18393 ^ n18392 ;
  assign n18395 = n18394 ^ n6656 ;
  assign n18396 = n18395 ^ x11 ;
  assign n18397 = n18394 ^ x11 ;
  assign n18401 = n18397 ^ n6657 ;
  assign n18402 = ~x10 & ~n14580 ;
  assign n18403 = n18401 & n18402 ;
  assign n18399 = n6657 & ~n14581 ;
  assign n18398 = ~n12152 & n18397 ;
  assign n18400 = n18399 ^ n18398 ;
  assign n18404 = n18403 ^ n18400 ;
  assign n18405 = ~n18396 & ~n18404 ;
  assign n18407 = n18406 ^ n18405 ;
  assign n18417 = n6650 & n12163 ;
  assign n18410 = n12160 ^ x11 ;
  assign n18411 = n18410 ^ x10 ;
  assign n18412 = n18411 ^ n12160 ;
  assign n18413 = ~n14866 & n18412 ;
  assign n18414 = n18413 ^ n12160 ;
  assign n18415 = n6648 & n18414 ;
  assign n18416 = n18415 ^ x11 ;
  assign n18418 = n18417 ^ n18416 ;
  assign n18409 = n6655 & n12167 ;
  assign n18419 = n18418 ^ n18409 ;
  assign n18408 = n17997 ^ n17865 ;
  assign n18420 = n18419 ^ n18408 ;
  assign n18436 = n17994 ^ n17885 ;
  assign n18422 = n6655 & n12168 ;
  assign n18421 = n6650 & n12167 ;
  assign n18423 = n18422 ^ n18421 ;
  assign n18424 = n18423 ^ n6656 ;
  assign n18425 = n18424 ^ x11 ;
  assign n18426 = n18423 ^ x11 ;
  assign n18430 = n18426 ^ n6657 ;
  assign n18431 = ~x10 & ~n14880 ;
  assign n18432 = n18430 & n18431 ;
  assign n18428 = n6657 & ~n14890 ;
  assign n18427 = ~n12163 & n18426 ;
  assign n18429 = n18428 ^ n18427 ;
  assign n18433 = n18432 ^ n18429 ;
  assign n18434 = ~n18425 & ~n18433 ;
  assign n18437 = n18436 ^ n18434 ;
  assign n18528 = n17992 ^ n17904 ;
  assign n18484 = n17974 ^ n17966 ;
  assign n18470 = ~n12183 & n16372 ;
  assign n18464 = n17911 ^ n12182 ;
  assign n18465 = n12182 ^ x12 ;
  assign n18466 = n18465 ^ n12182 ;
  assign n18467 = ~n18464 & ~n18466 ;
  assign n18468 = n18467 ^ n12182 ;
  assign n18469 = n4897 & ~n18468 ;
  assign n18471 = n18470 ^ n18469 ;
  assign n18438 = n4897 & ~n12183 ;
  assign n18439 = ~n12184 & ~n16289 ;
  assign n18440 = n12187 ^ n12182 ;
  assign n18441 = n15413 & n18440 ;
  assign n18447 = n6658 & n12181 ;
  assign n18442 = n12181 ^ n6655 ;
  assign n18443 = n18442 ^ n6655 ;
  assign n18444 = n15413 & n18443 ;
  assign n18445 = n18444 ^ n6655 ;
  assign n18446 = ~n12183 & n18445 ;
  assign n18448 = n18447 ^ n18446 ;
  assign n18449 = n18441 & ~n18448 ;
  assign n18450 = n18449 ^ n18448 ;
  assign n18451 = x11 & ~n18450 ;
  assign n18452 = ~n18439 & n18451 ;
  assign n18453 = ~n18438 & ~n18452 ;
  assign n18457 = n6655 & ~n12182 ;
  assign n18456 = n6658 & n12180 ;
  assign n18458 = n18457 ^ n18456 ;
  assign n18459 = n18458 ^ x11 ;
  assign n18455 = ~n15151 & n15413 ;
  assign n18460 = n18459 ^ n18455 ;
  assign n18454 = n6650 & n12181 ;
  assign n18461 = n18460 ^ n18454 ;
  assign n18462 = n18453 & n18461 ;
  assign n18463 = n18462 ^ n18461 ;
  assign n18472 = n18471 ^ n18463 ;
  assign n18479 = ~n15128 & n15413 ;
  assign n18477 = n6655 & n12181 ;
  assign n18475 = n6658 & n12179 ;
  assign n18474 = n18471 ^ x11 ;
  assign n18476 = n18475 ^ n18474 ;
  assign n18478 = n18477 ^ n18476 ;
  assign n18480 = n18479 ^ n18478 ;
  assign n18473 = n6650 & n12180 ;
  assign n18481 = n18480 ^ n18473 ;
  assign n18482 = n18472 & n18481 ;
  assign n18483 = n18482 ^ n18471 ;
  assign n18485 = n18484 ^ n18483 ;
  assign n18493 = n6650 & n12179 ;
  assign n18490 = n6658 & n12175 ;
  assign n18488 = n6655 & n12180 ;
  assign n18487 = n18483 ^ x11 ;
  assign n18489 = n18488 ^ n18487 ;
  assign n18491 = n18490 ^ n18489 ;
  assign n18486 = ~n15049 & n15413 ;
  assign n18492 = n18491 ^ n18486 ;
  assign n18494 = n18493 ^ n18492 ;
  assign n18495 = ~n18485 & ~n18494 ;
  assign n18496 = n18495 ^ n18484 ;
  assign n18497 = n17975 ^ n17942 ;
  assign n18498 = n18497 ^ n17986 ;
  assign n18500 = n18496 & ~n18498 ;
  assign n18499 = n18498 ^ n18496 ;
  assign n18501 = n18500 ^ n18499 ;
  assign n18506 = n6655 & n12179 ;
  assign n18505 = n6658 & ~n12169 ;
  assign n18507 = n18506 ^ n18505 ;
  assign n18503 = n6650 & n12175 ;
  assign n18502 = n15035 & n15413 ;
  assign n18504 = n18503 ^ n18502 ;
  assign n18508 = n18507 ^ n18504 ;
  assign n18509 = n18508 ^ x11 ;
  assign n18516 = n6655 & n12175 ;
  assign n18515 = n6658 & n12168 ;
  assign n18517 = n18516 ^ n18515 ;
  assign n18513 = n6650 & ~n12169 ;
  assign n18512 = ~n14949 & n15413 ;
  assign n18514 = n18513 ^ n18512 ;
  assign n18518 = n18517 ^ n18514 ;
  assign n18510 = n17989 ^ n17924 ;
  assign n18511 = n18510 ^ n18508 ;
  assign n18519 = n18518 ^ n18511 ;
  assign n18520 = ~n18509 & ~n18519 ;
  assign n18521 = ~n18501 & n18520 ;
  assign n18522 = n18510 ^ n18500 ;
  assign n18523 = n18510 ^ x11 ;
  assign n18524 = n18523 ^ n18518 ;
  assign n18525 = n18522 & n18524 ;
  assign n18526 = n18525 ^ n18500 ;
  assign n18527 = ~n18521 & ~n18526 ;
  assign n18529 = n18528 ^ n18527 ;
  assign n18541 = n6655 & ~n12169 ;
  assign n18538 = n18527 ^ x11 ;
  assign n18533 = n12167 ^ n9154 ;
  assign n18534 = n18533 ^ n12167 ;
  assign n18535 = ~n14914 & n18534 ;
  assign n18536 = n18535 ^ n12167 ;
  assign n18537 = n6648 & n18536 ;
  assign n18539 = n18538 ^ n18537 ;
  assign n18530 = n6650 & n12168 ;
  assign n18540 = n18539 ^ n18530 ;
  assign n18542 = n18541 ^ n18540 ;
  assign n18543 = ~n18529 & ~n18542 ;
  assign n18544 = n18543 ^ n18528 ;
  assign n18545 = n18544 ^ n18434 ;
  assign n18546 = n18437 & n18545 ;
  assign n18435 = n18434 ^ n18408 ;
  assign n18547 = n18546 ^ n18435 ;
  assign n18548 = ~n18420 & ~n18547 ;
  assign n18549 = n18548 ^ n18419 ;
  assign n18550 = n18549 ^ n18405 ;
  assign n18551 = ~n18407 & n18550 ;
  assign n18552 = n18551 ^ n18406 ;
  assign n18553 = n18552 ^ n18389 ;
  assign n18554 = n18391 & n18553 ;
  assign n18555 = n18554 ^ n18389 ;
  assign n18556 = n18555 ^ n18377 ;
  assign n18557 = n18379 & n18556 ;
  assign n18558 = n18557 ^ n18377 ;
  assign n18559 = n18558 ^ n18364 ;
  assign n18560 = ~n18366 & n18559 ;
  assign n18561 = n18560 ^ n18364 ;
  assign n18562 = n18561 ^ n18354 ;
  assign n18563 = ~n18356 & n18562 ;
  assign n18564 = n18563 ^ n18354 ;
  assign n18565 = n18564 ^ n18344 ;
  assign n18566 = ~n18346 & n18565 ;
  assign n18567 = n18566 ^ n18344 ;
  assign n18568 = n18567 ^ n18334 ;
  assign n18569 = n18336 & n18568 ;
  assign n18570 = n18569 ^ n18334 ;
  assign n18571 = n18570 ^ n18324 ;
  assign n18572 = ~n18326 & n18571 ;
  assign n18573 = n18572 ^ n18324 ;
  assign n18574 = n18573 ^ n18314 ;
  assign n18575 = n18316 & n18574 ;
  assign n18576 = n18575 ^ n18314 ;
  assign n18577 = n18576 ^ n18298 ;
  assign n18578 = n18306 & n18577 ;
  assign n18579 = n18578 ^ n18298 ;
  assign n18580 = n18579 ^ n18294 ;
  assign n18581 = n18296 & n18580 ;
  assign n18582 = n18581 ^ n18294 ;
  assign n18583 = n18582 ^ n18284 ;
  assign n18584 = n18286 & n18583 ;
  assign n18585 = n18584 ^ n18284 ;
  assign n18586 = n18585 ^ n18274 ;
  assign n18587 = n18276 & n18586 ;
  assign n18588 = n18587 ^ n18274 ;
  assign n18589 = n18588 ^ n18258 ;
  assign n18590 = ~n18266 & ~n18589 ;
  assign n18591 = n18590 ^ n18258 ;
  assign n18592 = n18591 ^ n18254 ;
  assign n18593 = ~n18256 & ~n18592 ;
  assign n18594 = n18593 ^ n18254 ;
  assign n18595 = n18594 ^ n18238 ;
  assign n18596 = ~n18246 & ~n18595 ;
  assign n18597 = n18596 ^ n18238 ;
  assign n18599 = n18598 ^ n18597 ;
  assign n18606 = ~n13283 & n15413 ;
  assign n18604 = n6655 & ~n12220 ;
  assign n18602 = n6658 & ~n12256 ;
  assign n18601 = n18598 ^ x11 ;
  assign n18603 = n18602 ^ n18601 ;
  assign n18605 = n18604 ^ n18603 ;
  assign n18607 = n18606 ^ n18605 ;
  assign n18600 = n6650 & ~n12262 ;
  assign n18608 = n18607 ^ n18600 ;
  assign n18609 = n18599 & ~n18608 ;
  assign n18610 = n18609 ^ n18598 ;
  assign n18611 = n18610 ^ n18235 ;
  assign n18612 = ~n18236 & n18611 ;
  assign n18613 = n18612 ^ n18235 ;
  assign n18614 = n18613 ^ n18215 ;
  assign n18615 = n18220 & ~n18614 ;
  assign n18616 = n18615 ^ n18215 ;
  assign n18617 = n18616 ^ n18202 ;
  assign n18618 = ~n18210 & ~n18617 ;
  assign n18619 = n18618 ^ n18202 ;
  assign n18620 = n18619 ^ n18192 ;
  assign n18621 = n18200 & ~n18620 ;
  assign n18622 = n18621 ^ n18192 ;
  assign n18623 = n18622 ^ n18188 ;
  assign n18624 = n18190 & ~n18623 ;
  assign n18625 = n18624 ^ n18188 ;
  assign n18628 = n18627 ^ x5 ;
  assign n18629 = n18628 ^ x4 ;
  assign n18630 = ~n12855 & n18627 ;
  assign n18631 = ~n18629 & n18630 ;
  assign n18632 = n18631 ^ n18628 ;
  assign n18626 = n18087 ^ n18079 ;
  assign n18633 = n18632 ^ n18626 ;
  assign n18634 = n18626 ^ n18625 ;
  assign n18635 = ~n18633 & ~n18634 ;
  assign n18636 = ~n18625 & n18635 ;
  assign n19664 = n10854 & n12855 ;
  assign n19659 = n9081 & ~n12972 ;
  assign n19137 = n7135 & ~n12872 ;
  assign n19135 = n7146 & ~n12367 ;
  assign n19133 = n8054 & n12656 ;
  assign n19129 = n18616 ^ n18210 ;
  assign n19132 = n19129 ^ x8 ;
  assign n19134 = n19133 ^ n19132 ;
  assign n19136 = n19135 ^ n19134 ;
  assign n19138 = n19137 ^ n19136 ;
  assign n19131 = n7141 & ~n12613 ;
  assign n19139 = n19138 ^ n19131 ;
  assign n18646 = n7135 & n13110 ;
  assign n18644 = n7146 & ~n12108 ;
  assign n18642 = n8054 & ~n12613 ;
  assign n18640 = n18613 ^ n18220 ;
  assign n18641 = n18640 ^ x8 ;
  assign n18643 = n18642 ^ n18641 ;
  assign n18645 = n18644 ^ n18643 ;
  assign n18647 = n18646 ^ n18645 ;
  assign n18639 = n7141 & ~n12367 ;
  assign n18648 = n18647 ^ n18639 ;
  assign n18660 = n18610 ^ n18236 ;
  assign n18657 = n7141 & ~n12108 ;
  assign n18650 = n12367 ^ x8 ;
  assign n18651 = n18650 ^ x7 ;
  assign n18652 = n18651 ^ n12367 ;
  assign n18653 = ~n12369 & n18652 ;
  assign n18654 = n18653 ^ n12367 ;
  assign n18655 = n7128 & ~n18654 ;
  assign n18656 = n18655 ^ x8 ;
  assign n18658 = n18657 ^ n18656 ;
  assign n18649 = n7146 & n11972 ;
  assign n18659 = n18658 ^ n18649 ;
  assign n18661 = n18660 ^ n18659 ;
  assign n19110 = n18608 ^ n18597 ;
  assign n18681 = n18594 ^ n18246 ;
  assign n18663 = n7146 & ~n12256 ;
  assign n18662 = n7141 & n12260 ;
  assign n18664 = n18663 ^ n18662 ;
  assign n18665 = n18664 ^ n7129 ;
  assign n18666 = n18665 ^ x8 ;
  assign n18667 = n18664 ^ x8 ;
  assign n18668 = n18667 ^ n7130 ;
  assign n18669 = n14078 & n18668 ;
  assign n18670 = n18669 ^ n7130 ;
  assign n18671 = n18670 ^ x7 ;
  assign n18672 = n18671 ^ n11972 ;
  assign n18673 = n18672 ^ n18670 ;
  assign n18674 = n18670 ^ n18668 ;
  assign n18675 = n18674 ^ n18670 ;
  assign n18676 = n18673 & n18675 ;
  assign n18677 = n18676 ^ n18670 ;
  assign n18678 = ~n12270 & n18677 ;
  assign n18679 = n18678 ^ n18670 ;
  assign n18680 = ~n18666 & ~n18679 ;
  assign n18682 = n18681 ^ n18680 ;
  assign n18690 = n7135 & n13054 ;
  assign n18688 = n7146 & ~n12262 ;
  assign n18686 = n8054 & n12260 ;
  assign n18684 = n18591 ^ n18256 ;
  assign n18685 = n18684 ^ x8 ;
  assign n18687 = n18686 ^ n18685 ;
  assign n18689 = n18688 ^ n18687 ;
  assign n18691 = n18690 ^ n18689 ;
  assign n18683 = n7141 & ~n12256 ;
  assign n18692 = n18691 ^ n18683 ;
  assign n18700 = n7135 & ~n13283 ;
  assign n18696 = n18588 ^ n18266 ;
  assign n18697 = n18696 ^ x8 ;
  assign n18695 = n8054 & ~n12256 ;
  assign n18698 = n18697 ^ n18695 ;
  assign n18694 = n7146 & ~n12220 ;
  assign n18699 = n18698 ^ n18694 ;
  assign n18701 = n18700 ^ n18699 ;
  assign n18693 = n7141 & ~n12262 ;
  assign n18702 = n18701 ^ n18693 ;
  assign n18711 = n18585 ^ n18276 ;
  assign n18709 = n7141 & ~n12220 ;
  assign n18707 = n7135 & n13712 ;
  assign n18704 = n7146 & ~n12110 ;
  assign n18703 = n8054 & ~n12262 ;
  assign n18705 = n18704 ^ n18703 ;
  assign n18706 = n18705 ^ x8 ;
  assign n18708 = n18707 ^ n18706 ;
  assign n18710 = n18709 ^ n18708 ;
  assign n18712 = n18711 ^ n18710 ;
  assign n18721 = n18582 ^ n18286 ;
  assign n18716 = n7146 & n12117 ;
  assign n18715 = n8054 & ~n12220 ;
  assign n18717 = n18716 ^ n18715 ;
  assign n18718 = n18717 ^ x8 ;
  assign n18714 = n7135 & n14047 ;
  assign n18719 = n18718 ^ n18714 ;
  assign n18713 = n7141 & ~n12110 ;
  assign n18720 = n18719 ^ n18713 ;
  assign n18722 = n18721 ^ n18720 ;
  assign n18731 = n18579 ^ n18296 ;
  assign n18729 = n7141 & n12117 ;
  assign n18727 = n7135 & n13196 ;
  assign n18724 = n7146 & n12121 ;
  assign n18723 = n8054 & ~n12110 ;
  assign n18725 = n18724 ^ n18723 ;
  assign n18726 = n18725 ^ x8 ;
  assign n18728 = n18727 ^ n18726 ;
  assign n18730 = n18729 ^ n18728 ;
  assign n18732 = n18731 ^ n18730 ;
  assign n18744 = n18576 ^ n18306 ;
  assign n18741 = n7141 & n12121 ;
  assign n18734 = n12117 ^ x8 ;
  assign n18735 = n18734 ^ x7 ;
  assign n18736 = n18735 ^ n12117 ;
  assign n18737 = ~n13586 & n18736 ;
  assign n18738 = n18737 ^ n12117 ;
  assign n18739 = n7128 & n18738 ;
  assign n18740 = n18739 ^ x8 ;
  assign n18742 = n18741 ^ n18740 ;
  assign n18733 = n7146 & ~n12129 ;
  assign n18743 = n18742 ^ n18733 ;
  assign n18745 = n18744 ^ n18743 ;
  assign n18748 = n7146 & n12130 ;
  assign n18747 = n7141 & ~n12129 ;
  assign n18749 = n18748 ^ n18747 ;
  assign n18750 = n18749 ^ n7129 ;
  assign n18751 = n18750 ^ x8 ;
  assign n18753 = n18749 ^ x8 ;
  assign n18756 = n18753 ^ n7130 ;
  assign n18757 = ~x7 & ~n13605 ;
  assign n18758 = n18756 & n18757 ;
  assign n18754 = ~n12121 & n18753 ;
  assign n18752 = n7130 & ~n13606 ;
  assign n18755 = n18754 ^ n18752 ;
  assign n18759 = n18758 ^ n18755 ;
  assign n18760 = ~n18751 & ~n18759 ;
  assign n18746 = n18573 ^ n18316 ;
  assign n18761 = n18760 ^ n18746 ;
  assign n18773 = n18570 ^ n18326 ;
  assign n18770 = n7141 & n12130 ;
  assign n18763 = n12129 ^ x8 ;
  assign n18764 = n18763 ^ x7 ;
  assign n18765 = n18764 ^ n12129 ;
  assign n18766 = ~n14271 & n18765 ;
  assign n18767 = n18766 ^ n12129 ;
  assign n18768 = n7128 & ~n18767 ;
  assign n18769 = n18768 ^ x8 ;
  assign n18771 = n18770 ^ n18769 ;
  assign n18762 = n7146 & ~n12136 ;
  assign n18772 = n18771 ^ n18762 ;
  assign n18774 = n18773 ^ n18772 ;
  assign n18789 = n18567 ^ n18336 ;
  assign n18776 = n7146 & n12137 ;
  assign n18775 = n7141 & ~n12136 ;
  assign n18777 = n18776 ^ n18775 ;
  assign n18778 = n18777 ^ n7129 ;
  assign n18779 = n18778 ^ x8 ;
  assign n18780 = n18777 ^ x8 ;
  assign n18784 = n18780 ^ n7130 ;
  assign n18785 = ~x7 & ~n13817 ;
  assign n18786 = n18784 & n18785 ;
  assign n18782 = n7130 & ~n13818 ;
  assign n18781 = ~n12130 & n18780 ;
  assign n18783 = n18782 ^ n18781 ;
  assign n18787 = n18786 ^ n18783 ;
  assign n18788 = ~n18779 & ~n18787 ;
  assign n18790 = n18789 ^ n18788 ;
  assign n18799 = n18564 ^ n18346 ;
  assign n18794 = n7146 & ~n12138 ;
  assign n18793 = n8054 & ~n12136 ;
  assign n18795 = n18794 ^ n18793 ;
  assign n18796 = n18795 ^ x8 ;
  assign n18792 = n7135 & n14129 ;
  assign n18797 = n18796 ^ n18792 ;
  assign n18791 = n7141 & n12137 ;
  assign n18798 = n18797 ^ n18791 ;
  assign n18800 = n18799 ^ n18798 ;
  assign n18812 = n18561 ^ n18356 ;
  assign n18809 = n7141 & ~n12138 ;
  assign n18802 = n12137 ^ x8 ;
  assign n18803 = n18802 ^ x7 ;
  assign n18804 = n18803 ^ n12137 ;
  assign n18805 = ~n13936 & n18804 ;
  assign n18806 = n18805 ^ n12137 ;
  assign n18807 = n7128 & n18806 ;
  assign n18808 = n18807 ^ x8 ;
  assign n18810 = n18809 ^ n18808 ;
  assign n18801 = n7146 & n12207 ;
  assign n18811 = n18810 ^ n18801 ;
  assign n18813 = n18812 ^ n18811 ;
  assign n18822 = n18558 ^ n18366 ;
  assign n18820 = n7141 & n12207 ;
  assign n18818 = n7135 & n14832 ;
  assign n18815 = n7146 & ~n12142 ;
  assign n18814 = n8054 & ~n12138 ;
  assign n18816 = n18815 ^ n18814 ;
  assign n18817 = n18816 ^ x8 ;
  assign n18819 = n18818 ^ n18817 ;
  assign n18821 = n18820 ^ n18819 ;
  assign n18823 = n18822 ^ n18821 ;
  assign n18838 = n18555 ^ n18379 ;
  assign n18825 = n7146 & n12143 ;
  assign n18824 = n7141 & ~n12142 ;
  assign n18826 = n18825 ^ n18824 ;
  assign n18827 = n18826 ^ n7129 ;
  assign n18828 = n18827 ^ x8 ;
  assign n18829 = n18826 ^ x8 ;
  assign n18833 = n18829 ^ n7130 ;
  assign n18834 = x7 & ~n14476 ;
  assign n18835 = n18833 & n18834 ;
  assign n18831 = n7130 & n12207 ;
  assign n18830 = n15500 & n18829 ;
  assign n18832 = n18831 ^ n18830 ;
  assign n18836 = n18835 ^ n18832 ;
  assign n18837 = ~n18828 & ~n18836 ;
  assign n18839 = n18838 ^ n18837 ;
  assign n19048 = n7146 & ~n12151 ;
  assign n19047 = n8054 & n12143 ;
  assign n19049 = n19048 ^ n19047 ;
  assign n19045 = n7141 & n12149 ;
  assign n19044 = n7135 & ~n14498 ;
  assign n19046 = n19045 ^ n19044 ;
  assign n19050 = n19049 ^ n19046 ;
  assign n18845 = n7146 & n12149 ;
  assign n18844 = n8054 & ~n12142 ;
  assign n18846 = n18845 ^ n18844 ;
  assign n18842 = n7141 & n12143 ;
  assign n18841 = n7135 & n14299 ;
  assign n18843 = n18842 ^ n18841 ;
  assign n18847 = n18846 ^ n18843 ;
  assign n19051 = n19050 ^ n18847 ;
  assign n19042 = n18549 ^ n18407 ;
  assign n19030 = n7146 & n12160 ;
  assign n19029 = n8054 & ~n12151 ;
  assign n19031 = n19030 ^ n19029 ;
  assign n19027 = n7141 & n12152 ;
  assign n19026 = n7135 & n15300 ;
  assign n19028 = n19027 ^ n19026 ;
  assign n19032 = n19031 ^ n19028 ;
  assign n19033 = n19032 ^ x8 ;
  assign n19013 = n18547 ^ n18419 ;
  assign n19034 = n19032 ^ n19013 ;
  assign n19020 = n7146 & n12152 ;
  assign n19019 = n8054 & n12149 ;
  assign n19021 = n19020 ^ n19019 ;
  assign n19017 = n7141 & ~n12151 ;
  assign n19016 = n7135 & ~n15312 ;
  assign n19018 = n19017 ^ n19016 ;
  assign n19022 = n19021 ^ n19018 ;
  assign n19035 = n19034 ^ n19022 ;
  assign n19036 = n19033 & ~n19035 ;
  assign n18857 = n18542 ^ n18528 ;
  assign n18855 = n7141 & n12160 ;
  assign n18853 = n7135 & ~n14581 ;
  assign n18850 = n7146 & n12163 ;
  assign n18849 = n8054 & n12152 ;
  assign n18851 = n18850 ^ n18849 ;
  assign n18852 = n18851 ^ x8 ;
  assign n18854 = n18853 ^ n18852 ;
  assign n18856 = n18855 ^ n18854 ;
  assign n18858 = n18857 ^ n18856 ;
  assign n18872 = n18509 ^ n18496 ;
  assign n18873 = n18499 & ~n18872 ;
  assign n18870 = n18518 ^ n18510 ;
  assign n18871 = n18870 ^ n18508 ;
  assign n18874 = n18873 ^ n18871 ;
  assign n18867 = n7141 & n12163 ;
  assign n18860 = n12160 ^ x8 ;
  assign n18861 = n18860 ^ x7 ;
  assign n18862 = n18861 ^ n12160 ;
  assign n18863 = ~n14866 & n18862 ;
  assign n18864 = n18863 ^ n12160 ;
  assign n18865 = n7128 & n18864 ;
  assign n18866 = n18865 ^ x8 ;
  assign n18868 = n18867 ^ n18866 ;
  assign n18859 = n7146 & n12167 ;
  assign n18869 = n18868 ^ n18859 ;
  assign n18875 = n18874 ^ n18869 ;
  assign n18883 = n7141 & n12167 ;
  assign n18881 = n7135 & ~n14890 ;
  assign n18878 = n7146 & n12168 ;
  assign n18877 = n8054 & n12163 ;
  assign n18879 = n18878 ^ n18877 ;
  assign n18880 = n18879 ^ x8 ;
  assign n18882 = n18881 ^ n18880 ;
  assign n18884 = n18883 ^ n18882 ;
  assign n19004 = n18884 ^ n18874 ;
  assign n18876 = n18509 ^ n18499 ;
  assign n18885 = n18884 ^ n18876 ;
  assign n18894 = n18494 ^ n18484 ;
  assign n18889 = n7146 & ~n12169 ;
  assign n18888 = n8054 & n12167 ;
  assign n18890 = n18889 ^ n18888 ;
  assign n18891 = n18890 ^ x8 ;
  assign n18887 = n7135 & ~n14915 ;
  assign n18892 = n18891 ^ n18887 ;
  assign n18886 = n7141 & n12168 ;
  assign n18893 = n18892 ^ n18886 ;
  assign n18895 = n18894 ^ n18893 ;
  assign n18904 = n18481 ^ n18463 ;
  assign n18902 = n7141 & ~n12169 ;
  assign n18900 = n7135 & ~n14949 ;
  assign n18897 = n7146 & n12175 ;
  assign n18896 = n8054 & n12168 ;
  assign n18898 = n18897 ^ n18896 ;
  assign n18899 = n18898 ^ x8 ;
  assign n18901 = n18900 ^ n18899 ;
  assign n18903 = n18902 ^ n18901 ;
  assign n18905 = n18904 ^ n18903 ;
  assign n18914 = n18452 ^ n18438 ;
  assign n18915 = n18914 ^ n18461 ;
  assign n18912 = n7141 & n12175 ;
  assign n18910 = n7135 & n15035 ;
  assign n18907 = n7146 & n12179 ;
  assign n18906 = n8054 & ~n12169 ;
  assign n18908 = n18907 ^ n18906 ;
  assign n18909 = n18908 ^ x8 ;
  assign n18911 = n18910 ^ n18909 ;
  assign n18913 = n18912 ^ n18911 ;
  assign n18916 = n18915 ^ n18913 ;
  assign n18971 = n7141 & n12179 ;
  assign n18964 = n12175 ^ x8 ;
  assign n18965 = n18964 ^ x7 ;
  assign n18966 = n18965 ^ n12175 ;
  assign n18967 = ~n15048 & n18966 ;
  assign n18968 = n18967 ^ n12175 ;
  assign n18969 = n7128 & n18968 ;
  assign n18970 = n18969 ^ x8 ;
  assign n18972 = n18971 ^ n18970 ;
  assign n18963 = n7146 & n12180 ;
  assign n18973 = n18972 ^ n18963 ;
  assign n18950 = n7141 & n12180 ;
  assign n18948 = n7135 & ~n15128 ;
  assign n18945 = n7146 & n12181 ;
  assign n18944 = n8054 & n12179 ;
  assign n18946 = n18945 ^ n18944 ;
  assign n18947 = n18946 ^ x8 ;
  assign n18949 = n18948 ^ n18947 ;
  assign n18951 = n18950 ^ n18949 ;
  assign n18917 = n6648 & ~n12183 ;
  assign n18918 = ~n12182 & ~n18156 ;
  assign n18919 = ~n12183 & ~n18156 ;
  assign n18920 = n7135 & n18440 ;
  assign n18926 = n8054 & n12181 ;
  assign n18923 = n7135 & n12181 ;
  assign n18924 = n18923 ^ n7146 ;
  assign n18925 = ~n12183 & n18924 ;
  assign n18927 = n18926 ^ n18925 ;
  assign n18928 = n18920 & ~n18927 ;
  assign n18929 = n18928 ^ n18927 ;
  assign n18930 = x8 & ~n18929 ;
  assign n18931 = ~n18919 & n18930 ;
  assign n18932 = ~n18918 & n18931 ;
  assign n18933 = ~n18917 & ~n18932 ;
  assign n18937 = n7146 & ~n12182 ;
  assign n18936 = n8054 & n12180 ;
  assign n18938 = n18937 ^ n18936 ;
  assign n18939 = n18938 ^ x8 ;
  assign n18935 = n7135 & ~n15151 ;
  assign n18940 = n18939 ^ n18935 ;
  assign n18934 = n7141 & n12181 ;
  assign n18941 = n18940 ^ n18934 ;
  assign n18942 = n18933 & n18941 ;
  assign n18943 = n18942 ^ n18941 ;
  assign n18952 = n18951 ^ n18943 ;
  assign n18957 = n18951 ^ n12182 ;
  assign n18956 = ~n6648 & ~n12182 ;
  assign n18958 = n18957 ^ n18956 ;
  assign n18955 = ~x9 & n18917 ;
  assign n18959 = n18958 ^ n18955 ;
  assign n18953 = x10 ^ x8 ;
  assign n18954 = ~n12183 & n18953 ;
  assign n18960 = n18959 ^ n18954 ;
  assign n18961 = n18952 & ~n18960 ;
  assign n18962 = n18961 ^ n18951 ;
  assign n18974 = n18973 ^ n18962 ;
  assign n18975 = n18439 & n18451 ;
  assign n18985 = n6656 & ~n12184 ;
  assign n18979 = n6657 ^ n6652 ;
  assign n18980 = n12182 ^ x11 ;
  assign n18981 = n18979 & ~n18980 ;
  assign n18982 = n18981 ^ n6650 ;
  assign n18983 = ~n12185 & n18982 ;
  assign n18976 = n18450 ^ n6650 ;
  assign n18977 = n18976 ^ n18962 ;
  assign n18984 = n18983 ^ n18977 ;
  assign n18986 = n18985 ^ n18984 ;
  assign n18987 = n18986 ^ n18962 ;
  assign n18988 = ~n18956 & ~n18987 ;
  assign n18989 = n18975 & n18988 ;
  assign n18990 = n18989 ^ n18986 ;
  assign n18991 = n18974 & ~n18990 ;
  assign n18992 = n18991 ^ n18973 ;
  assign n18993 = n18992 ^ n18913 ;
  assign n18994 = n18916 & n18993 ;
  assign n18995 = n18994 ^ n18913 ;
  assign n18996 = n18995 ^ n18903 ;
  assign n18997 = n18905 & n18996 ;
  assign n18998 = n18997 ^ n18903 ;
  assign n18999 = n18998 ^ n18893 ;
  assign n19000 = ~n18895 & n18999 ;
  assign n19001 = n19000 ^ n18893 ;
  assign n19002 = n19001 ^ n18884 ;
  assign n19003 = ~n18885 & n19002 ;
  assign n19005 = n19004 ^ n19003 ;
  assign n19006 = ~n18875 & ~n19005 ;
  assign n19007 = n19006 ^ n18874 ;
  assign n19008 = n19007 ^ n18856 ;
  assign n19009 = ~n18858 & ~n19008 ;
  assign n19010 = n19009 ^ n18856 ;
  assign n19011 = n18544 ^ n18437 ;
  assign n19012 = n19010 & ~n19011 ;
  assign n19014 = n19013 ^ n19012 ;
  assign n19015 = n19012 ^ x8 ;
  assign n19023 = n19022 ^ n19015 ;
  assign n19024 = n19014 & ~n19023 ;
  assign n19025 = n19024 ^ n19013 ;
  assign n19037 = n19011 ^ n19010 ;
  assign n19038 = n19037 ^ n19012 ;
  assign n19039 = ~n19025 & ~n19038 ;
  assign n19040 = n19036 & n19039 ;
  assign n19041 = n19040 ^ n19025 ;
  assign n19043 = n19042 ^ n19041 ;
  assign n19052 = n19051 ^ n19043 ;
  assign n19053 = n19052 ^ n19051 ;
  assign n19060 = n19050 ^ n19042 ;
  assign n19061 = n19060 ^ n19051 ;
  assign n18840 = n18552 ^ n18391 ;
  assign n18848 = n18847 ^ n18840 ;
  assign n19062 = n19061 ^ n18848 ;
  assign n19063 = n19062 ^ n19051 ;
  assign n19064 = n19053 & n19063 ;
  assign n19065 = n19064 ^ n19051 ;
  assign n19066 = x8 & ~n19065 ;
  assign n19054 = n19041 ^ n18847 ;
  assign n19055 = n19054 ^ n19051 ;
  assign n19056 = n19053 & n19055 ;
  assign n19057 = n19056 ^ n19051 ;
  assign n19058 = n18848 & n19057 ;
  assign n19059 = n19058 ^ n18847 ;
  assign n19067 = n19066 ^ n19059 ;
  assign n19068 = n19067 ^ n18837 ;
  assign n19069 = ~n18839 & ~n19068 ;
  assign n19070 = n19069 ^ n18837 ;
  assign n19071 = n19070 ^ n18821 ;
  assign n19072 = ~n18823 & ~n19071 ;
  assign n19073 = n19072 ^ n18821 ;
  assign n19074 = n19073 ^ n18811 ;
  assign n19075 = ~n18813 & n19074 ;
  assign n19076 = n19075 ^ n18811 ;
  assign n19077 = n19076 ^ n18798 ;
  assign n19078 = ~n18800 & n19077 ;
  assign n19079 = n19078 ^ n18798 ;
  assign n19080 = n19079 ^ n18788 ;
  assign n19081 = ~n18790 & ~n19080 ;
  assign n19082 = n19081 ^ n18788 ;
  assign n19083 = n19082 ^ n18772 ;
  assign n19084 = ~n18774 & ~n19083 ;
  assign n19085 = n19084 ^ n18772 ;
  assign n19086 = n19085 ^ n18760 ;
  assign n19087 = ~n18761 & ~n19086 ;
  assign n19088 = n19087 ^ n18760 ;
  assign n19089 = n19088 ^ n18743 ;
  assign n19090 = n18745 & ~n19089 ;
  assign n19091 = n19090 ^ n18743 ;
  assign n19092 = n19091 ^ n18730 ;
  assign n19093 = n18732 & n19092 ;
  assign n19094 = n19093 ^ n18730 ;
  assign n19095 = n19094 ^ n18720 ;
  assign n19096 = n18722 & n19095 ;
  assign n19097 = n19096 ^ n18720 ;
  assign n19098 = n19097 ^ n18710 ;
  assign n19099 = n18712 & n19098 ;
  assign n19100 = n19099 ^ n18710 ;
  assign n19101 = n19100 ^ n18696 ;
  assign n19102 = ~n18702 & ~n19101 ;
  assign n19103 = n19102 ^ n18696 ;
  assign n19104 = n19103 ^ n18684 ;
  assign n19105 = n18692 & ~n19104 ;
  assign n19106 = n19105 ^ n18684 ;
  assign n19107 = n19106 ^ n18680 ;
  assign n19108 = n18682 & ~n19107 ;
  assign n19109 = n19108 ^ n18680 ;
  assign n19111 = n19110 ^ n19109 ;
  assign n19118 = n7135 & n12376 ;
  assign n19116 = n7146 & n12260 ;
  assign n19114 = n8054 & ~n12108 ;
  assign n19113 = n19110 ^ x8 ;
  assign n19115 = n19114 ^ n19113 ;
  assign n19117 = n19116 ^ n19115 ;
  assign n19119 = n19118 ^ n19117 ;
  assign n19112 = n7141 & n11972 ;
  assign n19120 = n19119 ^ n19112 ;
  assign n19121 = ~n19111 & n19120 ;
  assign n19122 = n19121 ^ n19110 ;
  assign n19123 = n19122 ^ n18659 ;
  assign n19124 = n18661 & n19123 ;
  assign n19125 = n19124 ^ n18659 ;
  assign n19126 = n19125 ^ n18640 ;
  assign n19127 = ~n18648 & ~n19126 ;
  assign n19128 = n19127 ^ n18640 ;
  assign n19655 = n19139 ^ n19128 ;
  assign n19656 = n19655 ^ x5 ;
  assign n19654 = n10131 & n12971 ;
  assign n19657 = n19656 ^ n19654 ;
  assign n19653 = n9085 & n12755 ;
  assign n19658 = n19657 ^ n19653 ;
  assign n19660 = n19659 ^ n19658 ;
  assign n19652 = ~n9092 & ~n12705 ;
  assign n19661 = n19660 ^ n19652 ;
  assign n19171 = n19125 ^ n18648 ;
  assign n19154 = ~n9092 & n12656 ;
  assign n19153 = n9085 & ~n12705 ;
  assign n19155 = n19154 ^ n19153 ;
  assign n9079 = x5 & ~n9077 ;
  assign n19156 = n19155 ^ n9079 ;
  assign n19158 = n25052 ^ n9077 ;
  assign n19157 = n19155 ^ x5 ;
  assign n19159 = n19158 ^ n19157 ;
  assign n19165 = ~x4 & n19159 ;
  assign n19166 = n19165 ^ n19158 ;
  assign n19167 = ~n12724 & n19166 ;
  assign n19168 = n19167 ^ n19158 ;
  assign n19160 = ~n12755 & n19159 ;
  assign n19169 = n19168 ^ n19160 ;
  assign n19170 = ~n19156 & ~n19169 ;
  assign n19172 = n19171 ^ n19170 ;
  assign n19180 = n9081 & n12706 ;
  assign n19176 = n19122 ^ n18661 ;
  assign n19177 = n19176 ^ x5 ;
  assign n19175 = n10131 & ~n12705 ;
  assign n19178 = n19177 ^ n19175 ;
  assign n19174 = n9085 & n12656 ;
  assign n19179 = n19178 ^ n19174 ;
  assign n19181 = n19180 ^ n19179 ;
  assign n19173 = ~n9092 & ~n12613 ;
  assign n19182 = n19181 ^ n19173 ;
  assign n19631 = n19120 ^ n19109 ;
  assign n19191 = ~n9092 & ~n12108 ;
  assign n19188 = n9085 & ~n12367 ;
  assign n19186 = n10131 & ~n12613 ;
  assign n19184 = n19106 ^ n18682 ;
  assign n19185 = n19184 ^ x5 ;
  assign n19187 = n19186 ^ n19185 ;
  assign n19189 = n19188 ^ n19187 ;
  assign n19183 = n9081 & n13110 ;
  assign n19190 = n19189 ^ n19183 ;
  assign n19192 = n19191 ^ n19190 ;
  assign n19201 = n19103 ^ n18692 ;
  assign n19196 = n9085 & ~n12108 ;
  assign n19195 = n10131 & ~n12367 ;
  assign n19197 = n19196 ^ n19195 ;
  assign n19198 = n19197 ^ x5 ;
  assign n19194 = n9081 & n12368 ;
  assign n19199 = n19198 ^ n19194 ;
  assign n19193 = ~n9092 & n11972 ;
  assign n19200 = n19199 ^ n19193 ;
  assign n19202 = n19201 ^ n19200 ;
  assign n19210 = n9081 & n12376 ;
  assign n19206 = n19100 ^ n18702 ;
  assign n19207 = n19206 ^ x5 ;
  assign n19205 = n10131 & ~n12108 ;
  assign n19208 = n19207 ^ n19205 ;
  assign n19204 = n9085 & n11972 ;
  assign n19209 = n19208 ^ n19204 ;
  assign n19211 = n19210 ^ n19209 ;
  assign n19203 = ~n9092 & n12260 ;
  assign n19212 = n19211 ^ n19203 ;
  assign n19221 = n19097 ^ n18712 ;
  assign n19219 = ~n9092 & ~n12256 ;
  assign n19217 = n9081 & ~n14078 ;
  assign n19214 = n9085 & n12260 ;
  assign n19213 = n10131 & n11972 ;
  assign n19215 = n19214 ^ n19213 ;
  assign n19216 = n19215 ^ x5 ;
  assign n19218 = n19217 ^ n19216 ;
  assign n19220 = n19219 ^ n19218 ;
  assign n19222 = n19221 ^ n19220 ;
  assign n19606 = n19094 ^ n18722 ;
  assign n19593 = n19091 ^ n18732 ;
  assign n19228 = n9085 & ~n12220 ;
  assign n19227 = n10131 & ~n12262 ;
  assign n19229 = n19228 ^ n19227 ;
  assign n19225 = ~n9092 & ~n12110 ;
  assign n19224 = n9081 & n13712 ;
  assign n19226 = n19225 ^ n19224 ;
  assign n19230 = n19229 ^ n19226 ;
  assign n19231 = n19230 ^ x5 ;
  assign n19223 = n19088 ^ n18745 ;
  assign n19232 = n19231 ^ n19223 ;
  assign n19242 = n19082 ^ n18774 ;
  assign n19240 = ~n9092 & n12121 ;
  assign n19238 = n9081 & n13196 ;
  assign n19235 = n9085 & n12117 ;
  assign n19234 = n10131 & ~n12110 ;
  assign n19236 = n19235 ^ n19234 ;
  assign n19237 = n19236 ^ x5 ;
  assign n19239 = n19238 ^ n19237 ;
  assign n19241 = n19240 ^ n19239 ;
  assign n19243 = n19242 ^ n19241 ;
  assign n19252 = n19079 ^ n18790 ;
  assign n19247 = n9085 & n12121 ;
  assign n19246 = n10131 & n12117 ;
  assign n19248 = n19247 ^ n19246 ;
  assign n19249 = n19248 ^ x5 ;
  assign n19245 = n9081 & ~n13596 ;
  assign n19250 = n19249 ^ n19245 ;
  assign n19244 = ~n9092 & ~n12129 ;
  assign n19251 = n19250 ^ n19244 ;
  assign n19253 = n19252 ^ n19251 ;
  assign n19263 = n9085 & ~n12129 ;
  assign n19261 = ~n9092 & n12130 ;
  assign n19259 = n19076 ^ n18800 ;
  assign n19260 = n19259 ^ x5 ;
  assign n19262 = n19261 ^ n19260 ;
  assign n19264 = n19263 ^ n19262 ;
  assign n19254 = n12121 ^ n9089 ;
  assign n19255 = n19254 ^ n12121 ;
  assign n19256 = ~n13605 & n19255 ;
  assign n19257 = n19256 ^ n12121 ;
  assign n19258 = n9077 & n19257 ;
  assign n19265 = n19264 ^ n19258 ;
  assign n19277 = n19073 ^ n18813 ;
  assign n19274 = n9085 & n12130 ;
  assign n19267 = n12129 ^ x5 ;
  assign n19268 = n19267 ^ x4 ;
  assign n19269 = n19268 ^ n12129 ;
  assign n19270 = ~n14271 & n19269 ;
  assign n19271 = n19270 ^ n12129 ;
  assign n19272 = n9077 & ~n19271 ;
  assign n19273 = n19272 ^ x5 ;
  assign n19275 = n19274 ^ n19273 ;
  assign n19266 = ~n9092 & ~n12136 ;
  assign n19276 = n19275 ^ n19266 ;
  assign n19278 = n19277 ^ n19276 ;
  assign n19287 = n19070 ^ n18823 ;
  assign n19285 = ~n9092 & n12137 ;
  assign n19283 = n9081 & ~n13818 ;
  assign n19280 = n9085 & ~n12136 ;
  assign n19279 = n10131 & n12130 ;
  assign n19281 = n19280 ^ n19279 ;
  assign n19282 = n19281 ^ x5 ;
  assign n19284 = n19283 ^ n19282 ;
  assign n19286 = n19285 ^ n19284 ;
  assign n19288 = n19287 ^ n19286 ;
  assign n19297 = n19067 ^ n18839 ;
  assign n19292 = n9085 & n12137 ;
  assign n19291 = n10131 & ~n12136 ;
  assign n19293 = n19292 ^ n19291 ;
  assign n19294 = n19293 ^ x5 ;
  assign n19290 = n9081 & n14129 ;
  assign n19295 = n19294 ^ n19290 ;
  assign n19289 = ~n9092 & ~n12138 ;
  assign n19296 = n19295 ^ n19289 ;
  assign n19298 = n19297 ^ n19296 ;
  assign n19551 = ~n9092 & n12207 ;
  assign n19549 = n9081 & ~n13939 ;
  assign n19546 = n9085 & ~n12138 ;
  assign n19545 = n10131 & n12137 ;
  assign n19547 = n19546 ^ n19545 ;
  assign n19548 = n19547 ^ x5 ;
  assign n19550 = n19549 ^ n19548 ;
  assign n19552 = n19551 ^ n19550 ;
  assign n19307 = n19060 ^ x8 ;
  assign n19308 = n19307 ^ n19041 ;
  assign n19305 = ~n9092 & ~n12142 ;
  assign n19303 = n9081 & n14832 ;
  assign n19300 = n9085 & n12207 ;
  assign n19299 = n10131 & ~n12138 ;
  assign n19301 = n19300 ^ n19299 ;
  assign n19302 = n19301 ^ x5 ;
  assign n19304 = n19303 ^ n19302 ;
  assign n19306 = n19305 ^ n19304 ;
  assign n19309 = n19308 ^ n19306 ;
  assign n19530 = n9085 & ~n12142 ;
  assign n19529 = n10131 & n12207 ;
  assign n19531 = n19530 ^ n19529 ;
  assign n19532 = n19531 ^ x5 ;
  assign n19528 = n9081 & ~n15500 ;
  assign n19533 = n19532 ^ n19528 ;
  assign n19527 = ~n9092 & n12143 ;
  assign n19534 = n19533 ^ n19527 ;
  assign n19318 = n19037 ^ n19033 ;
  assign n19313 = n9085 & n12143 ;
  assign n19312 = n10131 & ~n12142 ;
  assign n19314 = n19313 ^ n19312 ;
  assign n19315 = n19314 ^ x5 ;
  assign n19311 = n9081 & n14299 ;
  assign n19316 = n19315 ^ n19311 ;
  assign n19310 = ~n9092 & n12149 ;
  assign n19317 = n19316 ^ n19310 ;
  assign n19319 = n19318 ^ n19317 ;
  assign n19328 = n19007 ^ n18858 ;
  assign n19323 = n9085 & n12149 ;
  assign n19322 = n10131 & n12143 ;
  assign n19324 = n19323 ^ n19322 ;
  assign n19325 = n19324 ^ x5 ;
  assign n19321 = n9081 & ~n14498 ;
  assign n19326 = n19325 ^ n19321 ;
  assign n19320 = ~n9092 & ~n12151 ;
  assign n19327 = n19326 ^ n19320 ;
  assign n19329 = n19328 ^ n19327 ;
  assign n19338 = n19005 ^ n18869 ;
  assign n19333 = n9085 & ~n12151 ;
  assign n19332 = n10131 & n12149 ;
  assign n19334 = n19333 ^ n19332 ;
  assign n19335 = n19334 ^ x5 ;
  assign n19331 = n9081 & ~n15312 ;
  assign n19336 = n19335 ^ n19331 ;
  assign n19330 = ~n9092 & n12152 ;
  assign n19337 = n19336 ^ n19330 ;
  assign n19339 = n19338 ^ n19337 ;
  assign n19348 = n19001 ^ n18885 ;
  assign n19346 = ~n9092 & n12160 ;
  assign n19344 = n9081 & n15300 ;
  assign n19341 = n9085 & n12152 ;
  assign n19340 = n10131 & ~n12151 ;
  assign n19342 = n19341 ^ n19340 ;
  assign n19343 = n19342 ^ x5 ;
  assign n19345 = n19344 ^ n19343 ;
  assign n19347 = n19346 ^ n19345 ;
  assign n19349 = n19348 ^ n19347 ;
  assign n19358 = n18998 ^ n18895 ;
  assign n19356 = ~n9092 & n12163 ;
  assign n19354 = n9081 & ~n14581 ;
  assign n19351 = n10131 & n12152 ;
  assign n19350 = n9085 & n12160 ;
  assign n19352 = n19351 ^ n19350 ;
  assign n19353 = n19352 ^ x5 ;
  assign n19355 = n19354 ^ n19353 ;
  assign n19357 = n19356 ^ n19355 ;
  assign n19359 = n19358 ^ n19357 ;
  assign n19499 = n18995 ^ n18905 ;
  assign n19360 = n18992 ^ n18916 ;
  assign n19365 = n9085 & n12167 ;
  assign n19364 = n10131 & n12163 ;
  assign n19366 = n19365 ^ n19364 ;
  assign n19362 = ~n9092 & n12168 ;
  assign n19361 = n9081 & ~n14890 ;
  assign n19363 = n19362 ^ n19361 ;
  assign n19367 = n19366 ^ n19363 ;
  assign n19368 = n19360 & ~n19367 ;
  assign n19379 = n19368 ^ n19360 ;
  assign n19492 = ~x5 & ~n19379 ;
  assign n19390 = n18960 ^ n18943 ;
  assign n19388 = ~n9092 & n12175 ;
  assign n19386 = n9081 & ~n14949 ;
  assign n19383 = n9085 & ~n12169 ;
  assign n19382 = n10131 & n12168 ;
  assign n19384 = n19383 ^ n19382 ;
  assign n19385 = n19384 ^ x5 ;
  assign n19387 = n19386 ^ n19385 ;
  assign n19389 = n19388 ^ n19387 ;
  assign n19391 = n19390 ^ n19389 ;
  assign n19400 = n18932 ^ n18917 ;
  assign n19401 = n19400 ^ n18941 ;
  assign n19398 = ~n9092 & n12179 ;
  assign n19396 = n9081 & n15035 ;
  assign n19393 = n10131 & ~n12169 ;
  assign n19392 = n9085 & n12175 ;
  assign n19394 = n19393 ^ n19392 ;
  assign n19395 = n19394 ^ x5 ;
  assign n19397 = n19396 ^ n19395 ;
  assign n19399 = n19398 ^ n19397 ;
  assign n19402 = n19401 ^ n19399 ;
  assign n19425 = n9085 & n12179 ;
  assign n19424 = n10131 & n12175 ;
  assign n19426 = n19425 ^ n19424 ;
  assign n19427 = n19426 ^ x5 ;
  assign n19423 = n9081 & ~n15049 ;
  assign n19428 = n19427 ^ n19423 ;
  assign n19422 = ~n9092 & n12180 ;
  assign n19429 = n19428 ^ n19422 ;
  assign n19409 = n13899 ^ n7130 ;
  assign n19410 = ~n12182 & n19409 ;
  assign n19403 = n18919 ^ n7128 ;
  assign n19404 = n18919 ^ n12182 ;
  assign n19405 = n19404 ^ n18919 ;
  assign n19406 = n19403 & ~n19405 ;
  assign n19407 = n19406 ^ n18919 ;
  assign n19408 = n18930 & n19407 ;
  assign n19411 = n19410 ^ n19408 ;
  assign n19414 = n7141 ^ n7129 ;
  assign n19417 = n12182 & n19414 ;
  assign n19418 = n19417 ^ n7141 ;
  assign n19419 = n12183 & n19418 ;
  assign n19412 = n18929 ^ n7129 ;
  assign n19420 = n19419 ^ n19412 ;
  assign n19421 = ~n19411 & ~n19420 ;
  assign n19430 = n19429 ^ n19421 ;
  assign n19462 = n7128 & n12183 ;
  assign n19463 = n19462 ^ n7128 ;
  assign n19466 = x5 & n19463 ;
  assign n19446 = n9077 & ~n12182 ;
  assign n19447 = x5 & ~n19446 ;
  assign n19448 = ~n12183 & n19447 ;
  assign n19449 = ~n18627 & n19448 ;
  assign n19450 = n19449 ^ n19447 ;
  assign n19457 = n9081 & n12185 ;
  assign n19456 = ~n9092 & ~n12183 ;
  assign n19458 = n19457 ^ n19456 ;
  assign n19454 = n9085 & ~n12182 ;
  assign n19453 = n9077 & n12181 ;
  assign n19455 = n19454 ^ n19453 ;
  assign n19459 = n19458 ^ n19455 ;
  assign n19460 = n19450 & ~n19459 ;
  assign n19443 = n9085 & n12181 ;
  assign n19442 = n10131 & n12180 ;
  assign n19444 = n19443 ^ n19442 ;
  assign n19440 = ~n9092 & ~n12182 ;
  assign n19439 = n9081 & ~n15151 ;
  assign n19441 = n19440 ^ n19439 ;
  assign n19445 = n19444 ^ n19441 ;
  assign n19461 = n19460 ^ n19445 ;
  assign n19464 = n19463 ^ n19460 ;
  assign n19465 = n19461 & n19464 ;
  assign n19467 = n19466 ^ n19465 ;
  assign n19437 = ~n9092 & n12181 ;
  assign n19435 = n9081 & ~n15128 ;
  assign n19432 = n9085 & n12180 ;
  assign n19431 = n10131 & n12179 ;
  assign n19433 = n19432 ^ n19431 ;
  assign n19434 = n19433 ^ x5 ;
  assign n19436 = n19435 ^ n19434 ;
  assign n19438 = n19437 ^ n19436 ;
  assign n19468 = n19467 ^ n19438 ;
  assign n19472 = n19466 ^ n19438 ;
  assign n19470 = x7 ^ x5 ;
  assign n19471 = ~n12183 & n19470 ;
  assign n19473 = n19472 ^ n19471 ;
  assign n19469 = n7128 & ~n12182 ;
  assign n19474 = n19473 ^ n19469 ;
  assign n19475 = n19468 & ~n19474 ;
  assign n19476 = n19475 ^ n19467 ;
  assign n19477 = n19476 ^ n19421 ;
  assign n19478 = ~n19430 & n19477 ;
  assign n19479 = n19478 ^ n19429 ;
  assign n19480 = n19479 ^ n19399 ;
  assign n19481 = n19402 & ~n19480 ;
  assign n19482 = n19481 ^ n19401 ;
  assign n19483 = n19482 ^ n19389 ;
  assign n19484 = ~n19391 & n19483 ;
  assign n19485 = n19484 ^ n19389 ;
  assign n19370 = n18990 ^ n18973 ;
  assign n19375 = n9085 & n12168 ;
  assign n19374 = n10131 & n12167 ;
  assign n19376 = n19375 ^ n19374 ;
  assign n19372 = ~n9092 & ~n12169 ;
  assign n19371 = n9081 & ~n14915 ;
  assign n19373 = n19372 ^ n19371 ;
  assign n19377 = n19376 ^ n19373 ;
  assign n19486 = n19377 ^ x5 ;
  assign n19487 = n19370 & n19486 ;
  assign n19488 = ~n19485 & n19487 ;
  assign n19489 = n19488 ^ n19485 ;
  assign n19378 = ~n19370 & n19377 ;
  assign n19493 = n19378 ^ n19370 ;
  assign n19380 = n19379 ^ n19367 ;
  assign n19494 = n19380 ^ n19360 ;
  assign n19495 = n19493 & n19494 ;
  assign n19496 = n19489 & n19495 ;
  assign n19497 = n19492 & ~n19496 ;
  assign n19369 = x5 & ~n19368 ;
  assign n19381 = ~n19378 & ~n19380 ;
  assign n19490 = n19381 & n19489 ;
  assign n19491 = n19369 & ~n19490 ;
  assign n19498 = n19497 ^ n19491 ;
  assign n19500 = n19499 ^ n19498 ;
  assign n19504 = n9085 & n12163 ;
  assign n19503 = n10131 & n12160 ;
  assign n19505 = n19504 ^ n19503 ;
  assign n19506 = n19505 ^ x5 ;
  assign n19502 = n9081 & ~n14867 ;
  assign n19507 = n19506 ^ n19502 ;
  assign n19501 = ~n9092 & n12167 ;
  assign n19508 = n19507 ^ n19501 ;
  assign n19509 = n19508 ^ n19498 ;
  assign n19510 = ~n19500 & n19509 ;
  assign n19511 = n19510 ^ n19499 ;
  assign n19512 = n19511 ^ n19357 ;
  assign n19513 = ~n19359 & ~n19512 ;
  assign n19514 = n19513 ^ n19358 ;
  assign n19515 = n19514 ^ n19347 ;
  assign n19516 = ~n19349 & ~n19515 ;
  assign n19517 = n19516 ^ n19347 ;
  assign n19518 = n19517 ^ n19337 ;
  assign n19519 = ~n19339 & ~n19518 ;
  assign n19520 = n19519 ^ n19338 ;
  assign n19521 = n19520 ^ n19327 ;
  assign n19522 = n19329 & n19521 ;
  assign n19523 = n19522 ^ n19328 ;
  assign n19524 = n19523 ^ n19317 ;
  assign n19525 = ~n19319 & n19524 ;
  assign n19526 = n19525 ^ n19317 ;
  assign n19535 = n19534 ^ n19526 ;
  assign n19537 = n19033 ^ n19011 ;
  assign n19538 = n19037 & ~n19537 ;
  assign n19536 = n19534 ^ n19035 ;
  assign n19539 = n19538 ^ n19536 ;
  assign n19540 = n19535 & n19539 ;
  assign n19541 = n19540 ^ n19534 ;
  assign n19542 = n19541 ^ n19306 ;
  assign n19543 = ~n19309 & n19542 ;
  assign n19544 = n19543 ^ n19306 ;
  assign n19553 = n19552 ^ n19544 ;
  assign n19556 = n19043 & ~n19307 ;
  assign n19554 = n19050 ^ n18848 ;
  assign n19555 = n19554 ^ n19552 ;
  assign n19557 = n19556 ^ n19555 ;
  assign n19558 = n19553 & n19557 ;
  assign n19559 = n19558 ^ n19552 ;
  assign n19560 = n19559 ^ n19296 ;
  assign n19561 = ~n19298 & n19560 ;
  assign n19562 = n19561 ^ n19296 ;
  assign n19563 = n19562 ^ n19286 ;
  assign n19564 = n19288 & n19563 ;
  assign n19565 = n19564 ^ n19286 ;
  assign n19566 = n19565 ^ n19276 ;
  assign n19567 = ~n19278 & ~n19566 ;
  assign n19568 = n19567 ^ n19277 ;
  assign n19569 = n19568 ^ n19259 ;
  assign n19570 = ~n19265 & n19569 ;
  assign n19571 = n19570 ^ n19259 ;
  assign n19572 = n19571 ^ n19251 ;
  assign n19573 = ~n19253 & ~n19572 ;
  assign n19574 = n19573 ^ n19251 ;
  assign n19575 = n19574 ^ n19241 ;
  assign n19576 = n19243 & n19575 ;
  assign n19577 = n19576 ^ n19241 ;
  assign n19589 = n19577 ^ n19223 ;
  assign n19233 = n19085 ^ n18761 ;
  assign n19578 = n19577 ^ n19233 ;
  assign n19585 = n9081 & n14047 ;
  assign n19583 = n9085 & ~n12110 ;
  assign n19581 = n10131 & ~n12220 ;
  assign n19580 = n19233 ^ x5 ;
  assign n19582 = n19581 ^ n19580 ;
  assign n19584 = n19583 ^ n19582 ;
  assign n19586 = n19585 ^ n19584 ;
  assign n19579 = ~n9092 & n12117 ;
  assign n19587 = n19586 ^ n19579 ;
  assign n19588 = ~n19578 & n19587 ;
  assign n19590 = n19589 ^ n19588 ;
  assign n19591 = ~n19232 & n19590 ;
  assign n19592 = n19591 ^ n19231 ;
  assign n19594 = n19593 ^ n19592 ;
  assign n19599 = n9085 & ~n12262 ;
  assign n19598 = n10131 & ~n12256 ;
  assign n19600 = n19599 ^ n19598 ;
  assign n19596 = ~n9092 & ~n12220 ;
  assign n19595 = n9081 & ~n13283 ;
  assign n19597 = n19596 ^ n19595 ;
  assign n19601 = n19600 ^ n19597 ;
  assign n19602 = n19601 ^ x5 ;
  assign n19603 = n19602 ^ n19592 ;
  assign n19604 = n19594 & ~n19603 ;
  assign n19605 = n19604 ^ n19593 ;
  assign n19607 = n19606 ^ n19605 ;
  assign n19614 = n9081 & n13054 ;
  assign n19612 = n9085 & ~n12256 ;
  assign n19610 = n10131 & n12260 ;
  assign n19609 = n19606 ^ x5 ;
  assign n19611 = n19610 ^ n19609 ;
  assign n19613 = n19612 ^ n19611 ;
  assign n19615 = n19614 ^ n19613 ;
  assign n19608 = ~n9092 & ~n12262 ;
  assign n19616 = n19615 ^ n19608 ;
  assign n19617 = n19607 & n19616 ;
  assign n19618 = n19617 ^ n19606 ;
  assign n19619 = n19618 ^ n19220 ;
  assign n19620 = n19222 & ~n19619 ;
  assign n19621 = n19620 ^ n19221 ;
  assign n19622 = n19621 ^ n19206 ;
  assign n19623 = ~n19212 & ~n19622 ;
  assign n19624 = n19623 ^ n19206 ;
  assign n19625 = n19624 ^ n19200 ;
  assign n19626 = ~n19202 & n19625 ;
  assign n19627 = n19626 ^ n19201 ;
  assign n19628 = n19627 ^ n19184 ;
  assign n19629 = n19192 & ~n19628 ;
  assign n19630 = n19629 ^ n19184 ;
  assign n19632 = n19631 ^ n19630 ;
  assign n19640 = n19631 ^ x5 ;
  assign n19639 = n9085 & ~n12613 ;
  assign n19641 = n19640 ^ n19639 ;
  assign n19638 = ~n9092 & ~n12367 ;
  assign n19642 = n19641 ^ n19638 ;
  assign n19633 = n12656 ^ n9089 ;
  assign n19634 = n19633 ^ n12656 ;
  assign n19635 = ~n12871 & n19634 ;
  assign n19636 = n19635 ^ n12656 ;
  assign n19637 = n9077 & n19636 ;
  assign n19643 = n19642 ^ n19637 ;
  assign n19644 = ~n19632 & ~n19643 ;
  assign n19645 = n19644 ^ n19631 ;
  assign n19646 = n19645 ^ n19176 ;
  assign n19647 = n19182 & ~n19646 ;
  assign n19648 = n19647 ^ n19176 ;
  assign n19649 = n19648 ^ n19171 ;
  assign n19650 = n19172 & ~n19649 ;
  assign n19651 = n19650 ^ n19171 ;
  assign n19662 = n19661 ^ n19651 ;
  assign n19663 = n19662 ^ n14315 ;
  assign n19665 = n19664 ^ n19663 ;
  assign n19672 = n12855 ^ x2 ;
  assign n19667 = n10828 & n14221 ;
  assign n19668 = n19667 ^ x1 ;
  assign n19673 = n19672 ^ n19668 ;
  assign n19674 = n19673 ^ n19668 ;
  assign n19675 = n19674 ^ n12855 ;
  assign n19676 = n12971 & n19675 ;
  assign n19677 = n19676 ^ n12855 ;
  assign n19678 = ~x1 & ~n19677 ;
  assign n19679 = n19678 ^ n19673 ;
  assign n19680 = ~x0 & n19679 ;
  assign n19666 = n19648 ^ n19172 ;
  assign n19669 = n19668 ^ n19666 ;
  assign n19681 = n19680 ^ n19669 ;
  assign n19698 = n19645 ^ n19182 ;
  assign n19682 = n12971 ^ n12755 ;
  assign n19683 = n19682 ^ n12971 ;
  assign n19688 = n12971 ^ x2 ;
  assign n19691 = n19688 ^ n12971 ;
  assign n19692 = n19683 & n19691 ;
  assign n19693 = n19692 ^ n12971 ;
  assign n19694 = ~x1 & n19693 ;
  assign n19684 = n19672 ^ x1 ;
  assign n19685 = ~n12855 & ~n13007 ;
  assign n19686 = n19684 & n19685 ;
  assign n19687 = n19686 ^ n19672 ;
  assign n19689 = n19688 ^ n19687 ;
  assign n19695 = n19694 ^ n19689 ;
  assign n19696 = ~x0 & ~n19695 ;
  assign n19697 = n19696 ^ n19687 ;
  assign n19699 = n19698 ^ n19697 ;
  assign n20481 = n10828 & ~n12918 ;
  assign n20482 = n20481 ^ n12971 ;
  assign n20483 = n20482 ^ n12755 ;
  assign n20484 = n20483 ^ n20482 ;
  assign n20485 = n20484 ^ n12705 ;
  assign n20486 = n20485 ^ n20484 ;
  assign n20489 = x2 & ~n20486 ;
  assign n20490 = n20489 ^ n20484 ;
  assign n20491 = ~x1 & n20490 ;
  assign n20492 = n20491 ^ n20483 ;
  assign n20493 = ~x0 & n20492 ;
  assign n20494 = n20493 ^ n20482 ;
  assign n19712 = n12656 ^ x2 ;
  assign n19715 = n19712 ^ n12656 ;
  assign n19716 = ~n19711 & n19715 ;
  assign n19717 = n19716 ^ n12656 ;
  assign n19718 = ~x1 & n19717 ;
  assign n19706 = n12705 ^ x1 ;
  assign n19705 = n12705 ^ x2 ;
  assign n19707 = n19706 ^ n19705 ;
  assign n19708 = n12663 & n19707 ;
  assign n19709 = n19708 ^ n19706 ;
  assign n19713 = n19712 ^ n19709 ;
  assign n19719 = n19718 ^ n19713 ;
  assign n19720 = ~x0 & ~n19719 ;
  assign n19721 = n19720 ^ n19709 ;
  assign n19738 = n19621 ^ n19212 ;
  assign n19726 = n12613 ^ n12367 ;
  assign n19727 = n19726 ^ n12613 ;
  assign n19728 = n12613 ^ x2 ;
  assign n19731 = n19728 ^ n12613 ;
  assign n19732 = ~n19727 & n19731 ;
  assign n19733 = n19732 ^ n12613 ;
  assign n19734 = ~x1 & ~n19733 ;
  assign n19722 = n12656 ^ x1 ;
  assign n19723 = n19722 ^ n19712 ;
  assign n19724 = n12871 & n19723 ;
  assign n19725 = n19724 ^ n19722 ;
  assign n19729 = n19728 ^ n19725 ;
  assign n19735 = n19734 ^ n19729 ;
  assign n19736 = ~x0 & ~n19735 ;
  assign n19737 = n19736 ^ n19725 ;
  assign n19739 = n19738 ^ n19737 ;
  assign n19745 = n16351 ^ n12367 ;
  assign n19746 = n12367 ^ x2 ;
  assign n19749 = n19746 ^ n12367 ;
  assign n19750 = ~n19745 & n19749 ;
  assign n19751 = n19750 ^ n12367 ;
  assign n19752 = ~x1 & ~n19751 ;
  assign n19741 = n12613 ^ x1 ;
  assign n19742 = n19741 ^ n19728 ;
  assign n19743 = n12777 & n19742 ;
  assign n19744 = n19743 ^ n19741 ;
  assign n19747 = n19746 ^ n19744 ;
  assign n19753 = n19752 ^ n19747 ;
  assign n19754 = ~x0 & n19753 ;
  assign n19755 = n19754 ^ n19744 ;
  assign n20427 = n19755 ^ n19737 ;
  assign n19740 = n19618 ^ n19222 ;
  assign n19756 = n19755 ^ n19740 ;
  assign n19773 = n19616 ^ n19605 ;
  assign n19761 = n12108 ^ n11972 ;
  assign n19762 = n19761 ^ n12108 ;
  assign n19763 = n12108 ^ x2 ;
  assign n19766 = n19763 ^ n12108 ;
  assign n19767 = n19762 & n19766 ;
  assign n19768 = n19767 ^ n12108 ;
  assign n19769 = ~x1 & ~n19768 ;
  assign n19757 = n12367 ^ x1 ;
  assign n19758 = n19757 ^ n19746 ;
  assign n19759 = n12277 & n19758 ;
  assign n19760 = n19759 ^ n19757 ;
  assign n19764 = n19763 ^ n19760 ;
  assign n19770 = n19769 ^ n19764 ;
  assign n19771 = ~x0 & n19770 ;
  assign n19772 = n19771 ^ n19760 ;
  assign n19774 = n19773 ^ n19772 ;
  assign n19792 = n19601 ^ n19593 ;
  assign n19791 = n19591 ^ n19230 ;
  assign n19793 = n19792 ^ n19791 ;
  assign n19777 = n12108 ^ x1 ;
  assign n19778 = n19777 ^ n19763 ;
  assign n19779 = n12375 & n19778 ;
  assign n19780 = n19779 ^ n19777 ;
  assign n19794 = n19793 ^ n19780 ;
  assign n19781 = n11972 ^ x2 ;
  assign n19784 = n19781 ^ n11972 ;
  assign n19785 = n12260 & n19784 ;
  assign n19786 = n19785 ^ n11972 ;
  assign n19787 = ~x1 & n19786 ;
  assign n19782 = n19781 ^ n19780 ;
  assign n19788 = n19787 ^ n19782 ;
  assign n19789 = ~x0 & ~n19788 ;
  assign n19795 = n19794 ^ n19789 ;
  assign n20404 = n12261 ^ n12260 ;
  assign n20400 = n11972 ^ x1 ;
  assign n20401 = n20400 ^ n19781 ;
  assign n20402 = n12270 & n20401 ;
  assign n20403 = n20402 ^ n20400 ;
  assign n20382 = n12260 ^ x2 ;
  assign n20405 = n20403 ^ n20382 ;
  assign n20406 = n20405 ^ n20403 ;
  assign n20407 = n20406 ^ n12260 ;
  assign n20408 = ~n20404 & n20407 ;
  assign n20409 = n20408 ^ n12260 ;
  assign n20410 = ~x1 & n20409 ;
  assign n20411 = n20410 ^ n20405 ;
  assign n20412 = ~x0 & n20411 ;
  assign n20413 = n20412 ^ n20403 ;
  assign n20414 = n20413 ^ n19793 ;
  assign n19797 = n19587 ^ n19577 ;
  assign n20398 = n19797 ^ n19793 ;
  assign n19800 = n12262 ^ n12220 ;
  assign n19801 = n19800 ^ n12262 ;
  assign n19802 = n12262 ^ x2 ;
  assign n19803 = n19802 ^ n12262 ;
  assign n19804 = ~n19801 & n19803 ;
  assign n19805 = n19804 ^ n12262 ;
  assign n19806 = ~x1 & ~n19805 ;
  assign n19807 = n19806 ^ n19802 ;
  assign n19796 = n19574 ^ n19243 ;
  assign n19817 = n19807 ^ n19796 ;
  assign n19799 = n12256 ^ x1 ;
  assign n19808 = n19807 ^ n19799 ;
  assign n19809 = n19808 ^ x2 ;
  assign n19810 = n19809 ^ x1 ;
  assign n19811 = n19810 ^ n19808 ;
  assign n19812 = n19808 ^ n13052 ;
  assign n19813 = n19812 ^ n19808 ;
  assign n19814 = n19811 & ~n19813 ;
  assign n19815 = n19814 ^ n19808 ;
  assign n19816 = x0 & n19815 ;
  assign n19818 = n19817 ^ n19816 ;
  assign n20331 = n19565 ^ n19278 ;
  assign n20332 = n20331 ^ n19265 ;
  assign n20284 = n12129 ^ x1 ;
  assign n20267 = n12129 ^ x2 ;
  assign n20285 = n20284 ^ n20267 ;
  assign n20286 = n13736 & n20285 ;
  assign n20287 = n20286 ^ n20284 ;
  assign n20238 = n12130 ^ x2 ;
  assign n20288 = n20287 ^ n20238 ;
  assign n20289 = n20288 ^ n20287 ;
  assign n20290 = n20289 ^ n12130 ;
  assign n20291 = ~n12136 & n20290 ;
  assign n20292 = n20291 ^ n12130 ;
  assign n20293 = ~x1 & n20292 ;
  assign n20294 = n20293 ^ n20288 ;
  assign n20295 = ~x0 & ~n20294 ;
  assign n20296 = n20295 ^ n20287 ;
  assign n20283 = n19557 ^ n19544 ;
  assign n20297 = n20296 ^ n20283 ;
  assign n20265 = n12130 ^ n12129 ;
  assign n20266 = n20265 ^ n12129 ;
  assign n20270 = n20267 ^ n12129 ;
  assign n20271 = n20266 & n20270 ;
  assign n20272 = n20271 ^ n12129 ;
  assign n20273 = ~x1 & ~n20272 ;
  assign n20261 = n12121 ^ x2 ;
  assign n20260 = n12121 ^ x1 ;
  assign n20262 = n20261 ^ n20260 ;
  assign n20263 = n13605 & n20262 ;
  assign n20264 = n20263 ^ n20260 ;
  assign n20268 = n20267 ^ n20264 ;
  assign n20274 = n20273 ^ n20268 ;
  assign n20275 = ~x0 & ~n20274 ;
  assign n20276 = n20275 ^ n20264 ;
  assign n20298 = n20296 ^ n20276 ;
  assign n20215 = n12136 ^ x1 ;
  assign n20214 = n12136 ^ x2 ;
  assign n20216 = n20215 ^ n20214 ;
  assign n20217 = n14128 & n20216 ;
  assign n20218 = n20217 ^ n20215 ;
  assign n20201 = n12137 ^ x2 ;
  assign n20221 = n20218 ^ n20201 ;
  assign n20222 = n20221 ^ n20218 ;
  assign n20223 = n20222 ^ n12137 ;
  assign n20224 = ~n12138 & n20223 ;
  assign n20225 = n20224 ^ n12137 ;
  assign n20226 = ~x1 & n20225 ;
  assign n20227 = n20226 ^ n20221 ;
  assign n20228 = ~x0 & ~n20227 ;
  assign n20229 = n20228 ^ n20218 ;
  assign n20202 = n12137 ^ x1 ;
  assign n20203 = n20202 ^ n20201 ;
  assign n20204 = n13936 & n20203 ;
  assign n20205 = n20204 ^ n20202 ;
  assign n20230 = n20229 ^ n20205 ;
  assign n20178 = n12138 ^ x2 ;
  assign n20206 = n20205 ^ n20178 ;
  assign n20207 = n20206 ^ n20205 ;
  assign n20208 = n20207 ^ n12138 ;
  assign n20209 = n12207 & n20208 ;
  assign n20210 = n20209 ^ n12138 ;
  assign n20211 = ~x1 & ~n20210 ;
  assign n20212 = n20211 ^ n20206 ;
  assign n20213 = ~x0 & ~n20212 ;
  assign n20231 = n20230 ^ n20213 ;
  assign n20232 = n20231 ^ n20229 ;
  assign n20183 = n12207 ^ n12142 ;
  assign n20184 = n20183 ^ n12207 ;
  assign n20179 = n12138 ^ x1 ;
  assign n20180 = n20179 ^ n20178 ;
  assign n20181 = n14370 & n20180 ;
  assign n20182 = n20181 ^ n20179 ;
  assign n20157 = n12207 ^ x2 ;
  assign n20185 = n20182 ^ n20157 ;
  assign n20186 = n20185 ^ n20182 ;
  assign n20187 = n20186 ^ n12207 ;
  assign n20188 = ~n20184 & n20187 ;
  assign n20189 = n20188 ^ n12207 ;
  assign n20190 = ~x1 & n20189 ;
  assign n20191 = n20190 ^ n20185 ;
  assign n20192 = ~x0 & ~n20191 ;
  assign n20193 = n20192 ^ n20182 ;
  assign n20162 = ~x2 & n14476 ;
  assign n20167 = n20162 ^ n14476 ;
  assign n20168 = n20167 ^ n12207 ;
  assign n20135 = n12142 ^ x2 ;
  assign n20163 = n20162 ^ n20135 ;
  assign n20164 = n20163 ^ n12207 ;
  assign n20165 = x0 & n20164 ;
  assign n20166 = n20165 ^ n20135 ;
  assign n20169 = n20168 ^ n20166 ;
  assign n20155 = n15500 ^ n12143 ;
  assign n20156 = n20155 ^ n12207 ;
  assign n20158 = n20157 ^ n12207 ;
  assign n20159 = ~n20156 & n20158 ;
  assign n20160 = n20159 ^ n12207 ;
  assign n20161 = ~x0 & n20160 ;
  assign n20170 = n20169 ^ n20161 ;
  assign n20171 = ~x1 & ~n20170 ;
  assign n20172 = n20171 ^ n20166 ;
  assign n20139 = n12149 ^ n12143 ;
  assign n20140 = n20139 ^ n12143 ;
  assign n20134 = n12142 ^ x1 ;
  assign n20136 = n20135 ^ n20134 ;
  assign n20137 = n14298 & n20136 ;
  assign n20138 = n20137 ^ n20134 ;
  assign n19838 = n12143 ^ x2 ;
  assign n20141 = n20138 ^ n19838 ;
  assign n20142 = n20141 ^ n20138 ;
  assign n20143 = n20142 ^ n12143 ;
  assign n20144 = n20140 & n20143 ;
  assign n20145 = n20144 ^ n12143 ;
  assign n20146 = ~x1 & n20145 ;
  assign n20147 = n20146 ^ n20141 ;
  assign n20148 = ~x0 & ~n20147 ;
  assign n20149 = n20148 ^ n20138 ;
  assign n19851 = n19511 ^ n19359 ;
  assign n19837 = n12143 ^ x1 ;
  assign n19839 = n19838 ^ n19837 ;
  assign n19840 = n14497 & n19839 ;
  assign n19841 = n19840 ^ n19837 ;
  assign n19852 = n19851 ^ n19841 ;
  assign n19842 = n12149 ^ x2 ;
  assign n19845 = n19842 ^ n12149 ;
  assign n19846 = ~n12151 & n19845 ;
  assign n19847 = n19846 ^ n12149 ;
  assign n19848 = ~x1 & n19847 ;
  assign n19843 = n19842 ^ n19841 ;
  assign n19849 = n19848 ^ n19843 ;
  assign n19850 = ~x0 & n19849 ;
  assign n19853 = n19852 ^ n19850 ;
  assign n19865 = x2 & n12152 ;
  assign n19866 = n19865 ^ n12151 ;
  assign n19867 = ~x1 & ~n19866 ;
  assign n19861 = n12151 ^ x2 ;
  assign n19855 = n12149 ^ x1 ;
  assign n19856 = n19855 ^ n19842 ;
  assign n19857 = n15311 & n19856 ;
  assign n19858 = n19857 ^ n19855 ;
  assign n19862 = n19861 ^ n19858 ;
  assign n19868 = n19867 ^ n19862 ;
  assign n19869 = ~x0 & ~n19868 ;
  assign n19870 = n19869 ^ n19858 ;
  assign n19854 = n19508 ^ n19500 ;
  assign n19871 = n19870 ^ n19854 ;
  assign n20128 = n19870 ^ n19851 ;
  assign n20101 = n12151 ^ x1 ;
  assign n20102 = n20101 ^ n19861 ;
  assign n20103 = n15299 & n20102 ;
  assign n20104 = n20103 ^ n20101 ;
  assign n19875 = n12152 ^ x2 ;
  assign n20107 = n20104 ^ n19875 ;
  assign n20108 = n20107 ^ n20104 ;
  assign n20109 = n20108 ^ n12152 ;
  assign n20110 = n12160 & n20109 ;
  assign n20111 = n20110 ^ n12152 ;
  assign n20112 = ~x1 & n20111 ;
  assign n20113 = n20112 ^ n20107 ;
  assign n20114 = ~x0 & ~n20113 ;
  assign n20115 = n20114 ^ n20104 ;
  assign n20126 = n20115 ^ n19851 ;
  assign n19888 = n19485 ^ n19370 ;
  assign n19889 = n19888 ^ n19486 ;
  assign n20116 = n20115 ^ n19889 ;
  assign n19874 = n12152 ^ x1 ;
  assign n19876 = n19875 ^ n19874 ;
  assign n19877 = n14580 & n19876 ;
  assign n19878 = n19877 ^ n19874 ;
  assign n19890 = n19889 ^ n19878 ;
  assign n19879 = n12160 ^ x2 ;
  assign n19882 = n19879 ^ n12160 ;
  assign n19883 = n12163 & n19882 ;
  assign n19884 = n19883 ^ n12160 ;
  assign n19885 = ~x1 & n19884 ;
  assign n19880 = n19879 ^ n19878 ;
  assign n19886 = n19885 ^ n19880 ;
  assign n19887 = ~x0 & n19886 ;
  assign n19891 = n19890 ^ n19887 ;
  assign n19920 = n15032 ^ n12175 ;
  assign n19921 = ~x2 & n19920 ;
  assign n19922 = n19921 ^ x2 ;
  assign n19918 = ~x1 & n12169 ;
  assign n19919 = n19918 ^ x1 ;
  assign n19923 = n19922 ^ n19919 ;
  assign n19924 = ~n12168 & n19923 ;
  assign n19925 = n19924 ^ n19922 ;
  assign n19927 = n19925 ^ n19918 ;
  assign n19926 = n19925 ^ n19921 ;
  assign n19928 = n19927 ^ n19926 ;
  assign n19931 = ~n12168 & n19928 ;
  assign n19932 = n19931 ^ n19927 ;
  assign n19933 = ~n12175 & ~n19932 ;
  assign n19934 = n19933 ^ n19925 ;
  assign n19911 = n12169 ^ n12168 ;
  assign n19936 = n12169 ^ n10828 ;
  assign n19937 = n19936 ^ n19920 ;
  assign n19938 = n19937 ^ n10828 ;
  assign n19939 = ~x1 & n19938 ;
  assign n19940 = n19939 ^ n10828 ;
  assign n19941 = ~n19911 & n19940 ;
  assign n19942 = n19941 ^ x2 ;
  assign n19943 = n19934 & n19942 ;
  assign n19944 = n19943 ^ n12167 ;
  assign n19909 = n19476 ^ n19430 ;
  assign n19948 = n19944 ^ n19909 ;
  assign n19913 = n12168 ^ x2 ;
  assign n19945 = n19944 ^ n19913 ;
  assign n19914 = n19913 ^ n12168 ;
  assign n19915 = ~n12169 & n19914 ;
  assign n19916 = n19915 ^ n12168 ;
  assign n19917 = ~x1 & n19916 ;
  assign n19946 = n19945 ^ n19917 ;
  assign n19947 = ~x0 & n19946 ;
  assign n19949 = n19948 ^ n19947 ;
  assign n20052 = n12168 ^ x1 ;
  assign n20053 = n20052 ^ n19913 ;
  assign n20054 = n14948 & n20053 ;
  assign n20055 = n20054 ^ n20052 ;
  assign n20035 = n12169 ^ x2 ;
  assign n20059 = n20055 ^ n20035 ;
  assign n20060 = n20059 ^ n20055 ;
  assign n20061 = n20060 ^ n12169 ;
  assign n20062 = n12175 & n20061 ;
  assign n20063 = n20062 ^ n12169 ;
  assign n20064 = ~x1 & ~n20063 ;
  assign n20065 = n20064 ^ n20059 ;
  assign n20066 = ~x0 & ~n20065 ;
  assign n19958 = n12175 ^ x1 ;
  assign n19957 = n12175 ^ x2 ;
  assign n19959 = n19958 ^ n19957 ;
  assign n19960 = n15048 & n19959 ;
  assign n19961 = n19960 ^ n19958 ;
  assign n19451 = n19450 ^ x5 ;
  assign n19953 = n19459 ^ n19451 ;
  assign n19971 = n19961 ^ n19953 ;
  assign n19966 = x2 & n12180 ;
  assign n19967 = n19966 ^ n12179 ;
  assign n19968 = ~x1 & n19967 ;
  assign n19962 = n12179 ^ x2 ;
  assign n19963 = n19962 ^ n19961 ;
  assign n19969 = n19968 ^ n19963 ;
  assign n19970 = ~x0 & n19969 ;
  assign n19972 = n19971 ^ n19970 ;
  assign n19991 = n11206 & ~n12183 ;
  assign n19992 = n19991 ^ n19446 ;
  assign n19977 = x2 & n12181 ;
  assign n19978 = n19977 ^ n12180 ;
  assign n19979 = ~x1 & n19978 ;
  assign n19975 = n12180 ^ x2 ;
  assign n19980 = n19979 ^ n19975 ;
  assign n19993 = n19992 ^ n19980 ;
  assign n19981 = n12179 ^ x1 ;
  assign n19982 = n19981 ^ n19980 ;
  assign n19983 = n19982 ^ x2 ;
  assign n19984 = n19983 ^ x1 ;
  assign n19985 = n19984 ^ n19982 ;
  assign n19986 = n19982 ^ n15127 ;
  assign n19987 = n19986 ^ n19982 ;
  assign n19988 = n19985 & n19987 ;
  assign n19989 = n19988 ^ n19982 ;
  assign n19990 = x0 & n19989 ;
  assign n19994 = n19993 ^ n19990 ;
  assign n20026 = n19992 ^ n19953 ;
  assign n20003 = n11468 & ~n12182 ;
  assign n20004 = n20003 ^ n12181 ;
  assign n20005 = ~x1 & n20004 ;
  assign n19999 = n12181 ^ x2 ;
  assign n19995 = n12180 ^ x1 ;
  assign n19996 = n19995 ^ n19975 ;
  assign n19997 = n12225 & n19996 ;
  assign n19998 = n19997 ^ n19995 ;
  assign n20000 = n19999 ^ n19998 ;
  assign n20006 = n20005 ^ n20000 ;
  assign n20007 = ~x0 & n20006 ;
  assign n20008 = n20007 ^ n19998 ;
  assign n20009 = n10702 & n12181 ;
  assign n20010 = n20009 ^ x2 ;
  assign n20011 = n20010 ^ n9077 ;
  assign n20012 = n20011 ^ n12182 ;
  assign n20013 = n20012 ^ n20011 ;
  assign n20016 = n20011 ^ n11240 ;
  assign n20017 = n20016 ^ n20011 ;
  assign n20018 = n20010 & ~n20017 ;
  assign n20019 = ~n20013 & n20018 ;
  assign n20020 = n20019 ^ n20013 ;
  assign n20021 = n20020 ^ n20012 ;
  assign n20022 = n12183 & n20021 ;
  assign n20023 = n20022 ^ n9077 ;
  assign n20024 = n20008 & n20023 ;
  assign n20025 = n20024 ^ n19953 ;
  assign n20027 = n20026 ^ n20025 ;
  assign n20028 = ~n19994 & n20027 ;
  assign n20029 = n20028 ^ n20025 ;
  assign n20030 = n19972 & n20029 ;
  assign n19950 = n19460 ^ x6 ;
  assign n19951 = n19950 ^ n19462 ;
  assign n19952 = n19951 ^ n19445 ;
  assign n19954 = n19953 ^ n19952 ;
  assign n20031 = n20030 ^ n19954 ;
  assign n20034 = n12169 ^ x1 ;
  assign n20036 = n20035 ^ n20034 ;
  assign n20037 = n15032 & n20036 ;
  assign n20038 = n20037 ^ n20034 ;
  assign n20047 = n20038 ^ n19952 ;
  assign n20039 = n20038 ^ n19957 ;
  assign n20040 = n20039 ^ n20038 ;
  assign n20041 = n20040 ^ n12175 ;
  assign n20042 = n12179 & n20041 ;
  assign n20043 = n20042 ^ n12175 ;
  assign n20044 = ~x1 & n20043 ;
  assign n20045 = n20044 ^ n20039 ;
  assign n20046 = ~x0 & ~n20045 ;
  assign n20048 = n20047 ^ n20046 ;
  assign n20049 = n20031 & ~n20048 ;
  assign n20050 = n20049 ^ n19952 ;
  assign n20056 = n20055 ^ n20050 ;
  assign n20067 = n20066 ^ n20056 ;
  assign n20068 = n20050 ^ n19474 ;
  assign n20069 = n20068 ^ n19467 ;
  assign n20070 = n20067 & n20069 ;
  assign n20051 = n20050 ^ n19909 ;
  assign n20071 = n20070 ^ n20051 ;
  assign n20072 = ~n19949 & ~n20071 ;
  assign n19908 = n19479 ^ n19402 ;
  assign n19910 = n19909 ^ n19908 ;
  assign n20073 = n20072 ^ n19910 ;
  assign n20074 = n12167 ^ x2 ;
  assign n20075 = n20074 ^ n12167 ;
  assign n20076 = n12168 ^ n12167 ;
  assign n20077 = n20076 ^ n12167 ;
  assign n20078 = n20075 & n20077 ;
  assign n20079 = n20078 ^ n12167 ;
  assign n20080 = ~x1 & n20079 ;
  assign n20081 = n20080 ^ n20074 ;
  assign n20090 = n20081 ^ n19908 ;
  assign n19898 = n12163 ^ x2 ;
  assign n20082 = n20081 ^ n19898 ;
  assign n20083 = n20082 ^ n10828 ;
  assign n20084 = n20083 ^ n20082 ;
  assign n20085 = n20082 ^ n14880 ;
  assign n20086 = n20085 ^ n20082 ;
  assign n20087 = n20084 & ~n20086 ;
  assign n20088 = n20087 ^ n20082 ;
  assign n20089 = x0 & n20088 ;
  assign n20091 = n20090 ^ n20089 ;
  assign n20092 = ~n20073 & n20091 ;
  assign n20093 = n20092 ^ n19908 ;
  assign n20098 = n20093 ^ n19889 ;
  assign n19901 = n19898 ^ n12163 ;
  assign n19902 = n12167 & n19901 ;
  assign n19903 = n19902 ^ n12163 ;
  assign n19904 = ~x1 & n19903 ;
  assign n19892 = n12160 ^ x1 ;
  assign n19893 = n19892 ^ n19879 ;
  assign n19894 = n14866 & n19893 ;
  assign n19895 = n19894 ^ n19892 ;
  assign n19899 = n19898 ^ n19895 ;
  assign n19905 = n19904 ^ n19899 ;
  assign n19906 = ~x0 & n19905 ;
  assign n19907 = n19906 ^ n19895 ;
  assign n20094 = n20093 ^ n19907 ;
  assign n20095 = n19907 ^ n19391 ;
  assign n20096 = n20095 ^ n19482 ;
  assign n20097 = n20094 & n20096 ;
  assign n20099 = n20098 ^ n20097 ;
  assign n20100 = n19891 & n20099 ;
  assign n20117 = n20116 ^ n20100 ;
  assign n20121 = n19377 ^ n19360 ;
  assign n20122 = n20121 ^ n19367 ;
  assign n20123 = n20122 ^ n20115 ;
  assign n20118 = n19486 ^ n19485 ;
  assign n20119 = n19486 ^ n19370 ;
  assign n20120 = n20118 & n20119 ;
  assign n20124 = n20123 ^ n20120 ;
  assign n20125 = ~n20117 & ~n20124 ;
  assign n20127 = n20126 ^ n20125 ;
  assign n20129 = n20128 ^ n20127 ;
  assign n20130 = n19871 & ~n20129 ;
  assign n20131 = n20130 ^ n20127 ;
  assign n20132 = ~n19853 & n20131 ;
  assign n20133 = n20132 ^ n19851 ;
  assign n20150 = n20149 ^ n20133 ;
  assign n20151 = n20133 ^ n19349 ;
  assign n20152 = n20151 ^ n19514 ;
  assign n20153 = n20150 & n20152 ;
  assign n20154 = n20153 ^ n20149 ;
  assign n20173 = n20172 ^ n20154 ;
  assign n20174 = n19517 ^ n19339 ;
  assign n20175 = n20174 ^ n20154 ;
  assign n20176 = n20173 & ~n20175 ;
  assign n20177 = n20176 ^ n20172 ;
  assign n20194 = n20193 ^ n20177 ;
  assign n20195 = n20177 ^ n19329 ;
  assign n20196 = n20195 ^ n19520 ;
  assign n20197 = n20194 & ~n20196 ;
  assign n20198 = n20197 ^ n20193 ;
  assign n20233 = n20232 ^ n20198 ;
  assign n20234 = n19523 ^ n19319 ;
  assign n20235 = n20234 ^ n20198 ;
  assign n20236 = ~n20233 & ~n20235 ;
  assign n20237 = n20236 ^ n20231 ;
  assign n20239 = n12130 ^ x1 ;
  assign n20240 = n20239 ^ n20238 ;
  assign n20241 = n13817 & n20240 ;
  assign n20242 = n20241 ^ n20239 ;
  assign n20245 = n20242 ^ n20214 ;
  assign n20246 = n20245 ^ n20242 ;
  assign n20247 = n20246 ^ n12136 ;
  assign n20248 = n12137 & n20247 ;
  assign n20249 = n20248 ^ n12136 ;
  assign n20250 = ~x1 & ~n20249 ;
  assign n20251 = n20250 ^ n20245 ;
  assign n20252 = ~x0 & ~n20251 ;
  assign n20253 = n20252 ^ n20242 ;
  assign n20254 = n20253 ^ n20229 ;
  assign n20255 = n20254 ^ n19539 ;
  assign n20256 = n20255 ^ n19526 ;
  assign n20257 = n20256 ^ n20253 ;
  assign n20258 = ~n20237 & ~n20257 ;
  assign n20259 = n20258 ^ n20254 ;
  assign n20277 = n20276 ^ n20253 ;
  assign n20278 = n20277 ^ n20276 ;
  assign n20279 = n20278 ^ n19541 ;
  assign n20280 = n20279 ^ n19309 ;
  assign n20281 = ~n20259 & ~n20280 ;
  assign n20282 = n20281 ^ n20277 ;
  assign n20299 = n20298 ^ n20282 ;
  assign n20300 = n20297 & ~n20299 ;
  assign n20301 = n20300 ^ n20282 ;
  assign n20303 = n12117 ^ x2 ;
  assign n20302 = n12117 ^ x1 ;
  assign n20304 = n20303 ^ n20302 ;
  assign n20305 = n13586 & n20304 ;
  assign n20306 = n20305 ^ n20302 ;
  assign n20309 = n20306 ^ n20261 ;
  assign n20310 = n20309 ^ n20306 ;
  assign n20311 = n20310 ^ n12121 ;
  assign n20312 = ~n12129 & n20311 ;
  assign n20313 = n20312 ^ n12121 ;
  assign n20314 = ~x1 & n20313 ;
  assign n20315 = n20314 ^ n20309 ;
  assign n20316 = ~x0 & n20315 ;
  assign n20317 = n20316 ^ n20306 ;
  assign n20318 = n20317 ^ n20276 ;
  assign n20319 = n20318 ^ n19298 ;
  assign n20320 = n20319 ^ n20317 ;
  assign n20321 = n20320 ^ n19559 ;
  assign n20322 = n20301 & ~n20321 ;
  assign n20323 = n20322 ^ n20318 ;
  assign n20324 = n20317 ^ n19265 ;
  assign n20325 = n20324 ^ n19562 ;
  assign n20326 = n20325 ^ n19265 ;
  assign n20327 = n20326 ^ n19288 ;
  assign n20328 = n20323 & n20327 ;
  assign n20329 = n20328 ^ n20324 ;
  assign n20333 = n20332 ^ n20329 ;
  assign n20335 = n12110 ^ x2 ;
  assign n20334 = n12110 ^ x1 ;
  assign n20336 = n20335 ^ n20334 ;
  assign n20337 = n13195 & n20336 ;
  assign n20338 = n20337 ^ n20334 ;
  assign n20341 = n20338 ^ n20303 ;
  assign n20342 = n20341 ^ n20338 ;
  assign n20343 = n20342 ^ n12117 ;
  assign n20344 = n12121 & n20343 ;
  assign n20345 = n20344 ^ n12117 ;
  assign n20346 = ~x1 & n20345 ;
  assign n20347 = n20346 ^ n20341 ;
  assign n20348 = ~x0 & ~n20347 ;
  assign n20339 = n20338 ^ n20331 ;
  assign n20349 = n20348 ^ n20339 ;
  assign n20350 = ~n20333 & ~n20349 ;
  assign n20330 = n20329 ^ n19568 ;
  assign n20351 = n20350 ^ n20330 ;
  assign n20354 = n12220 ^ x1 ;
  assign n20355 = n20354 ^ x2 ;
  assign n20356 = n20355 ^ n12220 ;
  assign n20357 = n13172 & n20356 ;
  assign n20358 = n20357 ^ n20354 ;
  assign n19824 = n12220 ^ x2 ;
  assign n19819 = n12262 ^ x1 ;
  assign n19820 = n19819 ^ x2 ;
  assign n19821 = n19820 ^ n12262 ;
  assign n19822 = n12250 & n19821 ;
  assign n19823 = n19822 ^ n19819 ;
  assign n19825 = n19824 ^ n19823 ;
  assign n19826 = n19825 ^ n19823 ;
  assign n19827 = n19826 ^ n13165 ;
  assign n19828 = ~n13166 & ~n19827 ;
  assign n19829 = n19828 ^ n13165 ;
  assign n19830 = ~x1 & n19829 ;
  assign n19831 = n19830 ^ n19825 ;
  assign n19832 = ~x0 & n19831 ;
  assign n19833 = n19832 ^ n19823 ;
  assign n20367 = n20358 ^ n19833 ;
  assign n20359 = n20358 ^ n20335 ;
  assign n20360 = n20359 ^ n20358 ;
  assign n20361 = n20360 ^ n12110 ;
  assign n20362 = n12117 & n20361 ;
  assign n20363 = n20362 ^ n12110 ;
  assign n20364 = ~x1 & ~n20363 ;
  assign n20365 = n20364 ^ n20359 ;
  assign n20366 = ~x0 & n20365 ;
  assign n20368 = n20367 ^ n20366 ;
  assign n20369 = n20368 ^ n19265 ;
  assign n20370 = n20369 ^ n19568 ;
  assign n20371 = n20370 ^ n19833 ;
  assign n20372 = ~n20351 & ~n20371 ;
  assign n20373 = n20372 ^ n20368 ;
  assign n20374 = n19833 ^ n19571 ;
  assign n20375 = n20374 ^ n19253 ;
  assign n20376 = n20373 & ~n20375 ;
  assign n19834 = n19833 ^ n19796 ;
  assign n20377 = n20376 ^ n19834 ;
  assign n20378 = ~n19818 & ~n20377 ;
  assign n19798 = n19797 ^ n19796 ;
  assign n20379 = n20378 ^ n19798 ;
  assign n20381 = n12260 ^ x1 ;
  assign n20383 = n20382 ^ n20381 ;
  assign n20384 = ~n13053 & n20383 ;
  assign n20385 = n20384 ^ n20381 ;
  assign n20395 = n20385 ^ n19797 ;
  assign n20386 = n12256 ^ x2 ;
  assign n20387 = n20386 ^ n20385 ;
  assign n20388 = n20387 ^ n20385 ;
  assign n20389 = n20388 ^ n12256 ;
  assign n20390 = ~n12262 & n20389 ;
  assign n20391 = n20390 ^ n12256 ;
  assign n20392 = ~x1 & ~n20391 ;
  assign n20393 = n20392 ^ n20387 ;
  assign n20394 = ~x0 & ~n20393 ;
  assign n20396 = n20395 ^ n20394 ;
  assign n20397 = ~n20379 & ~n20396 ;
  assign n20399 = n20398 ^ n20397 ;
  assign n20415 = n20414 ^ n20399 ;
  assign n20416 = n20413 ^ n19231 ;
  assign n20417 = n20416 ^ n19590 ;
  assign n20418 = ~n20415 & n20417 ;
  assign n20419 = n20418 ^ n20399 ;
  assign n20420 = ~n19795 & ~n20419 ;
  assign n20421 = n20420 ^ n19793 ;
  assign n20422 = n20421 ^ n19772 ;
  assign n20423 = ~n19774 & ~n20422 ;
  assign n20424 = n20423 ^ n19772 ;
  assign n20425 = n20424 ^ n19740 ;
  assign n20426 = ~n19756 & n20425 ;
  assign n20428 = n20427 ^ n20426 ;
  assign n20429 = ~n19739 & n20428 ;
  assign n20430 = n20429 ^ n19738 ;
  assign n20445 = ~n19721 & ~n20430 ;
  assign n19700 = ~n19200 & n19624 ;
  assign n20446 = n19700 ^ n19627 ;
  assign n19701 = n19700 ^ n19192 ;
  assign n20447 = n19701 ^ n19700 ;
  assign n20448 = ~n20446 & ~n20447 ;
  assign n20449 = n20448 ^ n19700 ;
  assign n20450 = n20445 & ~n20449 ;
  assign n20460 = n20450 ^ n20445 ;
  assign n20439 = n20430 ^ n19721 ;
  assign n20451 = n20450 ^ n20439 ;
  assign n19702 = n19624 ^ n19201 ;
  assign n19703 = n19702 ^ n19200 ;
  assign n20452 = n19201 ^ n19192 ;
  assign n20453 = n20452 ^ n19192 ;
  assign n20454 = n19200 ^ n19192 ;
  assign n20455 = n20454 ^ n19192 ;
  assign n20456 = ~n20453 & n20455 ;
  assign n20457 = n20456 ^ n19192 ;
  assign n20458 = n19703 & n20457 ;
  assign n20459 = n20451 & n20458 ;
  assign n20461 = n20460 ^ n20459 ;
  assign n20431 = n19721 & n20430 ;
  assign n20432 = n19700 ^ n19625 ;
  assign n20433 = n20432 ^ n19627 ;
  assign n20434 = n20432 ^ n19192 ;
  assign n20435 = n20434 ^ n20432 ;
  assign n20436 = n20433 & ~n20435 ;
  assign n20437 = n20436 ^ n20432 ;
  assign n20438 = n20431 & ~n20437 ;
  assign n20442 = n20438 ^ n20431 ;
  assign n19704 = n19701 & ~n19703 ;
  assign n20440 = n20439 ^ n20438 ;
  assign n20441 = n19704 & n20440 ;
  assign n20443 = n20442 ^ n20441 ;
  assign n20462 = n20461 ^ n20443 ;
  assign n20473 = n11240 ^ x2 ;
  assign n20476 = n11240 & n12656 ;
  assign n20477 = ~n20473 & n20476 ;
  assign n20463 = n10828 & ~n12724 ;
  assign n20464 = n20463 ^ n12755 ;
  assign n20467 = n20464 ^ n12705 ;
  assign n20468 = n20467 ^ n20464 ;
  assign n20469 = x1 & n20468 ;
  assign n20470 = n20469 ^ n20464 ;
  assign n20471 = ~x0 & ~n20470 ;
  assign n20472 = n20471 ^ n20464 ;
  assign n20474 = n20473 ^ n20472 ;
  assign n20478 = n20477 ^ n20474 ;
  assign n20479 = ~n20462 & ~n20478 ;
  assign n20444 = n20443 ^ x2 ;
  assign n20480 = n20479 ^ n20444 ;
  assign n20495 = n20494 ^ n20480 ;
  assign n20497 = n19643 ^ n19630 ;
  assign n20498 = n20497 ^ n20494 ;
  assign n20499 = n20498 ^ n20480 ;
  assign n20496 = n20480 ^ x2 ;
  assign n20500 = n20499 ^ n20496 ;
  assign n20501 = n20495 & n20500 ;
  assign n20502 = n20501 ^ n20499 ;
  assign n20503 = n20502 ^ n19697 ;
  assign n20504 = n19699 & n20503 ;
  assign n20505 = n20504 ^ n19697 ;
  assign n20506 = n20505 ^ n19666 ;
  assign n20507 = ~n19681 & ~n20506 ;
  assign n20508 = n20507 ^ n19666 ;
  assign n20509 = n20508 ^ n19662 ;
  assign n20510 = ~n19665 & ~n20509 ;
  assign n20511 = n20510 ^ n19662 ;
  assign n19149 = n7135 & n12706 ;
  assign n19145 = n18619 ^ n18200 ;
  assign n19146 = n19145 ^ x8 ;
  assign n19144 = n8054 & ~n12705 ;
  assign n19147 = n19146 ^ n19144 ;
  assign n19143 = n7146 & ~n12613 ;
  assign n19148 = n19147 ^ n19143 ;
  assign n19150 = n19149 ^ n19148 ;
  assign n19142 = n7141 & n12656 ;
  assign n19151 = n19150 ^ n19142 ;
  assign n19130 = n19129 ^ n19128 ;
  assign n19140 = n19130 & ~n19139 ;
  assign n19141 = n19140 ^ n19129 ;
  assign n19152 = n19151 ^ n19141 ;
  assign n20550 = n20511 ^ n19152 ;
  assign n20512 = n19152 & ~n20511 ;
  assign n20551 = n20550 ^ n20512 ;
  assign n20523 = n18622 ^ n18190 ;
  assign n20520 = n9081 & ~n14221 ;
  assign n20518 = n9077 ^ x5 ;
  assign n20517 = ~n9092 & n12971 ;
  assign n20519 = n20518 ^ n20517 ;
  assign n20521 = n20520 ^ n20519 ;
  assign n20516 = n9085 & ~n12855 ;
  assign n20522 = n20521 ^ n20516 ;
  assign n20524 = n20523 ^ n20522 ;
  assign n20513 = n19145 ^ n19141 ;
  assign n20514 = ~n19151 & n20513 ;
  assign n20515 = n20514 ^ n19145 ;
  assign n20525 = n20524 ^ n20515 ;
  assign n20526 = n20525 ^ n20512 ;
  assign n20531 = n9089 & ~n13007 ;
  assign n20534 = ~n9092 & n12755 ;
  assign n20533 = n9085 & n12971 ;
  assign n20535 = n20534 ^ n20533 ;
  assign n20536 = n20535 ^ x5 ;
  assign n20532 = n9077 & ~n12855 ;
  assign n20537 = n20536 ^ n20532 ;
  assign n20538 = n20537 ^ n20536 ;
  assign n20539 = n20531 & n20538 ;
  assign n20540 = n20539 ^ n20537 ;
  assign n20528 = n19655 ^ n19651 ;
  assign n20529 = n19661 & ~n20528 ;
  assign n20530 = n20529 ^ n19655 ;
  assign n20541 = n20540 ^ n20530 ;
  assign n20544 = n20540 ^ n20512 ;
  assign n20527 = n20512 ^ n14315 ;
  assign n20545 = n20544 ^ n20527 ;
  assign n20546 = ~n20541 & n20545 ;
  assign n20547 = n20546 ^ n20527 ;
  assign n20548 = ~n20526 & ~n20547 ;
  assign n20549 = n20548 ^ n20525 ;
  assign n20552 = n20540 ^ n20525 ;
  assign n20553 = n20525 ^ n14315 ;
  assign n20554 = n20530 ^ n20525 ;
  assign n20555 = ~n20553 & ~n20554 ;
  assign n20556 = ~n20552 & n20555 ;
  assign n20557 = n20556 ^ n20552 ;
  assign n20558 = n20557 ^ n20540 ;
  assign n20559 = n20549 & ~n20558 ;
  assign n20560 = ~n20551 & n20559 ;
  assign n20561 = n20560 ^ n20549 ;
  assign n20562 = n20522 ^ n20515 ;
  assign n20563 = n20524 & ~n20562 ;
  assign n20564 = n20563 ^ n20522 ;
  assign n20565 = n20561 & ~n20564 ;
  assign n18637 = n18090 ^ n14314 ;
  assign n18638 = n18637 ^ n18121 ;
  assign n20566 = n20565 ^ n18638 ;
  assign n20568 = n18638 ^ n18626 ;
  assign n20567 = n18638 ^ n18625 ;
  assign n20569 = n20568 ^ n20567 ;
  assign n20570 = n20568 ^ n18633 ;
  assign n20571 = n20570 ^ n20568 ;
  assign n20572 = n20569 & n20571 ;
  assign n20573 = n20572 ^ n20568 ;
  assign n20574 = ~n20566 & n20573 ;
  assign n20575 = n20574 ^ n20565 ;
  assign n20576 = n20564 ^ n20561 ;
  assign n20577 = n20576 ^ n20565 ;
  assign n20578 = ~n20575 & ~n20577 ;
  assign n20579 = n18638 ^ n18635 ;
  assign n20580 = n20578 & ~n20579 ;
  assign n20581 = n20580 ^ n20575 ;
  assign n20582 = n20581 ^ n20575 ;
  assign n20583 = n18636 & n20582 ;
  assign n20584 = n20583 ^ n20581 ;
  assign n20585 = n20584 ^ n18154 ;
  assign n20586 = n20585 ^ n18173 ;
  assign n20587 = ~n18174 & n20586 ;
  assign n20589 = n20585 ^ n18172 ;
  assign n20588 = n18153 ^ n18138 ;
  assign n20590 = n20589 ^ n20588 ;
  assign n20591 = n20587 & ~n20590 ;
  assign n20592 = n20591 ^ n18174 ;
  assign n20593 = ~n18129 & n20592 ;
  assign n20594 = n20584 ^ n18169 ;
  assign n20595 = n20593 & n20594 ;
  assign n20596 = n20595 ^ n20592 ;
  assign n20597 = n20596 ^ n20592 ;
  assign n20598 = n20588 ^ n18154 ;
  assign n20599 = ~n20585 & ~n20598 ;
  assign n20600 = n20597 & n20599 ;
  assign n20601 = n20600 ^ n20596 ;
  assign n16707 = n16706 ^ n16339 ;
  assign n20602 = n20601 ^ n16707 ;
  assign n20604 = n18167 ^ n16707 ;
  assign n20603 = n18160 ^ n16707 ;
  assign n20605 = n20604 ^ n20603 ;
  assign n20606 = n18166 & n20605 ;
  assign n20607 = n20606 ^ n20604 ;
  assign n20608 = n20602 & n20607 ;
  assign n20609 = n20608 ^ n20601 ;
  assign n20613 = n20612 ^ n20609 ;
  assign n16336 = n16284 ^ n16250 ;
  assign n16337 = n16336 ^ n16233 ;
  assign n20614 = n20613 ^ n16337 ;
  assign n20615 = n20614 ^ n16337 ;
  assign n20616 = n20612 ^ n16233 ;
  assign n20617 = n20616 ^ n16337 ;
  assign n20618 = n20615 & ~n20617 ;
  assign n20619 = n20618 ^ n16337 ;
  assign n20620 = n16335 & n20619 ;
  assign n20621 = n20620 ^ n16334 ;
  assign n20622 = n16232 ^ n15419 ;
  assign n20623 = n20622 ^ n16233 ;
  assign n20624 = ~n20621 & n20623 ;
  assign n20625 = n20612 ^ n16336 ;
  assign n20626 = n20625 ^ n20609 ;
  assign n20631 = ~n20609 & n20612 ;
  assign n20632 = n20631 ^ n16334 ;
  assign n20633 = n20626 & n20632 ;
  assign n20634 = n20624 & n20633 ;
  assign n20635 = n20634 ^ n20621 ;
  assign n20666 = n20665 ^ n20635 ;
  assign n20669 = n20665 ^ n16327 ;
  assign n20667 = n16327 ^ n16287 ;
  assign n20668 = ~n16333 & ~n20667 ;
  assign n20670 = n20669 ^ n20668 ;
  assign n20671 = n20666 & n20670 ;
  assign n20672 = n20671 ^ n20665 ;
  assign n20694 = n20693 ^ n20672 ;
  assign n20695 = n20689 & ~n20694 ;
  assign n15408 = n15407 ^ n15406 ;
  assign n20677 = n20676 ^ n15407 ;
  assign n20673 = n20672 ^ n15406 ;
  assign n20678 = n20677 ^ n20673 ;
  assign n20682 = n20681 ^ n15406 ;
  assign n20683 = n20682 ^ n20677 ;
  assign n20684 = n20678 & n20683 ;
  assign n20685 = n20684 ^ n20677 ;
  assign n20686 = ~n15408 & n20685 ;
  assign n20687 = n20686 ^ n15407 ;
  assign n20696 = n20690 ^ n15407 ;
  assign n20697 = n20687 & ~n20696 ;
  assign n20698 = n20695 & n20697 ;
  assign n20699 = n20698 ^ n20687 ;
  assign n20700 = n14788 ^ n14698 ;
  assign n20701 = n14790 & n20700 ;
  assign n20702 = n20701 ^ n14788 ;
  assign n20703 = n20699 & n20702 ;
  assign n20704 = n20703 ^ n15396 ;
  assign n20705 = ~n15398 & ~n20704 ;
  assign n20706 = n20705 ^ n15396 ;
  assign n20707 = n15393 & ~n20706 ;
  assign n20708 = n20707 ^ n14686 ;
  assign n20709 = n14687 ^ n14686 ;
  assign n20710 = n14686 ^ n6070 ;
  assign n20711 = n15391 ^ n6070 ;
  assign n20712 = n20710 & n20711 ;
  assign n20713 = n20709 & n20712 ;
  assign n20718 = n20713 ^ n15396 ;
  assign n20714 = n20713 ^ n14686 ;
  assign n20715 = n20714 ^ n20699 ;
  assign n20716 = n20714 ^ n20702 ;
  assign n20717 = n20715 & n20716 ;
  assign n20719 = n20702 & n20717 ;
  assign n20720 = ~n20718 & n20719 ;
  assign n20721 = n20720 ^ n20717 ;
  assign n20722 = n20721 ^ n20714 ;
  assign n20723 = ~n20708 & ~n20722 ;
  assign n20757 = n20754 ^ n20723 ;
  assign n20758 = n20757 ^ n20754 ;
  assign n20759 = ~n20756 & n20758 ;
  assign n20760 = n20759 ^ n20754 ;
  assign n20761 = n20753 & ~n20760 ;
  assign n20762 = n20761 ^ n20723 ;
  assign n20724 = n20723 ^ n14423 ;
  assign n20739 = n20738 ^ n20733 ;
  assign n20741 = n20740 ^ n20733 ;
  assign n20742 = n20741 ^ n20740 ;
  assign n20743 = n20740 ^ n20734 ;
  assign n20744 = n20743 ^ n20740 ;
  assign n20745 = ~n20742 & n20744 ;
  assign n20746 = n20745 ^ n20740 ;
  assign n20747 = n20739 & n20746 ;
  assign n20748 = n20747 ^ n14423 ;
  assign n20749 = ~n20724 & n20748 ;
  assign n20763 = n20762 ^ n20749 ;
  assign n20765 = n20763 ^ n14036 ;
  assign n14224 = n4678 ^ x20 ;
  assign n14223 = n12971 & n14027 ;
  assign n14225 = n14224 ^ n14223 ;
  assign n14222 = n4684 & ~n14221 ;
  assign n14226 = n14225 ^ n14222 ;
  assign n14220 = n4916 & ~n12855 ;
  assign n14227 = n14226 ^ n14220 ;
  assign n20764 = n20763 ^ n14227 ;
  assign n20766 = n20765 ^ n20764 ;
  assign n20767 = n20766 ^ n20765 ;
  assign n20768 = n14212 ^ n14197 ;
  assign n20769 = ~n14202 & n20768 ;
  assign n20770 = n20769 ^ n14197 ;
  assign n20771 = n20770 ^ n14227 ;
  assign n20772 = n20771 ^ n20765 ;
  assign n20773 = n20772 ^ n20765 ;
  assign n20774 = ~n20767 & ~n20773 ;
  assign n20775 = n20774 ^ n20765 ;
  assign n20776 = ~n14219 & n20775 ;
  assign n20777 = n20776 ^ n14218 ;
  assign n20780 = n14227 ^ n14036 ;
  assign n20781 = n20770 ^ n14036 ;
  assign n20782 = ~n20765 & n20781 ;
  assign n20783 = n20780 & n20782 ;
  assign n20784 = n20783 ^ n20780 ;
  assign n20785 = n20784 ^ n14227 ;
  assign n20786 = ~n20777 & ~n20785 ;
  assign n20787 = n20779 & n20786 ;
  assign n20788 = n20787 ^ n20777 ;
  assign n20789 = ~n14035 & n20788 ;
  assign n20790 = n13698 ^ n13533 ;
  assign n20791 = n20790 ^ n13699 ;
  assign n20792 = ~n14033 & ~n20791 ;
  assign n20793 = ~n20789 & n20792 ;
  assign n20794 = n14035 ^ n13533 ;
  assign n20795 = ~n13697 & n20794 ;
  assign n20796 = n14033 ^ n13533 ;
  assign n20797 = n20796 ^ n20788 ;
  assign n20798 = n20795 & ~n20797 ;
  assign n20799 = ~n20793 & ~n20798 ;
  assign n20800 = ~n13699 & n20799 ;
  assign n13529 = n13528 ^ n13422 ;
  assign n13530 = n13426 & n13529 ;
  assign n13531 = n13530 ^ n13422 ;
  assign n20801 = n20800 ^ n13531 ;
  assign n20825 = n20801 ^ n13355 ;
  assign n20804 = n13419 ^ n13406 ;
  assign n20805 = n13421 & n20804 ;
  assign n20806 = n20805 ^ n13420 ;
  assign n20826 = n20825 ^ n20806 ;
  assign n20827 = ~n20809 & ~n20826 ;
  assign n20823 = n20806 ^ n13531 ;
  assign n20824 = n20801 & n20823 ;
  assign n20828 = n20827 ^ n20824 ;
  assign n20829 = n20822 & ~n20828 ;
  assign n13532 = n13531 ^ n13355 ;
  assign n20802 = ~n13532 & ~n20801 ;
  assign n20803 = n20802 ^ n13531 ;
  assign n20816 = n20801 ^ n13532 ;
  assign n20817 = n20816 ^ n13531 ;
  assign n20810 = n20809 ^ n13355 ;
  assign n20811 = n20810 ^ n20806 ;
  assign n20812 = n20806 ^ n20800 ;
  assign n20813 = n20812 ^ n13355 ;
  assign n20814 = n20813 ^ n13531 ;
  assign n20815 = ~n20811 & ~n20814 ;
  assign n20818 = n20817 ^ n20815 ;
  assign n20819 = ~n20803 & ~n20818 ;
  assign n20820 = n20819 ^ n13531 ;
  assign n20821 = n20820 ^ n13531 ;
  assign n20830 = n20829 ^ n20821 ;
  assign n20831 = n20830 ^ n13352 ;
  assign n20832 = n13354 & n20831 ;
  assign n20833 = n20832 ^ n20830 ;
  assign n24005 = n13104 ^ n12984 ;
  assign n24007 = n24006 ^ n24005 ;
  assign n24008 = ~n20833 & ~n24007 ;
  assign n24464 = ~n24006 & ~n24008 ;
  assign n12768 = n12767 ^ n12720 ;
  assign n12843 = n12842 ^ n12720 ;
  assign n12844 = ~n12768 & n12843 ;
  assign n12845 = n12844 ^ n12767 ;
  assign n12863 = n80 ^ n73 ;
  assign n12864 = n12863 ^ n114 ;
  assign n12862 = ~n12855 & n12861 ;
  assign n12865 = n12864 ^ n12862 ;
  assign n24469 = n12845 & n12865 ;
  assign n24470 = n24469 ^ n24007 ;
  assign n24074 = n24073 ^ n24062 ;
  assign n12866 = n12865 ^ n12845 ;
  assign n24009 = n24006 ^ n12865 ;
  assign n24010 = ~n12866 & n24009 ;
  assign n24011 = n24010 ^ n24006 ;
  assign n24466 = n24074 ^ n24011 ;
  assign n24471 = n24470 ^ n24466 ;
  assign n24584 = n24471 ^ n24007 ;
  assign n24585 = n24584 ^ n20833 ;
  assign n24586 = n24585 ^ n24011 ;
  assign n24590 = n24586 ^ n20833 ;
  assign n24593 = n24590 ^ n24471 ;
  assign n24587 = n24586 ^ n24466 ;
  assign n24594 = n24593 ^ n24587 ;
  assign n24595 = n24594 ^ n24011 ;
  assign n24597 = n24595 ^ n24593 ;
  assign n24478 = n24011 ^ n24007 ;
  assign n24482 = n24478 ^ n24469 ;
  assign n24483 = n24482 ^ n24011 ;
  assign n24567 = n24483 ^ n20833 ;
  assign n24479 = n24478 ^ n20833 ;
  assign n24480 = n24479 ^ n24011 ;
  assign n24564 = n24483 ^ n24480 ;
  assign n24565 = n24564 ^ n24483 ;
  assign n24566 = n24565 ^ n24466 ;
  assign n24573 = n24567 ^ n24566 ;
  assign n24577 = n24573 ^ n24478 ;
  assign n24568 = n24567 ^ n24466 ;
  assign n24569 = n24568 ^ n24566 ;
  assign n24473 = n24466 ^ n24007 ;
  assign n24555 = n24473 ^ n20833 ;
  assign n24556 = n24555 ^ n24466 ;
  assign n24490 = n24473 ^ n24469 ;
  assign n24557 = n24556 ^ n24490 ;
  assign n24494 = n24473 ^ n24466 ;
  assign n24558 = n24557 ^ n24494 ;
  assign n24560 = n24558 ^ n24074 ;
  assign n24561 = n24560 ^ n24557 ;
  assign n24465 = n24007 ^ n20833 ;
  assign n24491 = n24490 ^ n24465 ;
  assign n24502 = n24494 ^ n24491 ;
  assign n24503 = n24502 ^ n24074 ;
  assign n24504 = n24503 ^ n20833 ;
  assign n24543 = n24504 ^ n24494 ;
  assign n24539 = n24503 ^ n24011 ;
  assign n24544 = n24543 ^ n24539 ;
  assign n24545 = n24544 ^ n24074 ;
  assign n24547 = n24545 ^ n24543 ;
  assign n24540 = n24494 ^ n24011 ;
  assign n24521 = ~n24074 & ~n24466 ;
  assign n24505 = n24504 ^ n24011 ;
  assign n24506 = n24505 ^ n24007 ;
  assign n24507 = n24506 ^ n24465 ;
  assign n24508 = n24507 ^ n24466 ;
  assign n24522 = n24521 ^ n24508 ;
  assign n24467 = n24466 ^ n24465 ;
  assign n24523 = n24522 ^ n24467 ;
  assign n24516 = n24540 ^ n24494 ;
  assign n24524 = n24523 ^ n24516 ;
  assign n24526 = n24516 ^ n24473 ;
  assign n24527 = n24524 & n24526 ;
  assign n24510 = n24505 ^ n24466 ;
  assign n24528 = n24510 ^ n24494 ;
  assign n24529 = n24540 ^ n24528 ;
  assign n24530 = n24508 ^ n24494 ;
  assign n24531 = n24540 ^ n24530 ;
  assign n24532 = n24529 & ~n24531 ;
  assign n24533 = n24527 & n24532 ;
  assign n24534 = n24533 ^ n24521 ;
  assign n24517 = n24510 ^ n24508 ;
  assign n24535 = n24534 ^ n24517 ;
  assign n24513 = n24494 ^ n24467 ;
  assign n24515 = n24540 ^ n24513 ;
  assign n24536 = n24535 ^ n24515 ;
  assign n24537 = n24536 ^ n24506 ;
  assign n24538 = n24540 ^ n24537 ;
  assign n24548 = n24547 ^ n24538 ;
  assign n24549 = n24548 ^ n24502 ;
  assign n24550 = n24549 ^ n24545 ;
  assign n24497 = n24490 ^ n24466 ;
  assign n24492 = n24491 ^ n24074 ;
  assign n24493 = n24492 ^ n24466 ;
  assign n24496 = n24493 ^ n24473 ;
  assign n24498 = n24497 ^ n24496 ;
  assign n24500 = n24498 ^ n24074 ;
  assign n24499 = n24498 ^ n24497 ;
  assign n24501 = n24500 ^ n24499 ;
  assign n24551 = n24550 ^ n24501 ;
  assign n24552 = n24551 ^ n24491 ;
  assign n24553 = n24552 ^ n24500 ;
  assign n24562 = n24561 ^ n24553 ;
  assign n24563 = n24562 ^ n24560 ;
  assign n24570 = n24569 ^ n24563 ;
  assign n24578 = n24577 ^ n24570 ;
  assign n24598 = n24597 ^ n24578 ;
  assign n24602 = n24598 ^ n24074 ;
  assign n24468 = n24467 ^ n24466 ;
  assign n24472 = n24471 ^ n24468 ;
  assign n24474 = n24473 ^ n24472 ;
  assign n24476 = n24474 ^ n24011 ;
  assign n24603 = n24602 ^ n24476 ;
  assign n24604 = n24469 ^ n24074 ;
  assign n24605 = n24604 ^ n12866 ;
  assign n24606 = n24603 & ~n24605 ;
  assign n24607 = n24464 & n24606 ;
  assign n24608 = n24607 ^ n24603 ;
  assign n24700 = n24699 ^ n24608 ;
  assign n24702 = n24700 ^ x2 ;
  assign n24990 = n10850 & ~n24702 ;
  assign n24012 = n24008 & n24011 ;
  assign n24026 = n13104 ^ n12865 ;
  assign n24017 = n12984 ^ n12845 ;
  assign n24018 = ~n24005 & ~n24017 ;
  assign n24027 = n24026 ^ n24018 ;
  assign n24075 = n24074 ^ n24027 ;
  assign n24013 = n12984 ^ n12865 ;
  assign n24014 = n24013 ^ n12845 ;
  assign n24015 = n24014 ^ n13104 ;
  assign n24016 = n24014 ^ n12865 ;
  assign n24019 = n24018 ^ n24016 ;
  assign n24020 = n24019 ^ n12865 ;
  assign n24021 = n20833 ^ n12865 ;
  assign n24022 = n24021 ^ n12865 ;
  assign n24023 = n24020 & ~n24022 ;
  assign n24024 = n24023 ^ n12865 ;
  assign n24025 = ~n24015 & n24024 ;
  assign n24076 = n24075 ^ n24025 ;
  assign n24077 = n24076 ^ n24074 ;
  assign n24078 = n24012 & ~n24077 ;
  assign n24079 = n24078 ^ n24076 ;
  assign n24989 = n10854 & ~n24079 ;
  assign n24991 = n24990 ^ n24989 ;
  assign n24978 = n24611 ^ n24608 ;
  assign n24979 = ~n24699 & ~n24978 ;
  assign n24975 = n24696 ^ n24668 ;
  assign n24976 = n24697 & n24975 ;
  assign n24968 = n12912 ^ n12859 ;
  assign n24969 = n24681 & n24968 ;
  assign n24970 = n24969 ^ n12859 ;
  assign n24966 = n24676 ^ n3939 ;
  assign n24967 = n24966 ^ n334 ;
  assign n24971 = n24970 ^ n24967 ;
  assign n24963 = ~n13005 & ~n24053 ;
  assign n24964 = x31 & n24963 ;
  assign n24959 = ~n3733 & n12755 ;
  assign n24958 = n3726 & n12971 ;
  assign n24960 = n24959 ^ n24958 ;
  assign n24961 = n24960 ^ x31 ;
  assign n24965 = n24964 ^ n24961 ;
  assign n24972 = n24971 ^ n24965 ;
  assign n24950 = n24684 ^ n24681 ;
  assign n24952 = n24688 ^ n828 ;
  assign n24953 = n24952 ^ n24674 ;
  assign n24951 = n24681 ^ n12912 ;
  assign n24954 = n24953 ^ n24951 ;
  assign n24955 = n24954 ^ n24952 ;
  assign n24956 = n24950 & ~n24955 ;
  assign n24957 = n24956 ^ n24953 ;
  assign n24973 = n24972 ^ n24957 ;
  assign n24974 = n24973 ^ n24697 ;
  assign n24977 = n24976 ^ n24974 ;
  assign n24980 = n24979 ^ n24977 ;
  assign n24981 = n24980 ^ x2 ;
  assign n12985 = n12984 ^ n12866 ;
  assign n13105 = n13104 ^ n12985 ;
  assign n20834 = n20833 ^ n13105 ;
  assign n20837 = n20830 ^ n13354 ;
  assign n20836 = n20828 ^ n20822 ;
  assign n20850 = n20809 ^ n20806 ;
  assign n20851 = n20850 ^ n13531 ;
  assign n20852 = n20851 ^ n20800 ;
  assign n20857 = n20789 ^ n14033 ;
  assign n20858 = n20857 ^ n13697 ;
  assign n20859 = n20858 ^ n13533 ;
  assign n20854 = n14033 ^ n13696 ;
  assign n20855 = n20788 ^ n14033 ;
  assign n20856 = n20854 & ~n20855 ;
  assign n20860 = n20859 ^ n20856 ;
  assign n20853 = n13696 & n14035 ;
  assign n20861 = n20860 ^ n20853 ;
  assign n20862 = n13534 ^ n8212 ;
  assign n20863 = n20862 ^ n13695 ;
  assign n20864 = n20863 ^ n14032 ;
  assign n20865 = n20864 ^ n20788 ;
  assign n20869 = n20778 ^ n20771 ;
  assign n20870 = n20764 & n20869 ;
  assign n20871 = n20870 ^ n14036 ;
  assign n20866 = n20770 ^ n14037 ;
  assign n20867 = n20770 ^ n14217 ;
  assign n20868 = n20866 & n20867 ;
  assign n20872 = n20871 ^ n20868 ;
  assign n20873 = n14227 ^ n14037 ;
  assign n20874 = n20873 ^ n20770 ;
  assign n20875 = n20874 ^ n14217 ;
  assign n20876 = n20875 ^ n20763 ;
  assign n20880 = n20750 ^ n20740 ;
  assign n20881 = n20880 ^ n20751 ;
  assign n20877 = n20750 ^ n14423 ;
  assign n20878 = n20877 ^ n20737 ;
  assign n20879 = n20724 & ~n20878 ;
  assign n20882 = n20881 ^ n20879 ;
  assign n20883 = n20878 ^ n20723 ;
  assign n21020 = n20699 ^ n14687 ;
  assign n21021 = n20711 ^ n20699 ;
  assign n21022 = n21021 ^ n20702 ;
  assign n21023 = ~n21020 & ~n21022 ;
  assign n21024 = n21023 ^ n14686 ;
  assign n21018 = n20702 ^ n15391 ;
  assign n21019 = n20711 & n21018 ;
  assign n21025 = n21024 ^ n21019 ;
  assign n20884 = n14687 ^ n6070 ;
  assign n20885 = n20884 ^ n20702 ;
  assign n20886 = n20885 ^ n15391 ;
  assign n20887 = n20886 ^ n20699 ;
  assign n20888 = n20688 ^ n20681 ;
  assign n20891 = n20688 ^ n20672 ;
  assign n20892 = n20888 & n20891 ;
  assign n20889 = n20888 ^ n20672 ;
  assign n20890 = n20676 & n20889 ;
  assign n20893 = n20892 ^ n20890 ;
  assign n20894 = n20893 ^ n15408 ;
  assign n20895 = n20688 ^ n20676 ;
  assign n20896 = n20895 ^ n20681 ;
  assign n20897 = n20896 ^ n20672 ;
  assign n20898 = n20670 ^ n20635 ;
  assign n20899 = n16336 ^ n15419 ;
  assign n21006 = n20609 ^ n16232 ;
  assign n21007 = n21006 ^ n20625 ;
  assign n21010 = n20899 & n21007 ;
  assign n21008 = n21007 ^ n20625 ;
  assign n21009 = n20613 & n21008 ;
  assign n21011 = n21010 ^ n21009 ;
  assign n21012 = n21011 ^ n16334 ;
  assign n20900 = n20899 ^ n16232 ;
  assign n20901 = n20900 ^ n20612 ;
  assign n20902 = n20901 ^ n20609 ;
  assign n20903 = n20607 ^ n20601 ;
  assign n20906 = n18170 ^ n18153 ;
  assign n20907 = n20906 ^ n20584 ;
  assign n20908 = n20588 & n20907 ;
  assign n20909 = n20908 ^ n18168 ;
  assign n20904 = n20584 ^ n18125 ;
  assign n20905 = ~n18170 & ~n20904 ;
  assign n20910 = n20909 ^ n20905 ;
  assign n20911 = n20588 ^ n18128 ;
  assign n20912 = n20911 ^ n18125 ;
  assign n20913 = n20912 ^ n20584 ;
  assign n20917 = n20561 ^ n18626 ;
  assign n20914 = n18632 ^ n18625 ;
  assign n20918 = n20914 ^ n20561 ;
  assign n20919 = n20918 ^ n20564 ;
  assign n20920 = ~n20917 & ~n20919 ;
  assign n20921 = n20920 ^ n18638 ;
  assign n20915 = n20564 ^ n18632 ;
  assign n20916 = ~n20914 & n20915 ;
  assign n20922 = n20921 ^ n20916 ;
  assign n20923 = n20922 ^ n20913 ;
  assign n20966 = n20540 ^ n19152 ;
  assign n20967 = n20966 ^ n14315 ;
  assign n20968 = n20967 ^ n20530 ;
  assign n20969 = n20968 ^ n20511 ;
  assign n20970 = n20505 ^ n19681 ;
  assign n20971 = ~n20969 & n20970 ;
  assign n20924 = n20502 ^ n19699 ;
  assign n20925 = n20478 ^ n20462 ;
  assign n20940 = n19721 ^ n19703 ;
  assign n20941 = n20940 ^ n20430 ;
  assign n20926 = n20424 ^ n19756 ;
  assign n20939 = n20428 ^ n19738 ;
  assign n20948 = n20926 & n20939 ;
  assign n20949 = ~n20941 & n20948 ;
  assign n20950 = n20949 ^ n20941 ;
  assign n20951 = ~n20925 & n20950 ;
  assign n20952 = ~n20499 & ~n20951 ;
  assign n20953 = ~n20924 & ~n20952 ;
  assign n20927 = n20421 ^ n19774 ;
  assign n20928 = n20926 & n20927 ;
  assign n20930 = n19755 ^ n19220 ;
  assign n20934 = n19755 ^ n19618 ;
  assign n20935 = n20930 & n20934 ;
  assign n20931 = n20930 ^ n19618 ;
  assign n20932 = ~n19221 & ~n20931 ;
  assign n20929 = n19737 ^ n19212 ;
  assign n20933 = n20932 ^ n20929 ;
  assign n20936 = n20935 ^ n20933 ;
  assign n20937 = n20928 & ~n20936 ;
  assign n20938 = n20937 ^ n20926 ;
  assign n20942 = ~n20939 & n20941 ;
  assign n20943 = ~n20938 & n20942 ;
  assign n20944 = n20943 ^ n20941 ;
  assign n20945 = n20925 & ~n20944 ;
  assign n20946 = n20499 & ~n20945 ;
  assign n20947 = n20924 & ~n20946 ;
  assign n20954 = n20953 ^ n20947 ;
  assign n20955 = n20954 ^ n20924 ;
  assign n20960 = n20540 ^ n20511 ;
  assign n20961 = ~n20541 & n20960 ;
  assign n20956 = n19152 ^ n14315 ;
  assign n20957 = n20550 ^ n20541 ;
  assign n20958 = ~n20956 & ~n20957 ;
  assign n20959 = n20958 ^ n20525 ;
  assign n20962 = n20961 ^ n20959 ;
  assign n20963 = n20508 ^ n19665 ;
  assign n20964 = n20962 & ~n20963 ;
  assign n20965 = n20955 & n20964 ;
  assign n20972 = n20971 ^ n20965 ;
  assign n20973 = n20969 ^ n20962 ;
  assign n20974 = n20969 ^ n20963 ;
  assign n20975 = n20970 ^ n20969 ;
  assign n20976 = n20974 & n20975 ;
  assign n20977 = n20976 ^ n20974 ;
  assign n20978 = n20977 ^ n20963 ;
  assign n20981 = n20977 ^ n20955 ;
  assign n20982 = n20976 & ~n20981 ;
  assign n20983 = n20978 & n20982 ;
  assign n20984 = n20983 ^ n20978 ;
  assign n20985 = n20984 ^ n20963 ;
  assign n20986 = ~n20973 & ~n20985 ;
  assign n20987 = n20986 ^ n20962 ;
  assign n20988 = ~n20924 & ~n20987 ;
  assign n20989 = n20972 & n20988 ;
  assign n20990 = n20989 ^ n20987 ;
  assign n20991 = n20990 ^ n20962 ;
  assign n20992 = n18633 ^ n18625 ;
  assign n20993 = n20992 ^ n20564 ;
  assign n20994 = n20993 ^ n20561 ;
  assign n20995 = n20994 ^ n20922 ;
  assign n20996 = ~n20991 & ~n20995 ;
  assign n20997 = n20990 ^ n20922 ;
  assign n20998 = n20996 & n20997 ;
  assign n20999 = n20998 ^ n20995 ;
  assign n21000 = ~n20923 & n20999 ;
  assign n21001 = n21000 ^ n20913 ;
  assign n21002 = ~n20913 & ~n21001 ;
  assign n21036 = n21002 ^ n21000 ;
  assign n21037 = ~n20910 & n21036 ;
  assign n21038 = n20903 & ~n21037 ;
  assign n21039 = ~n20902 & ~n21038 ;
  assign n21040 = ~n21012 & ~n21039 ;
  assign n21041 = ~n20898 & ~n21040 ;
  assign n21042 = n20897 & ~n21041 ;
  assign n21043 = n20894 & ~n21042 ;
  assign n21044 = ~n20887 & ~n21043 ;
  assign n21045 = n21025 & ~n21044 ;
  assign n21046 = n20883 & ~n21045 ;
  assign n21047 = ~n20882 & ~n21046 ;
  assign n21048 = ~n20876 & ~n21047 ;
  assign n21049 = n20872 & ~n21048 ;
  assign n21050 = n20865 & ~n21049 ;
  assign n21051 = ~n20861 & ~n21050 ;
  assign n21052 = n20852 & ~n21051 ;
  assign n21053 = ~n20836 & ~n21052 ;
  assign n21054 = n20837 & ~n21053 ;
  assign n24003 = ~n20834 & ~n21054 ;
  assign n24462 = ~n24003 & n24079 ;
  assign n24948 = ~n24462 & n24700 ;
  assign n21003 = n20910 & ~n21002 ;
  assign n21004 = ~n20903 & ~n21003 ;
  assign n21005 = n20902 & ~n21004 ;
  assign n21013 = ~n21005 & n21012 ;
  assign n21014 = n20898 & ~n21013 ;
  assign n21015 = ~n20897 & ~n21014 ;
  assign n21016 = ~n20894 & ~n21015 ;
  assign n21017 = n20887 & ~n21016 ;
  assign n21026 = ~n21017 & ~n21025 ;
  assign n21027 = ~n20883 & ~n21026 ;
  assign n21028 = n20882 & ~n21027 ;
  assign n21029 = n20876 & ~n21028 ;
  assign n21030 = ~n20872 & ~n21029 ;
  assign n21031 = ~n20865 & ~n21030 ;
  assign n21032 = n20861 & ~n21031 ;
  assign n21033 = ~n20852 & ~n21032 ;
  assign n21034 = n20836 & ~n21033 ;
  assign n21035 = ~n20837 & ~n21034 ;
  assign n24002 = n20834 & ~n21035 ;
  assign n24461 = ~n24002 & ~n24079 ;
  assign n24947 = ~n24461 & ~n24700 ;
  assign n24949 = n24948 ^ n24947 ;
  assign n24982 = n24981 ^ n24949 ;
  assign n24983 = n24982 ^ n24981 ;
  assign n24984 = n24981 ^ n10828 ;
  assign n24985 = n24984 ^ n24981 ;
  assign n24986 = ~n24983 & n24985 ;
  assign n24987 = n24986 ^ n24981 ;
  assign n24988 = x0 & ~n24987 ;
  assign n24992 = n24991 ^ n24988 ;
  assign n24939 = n9085 & n20837 ;
  assign n24938 = n10131 & n20834 ;
  assign n24940 = n24939 ^ n24938 ;
  assign n24941 = n24940 ^ x5 ;
  assign n21055 = n21054 ^ n21035 ;
  assign n24936 = n21055 ^ n20834 ;
  assign n24937 = n9081 & ~n24936 ;
  assign n24942 = n24941 ^ n24937 ;
  assign n24935 = ~n9092 & n20836 ;
  assign n24943 = n24942 ^ n24935 ;
  assign n22414 = n21044 ^ n21017 ;
  assign n24294 = ~x13 & ~n22414 ;
  assign n24295 = n24294 ^ n21025 ;
  assign n24416 = n6060 & ~n24295 ;
  assign n24414 = ~n6072 & ~n20894 ;
  assign n24412 = ~n6074 & ~n20887 ;
  assign n24407 = n5696 & n20897 ;
  assign n23919 = ~n3520 & ~n20939 ;
  assign n24226 = n20939 ^ x31 ;
  assign n24227 = ~n23919 & n24226 ;
  assign n24222 = ~n35 & n20939 ;
  assign n24221 = n20939 ^ n3722 ;
  assign n24223 = n24222 ^ n24221 ;
  assign n24224 = n24223 ^ x31 ;
  assign n21170 = n20939 ^ n20938 ;
  assign n24218 = x31 & ~n21170 ;
  assign n24219 = n24218 ^ n20941 ;
  assign n24220 = n3520 & n24219 ;
  assign n24225 = n24224 ^ n24220 ;
  assign n24228 = n24227 ^ n24225 ;
  assign n24215 = ~n20926 & n24214 ;
  assign n24229 = n24228 ^ n24215 ;
  assign n24207 = n5115 ^ n4185 ;
  assign n24205 = n768 ^ n540 ;
  assign n24206 = n24205 ^ n2260 ;
  assign n24208 = n24207 ^ n24206 ;
  assign n24202 = n3692 ^ n283 ;
  assign n24201 = n1444 ^ n495 ;
  assign n24203 = n24202 ^ n24201 ;
  assign n24199 = n779 ^ n370 ;
  assign n24196 = n2764 ^ n431 ;
  assign n24197 = n24196 ^ n363 ;
  assign n24198 = n24197 ^ n391 ;
  assign n24200 = n24199 ^ n24198 ;
  assign n24204 = n24203 ^ n24200 ;
  assign n24209 = n24208 ^ n24204 ;
  assign n24210 = n24209 ^ n3789 ;
  assign n24211 = n24210 ^ n5053 ;
  assign n24212 = ~n1112 & ~n1702 ;
  assign n24213 = ~n24211 & n24212 ;
  assign n24230 = n24229 ^ n24213 ;
  assign n23904 = n12797 ^ n2693 ;
  assign n23903 = n865 ^ n131 ;
  assign n23905 = n23904 ^ n23903 ;
  assign n23901 = n1172 ^ n759 ;
  assign n23899 = n790 ^ n356 ;
  assign n23898 = n1001 ^ n143 ;
  assign n23900 = n23899 ^ n23898 ;
  assign n23902 = n23901 ^ n23900 ;
  assign n23906 = n23905 ^ n23902 ;
  assign n23907 = n23906 ^ n3758 ;
  assign n23894 = n13259 ^ n2157 ;
  assign n23895 = n23894 ^ n3768 ;
  assign n23896 = n23895 ^ n4967 ;
  assign n23897 = n23896 ^ n1627 ;
  assign n23908 = n23907 ^ n23897 ;
  assign n23909 = n23908 ^ n6339 ;
  assign n23910 = ~n15028 & ~n23909 ;
  assign n23721 = ~n3720 & ~n20927 ;
  assign n23719 = ~n3520 & ~n20926 ;
  assign n23718 = n20926 ^ n3520 ;
  assign n23720 = n23719 ^ n23718 ;
  assign n23722 = n23721 ^ n23720 ;
  assign n23751 = n2308 ^ n228 ;
  assign n23750 = n3692 ^ n982 ;
  assign n23752 = n23751 ^ n23750 ;
  assign n23748 = n4181 ^ n239 ;
  assign n23746 = n14851 ^ n321 ;
  assign n23747 = n23746 ^ n1219 ;
  assign n23749 = n23748 ^ n23747 ;
  assign n23753 = n23752 ^ n23749 ;
  assign n23742 = n13847 ^ n5354 ;
  assign n23743 = n23742 ^ n3678 ;
  assign n23740 = n2195 ^ n1250 ;
  assign n23739 = n1731 ^ n1722 ;
  assign n23741 = n23740 ^ n23739 ;
  assign n23744 = n23743 ^ n23741 ;
  assign n23735 = n1798 ^ n269 ;
  assign n23736 = n23735 ^ n361 ;
  assign n23737 = n23736 ^ n1611 ;
  assign n23738 = n23737 ^ n15122 ;
  assign n23745 = n23744 ^ n23738 ;
  assign n23754 = n23753 ^ n23745 ;
  assign n23732 = n2506 ^ n1893 ;
  assign n23731 = n3984 ^ n3961 ;
  assign n23733 = n23732 ^ n23731 ;
  assign n23729 = n13631 ^ n4139 ;
  assign n23726 = n1355 ^ n511 ;
  assign n23725 = n550 ^ n450 ;
  assign n23727 = n23726 ^ n23725 ;
  assign n23723 = n13775 ^ n1282 ;
  assign n23724 = n23723 ^ n3331 ;
  assign n23728 = n23727 ^ n23724 ;
  assign n23730 = n23729 ^ n23728 ;
  assign n23734 = n23733 ^ n23730 ;
  assign n23755 = n23754 ^ n23734 ;
  assign n23756 = ~n15027 & ~n23755 ;
  assign n23893 = ~n23722 & ~n23756 ;
  assign n23911 = n23910 ^ n23893 ;
  assign n23922 = ~n3721 & ~n23719 ;
  assign n23918 = n24214 ^ n20939 ;
  assign n23920 = n23919 ^ n23918 ;
  assign n23913 = n20926 ^ n4851 ;
  assign n23914 = n23913 ^ n4851 ;
  assign n23915 = n23912 & ~n23914 ;
  assign n23916 = n23915 ^ n4851 ;
  assign n23917 = n20927 & n23916 ;
  assign n23921 = n23920 ^ n23917 ;
  assign n23923 = n23922 ^ n23921 ;
  assign n24193 = n23923 ^ n23893 ;
  assign n24194 = n23911 & ~n24193 ;
  assign n24195 = n24194 ^ n23923 ;
  assign n24231 = n24230 ^ n24195 ;
  assign n24190 = n3484 & n20499 ;
  assign n21210 = n20952 ^ n20946 ;
  assign n24183 = n20924 ^ x29 ;
  assign n24184 = n24183 ^ x28 ;
  assign n24185 = n24184 ^ n20924 ;
  assign n24186 = ~n21210 & n24185 ;
  assign n24187 = n24186 ^ n20924 ;
  assign n24188 = n650 & ~n24187 ;
  assign n24189 = n24188 ^ x29 ;
  assign n24191 = n24190 ^ n24189 ;
  assign n24182 = n831 & ~n20925 ;
  assign n24192 = n24191 ^ n24182 ;
  assign n24232 = n24231 ^ n24192 ;
  assign n23927 = n3484 & ~n20925 ;
  assign n23924 = n23923 ^ n23911 ;
  assign n23925 = n23924 ^ x29 ;
  assign n21123 = n20951 ^ n20945 ;
  assign n23888 = n20499 ^ n4536 ;
  assign n23889 = n23888 ^ n20499 ;
  assign n23890 = ~n21123 & n23889 ;
  assign n23891 = n23890 ^ n20499 ;
  assign n23892 = n650 & n23891 ;
  assign n23926 = n23925 ^ n23892 ;
  assign n23928 = n23927 ^ n23926 ;
  assign n23887 = n831 & n20941 ;
  assign n23929 = n23928 ^ n23887 ;
  assign n23757 = n23756 ^ n23722 ;
  assign n22617 = n3484 & n20939 ;
  assign n22610 = n20941 ^ x29 ;
  assign n22611 = n22610 ^ x28 ;
  assign n22612 = n22611 ^ n20941 ;
  assign n22613 = n21170 & n22612 ;
  assign n22614 = n22613 ^ n20941 ;
  assign n22615 = n650 & n22614 ;
  assign n22616 = n22615 ^ x29 ;
  assign n22618 = n22617 ^ n22616 ;
  assign n22609 = n831 & n20926 ;
  assign n22619 = n22618 ^ n22609 ;
  assign n21142 = ~n20926 & n20927 ;
  assign n21143 = n21142 ^ n20927 ;
  assign n21144 = n21143 ^ n20939 ;
  assign n22500 = n3481 & n21144 ;
  assign n22499 = n656 & n20939 ;
  assign n22501 = n22500 ^ n22499 ;
  assign n22497 = n831 & ~n20927 ;
  assign n22496 = n3484 & n20926 ;
  assign n22498 = n22497 ^ n22496 ;
  assign n22502 = n22501 ^ n22498 ;
  assign n22390 = n650 & n20926 ;
  assign n22503 = x29 & ~n22390 ;
  assign n22504 = n827 & ~n20927 ;
  assign n22505 = n22503 & n22504 ;
  assign n22506 = n22505 ^ n22503 ;
  assign n22620 = ~n22502 & n22506 ;
  assign n22622 = n3520 & ~n20927 ;
  assign n23715 = ~n22620 & ~n22622 ;
  assign n23716 = n22619 & n23715 ;
  assign n23717 = n23716 ^ n22619 ;
  assign n23758 = n23757 ^ n23717 ;
  assign n23711 = n831 & n20939 ;
  assign n23710 = n3484 & n20941 ;
  assign n23712 = n23711 ^ n23710 ;
  assign n23713 = n23712 ^ n651 ;
  assign n23703 = n20925 ^ x29 ;
  assign n23702 = n20925 ^ x28 ;
  assign n23704 = n23703 ^ n23702 ;
  assign n21187 = n20950 ^ n20944 ;
  assign n23705 = n23703 ^ n21187 ;
  assign n23706 = n23705 ^ n23703 ;
  assign n23707 = n23704 & n23706 ;
  assign n23708 = n23707 ^ n23703 ;
  assign n23709 = n650 & ~n23708 ;
  assign n23714 = n23713 ^ n23709 ;
  assign n23930 = n23717 ^ n23714 ;
  assign n23931 = ~n23758 & n23930 ;
  assign n23932 = n23931 ^ n23714 ;
  assign n24179 = n23932 ^ n23924 ;
  assign n24180 = ~n23929 & n24179 ;
  assign n24181 = n24180 ^ n23932 ;
  assign n24233 = n24232 ^ n24181 ;
  assign n24174 = n12861 & n20970 ;
  assign n24173 = n446 & ~n20963 ;
  assign n24175 = n24174 ^ n24173 ;
  assign n24176 = n24175 ^ x26 ;
  assign n24172 = ~n487 & ~n20969 ;
  assign n24177 = n24176 ^ n24172 ;
  assign n21104 = ~n20953 & ~n20970 ;
  assign n21105 = ~n20963 & ~n21104 ;
  assign n21102 = ~n20947 & n20970 ;
  assign n21103 = n20963 & ~n21102 ;
  assign n21106 = n21105 ^ n21103 ;
  assign n21114 = n21106 ^ n20969 ;
  assign n24171 = ~n3501 & n21114 ;
  assign n24178 = n24177 ^ n24171 ;
  assign n24234 = n24233 ^ n24178 ;
  assign n23933 = n23932 ^ n23929 ;
  assign n23882 = n12861 & ~n20924 ;
  assign n23881 = n446 & n20970 ;
  assign n23883 = n23882 ^ n23881 ;
  assign n23884 = n23883 ^ x26 ;
  assign n23880 = ~n487 & ~n20963 ;
  assign n23885 = n23884 ^ n23880 ;
  assign n21239 = n21104 ^ n21102 ;
  assign n21240 = n21239 ^ n20963 ;
  assign n23879 = ~n3501 & n21240 ;
  assign n23886 = n23885 ^ n23879 ;
  assign n23934 = n23933 ^ n23886 ;
  assign n23759 = n23758 ^ n23714 ;
  assign n23697 = n12861 & n20499 ;
  assign n23696 = n446 & ~n20924 ;
  assign n23698 = n23697 ^ n23696 ;
  assign n23699 = n23698 ^ x26 ;
  assign n23695 = ~n487 & n20970 ;
  assign n23700 = n23699 ^ n23695 ;
  assign n21251 = n20970 ^ n20954 ;
  assign n23694 = ~n3501 & ~n21251 ;
  assign n23701 = n23700 ^ n23694 ;
  assign n23760 = n23759 ^ n23701 ;
  assign n22621 = n22620 ^ n22619 ;
  assign n22623 = n22622 ^ n22621 ;
  assign n22604 = n12861 & ~n20925 ;
  assign n22603 = n446 & n20499 ;
  assign n22605 = n22604 ^ n22603 ;
  assign n22606 = n22605 ^ x26 ;
  assign n22602 = ~n487 & ~n20924 ;
  assign n22607 = n22606 ^ n22602 ;
  assign n21211 = n21210 ^ n20924 ;
  assign n22601 = ~n3501 & n21211 ;
  assign n22608 = n22607 ^ n22601 ;
  assign n22624 = n22623 ^ n22608 ;
  assign n22514 = ~n487 & n20499 ;
  assign n22512 = n12861 & n20941 ;
  assign n22510 = n446 & ~n20925 ;
  assign n22507 = n22506 ^ x29 ;
  assign n22508 = n22507 ^ n22502 ;
  assign n22509 = n22508 ^ x26 ;
  assign n22511 = n22510 ^ n22509 ;
  assign n22513 = n22512 ^ n22511 ;
  assign n22515 = n22514 ^ n22513 ;
  assign n21124 = n21123 ^ n20499 ;
  assign n22495 = ~n3501 & ~n21124 ;
  assign n22516 = n22515 ^ n22495 ;
  assign n22392 = n826 & ~n20927 ;
  assign n22274 = n650 & ~n20927 ;
  assign n21385 = n64 & n20926 ;
  assign n21697 = x26 & ~n21385 ;
  assign n21698 = n7214 & ~n20927 ;
  assign n21699 = n21697 & n21698 ;
  assign n21700 = n21699 ^ n21697 ;
  assign n21707 = ~n3501 & n21144 ;
  assign n21704 = n12861 & ~n20927 ;
  assign n21703 = n446 & n20926 ;
  assign n21705 = n21704 ^ n21703 ;
  assign n21702 = ~n487 & n20939 ;
  assign n21706 = n21705 ^ n21702 ;
  assign n21708 = n21707 ^ n21706 ;
  assign n22275 = n21700 & ~n21708 ;
  assign n22280 = n12861 & n20926 ;
  assign n22279 = n446 & n20939 ;
  assign n22281 = n22280 ^ n22279 ;
  assign n22282 = n22281 ^ x26 ;
  assign n22278 = ~n487 & n20941 ;
  assign n22283 = n22282 ^ n22278 ;
  assign n21172 = n21170 ^ n20941 ;
  assign n22277 = ~n3501 & n21172 ;
  assign n22284 = n22283 ^ n22277 ;
  assign n22387 = ~n22275 & n22284 ;
  assign n22388 = ~n22274 & n22387 ;
  assign n22389 = n22388 ^ n22284 ;
  assign n22391 = n22390 ^ n22389 ;
  assign n22393 = n22392 ^ n22391 ;
  assign n22382 = n12861 & n20939 ;
  assign n22381 = n446 & n20941 ;
  assign n22383 = n22382 ^ n22381 ;
  assign n22384 = n22383 ^ x26 ;
  assign n22380 = ~n487 & ~n20925 ;
  assign n22385 = n22384 ^ n22380 ;
  assign n21188 = n21187 ^ n20925 ;
  assign n22379 = ~n3501 & ~n21188 ;
  assign n22386 = n22385 ^ n22379 ;
  assign n22492 = n22389 ^ n22386 ;
  assign n22493 = ~n22393 & n22492 ;
  assign n22494 = n22493 ^ n22386 ;
  assign n22598 = n22508 ^ n22494 ;
  assign n22599 = n22516 & n22598 ;
  assign n22600 = n22599 ^ n22508 ;
  assign n23761 = n22608 ^ n22600 ;
  assign n23762 = n22624 & n23761 ;
  assign n23763 = n23762 ^ n22608 ;
  assign n23876 = n23763 ^ n23701 ;
  assign n23877 = ~n23760 & n23876 ;
  assign n23878 = n23877 ^ n23763 ;
  assign n24168 = n23886 ^ n23878 ;
  assign n24169 = n23934 & n24168 ;
  assign n24170 = n24169 ^ n23886 ;
  assign n24235 = n24234 ^ n24170 ;
  assign n23775 = ~n4496 & ~n20969 ;
  assign n23772 = n4491 & n20962 ;
  assign n23770 = n4504 & ~n20963 ;
  assign n22625 = n22624 ^ n22600 ;
  assign n22593 = n4504 & n20970 ;
  assign n22592 = n4491 & ~n20969 ;
  assign n22594 = n22593 ^ n22592 ;
  assign n22595 = n22594 ^ x23 ;
  assign n22591 = n4492 & n21114 ;
  assign n22596 = n22595 ^ n22591 ;
  assign n22590 = ~n4496 & ~n20963 ;
  assign n22597 = n22596 ^ n22590 ;
  assign n22626 = n22625 ^ n22597 ;
  assign n22517 = n22516 ^ n22494 ;
  assign n22487 = n4504 & ~n20924 ;
  assign n22486 = n4491 & ~n20963 ;
  assign n22488 = n22487 ^ n22486 ;
  assign n22489 = n22488 ^ x23 ;
  assign n22485 = n4492 & n21240 ;
  assign n22490 = n22489 ^ n22485 ;
  assign n22484 = ~n4496 & n20970 ;
  assign n22491 = n22490 ^ n22484 ;
  assign n22518 = n22517 ^ n22491 ;
  assign n22394 = n22393 ^ n22386 ;
  assign n22374 = n4504 & n20499 ;
  assign n22373 = n4491 & n20970 ;
  assign n22375 = n22374 ^ n22373 ;
  assign n22376 = n22375 ^ x23 ;
  assign n22372 = n4492 & ~n21251 ;
  assign n22377 = n22376 ^ n22372 ;
  assign n22371 = ~n4496 & ~n20924 ;
  assign n22378 = n22377 ^ n22371 ;
  assign n22395 = n22394 ^ n22378 ;
  assign n22276 = n22275 ^ n22274 ;
  assign n22285 = n22284 ^ n22276 ;
  assign n22269 = n4504 & ~n20925 ;
  assign n22268 = n4491 & ~n20924 ;
  assign n22270 = n22269 ^ n22268 ;
  assign n22271 = n22270 ^ x23 ;
  assign n22267 = n4492 & n21211 ;
  assign n22272 = n22271 ^ n22267 ;
  assign n22266 = ~n4496 & n20499 ;
  assign n22273 = n22272 ^ n22266 ;
  assign n22286 = n22285 ^ n22273 ;
  assign n21720 = ~n4496 & ~n20925 ;
  assign n21387 = ~n7434 & ~n20927 ;
  assign n21223 = n64 & ~n20927 ;
  assign n21136 = n4488 & n20926 ;
  assign n21137 = x23 & ~n21136 ;
  assign n21138 = ~n4500 & ~n20927 ;
  assign n21139 = n21137 & n21138 ;
  assign n21140 = n21139 ^ n21137 ;
  assign n21149 = ~n4496 & n20926 ;
  assign n21148 = n4491 & n20939 ;
  assign n21150 = n21149 ^ n21148 ;
  assign n21146 = n4504 & ~n20927 ;
  assign n21145 = n4492 & n21144 ;
  assign n21147 = n21146 ^ n21145 ;
  assign n21151 = n21150 ^ n21147 ;
  assign n21224 = n21140 & ~n21151 ;
  assign n21229 = n4504 & n20926 ;
  assign n21228 = n4491 & n20941 ;
  assign n21230 = n21229 ^ n21228 ;
  assign n21231 = n21230 ^ x23 ;
  assign n21227 = n4492 & n21172 ;
  assign n21232 = n21231 ^ n21227 ;
  assign n21226 = ~n4496 & n20939 ;
  assign n21233 = n21232 ^ n21226 ;
  assign n21382 = ~n21224 & n21233 ;
  assign n21383 = ~n21223 & n21382 ;
  assign n21384 = n21383 ^ n21233 ;
  assign n21386 = n21385 ^ n21384 ;
  assign n21388 = n21387 ^ n21386 ;
  assign n21377 = n4504 & n20939 ;
  assign n21376 = n4491 & ~n20925 ;
  assign n21378 = n21377 ^ n21376 ;
  assign n21379 = n21378 ^ x23 ;
  assign n21375 = n4492 & ~n21188 ;
  assign n21380 = n21379 ^ n21375 ;
  assign n21374 = ~n4496 & n20941 ;
  assign n21381 = n21380 ^ n21374 ;
  assign n21713 = n21384 ^ n21381 ;
  assign n21714 = ~n21388 & n21713 ;
  assign n21715 = n21714 ^ n21381 ;
  assign n21716 = n21715 ^ x23 ;
  assign n21712 = n4504 & n20941 ;
  assign n21717 = n21716 ^ n21712 ;
  assign n21711 = n4491 & n20499 ;
  assign n21718 = n21717 ^ n21711 ;
  assign n21710 = n4492 & ~n21124 ;
  assign n21719 = n21718 ^ n21710 ;
  assign n21721 = n21720 ^ n21719 ;
  assign n21701 = n21700 ^ x26 ;
  assign n21709 = n21708 ^ n21701 ;
  assign n22263 = n21715 ^ n21709 ;
  assign n22264 = n21721 & n22263 ;
  assign n22265 = n22264 ^ n21715 ;
  assign n22368 = n22273 ^ n22265 ;
  assign n22369 = n22286 & n22368 ;
  assign n22370 = n22369 ^ n22273 ;
  assign n22481 = n22378 ^ n22370 ;
  assign n22482 = n22395 & n22481 ;
  assign n22483 = n22482 ^ n22378 ;
  assign n22587 = n22491 ^ n22483 ;
  assign n22588 = n22518 & n22587 ;
  assign n22589 = n22588 ^ n22491 ;
  assign n23766 = n22597 ^ n22589 ;
  assign n23767 = n22626 & n23766 ;
  assign n23768 = n23767 ^ n22597 ;
  assign n23769 = n23768 ^ x23 ;
  assign n23771 = n23770 ^ n23769 ;
  assign n23773 = n23772 ^ n23771 ;
  assign n21107 = n20969 & n21106 ;
  assign n21108 = n21107 ^ n21103 ;
  assign n21109 = n21108 ^ n20962 ;
  assign n23765 = n4492 & n21109 ;
  assign n23774 = n23773 ^ n23765 ;
  assign n23776 = n23775 ^ n23774 ;
  assign n23764 = n23763 ^ n23760 ;
  assign n23936 = n23768 ^ n23764 ;
  assign n23937 = ~n23776 & n23936 ;
  assign n23938 = n23937 ^ n23764 ;
  assign n23935 = n23934 ^ n23878 ;
  assign n23939 = n23938 ^ n23935 ;
  assign n23874 = ~n4496 & n20962 ;
  assign n21394 = n20994 ^ n20962 ;
  assign n21630 = n21394 ^ n20990 ;
  assign n23872 = n4492 & n21630 ;
  assign n23869 = n4504 & ~n20969 ;
  assign n23868 = n4491 & n20994 ;
  assign n23870 = n23869 ^ n23868 ;
  assign n23871 = n23870 ^ x23 ;
  assign n23873 = n23872 ^ n23871 ;
  assign n23875 = n23874 ^ n23873 ;
  assign n24165 = n23938 ^ n23875 ;
  assign n24166 = n23939 & n24165 ;
  assign n24167 = n24166 ^ n23938 ;
  assign n24236 = n24235 ^ n24167 ;
  assign n24162 = ~n4496 & n20994 ;
  assign n21395 = ~n20991 & n21394 ;
  assign n24155 = n20922 ^ x23 ;
  assign n24156 = n24155 ^ x22 ;
  assign n24157 = n24156 ^ n20922 ;
  assign n24158 = n21395 & n24157 ;
  assign n24159 = n24158 ^ n20922 ;
  assign n24160 = n4488 & ~n24159 ;
  assign n24161 = n24160 ^ x23 ;
  assign n24163 = n24162 ^ n24161 ;
  assign n24154 = n4504 & n20962 ;
  assign n24164 = n24163 ^ n24154 ;
  assign n24397 = n24167 ^ n24164 ;
  assign n24398 = ~n24236 & n24397 ;
  assign n24399 = n24398 ^ n24164 ;
  assign n24389 = n24229 ^ n24195 ;
  assign n24390 = ~n24230 & ~n24389 ;
  assign n24391 = n24390 ^ n24229 ;
  assign n24383 = ~n35 & n20941 ;
  assign n24382 = n20941 ^ n3726 ;
  assign n24384 = n24383 ^ n24382 ;
  assign n24378 = n21188 ^ n21187 ;
  assign n24379 = ~n3726 & n24378 ;
  assign n24380 = n24379 ^ n21187 ;
  assign n24381 = ~x31 & ~n24380 ;
  assign n24385 = n24384 ^ n24381 ;
  assign n24371 = n14963 ^ n12458 ;
  assign n24367 = n848 ^ n725 ;
  assign n24368 = n24367 ^ n614 ;
  assign n24365 = n3192 ^ n745 ;
  assign n24366 = n24365 ^ n589 ;
  assign n24369 = n24368 ^ n24366 ;
  assign n24363 = n2262 ^ n1122 ;
  assign n24361 = n13880 ^ n1116 ;
  assign n24362 = n24361 ^ n91 ;
  assign n24364 = n24363 ^ n24362 ;
  assign n24370 = n24369 ^ n24364 ;
  assign n24372 = n24371 ^ n24370 ;
  assign n24373 = n24372 ^ n12441 ;
  assign n24374 = n24373 ^ n12515 ;
  assign n24375 = ~n15077 & ~n24374 ;
  assign n24386 = n24385 ^ n24375 ;
  assign n24359 = n21188 ^ n20941 ;
  assign n24360 = ~n12015 & ~n24359 ;
  assign n24387 = n24386 ^ n24360 ;
  assign n24358 = x31 & n24222 ;
  assign n24388 = n24387 ^ n24358 ;
  assign n24392 = n24391 ^ n24388 ;
  assign n24355 = n3484 & ~n20924 ;
  assign n21456 = n21251 ^ n20970 ;
  assign n24348 = n20970 ^ x29 ;
  assign n24349 = n24348 ^ x28 ;
  assign n24350 = n24349 ^ n20970 ;
  assign n24351 = ~n21456 & n24350 ;
  assign n24352 = n24351 ^ n20970 ;
  assign n24353 = n650 & n24352 ;
  assign n24354 = n24353 ^ x29 ;
  assign n24356 = n24355 ^ n24354 ;
  assign n24347 = n831 & n20499 ;
  assign n24357 = n24356 ^ n24347 ;
  assign n24393 = n24392 ^ n24357 ;
  assign n24344 = n24192 ^ n24181 ;
  assign n24345 = n24232 & n24344 ;
  assign n24346 = n24345 ^ n24192 ;
  assign n24394 = n24393 ^ n24346 ;
  assign n24340 = n24178 ^ n24170 ;
  assign n24341 = n24234 & n24340 ;
  assign n24342 = n24341 ^ n24178 ;
  assign n24335 = n12861 & ~n20963 ;
  assign n24334 = n446 & ~n20969 ;
  assign n24336 = n24335 ^ n24334 ;
  assign n24337 = n24336 ^ x26 ;
  assign n24333 = ~n487 & n20962 ;
  assign n24338 = n24337 ^ n24333 ;
  assign n24332 = ~n3501 & n21109 ;
  assign n24339 = n24338 ^ n24332 ;
  assign n24343 = n24342 ^ n24339 ;
  assign n24395 = n24394 ^ n24343 ;
  assign n24329 = ~n4496 & ~n20922 ;
  assign n21087 = n20999 ^ n20913 ;
  assign n21088 = n21087 ^ n20913 ;
  assign n24322 = n20913 ^ x23 ;
  assign n24323 = n24322 ^ x22 ;
  assign n24324 = n24323 ^ n20913 ;
  assign n24325 = ~n21088 & n24324 ;
  assign n24326 = n24325 ^ n20913 ;
  assign n24327 = n4488 & n24326 ;
  assign n24328 = n24327 ^ x23 ;
  assign n24330 = n24329 ^ n24328 ;
  assign n24321 = n4504 & n20994 ;
  assign n24331 = n24330 ^ n24321 ;
  assign n24396 = n24395 ^ n24331 ;
  assign n24400 = n24399 ^ n24396 ;
  assign n24318 = n14027 & n20910 ;
  assign n21743 = n21038 ^ n21004 ;
  assign n24311 = n20902 ^ x20 ;
  assign n24312 = n24311 ^ x19 ;
  assign n24313 = n24312 ^ n20902 ;
  assign n24314 = ~n21743 & n24313 ;
  assign n24315 = n24314 ^ n20902 ;
  assign n24316 = n4678 & n24315 ;
  assign n24317 = n24316 ^ x20 ;
  assign n24319 = n24318 ^ n24317 ;
  assign n24309 = n4916 & n20903 ;
  assign n24320 = n24319 ^ n24309 ;
  assign n24401 = n24400 ^ n24320 ;
  assign n24237 = n24236 ^ n24164 ;
  assign n24149 = n14027 & n20913 ;
  assign n21755 = n21037 ^ n21003 ;
  assign n21756 = n21755 ^ n20903 ;
  assign n24148 = n4684 & ~n21756 ;
  assign n24150 = n24149 ^ n24148 ;
  assign n24151 = n24150 ^ x20 ;
  assign n24147 = n4683 & n20903 ;
  assign n24152 = n24151 ^ n24147 ;
  assign n24146 = n4916 & n20910 ;
  assign n24153 = n24152 ^ n24146 ;
  assign n24238 = n24237 ^ n24153 ;
  assign n23940 = n23939 ^ n23875 ;
  assign n23865 = n14027 & ~n20922 ;
  assign n21667 = n21000 ^ n20910 ;
  assign n22951 = n21667 ^ n20910 ;
  assign n23858 = n20910 ^ x20 ;
  assign n23859 = n23858 ^ x19 ;
  assign n23860 = n23859 ^ n20910 ;
  assign n23861 = n22951 & n23860 ;
  assign n23862 = n23861 ^ n20910 ;
  assign n23863 = n4678 & n23862 ;
  assign n23864 = n23863 ^ x20 ;
  assign n23866 = n23865 ^ n23864 ;
  assign n23857 = n4916 & n20913 ;
  assign n23867 = n23866 ^ n23857 ;
  assign n23941 = n23940 ^ n23867 ;
  assign n23777 = n23776 ^ n23764 ;
  assign n22581 = n4916 & n20994 ;
  assign n22574 = n20922 ^ x20 ;
  assign n22575 = n22574 ^ x19 ;
  assign n22576 = n22575 ^ n20922 ;
  assign n22577 = n21395 & n22576 ;
  assign n22578 = n22577 ^ n20922 ;
  assign n22579 = n4678 & ~n22578 ;
  assign n22580 = n22579 ^ x20 ;
  assign n22582 = n22581 ^ n22580 ;
  assign n22573 = n14027 & n20962 ;
  assign n22583 = n22582 ^ n22573 ;
  assign n23778 = n23777 ^ n22583 ;
  assign n22627 = n22626 ^ n22589 ;
  assign n22396 = n22395 ^ n22370 ;
  assign n22287 = n22286 ^ n22265 ;
  assign n22260 = n4916 & ~n20963 ;
  assign n22253 = n20969 ^ x20 ;
  assign n22254 = n22253 ^ x19 ;
  assign n22255 = n22254 ^ n20969 ;
  assign n22256 = ~n21106 & n22255 ;
  assign n22257 = n22256 ^ n20969 ;
  assign n22258 = n4678 & ~n22257 ;
  assign n22259 = n22258 ^ x20 ;
  assign n22261 = n22260 ^ n22259 ;
  assign n22252 = n14027 & n20970 ;
  assign n22262 = n22261 ^ n22252 ;
  assign n22288 = n22287 ^ n22262 ;
  assign n21722 = n21721 ^ n21709 ;
  assign n21694 = n4916 & n20970 ;
  assign n21686 = n21240 ^ n20963 ;
  assign n21687 = n20963 ^ x20 ;
  assign n21688 = n21687 ^ x19 ;
  assign n21689 = n21688 ^ n20963 ;
  assign n21690 = ~n21686 & n21689 ;
  assign n21691 = n21690 ^ n20963 ;
  assign n21692 = n4678 & ~n21691 ;
  assign n21693 = n21692 ^ x20 ;
  assign n21695 = n21694 ^ n21693 ;
  assign n21685 = n14027 & ~n20924 ;
  assign n21696 = n21695 ^ n21685 ;
  assign n21723 = n21722 ^ n21696 ;
  assign n21389 = n21388 ^ n21381 ;
  assign n21369 = n14027 & n20499 ;
  assign n21368 = n4684 & ~n21251 ;
  assign n21370 = n21369 ^ n21368 ;
  assign n21371 = n21370 ^ x20 ;
  assign n21367 = n4683 & n20970 ;
  assign n21372 = n21371 ^ n21367 ;
  assign n21366 = n4916 & ~n20924 ;
  assign n21373 = n21372 ^ n21366 ;
  assign n21390 = n21389 ^ n21373 ;
  assign n21225 = n21224 ^ n21223 ;
  assign n21234 = n21233 ^ n21225 ;
  assign n21220 = n4916 & n20499 ;
  assign n21213 = n20924 ^ x20 ;
  assign n21214 = n21213 ^ x19 ;
  assign n21215 = n21214 ^ n20924 ;
  assign n21216 = ~n21210 & n21215 ;
  assign n21217 = n21216 ^ n20924 ;
  assign n21218 = n4678 & ~n21217 ;
  assign n21219 = n21218 ^ x20 ;
  assign n21221 = n21220 ^ n21219 ;
  assign n21209 = n14027 & ~n20925 ;
  assign n21222 = n21221 ^ n21209 ;
  assign n21235 = n21234 ^ n21222 ;
  assign n21141 = n21140 ^ x23 ;
  assign n21152 = n21151 ^ n21141 ;
  assign n21133 = n4916 & ~n20925 ;
  assign n21126 = n20499 ^ x20 ;
  assign n21127 = n21126 ^ x19 ;
  assign n21128 = n21127 ^ n20499 ;
  assign n21129 = ~n21123 & n21128 ;
  assign n21130 = n21129 ^ n20499 ;
  assign n21131 = n4678 & n21130 ;
  assign n21132 = n21131 ^ x20 ;
  assign n21134 = n21133 ^ n21132 ;
  assign n21122 = n14027 & n20941 ;
  assign n21135 = n21134 ^ n21122 ;
  assign n21153 = n21152 ^ n21135 ;
  assign n21197 = n4916 & n20941 ;
  assign n21190 = n20925 ^ x20 ;
  assign n21191 = n21190 ^ x19 ;
  assign n21192 = n21191 ^ n20925 ;
  assign n21193 = n21187 & n21192 ;
  assign n21194 = n21193 ^ n20925 ;
  assign n21195 = n4678 & ~n21194 ;
  assign n21196 = n21195 ^ x20 ;
  assign n21198 = n21197 ^ n21196 ;
  assign n21186 = n14027 & n20939 ;
  assign n21199 = n21198 ^ n21186 ;
  assign n21205 = n21199 ^ n21152 ;
  assign n21154 = n7824 & ~n21142 ;
  assign n21155 = n21143 ^ n20926 ;
  assign n21156 = ~n20939 & ~n21155 ;
  assign n21157 = n21156 ^ n20926 ;
  assign n21158 = n4684 & ~n21157 ;
  assign n21164 = n4683 & n20939 ;
  assign n21161 = n4684 & n20939 ;
  assign n21162 = n21161 ^ n14027 ;
  assign n21163 = ~n20927 & n21162 ;
  assign n21165 = n21164 ^ n21163 ;
  assign n21166 = n21158 & ~n21165 ;
  assign n21167 = n21166 ^ n21165 ;
  assign n21168 = n21154 & ~n21167 ;
  assign n21169 = n21168 ^ n21167 ;
  assign n21176 = n14027 & n20926 ;
  assign n21175 = n4916 & n20939 ;
  assign n21177 = n21176 ^ n21175 ;
  assign n21173 = n4678 & n21172 ;
  assign n21171 = n4683 & n21170 ;
  assign n21174 = n21173 ^ n21171 ;
  assign n21178 = n21177 ^ n21174 ;
  assign n21179 = n4488 & ~n20927 ;
  assign n21180 = n21178 ^ x20 ;
  assign n21181 = ~n21179 & n21180 ;
  assign n21182 = ~n21178 & n21181 ;
  assign n21183 = ~n21169 & n21182 ;
  assign n21184 = n21183 ^ n21181 ;
  assign n21185 = n21184 ^ n21180 ;
  assign n21200 = n21199 ^ n21185 ;
  assign n21202 = ~n7810 & ~n20927 ;
  assign n21201 = n21185 ^ n21136 ;
  assign n21203 = n21202 ^ n21201 ;
  assign n21204 = n21200 & ~n21203 ;
  assign n21206 = n21205 ^ n21204 ;
  assign n21207 = n21153 & n21206 ;
  assign n21208 = n21207 ^ n21152 ;
  assign n21363 = n21222 ^ n21208 ;
  assign n21364 = n21235 & n21363 ;
  assign n21365 = n21364 ^ n21222 ;
  assign n21682 = n21373 ^ n21365 ;
  assign n21683 = n21390 & n21682 ;
  assign n21684 = n21683 ^ n21373 ;
  assign n22249 = n21696 ^ n21684 ;
  assign n22250 = n21723 & n22249 ;
  assign n22251 = n22250 ^ n21696 ;
  assign n22365 = n22262 ^ n22251 ;
  assign n22366 = n22288 & n22365 ;
  assign n22367 = n22366 ^ n22262 ;
  assign n22397 = n22396 ^ n22367 ;
  assign n22362 = n4916 & ~n20969 ;
  assign n21596 = n21109 ^ n20962 ;
  assign n22355 = n20962 ^ x20 ;
  assign n22356 = n22355 ^ x19 ;
  assign n22357 = n22356 ^ n20962 ;
  assign n22358 = n21596 & n22357 ;
  assign n22359 = n22358 ^ n20962 ;
  assign n22360 = n4678 & n22359 ;
  assign n22361 = n22360 ^ x20 ;
  assign n22363 = n22362 ^ n22361 ;
  assign n22354 = n14027 & ~n20963 ;
  assign n22364 = n22363 ^ n22354 ;
  assign n22520 = n22367 ^ n22364 ;
  assign n22521 = ~n22397 & n22520 ;
  assign n22522 = n22521 ^ n22364 ;
  assign n22519 = n22518 ^ n22483 ;
  assign n22523 = n22522 ^ n22519 ;
  assign n22478 = n4916 & n20962 ;
  assign n21631 = n21630 ^ n20994 ;
  assign n22471 = n20994 ^ x20 ;
  assign n22472 = n22471 ^ x19 ;
  assign n22473 = n22472 ^ n20994 ;
  assign n22474 = n21631 & n22473 ;
  assign n22475 = n22474 ^ n20994 ;
  assign n22476 = n4678 & n22475 ;
  assign n22477 = n22476 ^ x20 ;
  assign n22479 = n22478 ^ n22477 ;
  assign n22470 = n14027 & ~n20969 ;
  assign n22480 = n22479 ^ n22470 ;
  assign n22584 = n22522 ^ n22480 ;
  assign n22585 = n22523 & n22584 ;
  assign n22586 = n22585 ^ n22522 ;
  assign n22628 = n22627 ^ n22586 ;
  assign n23692 = n22586 ^ n22583 ;
  assign n23693 = ~n22628 & n23692 ;
  assign n23779 = n23778 ^ n23693 ;
  assign n23788 = n4916 & ~n20922 ;
  assign n23781 = n20913 ^ x20 ;
  assign n23782 = n23781 ^ x19 ;
  assign n23783 = n23782 ^ n20913 ;
  assign n23784 = ~n21088 & n23783 ;
  assign n23785 = n23784 ^ n20913 ;
  assign n23786 = n4678 & n23785 ;
  assign n23787 = n23786 ^ x20 ;
  assign n23789 = n23788 ^ n23787 ;
  assign n23780 = n14027 & n20994 ;
  assign n23790 = n23789 ^ n23780 ;
  assign n23854 = n23790 ^ n23777 ;
  assign n23855 = ~n23779 & n23854 ;
  assign n23856 = n23855 ^ n23790 ;
  assign n24143 = n23867 ^ n23856 ;
  assign n24144 = n23941 & n24143 ;
  assign n24145 = n24144 ^ n23867 ;
  assign n24306 = n24153 ^ n24145 ;
  assign n24307 = n24238 & n24306 ;
  assign n24308 = n24307 ^ n24153 ;
  assign n24402 = n24401 ^ n24308 ;
  assign n24403 = n24402 ^ x17 ;
  assign n21965 = n21041 ^ n21014 ;
  assign n24305 = ~n21965 & n24304 ;
  assign n24404 = n24403 ^ n24305 ;
  assign n21966 = n21965 ^ n20897 ;
  assign n24303 = n17163 & ~n21966 ;
  assign n24405 = n24404 ^ n24303 ;
  assign n24302 = n20731 & ~n21012 ;
  assign n24406 = n24405 ^ n24302 ;
  assign n24408 = n24407 ^ n24406 ;
  assign n24301 = n5700 & n20898 ;
  assign n24409 = n24408 ^ n24301 ;
  assign n24239 = n24238 ^ n24145 ;
  assign n24141 = n20731 & n20902 ;
  assign n21971 = n21040 ^ n21013 ;
  assign n21972 = n21971 ^ n20898 ;
  assign n24139 = n5703 & ~n21972 ;
  assign n24136 = n5700 & ~n21012 ;
  assign n24135 = n5702 & n20898 ;
  assign n24137 = n24136 ^ n24135 ;
  assign n24138 = n24137 ^ x17 ;
  assign n24140 = n24139 ^ n24138 ;
  assign n24142 = n24141 ^ n24140 ;
  assign n24240 = n24239 ^ n24142 ;
  assign n23942 = n23941 ^ n23856 ;
  assign n23852 = n20731 & n20903 ;
  assign n21734 = n21039 ^ n21005 ;
  assign n21735 = n21734 ^ n21012 ;
  assign n23850 = n5703 & n21735 ;
  assign n23847 = n5700 & n20902 ;
  assign n23846 = n5702 & ~n21012 ;
  assign n23848 = n23847 ^ n23846 ;
  assign n23849 = n23848 ^ x17 ;
  assign n23851 = n23850 ^ n23849 ;
  assign n23853 = n23852 ^ n23851 ;
  assign n23943 = n23942 ^ n23853 ;
  assign n23791 = n23790 ^ n23779 ;
  assign n23690 = n20731 & n20910 ;
  assign n21744 = n21743 ^ n20902 ;
  assign n23688 = n5703 & ~n21744 ;
  assign n23685 = n5700 & n20903 ;
  assign n23684 = n5702 & n20902 ;
  assign n23686 = n23685 ^ n23684 ;
  assign n23687 = n23686 ^ x17 ;
  assign n23689 = n23688 ^ n23687 ;
  assign n23691 = n23690 ^ n23689 ;
  assign n23792 = n23791 ^ n23691 ;
  assign n22629 = n22628 ^ n22583 ;
  assign n22571 = n20731 & n20913 ;
  assign n22569 = n5703 & ~n21756 ;
  assign n22566 = n5702 & n20903 ;
  assign n22565 = n5700 & n20910 ;
  assign n22567 = n22566 ^ n22565 ;
  assign n22568 = n22567 ^ x17 ;
  assign n22570 = n22569 ^ n22568 ;
  assign n22572 = n22571 ^ n22570 ;
  assign n22630 = n22629 ^ n22572 ;
  assign n22524 = n22523 ^ n22480 ;
  assign n22468 = n20731 & ~n20922 ;
  assign n22466 = n5703 & n21667 ;
  assign n22463 = n5700 & n20913 ;
  assign n22462 = n5702 & n20910 ;
  assign n22464 = n22463 ^ n22462 ;
  assign n22465 = n22464 ^ x17 ;
  assign n22467 = n22466 ^ n22465 ;
  assign n22469 = n22468 ^ n22467 ;
  assign n22525 = n22524 ^ n22469 ;
  assign n22398 = n22397 ^ n22364 ;
  assign n22351 = n5700 & ~n20922 ;
  assign n22344 = n20913 ^ x17 ;
  assign n22345 = n22344 ^ x16 ;
  assign n22346 = n22345 ^ n20913 ;
  assign n22347 = ~n21088 & n22346 ;
  assign n22348 = n22347 ^ n20913 ;
  assign n22349 = n5693 & n22348 ;
  assign n22350 = n22349 ^ x17 ;
  assign n22352 = n22351 ^ n22350 ;
  assign n22343 = n20731 & n20994 ;
  assign n22353 = n22352 ^ n22343 ;
  assign n22399 = n22398 ^ n22353 ;
  assign n22289 = n22288 ^ n22251 ;
  assign n21724 = n21723 ^ n21684 ;
  assign n21361 = n20731 & ~n20963 ;
  assign n21236 = n21235 ^ n21208 ;
  assign n21117 = n5700 & ~n20963 ;
  assign n21116 = n5702 & ~n20969 ;
  assign n21118 = n21117 ^ n21116 ;
  assign n21119 = n21118 ^ x17 ;
  assign n21115 = n5703 & n21114 ;
  assign n21120 = n21119 ^ n21115 ;
  assign n21113 = n20731 & n20970 ;
  assign n21121 = n21120 ^ n21113 ;
  assign n21237 = n21236 ^ n21121 ;
  assign n21248 = n21206 ^ n21135 ;
  assign n21243 = n5700 & n20970 ;
  assign n21242 = n5702 & ~n20963 ;
  assign n21244 = n21243 ^ n21242 ;
  assign n21245 = n21244 ^ x17 ;
  assign n21241 = n5703 & n21240 ;
  assign n21246 = n21245 ^ n21241 ;
  assign n21238 = n20731 & ~n20924 ;
  assign n21247 = n21246 ^ n21238 ;
  assign n21249 = n21248 ^ n21247 ;
  assign n21259 = n21203 ^ n21199 ;
  assign n21254 = n5700 & ~n20924 ;
  assign n21253 = n5702 & n20970 ;
  assign n21255 = n21254 ^ n21253 ;
  assign n21256 = n21255 ^ x17 ;
  assign n21252 = n5703 & ~n21251 ;
  assign n21257 = n21256 ^ n21252 ;
  assign n21250 = n20499 & n20731 ;
  assign n21258 = n21257 ^ n21250 ;
  assign n21260 = n21259 ^ n21258 ;
  assign n21336 = n5700 & n20499 ;
  assign n21335 = n5702 & ~n20924 ;
  assign n21337 = n21336 ^ n21335 ;
  assign n21338 = n21337 ^ x17 ;
  assign n21334 = n5703 & n21211 ;
  assign n21339 = n21338 ^ n21334 ;
  assign n21333 = n20731 & ~n20925 ;
  assign n21340 = n21339 ^ n21333 ;
  assign n21306 = n5700 & ~n20925 ;
  assign n21305 = n5702 & n20499 ;
  assign n21307 = n21306 ^ n21305 ;
  assign n21308 = n21307 ^ x17 ;
  assign n21304 = n5703 & ~n21124 ;
  assign n21309 = n21308 ^ n21304 ;
  assign n21303 = n20731 & n20941 ;
  assign n21310 = n21309 ^ n21303 ;
  assign n21289 = n8156 & ~n20927 ;
  assign n21288 = n4678 & n20926 ;
  assign n21290 = n21289 ^ n21288 ;
  assign n21261 = n4678 & ~n20927 ;
  assign n21262 = n5693 & n20926 ;
  assign n21263 = x17 & ~n21262 ;
  assign n21264 = ~n20927 & n21263 ;
  assign n21265 = n5705 & n21264 ;
  assign n21266 = n21265 ^ n21263 ;
  assign n21273 = n5700 & n20926 ;
  assign n21272 = n5702 & n20939 ;
  assign n21274 = n21273 ^ n21272 ;
  assign n21270 = n20731 & ~n20927 ;
  assign n21269 = n5703 & n21144 ;
  assign n21271 = n21270 ^ n21269 ;
  assign n21275 = n21274 ^ n21271 ;
  assign n21276 = n21266 & ~n21275 ;
  assign n21277 = ~n21261 & ~n21276 ;
  assign n21281 = n5700 & n20939 ;
  assign n21280 = n5702 & n20941 ;
  assign n21282 = n21281 ^ n21280 ;
  assign n21283 = n21282 ^ x17 ;
  assign n21279 = n5703 & n21172 ;
  assign n21284 = n21283 ^ n21279 ;
  assign n21278 = n20731 & n20926 ;
  assign n21285 = n21284 ^ n21278 ;
  assign n21286 = n21277 & n21285 ;
  assign n21287 = n21286 ^ n21285 ;
  assign n21291 = n21290 ^ n21287 ;
  assign n21295 = n5700 & n20941 ;
  assign n21294 = n5702 & ~n20925 ;
  assign n21296 = n21295 ^ n21294 ;
  assign n21297 = n21296 ^ x17 ;
  assign n21293 = n5703 & ~n21188 ;
  assign n21298 = n21297 ^ n21293 ;
  assign n21292 = n20731 & n20939 ;
  assign n21299 = n21298 ^ n21292 ;
  assign n21300 = n21299 ^ n21287 ;
  assign n21301 = n21291 & n21300 ;
  assign n21302 = n21301 ^ n21287 ;
  assign n21311 = n21310 ^ n21302 ;
  assign n21328 = n21310 ^ n21167 ;
  assign n21312 = n20927 ^ n20926 ;
  assign n21313 = n8214 ^ n4916 ;
  assign n21318 = ~n20927 & ~n21313 ;
  assign n21319 = n21318 ^ n4916 ;
  assign n21320 = ~n21312 & n21319 ;
  assign n21329 = n21328 ^ n21320 ;
  assign n21323 = n21167 ^ n4916 ;
  assign n21324 = n21323 ^ n21313 ;
  assign n21325 = n21320 & n21324 ;
  assign n21326 = n21325 ^ n21313 ;
  assign n21327 = n20926 & ~n21326 ;
  assign n21330 = n21329 ^ n21327 ;
  assign n21331 = n21311 & n21330 ;
  assign n21332 = n21331 ^ n21310 ;
  assign n21341 = n21340 ^ n21332 ;
  assign n21344 = x20 & n21169 ;
  assign n21342 = n21179 ^ n21178 ;
  assign n21343 = n21342 ^ n21340 ;
  assign n21345 = n21344 ^ n21343 ;
  assign n21346 = n21341 & n21345 ;
  assign n21347 = n21346 ^ n21340 ;
  assign n21348 = n21347 ^ n21258 ;
  assign n21349 = n21260 & n21348 ;
  assign n21350 = n21349 ^ n21258 ;
  assign n21351 = n21350 ^ n21247 ;
  assign n21352 = n21249 & n21351 ;
  assign n21353 = n21352 ^ n21247 ;
  assign n21354 = n21353 ^ n21121 ;
  assign n21355 = n21237 & n21354 ;
  assign n21356 = n21355 ^ n21121 ;
  assign n21357 = n21356 ^ x17 ;
  assign n21112 = n5700 & ~n20969 ;
  assign n21358 = n21357 ^ n21112 ;
  assign n21111 = n5702 & n20962 ;
  assign n21359 = n21358 ^ n21111 ;
  assign n21110 = n5703 & n21109 ;
  assign n21360 = n21359 ^ n21110 ;
  assign n21362 = n21361 ^ n21360 ;
  assign n21391 = n21390 ^ n21365 ;
  assign n21679 = n21391 ^ n21356 ;
  assign n21680 = n21362 & n21679 ;
  assign n21681 = n21680 ^ n21356 ;
  assign n21725 = n21724 ^ n21681 ;
  assign n21677 = n20731 & ~n20969 ;
  assign n21675 = n5703 & n21630 ;
  assign n21672 = n5700 & n20962 ;
  assign n21671 = n5702 & n20994 ;
  assign n21673 = n21672 ^ n21671 ;
  assign n21674 = n21673 ^ x17 ;
  assign n21676 = n21675 ^ n21674 ;
  assign n21678 = n21677 ^ n21676 ;
  assign n22246 = n21681 ^ n21678 ;
  assign n22247 = ~n21725 & n22246 ;
  assign n22248 = n22247 ^ n21678 ;
  assign n22290 = n22289 ^ n22248 ;
  assign n22243 = n5700 & n20994 ;
  assign n22236 = n20922 ^ x17 ;
  assign n22237 = n22236 ^ x16 ;
  assign n22238 = n22237 ^ n20922 ;
  assign n22239 = n21395 & n22238 ;
  assign n22240 = n22239 ^ n20922 ;
  assign n22241 = n5693 & ~n22240 ;
  assign n22242 = n22241 ^ x17 ;
  assign n22244 = n22243 ^ n22242 ;
  assign n22235 = n20731 & n20962 ;
  assign n22245 = n22244 ^ n22235 ;
  assign n22340 = n22248 ^ n22245 ;
  assign n22341 = n22290 & n22340 ;
  assign n22342 = n22341 ^ n22248 ;
  assign n22459 = n22353 ^ n22342 ;
  assign n22460 = n22399 & n22459 ;
  assign n22461 = n22460 ^ n22353 ;
  assign n22562 = n22469 ^ n22461 ;
  assign n22563 = n22525 & n22562 ;
  assign n22564 = n22563 ^ n22469 ;
  assign n23681 = n22572 ^ n22564 ;
  assign n23682 = n22630 & n23681 ;
  assign n23683 = n23682 ^ n22572 ;
  assign n23843 = n23691 ^ n23683 ;
  assign n23844 = n23792 & n23843 ;
  assign n23845 = n23844 ^ n23691 ;
  assign n24132 = n23853 ^ n23845 ;
  assign n24133 = n23943 & n24132 ;
  assign n24134 = n24133 ^ n23853 ;
  assign n24298 = n24142 ^ n24134 ;
  assign n24299 = n24240 & n24298 ;
  assign n24300 = n24299 ^ n24142 ;
  assign n24410 = n24409 ^ n24300 ;
  assign n24411 = n24410 ^ x14 ;
  assign n24413 = n24412 ^ n24411 ;
  assign n24415 = n24414 ^ n24413 ;
  assign n24417 = n24416 ^ n24415 ;
  assign n24296 = n24295 ^ n22414 ;
  assign n24297 = n6063 & n24296 ;
  assign n24418 = n24417 ^ n24297 ;
  assign n24241 = n24240 ^ n24134 ;
  assign n24113 = ~n6072 & n20897 ;
  assign n24112 = ~n6074 & ~n20894 ;
  assign n24114 = n24113 ^ n24112 ;
  assign n24115 = n24114 ^ n6060 ;
  assign n24116 = n24115 ^ x14 ;
  assign n24127 = n8465 & ~n20887 ;
  assign n22306 = n21043 ^ n21016 ;
  assign n22307 = n22306 ^ n20887 ;
  assign n24126 = x13 & ~n22307 ;
  assign n24128 = n24127 ^ n24126 ;
  assign n24129 = ~n6063 & n24128 ;
  assign n24124 = n22306 ^ n8465 ;
  assign n24117 = n24114 ^ x14 ;
  assign n24119 = n20887 ^ x13 ;
  assign n24120 = n24119 ^ n20887 ;
  assign n24121 = ~n22306 & ~n24120 ;
  assign n24122 = n24121 ^ n20887 ;
  assign n24123 = ~n24117 & n24122 ;
  assign n24125 = n24124 ^ n24123 ;
  assign n24130 = n24129 ^ n24125 ;
  assign n24131 = ~n24116 & n24130 ;
  assign n24242 = n24241 ^ n24131 ;
  assign n23946 = ~n6072 & n20898 ;
  assign n23945 = ~n6074 & n20897 ;
  assign n23947 = n23946 ^ n23945 ;
  assign n23948 = n23947 ^ n6060 ;
  assign n23949 = n23948 ^ x14 ;
  assign n23966 = n20894 ^ n6063 ;
  assign n23952 = n23947 ^ n6062 ;
  assign n21953 = n21042 ^ n21015 ;
  assign n23956 = n20894 ^ n17542 ;
  assign n23957 = n23956 ^ n20894 ;
  assign n23958 = ~n21953 & ~n23957 ;
  assign n23959 = n23958 ^ n20894 ;
  assign n23960 = ~n23952 & n23959 ;
  assign n23967 = n23966 ^ n23960 ;
  assign n23965 = ~n17542 & ~n21953 ;
  assign n23968 = n23967 ^ n23965 ;
  assign n23969 = ~n23949 & ~n23968 ;
  assign n23944 = n23943 ^ n23845 ;
  assign n23970 = n23969 ^ n23944 ;
  assign n22633 = ~n6072 & n20902 ;
  assign n22632 = ~n6074 & ~n21012 ;
  assign n22634 = n22633 ^ n22632 ;
  assign n22635 = n22634 ^ n6060 ;
  assign n22636 = n22635 ^ x14 ;
  assign n22653 = n20898 ^ n6063 ;
  assign n22640 = n22634 ^ n6062 ;
  assign n22642 = n21972 ^ n20898 ;
  assign n22643 = n20898 ^ n17542 ;
  assign n22644 = n22643 ^ n20898 ;
  assign n22645 = ~n22642 & ~n22644 ;
  assign n22646 = n22645 ^ n20898 ;
  assign n22647 = ~n22640 & ~n22646 ;
  assign n22654 = n22653 ^ n22647 ;
  assign n22652 = ~n17542 & ~n21971 ;
  assign n22655 = n22654 ^ n22652 ;
  assign n22656 = ~n22636 & n22655 ;
  assign n22631 = n22630 ^ n22564 ;
  assign n22657 = n22656 ^ n22631 ;
  assign n23672 = ~n6072 & ~n21012 ;
  assign n23671 = ~n6074 & n20898 ;
  assign n23673 = n23672 ^ n23671 ;
  assign n23674 = n23673 ^ x14 ;
  assign n23665 = n21966 ^ n20897 ;
  assign n23666 = n20897 ^ n4899 ;
  assign n23667 = n23666 ^ n20897 ;
  assign n23668 = ~n23665 & n23667 ;
  assign n23669 = n23668 ^ n20897 ;
  assign n23670 = n4897 & n23669 ;
  assign n23675 = n23674 ^ n23670 ;
  assign n23676 = n23675 ^ n22631 ;
  assign n23677 = n23676 ^ n23675 ;
  assign n22526 = n22525 ^ n22461 ;
  assign n22440 = ~n6072 & n20903 ;
  assign n22439 = ~n6074 & n20902 ;
  assign n22441 = n22440 ^ n22439 ;
  assign n22442 = n22441 ^ n6060 ;
  assign n22443 = n22442 ^ x14 ;
  assign n22455 = n21734 ^ n8465 ;
  assign n22448 = n22441 ^ x14 ;
  assign n22450 = n21012 ^ x13 ;
  assign n22451 = n22450 ^ n21012 ;
  assign n22452 = ~n21734 & ~n22451 ;
  assign n22453 = n22452 ^ n21012 ;
  assign n22454 = ~n22448 & n22453 ;
  assign n22456 = n22455 ^ n22454 ;
  assign n22445 = n8465 & ~n21012 ;
  assign n22444 = x13 & ~n21735 ;
  assign n22446 = n22445 ^ n22444 ;
  assign n22447 = ~n6063 & n22446 ;
  assign n22457 = n22456 ^ n22447 ;
  assign n22458 = ~n22443 & n22457 ;
  assign n22527 = n22526 ^ n22458 ;
  assign n22400 = n22399 ^ n22342 ;
  assign n22325 = ~n6074 & n20903 ;
  assign n22324 = ~n6072 & n20910 ;
  assign n22326 = n22325 ^ n22324 ;
  assign n22327 = n22326 ^ n6060 ;
  assign n22328 = n22327 ^ x14 ;
  assign n22329 = n22326 ^ x14 ;
  assign n22330 = n22329 ^ n6063 ;
  assign n22337 = ~n20902 & n22330 ;
  assign n22333 = ~x13 & ~n22330 ;
  assign n22334 = n22333 ^ n17542 ;
  assign n22335 = ~n21743 & ~n22334 ;
  assign n22336 = n22335 ^ n6063 ;
  assign n22338 = n22337 ^ n22336 ;
  assign n22339 = ~n22328 & ~n22338 ;
  assign n22401 = n22400 ^ n22339 ;
  assign n22291 = n22290 ^ n22245 ;
  assign n22220 = ~n6072 & n20913 ;
  assign n22219 = ~n6074 & n20910 ;
  assign n22221 = n22220 ^ n22219 ;
  assign n22222 = n22221 ^ n6060 ;
  assign n22223 = n22222 ^ x14 ;
  assign n22224 = n22221 ^ x14 ;
  assign n22225 = n22224 ^ n6063 ;
  assign n22232 = ~n20903 & n22225 ;
  assign n22228 = ~x13 & ~n22225 ;
  assign n22229 = n22228 ^ n17542 ;
  assign n22230 = ~n21755 & ~n22229 ;
  assign n22231 = n22230 ^ n6063 ;
  assign n22233 = n22232 ^ n22231 ;
  assign n22234 = ~n22223 & ~n22233 ;
  assign n22292 = n22291 ^ n22234 ;
  assign n21726 = n21725 ^ n21678 ;
  assign n21668 = n21667 ^ x13 ;
  assign n21656 = n21000 ^ n4899 ;
  assign n21657 = n21656 ^ n21000 ;
  assign n21658 = n21656 ^ n6066 ;
  assign n21659 = n21658 ^ n21656 ;
  assign n21660 = n21656 ^ n20922 ;
  assign n21661 = n21660 ^ n21656 ;
  assign n21662 = ~n21659 & ~n21661 ;
  assign n21663 = n21657 & n21662 ;
  assign n21664 = n21663 ^ n21657 ;
  assign n21665 = n21664 ^ n21000 ;
  assign n21666 = ~n8435 & ~n21665 ;
  assign n21669 = n21668 ^ n21666 ;
  assign n21651 = n20910 ^ n6066 ;
  assign n21652 = n21651 ^ n20910 ;
  assign n21653 = n20913 & n21652 ;
  assign n21654 = n21653 ^ n20910 ;
  assign n21655 = ~n4897 & n21654 ;
  assign n21670 = n21669 ^ n21655 ;
  assign n21727 = n21726 ^ n21670 ;
  assign n21392 = n21391 ^ n21362 ;
  assign n21082 = ~n6072 & n20994 ;
  assign n21081 = ~n6074 & ~n20922 ;
  assign n21083 = n21082 ^ n21081 ;
  assign n21084 = n21083 ^ n6060 ;
  assign n21085 = n21084 ^ x14 ;
  assign n21097 = n8465 & n20913 ;
  assign n21096 = x13 & n21087 ;
  assign n21098 = n21097 ^ n21096 ;
  assign n21099 = ~n6063 & n21098 ;
  assign n21094 = n20999 ^ n8465 ;
  assign n21086 = n21083 ^ x14 ;
  assign n21091 = ~x13 & ~n21088 ;
  assign n21092 = n21091 ^ n20913 ;
  assign n21093 = ~n21086 & ~n21092 ;
  assign n21095 = n21094 ^ n21093 ;
  assign n21100 = n21099 ^ n21095 ;
  assign n21101 = ~n21085 & n21100 ;
  assign n21393 = n21392 ^ n21101 ;
  assign n21407 = n21353 ^ n21237 ;
  assign n21396 = ~x13 & n21395 ;
  assign n21397 = n21396 ^ n20922 ;
  assign n21404 = n21397 ^ n21395 ;
  assign n21405 = n6063 & ~n21404 ;
  assign n21400 = ~n6072 & n20962 ;
  assign n21399 = ~n6074 & n20994 ;
  assign n21401 = n21400 ^ n21399 ;
  assign n21402 = n21401 ^ x14 ;
  assign n21398 = n6060 & ~n21397 ;
  assign n21403 = n21402 ^ n21398 ;
  assign n21406 = n21405 ^ n21403 ;
  assign n21408 = n21407 ^ n21406 ;
  assign n21594 = n21347 ^ n21260 ;
  assign n21430 = n21345 ^ n21332 ;
  assign n21411 = ~n6072 & n20970 ;
  assign n21410 = ~n6074 & ~n20963 ;
  assign n21412 = n21411 ^ n21410 ;
  assign n21413 = n21412 ^ n6060 ;
  assign n21414 = n21413 ^ x14 ;
  assign n21425 = n8465 & ~n20969 ;
  assign n21424 = x13 & ~n21114 ;
  assign n21426 = n21425 ^ n21424 ;
  assign n21427 = ~n6063 & n21426 ;
  assign n21422 = n21106 ^ n8465 ;
  assign n21415 = n21412 ^ x14 ;
  assign n21417 = n20969 ^ x13 ;
  assign n21418 = n21417 ^ n20969 ;
  assign n21419 = ~n21106 & ~n21418 ;
  assign n21420 = n21419 ^ n20969 ;
  assign n21421 = ~n21415 & n21420 ;
  assign n21423 = n21422 ^ n21421 ;
  assign n21428 = n21427 ^ n21423 ;
  assign n21429 = ~n21414 & n21428 ;
  assign n21431 = n21430 ^ n21429 ;
  assign n21447 = n21330 ^ n21302 ;
  assign n21433 = ~n6072 & ~n20924 ;
  assign n21432 = ~n6074 & n20970 ;
  assign n21434 = n21433 ^ n21432 ;
  assign n21435 = n21434 ^ n6060 ;
  assign n21436 = n21435 ^ x14 ;
  assign n21437 = n21434 ^ n6062 ;
  assign n21444 = n20963 & n21437 ;
  assign n21440 = ~x13 & ~n21437 ;
  assign n21441 = n21440 ^ n17542 ;
  assign n21442 = ~n21239 & ~n21441 ;
  assign n21443 = n21442 ^ n6063 ;
  assign n21445 = n21444 ^ n21443 ;
  assign n21446 = ~n21436 & ~n21445 ;
  assign n21448 = n21447 ^ n21446 ;
  assign n21465 = n21299 ^ n21291 ;
  assign n21450 = ~n6072 & n20499 ;
  assign n21449 = ~n6074 & ~n20924 ;
  assign n21451 = n21450 ^ n21449 ;
  assign n21452 = n21451 ^ n6060 ;
  assign n21453 = n21452 ^ x14 ;
  assign n21454 = n21451 ^ x14 ;
  assign n21455 = n21454 ^ n6063 ;
  assign n21457 = n20970 ^ x13 ;
  assign n21458 = n21457 ^ n21454 ;
  assign n21459 = n21458 ^ n20970 ;
  assign n21460 = ~n21456 & n21459 ;
  assign n21461 = n21460 ^ n20970 ;
  assign n21462 = n21455 & ~n21461 ;
  assign n21463 = n21462 ^ n6063 ;
  assign n21464 = ~n21453 & ~n21463 ;
  assign n21466 = n21465 ^ n21464 ;
  assign n21479 = n21276 ^ n21261 ;
  assign n21480 = n21479 ^ n21285 ;
  assign n21474 = ~n6074 & n20499 ;
  assign n21473 = n6060 & ~n21210 ;
  assign n21475 = n21474 ^ n21473 ;
  assign n21476 = n21475 ^ x14 ;
  assign n21472 = ~n6072 & ~n20925 ;
  assign n21477 = n21476 ^ n21472 ;
  assign n21467 = n20924 ^ x13 ;
  assign n21468 = n21467 ^ n20924 ;
  assign n21469 = ~n21210 & n21468 ;
  assign n21470 = n21469 ^ n20924 ;
  assign n21471 = n4897 & ~n21470 ;
  assign n21478 = n21477 ^ n21471 ;
  assign n21481 = n21480 ^ n21478 ;
  assign n21267 = n21266 ^ x17 ;
  assign n21558 = n21275 ^ n21267 ;
  assign n21534 = n5698 & ~n20927 ;
  assign n21482 = n5693 & ~n20927 ;
  assign n21484 = ~n6072 & n20926 ;
  assign n21483 = ~n6074 & n20939 ;
  assign n21485 = n21484 ^ n21483 ;
  assign n21486 = n21485 ^ n6060 ;
  assign n21487 = n21486 ^ x14 ;
  assign n21497 = n6063 & ~n21170 ;
  assign n21488 = n21485 ^ n6062 ;
  assign n21492 = n20941 ^ x13 ;
  assign n21493 = n21492 ^ n20941 ;
  assign n21494 = n21170 & ~n21493 ;
  assign n21495 = n21494 ^ n20941 ;
  assign n21496 = n21488 & ~n21495 ;
  assign n21498 = n21497 ^ n21496 ;
  assign n21499 = ~n21487 & ~n21498 ;
  assign n21501 = ~n6072 & ~n20927 ;
  assign n21500 = ~n6074 & n20926 ;
  assign n21502 = n21501 ^ n21500 ;
  assign n21503 = n21502 ^ n6060 ;
  assign n21504 = n21503 ^ x14 ;
  assign n21520 = n20939 ^ n6063 ;
  assign n21508 = n21502 ^ n6062 ;
  assign n21509 = n21144 ^ n20939 ;
  assign n21510 = n20939 ^ n17542 ;
  assign n21511 = n21510 ^ n20939 ;
  assign n21512 = n21509 & ~n21511 ;
  assign n21513 = n21512 ^ n20939 ;
  assign n21514 = ~n21508 & ~n21513 ;
  assign n21521 = n21520 ^ n21514 ;
  assign n21519 = ~n17542 & n21143 ;
  assign n21522 = n21521 ^ n21519 ;
  assign n21523 = ~n21504 & n21522 ;
  assign n21524 = n4897 & n20926 ;
  assign n21525 = x14 & ~n21524 ;
  assign n21526 = ~n15382 & ~n20927 ;
  assign n21527 = n21525 & n21526 ;
  assign n21528 = n21527 ^ n21525 ;
  assign n21529 = ~n21523 & n21528 ;
  assign n21530 = ~n21499 & ~n21529 ;
  assign n21531 = ~n21482 & n21530 ;
  assign n21532 = n21531 ^ n21499 ;
  assign n21533 = n21532 ^ n21262 ;
  assign n21535 = n21534 ^ n21533 ;
  assign n21537 = ~n6072 & n20939 ;
  assign n21536 = ~n6074 & n20941 ;
  assign n21538 = n21537 ^ n21536 ;
  assign n21539 = n21538 ^ n6060 ;
  assign n21540 = n21539 ^ x14 ;
  assign n21550 = n8465 & ~n20925 ;
  assign n21549 = x13 & n21188 ;
  assign n21551 = n21550 ^ n21549 ;
  assign n21552 = ~n6063 & n21551 ;
  assign n21547 = n21187 ^ n8465 ;
  assign n21541 = n21538 ^ x14 ;
  assign n21542 = n20925 ^ x13 ;
  assign n21543 = n21542 ^ n20925 ;
  assign n21544 = n21187 & ~n21543 ;
  assign n21545 = n21544 ^ n20925 ;
  assign n21546 = ~n21541 & n21545 ;
  assign n21548 = n21547 ^ n21546 ;
  assign n21553 = n21552 ^ n21548 ;
  assign n21554 = ~n21540 & ~n21553 ;
  assign n21555 = n21554 ^ n21532 ;
  assign n21556 = n21535 & n21555 ;
  assign n21557 = n21556 ^ n21554 ;
  assign n21559 = n21558 ^ n21557 ;
  assign n21561 = ~n6072 & n20941 ;
  assign n21560 = ~n6074 & ~n20925 ;
  assign n21562 = n21561 ^ n21560 ;
  assign n21563 = n21562 ^ n6060 ;
  assign n21564 = n21563 ^ x14 ;
  assign n21574 = n8465 & n20499 ;
  assign n21573 = x13 & n21124 ;
  assign n21575 = n21574 ^ n21573 ;
  assign n21576 = ~n6063 & n21575 ;
  assign n21571 = n21123 ^ n8465 ;
  assign n21565 = n21562 ^ x14 ;
  assign n21566 = n20499 ^ x13 ;
  assign n21567 = n21566 ^ n20499 ;
  assign n21568 = ~n21123 & ~n21567 ;
  assign n21569 = n21568 ^ n20499 ;
  assign n21570 = ~n21565 & ~n21569 ;
  assign n21572 = n21571 ^ n21570 ;
  assign n21577 = n21576 ^ n21572 ;
  assign n21578 = ~n21564 & n21577 ;
  assign n21579 = n21578 ^ n21558 ;
  assign n21580 = ~n21559 & ~n21579 ;
  assign n21581 = n21580 ^ n21558 ;
  assign n21582 = n21581 ^ n21478 ;
  assign n21583 = n21481 & ~n21582 ;
  assign n21584 = n21583 ^ n21480 ;
  assign n21585 = n21584 ^ n21464 ;
  assign n21586 = ~n21466 & ~n21585 ;
  assign n21587 = n21586 ^ n21464 ;
  assign n21588 = n21587 ^ n21446 ;
  assign n21589 = ~n21448 & n21588 ;
  assign n21590 = n21589 ^ n21446 ;
  assign n21591 = n21590 ^ n21429 ;
  assign n21592 = ~n21431 & n21591 ;
  assign n21593 = n21592 ^ n21429 ;
  assign n21595 = n21594 ^ n21593 ;
  assign n21603 = ~n6072 & ~n20963 ;
  assign n21602 = ~n6074 & ~n20969 ;
  assign n21604 = n21603 ^ n21602 ;
  assign n21605 = n21604 ^ x14 ;
  assign n21606 = n21604 ^ n16242 ;
  assign n21607 = x14 & ~n21606 ;
  assign n21597 = n20962 ^ x13 ;
  assign n21598 = n21597 ^ n20962 ;
  assign n21608 = n21596 & ~n21598 ;
  assign n21609 = n21608 ^ n20962 ;
  assign n21610 = n21607 & ~n21609 ;
  assign n21611 = n21610 ^ n21606 ;
  assign n21612 = n21605 & n21611 ;
  assign n21599 = n21596 & n21598 ;
  assign n21600 = n21599 ^ n20962 ;
  assign n21601 = n6063 & n21600 ;
  assign n21613 = n21612 ^ n21601 ;
  assign n21614 = n21613 ^ n21593 ;
  assign n21615 = ~n21595 & ~n21614 ;
  assign n21616 = n21615 ^ n21593 ;
  assign n21409 = n21350 ^ n21249 ;
  assign n21617 = n21616 ^ n21409 ;
  assign n21626 = ~n6072 & ~n20969 ;
  assign n21625 = ~n6074 & n20962 ;
  assign n21627 = n21626 ^ n21625 ;
  assign n21628 = ~n6061 & ~n21627 ;
  assign n21629 = n21627 ^ x14 ;
  assign n21618 = n20994 ^ x13 ;
  assign n21619 = n21618 ^ n20994 ;
  assign n21634 = ~n21619 & n21631 ;
  assign n21635 = n21634 ^ n20994 ;
  assign n21636 = n21629 & n21635 ;
  assign n21637 = n21628 & n21636 ;
  assign n21638 = n21637 ^ n21629 ;
  assign n21620 = n20994 ^ n20991 ;
  assign n21621 = n21620 ^ n20994 ;
  assign n21622 = n21619 & n21621 ;
  assign n21623 = n21622 ^ n20994 ;
  assign n21624 = n6063 & n21623 ;
  assign n21639 = n21638 ^ n21624 ;
  assign n21640 = n21639 ^ n21616 ;
  assign n21641 = ~n21617 & ~n21640 ;
  assign n21642 = n21641 ^ n21616 ;
  assign n21643 = n21642 ^ n21406 ;
  assign n21644 = n21408 & n21643 ;
  assign n21645 = n21644 ^ n21407 ;
  assign n21646 = n21645 ^ n21101 ;
  assign n21647 = ~n21393 & ~n21646 ;
  assign n21648 = n21647 ^ n21101 ;
  assign n22216 = n21670 ^ n21648 ;
  assign n22217 = n21727 & n22216 ;
  assign n22218 = n22217 ^ n21648 ;
  assign n22321 = n22234 ^ n22218 ;
  assign n22322 = ~n22292 & n22321 ;
  assign n22323 = n22322 ^ n22234 ;
  assign n22436 = n22339 ^ n22323 ;
  assign n22437 = ~n22401 & n22436 ;
  assign n22438 = n22437 ^ n22339 ;
  assign n22559 = n22458 ^ n22438 ;
  assign n22560 = ~n22527 & n22559 ;
  assign n22561 = n22560 ^ n22458 ;
  assign n23678 = n23677 ^ n22561 ;
  assign n23679 = ~n22657 & ~n23678 ;
  assign n23680 = n23679 ^ n23676 ;
  assign n23793 = n23792 ^ n23683 ;
  assign n23840 = n23793 ^ n23675 ;
  assign n23841 = ~n23680 & n23840 ;
  assign n23842 = n23841 ^ n23793 ;
  assign n24109 = n23944 ^ n23842 ;
  assign n24110 = ~n23970 & n24109 ;
  assign n24111 = n24110 ^ n23944 ;
  assign n24291 = n24241 ^ n24111 ;
  assign n24292 = ~n24242 & n24291 ;
  assign n24293 = n24292 ^ n24241 ;
  assign n24419 = n24418 ^ n24293 ;
  assign n22671 = n21046 ^ n21027 ;
  assign n22672 = n22671 ^ n20882 ;
  assign n24247 = n15413 & ~n22672 ;
  assign n24243 = n24242 ^ n24111 ;
  assign n24244 = n24243 ^ x11 ;
  assign n24108 = n6658 & n20882 ;
  assign n24245 = n24244 ^ n24108 ;
  assign n24107 = n6655 & ~n21025 ;
  assign n24246 = n24245 ^ n24107 ;
  assign n24248 = n24247 ^ n24246 ;
  assign n24106 = n6650 & n20883 ;
  assign n24249 = n24248 ^ n24106 ;
  assign n24284 = n6650 & n20882 ;
  assign n23009 = n21047 ^ n21028 ;
  assign n23010 = n23009 ^ n20876 ;
  assign n24282 = n15413 & n23010 ;
  assign n24279 = n6655 & n20883 ;
  assign n24278 = n6658 & ~n20876 ;
  assign n24280 = n24279 ^ n24278 ;
  assign n24281 = n24280 ^ x11 ;
  assign n24283 = n24282 ^ n24281 ;
  assign n24285 = n24284 ^ n24283 ;
  assign n24286 = n24285 ^ n24243 ;
  assign n23973 = n6655 & ~n20887 ;
  assign n23972 = n6650 & ~n21025 ;
  assign n23974 = n23973 ^ n23972 ;
  assign n23975 = n23974 ^ n6656 ;
  assign n23976 = n23975 ^ x11 ;
  assign n23977 = n23974 ^ x11 ;
  assign n23981 = n23977 ^ n6657 ;
  assign n22545 = n21045 ^ n21026 ;
  assign n23982 = ~x10 & ~n22545 ;
  assign n23983 = n23981 & n23982 ;
  assign n22546 = n22545 ^ n20883 ;
  assign n23979 = n6657 & ~n22546 ;
  assign n23978 = ~n20883 & n23977 ;
  assign n23980 = n23979 ^ n23978 ;
  assign n23984 = n23983 ^ n23980 ;
  assign n23985 = ~n23976 & ~n23984 ;
  assign n23971 = n23970 ^ n23842 ;
  assign n23986 = n23985 ^ n23971 ;
  assign n23660 = n6650 & ~n20887 ;
  assign n22415 = n22414 ^ n21025 ;
  assign n23652 = n22415 ^ n21025 ;
  assign n23653 = n22415 ^ x11 ;
  assign n23654 = n23653 ^ x10 ;
  assign n23655 = n23654 ^ n22415 ;
  assign n23656 = ~n23652 & ~n23655 ;
  assign n23657 = n23656 ^ n22415 ;
  assign n23658 = n6648 & n23657 ;
  assign n23659 = n23658 ^ x11 ;
  assign n23661 = n23660 ^ n23659 ;
  assign n23651 = n6655 & ~n20894 ;
  assign n23662 = n23661 ^ n23651 ;
  assign n22658 = n22657 ^ n22561 ;
  assign n23663 = n23662 ^ n22658 ;
  assign n22662 = n15413 & n22307 ;
  assign n22659 = n22658 ^ x11 ;
  assign n22558 = n6658 & ~n20887 ;
  assign n22660 = n22659 ^ n22558 ;
  assign n22557 = n6655 & n20897 ;
  assign n22661 = n22660 ^ n22557 ;
  assign n22663 = n22662 ^ n22661 ;
  assign n22556 = n6650 & ~n20894 ;
  assign n22664 = n22663 ^ n22556 ;
  assign n21954 = n21953 ^ n20894 ;
  assign n22534 = n15413 & n21954 ;
  assign n22532 = n6655 & n20898 ;
  assign n22530 = n6658 & ~n20894 ;
  assign n22528 = n22527 ^ n22438 ;
  assign n22529 = n22528 ^ x11 ;
  assign n22531 = n22530 ^ n22529 ;
  assign n22533 = n22532 ^ n22531 ;
  assign n22535 = n22534 ^ n22533 ;
  assign n22435 = n6650 & n20897 ;
  assign n22536 = n22535 ^ n22435 ;
  assign n22410 = n6650 & n20898 ;
  assign n22407 = n6649 & ~n21965 ;
  assign n22406 = n6656 & ~n21966 ;
  assign n22408 = n22407 ^ n22406 ;
  assign n22402 = n22401 ^ n22323 ;
  assign n22403 = n22402 ^ x11 ;
  assign n22320 = n6655 & ~n21012 ;
  assign n22404 = n22403 ^ n22320 ;
  assign n22319 = n6657 & n20897 ;
  assign n22405 = n22404 ^ n22319 ;
  assign n22409 = n22408 ^ n22405 ;
  assign n22411 = n22410 ^ n22409 ;
  assign n22299 = n15413 & ~n21972 ;
  assign n22297 = n6655 & n20902 ;
  assign n22295 = n6658 & n20898 ;
  assign n22293 = n22292 ^ n22218 ;
  assign n22294 = n22293 ^ x11 ;
  assign n22296 = n22295 ^ n22294 ;
  assign n22298 = n22297 ^ n22296 ;
  assign n22300 = n22299 ^ n22298 ;
  assign n22215 = n6650 & ~n21012 ;
  assign n22301 = n22300 ^ n22215 ;
  assign n21736 = n15413 & n21735 ;
  assign n21732 = n6655 & n20903 ;
  assign n21730 = n6658 & ~n21012 ;
  assign n21728 = n21727 ^ n21648 ;
  assign n21729 = n21728 ^ x11 ;
  assign n21731 = n21730 ^ n21729 ;
  assign n21733 = n21732 ^ n21731 ;
  assign n21737 = n21736 ^ n21733 ;
  assign n21080 = n6650 & n20902 ;
  assign n21738 = n21737 ^ n21080 ;
  assign n21749 = n21645 ^ n21393 ;
  assign n21747 = n6650 & n20903 ;
  assign n21745 = n15413 & ~n21744 ;
  assign n21740 = n6655 & n20910 ;
  assign n21739 = n6658 & n20902 ;
  assign n21741 = n21740 ^ n21739 ;
  assign n21742 = n21741 ^ x11 ;
  assign n21746 = n21745 ^ n21742 ;
  assign n21748 = n21747 ^ n21746 ;
  assign n21750 = n21749 ^ n21748 ;
  assign n21761 = n21642 ^ n21408 ;
  assign n21759 = n6650 & n20910 ;
  assign n21757 = n15413 & ~n21756 ;
  assign n21752 = n6655 & n20913 ;
  assign n21751 = n6658 & n20903 ;
  assign n21753 = n21752 ^ n21751 ;
  assign n21754 = n21753 ^ x11 ;
  assign n21758 = n21757 ^ n21754 ;
  assign n21760 = n21759 ^ n21758 ;
  assign n21762 = n21761 ^ n21760 ;
  assign n21771 = n21639 ^ n21617 ;
  assign n21769 = n6650 & n20913 ;
  assign n21767 = n15413 & n21667 ;
  assign n21764 = n6655 & ~n20922 ;
  assign n21763 = n6658 & n20910 ;
  assign n21765 = n21764 ^ n21763 ;
  assign n21766 = n21765 ^ x11 ;
  assign n21768 = n21767 ^ n21766 ;
  assign n21770 = n21769 ^ n21768 ;
  assign n21772 = n21771 ^ n21770 ;
  assign n21781 = n21613 ^ n21595 ;
  assign n21779 = n6650 & ~n20922 ;
  assign n21777 = n15413 & ~n21087 ;
  assign n21774 = n6655 & n20994 ;
  assign n21773 = n6658 & n20913 ;
  assign n21775 = n21774 ^ n21773 ;
  assign n21776 = n21775 ^ x11 ;
  assign n21778 = n21777 ^ n21776 ;
  assign n21780 = n21779 ^ n21778 ;
  assign n21782 = n21781 ^ n21780 ;
  assign n21917 = n21590 ^ n21431 ;
  assign n21911 = n6650 & n20962 ;
  assign n21909 = n15413 & n21630 ;
  assign n21907 = n6658 & n20994 ;
  assign n21905 = n6655 & ~n20969 ;
  assign n21792 = n21581 ^ n21481 ;
  assign n21787 = n6655 & n20970 ;
  assign n21786 = n6658 & ~n20969 ;
  assign n21788 = n21787 ^ n21786 ;
  assign n21789 = n21788 ^ x11 ;
  assign n21785 = n15413 & n21114 ;
  assign n21790 = n21789 ^ n21785 ;
  assign n21784 = n6650 & ~n20963 ;
  assign n21791 = n21790 ^ n21784 ;
  assign n21793 = n21792 ^ n21791 ;
  assign n21802 = n21579 ^ n21557 ;
  assign n21797 = n6655 & ~n20924 ;
  assign n21796 = n6658 & ~n20963 ;
  assign n21798 = n21797 ^ n21796 ;
  assign n21799 = n21798 ^ x11 ;
  assign n21795 = n15413 & n21240 ;
  assign n21800 = n21799 ^ n21795 ;
  assign n21794 = n6650 & n20970 ;
  assign n21801 = n21800 ^ n21794 ;
  assign n21803 = n21802 ^ n21801 ;
  assign n21812 = n21554 ^ n21535 ;
  assign n21807 = n6655 & n20499 ;
  assign n21806 = n6658 & n20970 ;
  assign n21808 = n21807 ^ n21806 ;
  assign n21809 = n21808 ^ x11 ;
  assign n21805 = n15413 & ~n21251 ;
  assign n21810 = n21809 ^ n21805 ;
  assign n21804 = n6650 & ~n20924 ;
  assign n21811 = n21810 ^ n21804 ;
  assign n21813 = n21812 ^ n21811 ;
  assign n21822 = n21529 ^ n21482 ;
  assign n21823 = n21822 ^ n21499 ;
  assign n21817 = n6655 & ~n20925 ;
  assign n21816 = n6658 & ~n20924 ;
  assign n21818 = n21817 ^ n21816 ;
  assign n21819 = n21818 ^ x11 ;
  assign n21815 = n15413 & n21211 ;
  assign n21820 = n21819 ^ n21815 ;
  assign n21814 = n6650 & n20499 ;
  assign n21821 = n21820 ^ n21814 ;
  assign n21824 = n21823 ^ n21821 ;
  assign n21867 = n21528 ^ n21523 ;
  assign n21833 = n4897 & ~n20927 ;
  assign n21834 = ~n16289 & ~n21142 ;
  assign n21835 = n20939 ^ n6655 ;
  assign n21836 = n21835 ^ n6655 ;
  assign n21837 = n15413 & n21836 ;
  assign n21838 = n21837 ^ n6655 ;
  assign n21839 = ~n20927 & n21838 ;
  assign n21840 = n6648 & ~n21839 ;
  assign n21841 = n21157 ^ n20939 ;
  assign n21842 = n20939 ^ n9154 ;
  assign n21843 = n21842 ^ n20939 ;
  assign n21844 = ~n21841 & n21843 ;
  assign n21845 = n21844 ^ n20939 ;
  assign n21846 = n21840 & n21845 ;
  assign n21847 = n21846 ^ n21839 ;
  assign n21848 = x11 & ~n21847 ;
  assign n21849 = ~n21834 & n21848 ;
  assign n21850 = ~n21833 & ~n21849 ;
  assign n21854 = n6655 & n20926 ;
  assign n21853 = n6658 & n20941 ;
  assign n21855 = n21854 ^ n21853 ;
  assign n21856 = n21855 ^ x11 ;
  assign n21852 = n15413 & n21172 ;
  assign n21857 = n21856 ^ n21852 ;
  assign n21851 = n6650 & n20939 ;
  assign n21858 = n21857 ^ n21851 ;
  assign n21859 = n21850 & n21858 ;
  assign n21860 = n21859 ^ n21858 ;
  assign n21828 = n6655 & n20939 ;
  assign n21827 = n6658 & ~n20925 ;
  assign n21829 = n21828 ^ n21827 ;
  assign n21830 = n21829 ^ x11 ;
  assign n21826 = n15413 & ~n21188 ;
  assign n21831 = n21830 ^ n21826 ;
  assign n21825 = n6650 & n20941 ;
  assign n21832 = n21831 ^ n21825 ;
  assign n21861 = n21860 ^ n21832 ;
  assign n21863 = ~n6056 & ~n20927 ;
  assign n21862 = n21860 ^ n21524 ;
  assign n21864 = n21863 ^ n21862 ;
  assign n21865 = n21861 & n21864 ;
  assign n21866 = n21865 ^ n21860 ;
  assign n21868 = n21867 ^ n21866 ;
  assign n21872 = n6655 & n20941 ;
  assign n21871 = n6658 & n20499 ;
  assign n21873 = n21872 ^ n21871 ;
  assign n21874 = n21873 ^ x11 ;
  assign n21870 = n15413 & ~n21124 ;
  assign n21875 = n21874 ^ n21870 ;
  assign n21869 = n6650 & ~n20925 ;
  assign n21876 = n21875 ^ n21869 ;
  assign n21877 = n21876 ^ n21866 ;
  assign n21878 = n21868 & n21877 ;
  assign n21879 = n21878 ^ n21876 ;
  assign n21880 = n21879 ^ n21821 ;
  assign n21881 = ~n21824 & n21880 ;
  assign n21882 = n21881 ^ n21821 ;
  assign n21883 = n21882 ^ n21811 ;
  assign n21884 = n21813 & n21883 ;
  assign n21885 = n21884 ^ n21811 ;
  assign n21886 = n21885 ^ n21801 ;
  assign n21887 = n21803 & n21886 ;
  assign n21888 = n21887 ^ n21801 ;
  assign n21889 = n21888 ^ n21791 ;
  assign n21890 = n21793 & n21889 ;
  assign n21891 = n21890 ^ n21791 ;
  assign n21783 = n21584 ^ n21466 ;
  assign n21892 = n21891 ^ n21783 ;
  assign n21900 = n6650 & ~n20969 ;
  assign n21896 = n21891 ^ x11 ;
  assign n21895 = n6655 & ~n20963 ;
  assign n21897 = n21896 ^ n21895 ;
  assign n21894 = n6658 & n20962 ;
  assign n21898 = n21897 ^ n21894 ;
  assign n21893 = n15413 & n21109 ;
  assign n21899 = n21898 ^ n21893 ;
  assign n21901 = n21900 ^ n21899 ;
  assign n21902 = ~n21892 & n21901 ;
  assign n21903 = n21902 ^ n21891 ;
  assign n21904 = n21903 ^ x11 ;
  assign n21906 = n21905 ^ n21904 ;
  assign n21908 = n21907 ^ n21906 ;
  assign n21910 = n21909 ^ n21908 ;
  assign n21912 = n21911 ^ n21910 ;
  assign n21913 = n21587 ^ n21448 ;
  assign n21914 = n21913 ^ n21903 ;
  assign n21915 = ~n21912 & n21914 ;
  assign n21916 = n21915 ^ n21913 ;
  assign n21918 = n21917 ^ n21916 ;
  assign n21929 = n6650 & n20994 ;
  assign n21922 = n20922 ^ x11 ;
  assign n21923 = n21922 ^ x10 ;
  assign n21924 = n21923 ^ n20922 ;
  assign n21925 = n21395 & n21924 ;
  assign n21926 = n21925 ^ n20922 ;
  assign n21927 = n6648 & ~n21926 ;
  assign n21928 = n21927 ^ x11 ;
  assign n21930 = n21929 ^ n21928 ;
  assign n21919 = n6655 & n20962 ;
  assign n21931 = n21930 ^ n21919 ;
  assign n21932 = n21931 ^ n21916 ;
  assign n21933 = n21918 & n21932 ;
  assign n21934 = n21933 ^ n21916 ;
  assign n21935 = n21934 ^ n21780 ;
  assign n21936 = ~n21782 & n21935 ;
  assign n21937 = n21936 ^ n21780 ;
  assign n21938 = n21937 ^ n21770 ;
  assign n21939 = ~n21772 & n21938 ;
  assign n21940 = n21939 ^ n21770 ;
  assign n21941 = n21940 ^ n21760 ;
  assign n21942 = ~n21762 & n21941 ;
  assign n21943 = n21942 ^ n21760 ;
  assign n21944 = n21943 ^ n21748 ;
  assign n21945 = ~n21750 & n21944 ;
  assign n21946 = n21945 ^ n21748 ;
  assign n22212 = n21946 ^ n21728 ;
  assign n22213 = n21738 & n22212 ;
  assign n22214 = n22213 ^ n21728 ;
  assign n22316 = n22293 ^ n22214 ;
  assign n22317 = n22301 & n22316 ;
  assign n22318 = n22317 ^ n22293 ;
  assign n22432 = n22402 ^ n22318 ;
  assign n22433 = n22411 & n22432 ;
  assign n22434 = n22433 ^ n22402 ;
  assign n22553 = n22528 ^ n22434 ;
  assign n22554 = n22536 & n22553 ;
  assign n22555 = n22554 ^ n22528 ;
  assign n23649 = n22658 ^ n22555 ;
  assign n23650 = n22664 & n23649 ;
  assign n23664 = n23663 ^ n23650 ;
  assign n23794 = n23793 ^ n23680 ;
  assign n23837 = n23794 ^ n23662 ;
  assign n23838 = ~n23664 & n23837 ;
  assign n23839 = n23838 ^ n23794 ;
  assign n24103 = n23971 ^ n23839 ;
  assign n24104 = n23986 & ~n24103 ;
  assign n24105 = n24104 ^ n23971 ;
  assign n24287 = n24286 ^ n24105 ;
  assign n24288 = n24287 ^ n24285 ;
  assign n24289 = ~n24249 & n24288 ;
  assign n24290 = n24289 ^ n24286 ;
  assign n24420 = n24419 ^ n24290 ;
  assign n22682 = n21049 ^ n21030 ;
  assign n22683 = n22682 ^ n20865 ;
  assign n24256 = n7135 & ~n22683 ;
  assign n24254 = n7146 & ~n20876 ;
  assign n24252 = n8054 & n20865 ;
  assign n24250 = n24249 ^ n24105 ;
  assign n24251 = n24250 ^ x8 ;
  assign n24253 = n24252 ^ n24251 ;
  assign n24255 = n24254 ^ n24253 ;
  assign n24257 = n24256 ^ n24255 ;
  assign n24102 = n7141 & ~n20872 ;
  assign n24258 = n24257 ^ n24102 ;
  assign n23987 = n23986 ^ n23839 ;
  assign n23795 = n23794 ^ n23664 ;
  assign n23988 = n23987 ^ n23795 ;
  assign n22673 = n7135 & ~n22672 ;
  assign n22669 = n7146 & ~n21025 ;
  assign n22667 = n8054 & n20882 ;
  assign n22665 = n22664 ^ n22555 ;
  assign n22666 = n22665 ^ x8 ;
  assign n22668 = n22667 ^ n22666 ;
  assign n22670 = n22669 ^ n22668 ;
  assign n22674 = n22673 ^ n22670 ;
  assign n22552 = n7141 & n20883 ;
  assign n22675 = n22674 ^ n22552 ;
  assign n23796 = n23795 ^ n22665 ;
  assign n23797 = n23796 ^ n23795 ;
  assign n22537 = n22536 ^ n22434 ;
  assign n21955 = n7135 & n21954 ;
  assign n21951 = n7146 & n20898 ;
  assign n21949 = n8054 & ~n20894 ;
  assign n21947 = n21946 ^ n21738 ;
  assign n21948 = n21947 ^ x8 ;
  assign n21950 = n21949 ^ n21948 ;
  assign n21952 = n21951 ^ n21950 ;
  assign n21956 = n21955 ^ n21952 ;
  assign n21079 = n7141 & n20897 ;
  assign n21957 = n21956 ^ n21079 ;
  assign n21967 = n7135 & ~n21966 ;
  assign n21963 = n7146 & ~n21012 ;
  assign n21961 = n8054 & n20897 ;
  assign n21959 = n21943 ^ n21750 ;
  assign n21960 = n21959 ^ x8 ;
  assign n21962 = n21961 ^ n21960 ;
  assign n21964 = n21963 ^ n21962 ;
  assign n21968 = n21967 ^ n21964 ;
  assign n21958 = n7141 & n20898 ;
  assign n21969 = n21968 ^ n21958 ;
  assign n21982 = n7141 & ~n21012 ;
  assign n21979 = n21940 ^ n21762 ;
  assign n21980 = n21979 ^ x8 ;
  assign n21974 = n20898 ^ n9577 ;
  assign n21975 = n21974 ^ n20898 ;
  assign n21976 = ~n21971 & n21975 ;
  assign n21977 = n21976 ^ n20898 ;
  assign n21978 = n7128 & n21977 ;
  assign n21981 = n21980 ^ n21978 ;
  assign n21983 = n21982 ^ n21981 ;
  assign n21970 = n7146 & n20902 ;
  assign n21984 = n21983 ^ n21970 ;
  assign n21992 = n7135 & n21735 ;
  assign n21988 = n21937 ^ n21772 ;
  assign n21989 = n21988 ^ x8 ;
  assign n21987 = n8054 & ~n21012 ;
  assign n21990 = n21989 ^ n21987 ;
  assign n21986 = n7146 & n20903 ;
  assign n21991 = n21990 ^ n21986 ;
  assign n21993 = n21992 ^ n21991 ;
  assign n21985 = n7141 & n20902 ;
  assign n21994 = n21993 ^ n21985 ;
  assign n22187 = n21934 ^ n21782 ;
  assign n22003 = n21931 ^ n21918 ;
  assign n22001 = n7141 & n20910 ;
  assign n21999 = n7135 & ~n21756 ;
  assign n21996 = n7146 & n20913 ;
  assign n21995 = n8054 & n20903 ;
  assign n21997 = n21996 ^ n21995 ;
  assign n21998 = n21997 ^ x8 ;
  assign n22000 = n21999 ^ n21998 ;
  assign n22002 = n22001 ^ n22000 ;
  assign n22004 = n22003 ^ n22002 ;
  assign n22013 = n21913 ^ n21912 ;
  assign n22011 = n7141 & n20913 ;
  assign n22009 = n7135 & n21667 ;
  assign n22006 = n7146 & ~n20922 ;
  assign n22005 = n8054 & n20910 ;
  assign n22007 = n22006 ^ n22005 ;
  assign n22008 = n22007 ^ x8 ;
  assign n22010 = n22009 ^ n22008 ;
  assign n22012 = n22011 ^ n22010 ;
  assign n22014 = n22013 ^ n22012 ;
  assign n22023 = n21901 ^ n21783 ;
  assign n22021 = n7141 & ~n20922 ;
  assign n22019 = n7135 & ~n21087 ;
  assign n22016 = n7146 & n20994 ;
  assign n22015 = n8054 & n20913 ;
  assign n22017 = n22016 ^ n22015 ;
  assign n22018 = n22017 ^ x8 ;
  assign n22020 = n22019 ^ n22018 ;
  assign n22022 = n22021 ^ n22020 ;
  assign n22024 = n22023 ^ n22022 ;
  assign n22153 = n21885 ^ n21803 ;
  assign n22140 = n21882 ^ n21813 ;
  assign n22033 = n7135 & n21114 ;
  assign n22029 = n21879 ^ n21824 ;
  assign n22030 = n22029 ^ x8 ;
  assign n22028 = n8054 & ~n20969 ;
  assign n22031 = n22030 ^ n22028 ;
  assign n22027 = n7146 & n20970 ;
  assign n22032 = n22031 ^ n22027 ;
  assign n22034 = n22033 ^ n22032 ;
  assign n22026 = n7141 & ~n20963 ;
  assign n22035 = n22034 ^ n22026 ;
  assign n22124 = n21876 ^ n21868 ;
  assign n22044 = n21864 ^ n21832 ;
  assign n22039 = n7146 & n20499 ;
  assign n22038 = n8054 & n20970 ;
  assign n22040 = n22039 ^ n22038 ;
  assign n22041 = n22040 ^ x8 ;
  assign n22037 = n7135 & ~n21251 ;
  assign n22042 = n22041 ^ n22037 ;
  assign n22036 = n7141 & ~n20924 ;
  assign n22043 = n22042 ^ n22036 ;
  assign n22045 = n22044 ^ n22043 ;
  assign n22107 = n21858 ^ n21833 ;
  assign n22108 = n22107 ^ n21849 ;
  assign n22093 = x11 & n21834 ;
  assign n22086 = n21848 ^ n20926 ;
  assign n22087 = n22086 ^ n20926 ;
  assign n22088 = n21155 ^ n20926 ;
  assign n22089 = n22087 & n22088 ;
  assign n22090 = n22089 ^ n20926 ;
  assign n22091 = n6650 & n22090 ;
  assign n22092 = n22091 ^ n21847 ;
  assign n22094 = n22093 ^ n22092 ;
  assign n22072 = n6647 & ~n20927 ;
  assign n22071 = n6648 & n20926 ;
  assign n22073 = n22072 ^ n22071 ;
  assign n22046 = n6648 & ~n20927 ;
  assign n22047 = n7128 & n20926 ;
  assign n22048 = n7144 & n20927 ;
  assign n22049 = ~n22047 & n22048 ;
  assign n22050 = n22049 ^ n7144 ;
  assign n22051 = n22050 ^ x8 ;
  assign n22056 = n7141 & n20926 ;
  assign n22055 = n8054 & n20939 ;
  assign n22057 = n22056 ^ n22055 ;
  assign n22053 = n7146 & ~n20927 ;
  assign n22052 = n7135 & n21144 ;
  assign n22054 = n22053 ^ n22052 ;
  assign n22058 = n22057 ^ n22054 ;
  assign n22059 = n22051 & ~n22058 ;
  assign n22060 = ~n22046 & ~n22059 ;
  assign n22064 = n7146 & n20926 ;
  assign n22063 = n8054 & n20941 ;
  assign n22065 = n22064 ^ n22063 ;
  assign n22066 = n22065 ^ x8 ;
  assign n22062 = n7135 & n21172 ;
  assign n22067 = n22066 ^ n22062 ;
  assign n22061 = n7141 & n20939 ;
  assign n22068 = n22067 ^ n22061 ;
  assign n22069 = n22060 & n22068 ;
  assign n22070 = n22069 ^ n22068 ;
  assign n22074 = n22073 ^ n22070 ;
  assign n22078 = n7146 & n20939 ;
  assign n22077 = n8054 & ~n20925 ;
  assign n22079 = n22078 ^ n22077 ;
  assign n22080 = n22079 ^ x8 ;
  assign n22076 = n7135 & ~n21188 ;
  assign n22081 = n22080 ^ n22076 ;
  assign n22075 = n7141 & n20941 ;
  assign n22082 = n22081 ^ n22075 ;
  assign n22083 = n22082 ^ n22070 ;
  assign n22084 = n22074 & n22083 ;
  assign n22085 = n22084 ^ n22070 ;
  assign n22095 = n22094 ^ n22085 ;
  assign n22099 = n7146 & n20941 ;
  assign n22098 = n8054 & n20499 ;
  assign n22100 = n22099 ^ n22098 ;
  assign n22101 = n22100 ^ x8 ;
  assign n22097 = n7135 & ~n21124 ;
  assign n22102 = n22101 ^ n22097 ;
  assign n22096 = n7141 & ~n20925 ;
  assign n22103 = n22102 ^ n22096 ;
  assign n22104 = n22103 ^ n22085 ;
  assign n22105 = n22095 & ~n22104 ;
  assign n22106 = n22105 ^ n22094 ;
  assign n22109 = n22108 ^ n22106 ;
  assign n22117 = n7141 & n20499 ;
  assign n22114 = n8054 & ~n20924 ;
  assign n22112 = n7146 & ~n20925 ;
  assign n22111 = n22106 ^ x8 ;
  assign n22113 = n22112 ^ n22111 ;
  assign n22115 = n22114 ^ n22113 ;
  assign n22110 = n7135 & n21211 ;
  assign n22116 = n22115 ^ n22110 ;
  assign n22118 = n22117 ^ n22116 ;
  assign n22119 = n22109 & ~n22118 ;
  assign n22120 = n22119 ^ n22108 ;
  assign n22121 = n22120 ^ n22043 ;
  assign n22122 = n22045 & ~n22121 ;
  assign n22123 = n22122 ^ n22044 ;
  assign n22125 = n22124 ^ n22123 ;
  assign n22132 = n7135 & n21240 ;
  assign n22130 = n7146 & ~n20924 ;
  assign n22128 = n8054 & ~n20963 ;
  assign n22127 = n22124 ^ x8 ;
  assign n22129 = n22128 ^ n22127 ;
  assign n22131 = n22130 ^ n22129 ;
  assign n22133 = n22132 ^ n22131 ;
  assign n22126 = n7141 & n20970 ;
  assign n22134 = n22133 ^ n22126 ;
  assign n22135 = ~n22125 & ~n22134 ;
  assign n22136 = n22135 ^ n22124 ;
  assign n22137 = n22136 ^ n22029 ;
  assign n22138 = ~n22035 & n22137 ;
  assign n22139 = n22138 ^ n22029 ;
  assign n22141 = n22140 ^ n22139 ;
  assign n22145 = n7146 & ~n20963 ;
  assign n22144 = n8054 & n20962 ;
  assign n22146 = n22145 ^ n22144 ;
  assign n22147 = n22146 ^ x8 ;
  assign n22143 = n7135 & n21109 ;
  assign n22148 = n22147 ^ n22143 ;
  assign n22142 = n7141 & ~n20969 ;
  assign n22149 = n22148 ^ n22142 ;
  assign n22150 = n22149 ^ n22139 ;
  assign n22151 = ~n22141 & n22150 ;
  assign n22152 = n22151 ^ n22140 ;
  assign n22154 = n22153 ^ n22152 ;
  assign n22161 = n7141 & n20962 ;
  assign n22159 = n7135 & n21630 ;
  assign n22156 = n7146 & ~n20969 ;
  assign n22155 = n8054 & n20994 ;
  assign n22157 = n22156 ^ n22155 ;
  assign n22158 = n22157 ^ x8 ;
  assign n22160 = n22159 ^ n22158 ;
  assign n22162 = n22161 ^ n22160 ;
  assign n22163 = n22162 ^ n22152 ;
  assign n22164 = ~n22154 & n22163 ;
  assign n22165 = n22164 ^ n22162 ;
  assign n22025 = n21888 ^ n21793 ;
  assign n22166 = n22165 ^ n22025 ;
  assign n22174 = n7141 & n20994 ;
  assign n22170 = n22165 ^ x8 ;
  assign n22169 = n7146 & n20962 ;
  assign n22171 = n22170 ^ n22169 ;
  assign n22168 = n8054 & ~n20922 ;
  assign n22172 = n22171 ^ n22168 ;
  assign n21920 = n21395 ^ n20922 ;
  assign n22167 = n7135 & ~n21920 ;
  assign n22173 = n22172 ^ n22167 ;
  assign n22175 = n22174 ^ n22173 ;
  assign n22176 = n22166 & n22175 ;
  assign n22177 = n22176 ^ n22165 ;
  assign n22178 = n22177 ^ n22022 ;
  assign n22179 = ~n22024 & n22178 ;
  assign n22180 = n22179 ^ n22022 ;
  assign n22181 = n22180 ^ n22012 ;
  assign n22182 = n22014 & n22181 ;
  assign n22183 = n22182 ^ n22012 ;
  assign n22184 = n22183 ^ n22002 ;
  assign n22185 = n22004 & n22184 ;
  assign n22186 = n22185 ^ n22002 ;
  assign n22188 = n22187 ^ n22186 ;
  assign n22195 = n7135 & ~n21744 ;
  assign n22193 = n7146 & n20910 ;
  assign n22191 = n8054 & n20902 ;
  assign n22190 = n22187 ^ x8 ;
  assign n22192 = n22191 ^ n22190 ;
  assign n22194 = n22193 ^ n22192 ;
  assign n22196 = n22195 ^ n22194 ;
  assign n22189 = n7141 & n20903 ;
  assign n22197 = n22196 ^ n22189 ;
  assign n22198 = ~n22188 & ~n22197 ;
  assign n22199 = n22198 ^ n22187 ;
  assign n22200 = n22199 ^ n21988 ;
  assign n22201 = ~n21994 & n22200 ;
  assign n22202 = n22201 ^ n21988 ;
  assign n22203 = n22202 ^ n21979 ;
  assign n22204 = ~n21984 & n22203 ;
  assign n22205 = n22204 ^ n21979 ;
  assign n22206 = n22205 ^ n21959 ;
  assign n22207 = ~n21969 & n22206 ;
  assign n22208 = n22207 ^ n21959 ;
  assign n22209 = n22208 ^ n21947 ;
  assign n22210 = n21957 & ~n22209 ;
  assign n22211 = n22210 ^ n21947 ;
  assign n22302 = n22301 ^ n22214 ;
  assign n22304 = n22211 & n22302 ;
  assign n22303 = n22302 ^ n22211 ;
  assign n22305 = n22304 ^ n22303 ;
  assign n22312 = n7146 & n20897 ;
  assign n22311 = n8054 & ~n20887 ;
  assign n22313 = n22312 ^ n22311 ;
  assign n22309 = n7141 & ~n20894 ;
  assign n22308 = n7135 & n22307 ;
  assign n22310 = n22309 ^ n22308 ;
  assign n22314 = n22313 ^ n22310 ;
  assign n22315 = n22314 ^ x8 ;
  assign n22420 = n7146 & ~n20894 ;
  assign n22419 = n8054 & ~n21025 ;
  assign n22421 = n22420 ^ n22419 ;
  assign n22417 = n7141 & ~n20887 ;
  assign n22416 = n7135 & n22415 ;
  assign n22418 = n22417 ^ n22416 ;
  assign n22422 = n22421 ^ n22418 ;
  assign n22412 = n22411 ^ n22318 ;
  assign n22413 = n22412 ^ n22314 ;
  assign n22423 = n22422 ^ n22413 ;
  assign n22424 = n22315 & ~n22423 ;
  assign n22425 = n22305 & n22424 ;
  assign n22426 = n22412 ^ n22304 ;
  assign n22427 = n22412 ^ x8 ;
  assign n22428 = n22427 ^ n22422 ;
  assign n22429 = n22426 & ~n22428 ;
  assign n22430 = n22429 ^ n22304 ;
  assign n22431 = ~n22425 & ~n22430 ;
  assign n22538 = n22537 ^ n22431 ;
  assign n22547 = n7135 & ~n22546 ;
  assign n22543 = n7146 & ~n20887 ;
  assign n22541 = n8054 & n20883 ;
  assign n22540 = n22537 ^ x8 ;
  assign n22542 = n22541 ^ n22540 ;
  assign n22544 = n22543 ^ n22542 ;
  assign n22548 = n22547 ^ n22544 ;
  assign n22539 = n7141 & ~n21025 ;
  assign n22549 = n22548 ^ n22539 ;
  assign n22550 = ~n22538 & n22549 ;
  assign n22551 = n22550 ^ n22537 ;
  assign n23798 = n23797 ^ n22551 ;
  assign n23799 = n22675 & n23798 ;
  assign n23800 = n23799 ^ n23796 ;
  assign n23807 = n7141 & n20882 ;
  assign n23805 = n7135 & n23010 ;
  assign n23802 = n7146 & n20883 ;
  assign n23801 = n8054 & ~n20876 ;
  assign n23803 = n23802 ^ n23801 ;
  assign n23804 = n23803 ^ x8 ;
  assign n23806 = n23805 ^ n23804 ;
  assign n23808 = n23807 ^ n23806 ;
  assign n23835 = n23808 ^ n23795 ;
  assign n23836 = n23800 & n23835 ;
  assign n23989 = n23988 ^ n23836 ;
  assign n23993 = n7146 & n20882 ;
  assign n23992 = n8054 & ~n20872 ;
  assign n23994 = n23993 ^ n23992 ;
  assign n23995 = n23994 ^ x8 ;
  assign n23032 = n21048 ^ n21029 ;
  assign n23033 = n23032 ^ n20872 ;
  assign n23991 = n7135 & n23033 ;
  assign n23996 = n23995 ^ n23991 ;
  assign n23990 = n7141 & ~n20876 ;
  assign n23997 = n23996 ^ n23990 ;
  assign n24272 = n23997 ^ n23987 ;
  assign n24273 = ~n23989 & n24272 ;
  assign n24274 = n24273 ^ n23997 ;
  assign n23608 = n21050 ^ n21031 ;
  assign n24259 = ~x7 & ~n23608 ;
  assign n23640 = n23608 ^ n20861 ;
  assign n24267 = n24259 ^ n23640 ;
  assign n24268 = n7130 & ~n24267 ;
  assign n24263 = n7146 & ~n20872 ;
  assign n24262 = n7141 & n20865 ;
  assign n24264 = n24263 ^ n24262 ;
  assign n24265 = n24264 ^ x8 ;
  assign n24260 = n24259 ^ n20861 ;
  assign n24261 = n7129 & n24260 ;
  assign n24266 = n24265 ^ n24261 ;
  assign n24269 = n24268 ^ n24266 ;
  assign n24270 = n24269 ^ n24250 ;
  assign n24271 = n24270 ^ n24269 ;
  assign n24275 = n24274 ^ n24271 ;
  assign n24276 = n24258 & n24275 ;
  assign n24277 = n24276 ^ n24270 ;
  assign n24421 = n24420 ^ n24277 ;
  assign n24944 = n24943 ^ n24421 ;
  assign n21061 = n21053 ^ n21034 ;
  assign n24427 = n21061 ^ n20837 ;
  assign n24428 = n9081 & ~n24427 ;
  assign n24425 = n9085 & n20836 ;
  assign n24423 = n10131 & n20837 ;
  assign n24422 = n24421 ^ x5 ;
  assign n24424 = n24423 ^ n24422 ;
  assign n24426 = n24425 ^ n24424 ;
  assign n24429 = n24428 ^ n24426 ;
  assign n24101 = ~n9092 & n20852 ;
  assign n24430 = n24429 ^ n24101 ;
  assign n24436 = n9085 & n20852 ;
  assign n24435 = n10131 & n20836 ;
  assign n24437 = n24436 ^ n24435 ;
  assign n24438 = n24437 ^ x5 ;
  assign n23041 = n21052 ^ n21033 ;
  assign n24433 = n23041 ^ n20836 ;
  assign n24434 = n9081 & ~n24433 ;
  assign n24439 = n24438 ^ n24434 ;
  assign n24432 = ~n9092 & n20861 ;
  assign n24440 = n24439 ^ n24432 ;
  assign n24925 = n24440 ^ n24421 ;
  assign n24443 = n24274 ^ n24258 ;
  assign n24926 = n24925 ^ n24443 ;
  assign n23812 = n9085 & n20865 ;
  assign n23809 = n23808 ^ n23800 ;
  assign n23810 = n23809 ^ x5 ;
  assign n23644 = n20861 ^ n9089 ;
  assign n23645 = n23644 ^ n20861 ;
  assign n23646 = ~n23608 & n23645 ;
  assign n23647 = n23646 ^ n20861 ;
  assign n23648 = n9077 & n23647 ;
  assign n23811 = n23810 ^ n23648 ;
  assign n23813 = n23812 ^ n23811 ;
  assign n23639 = ~n9092 & ~n20872 ;
  assign n23814 = n23813 ^ n23639 ;
  assign n22684 = n9081 & ~n22683 ;
  assign n22680 = n9085 & ~n20872 ;
  assign n22678 = n10131 & n20865 ;
  assign n22676 = n22675 ^ n22551 ;
  assign n22677 = n22676 ^ x5 ;
  assign n22679 = n22678 ^ n22677 ;
  assign n22681 = n22680 ^ n22679 ;
  assign n22685 = n22684 ^ n22681 ;
  assign n21078 = ~n9092 & ~n20876 ;
  assign n22686 = n22685 ^ n21078 ;
  assign n23024 = n22549 ^ n22431 ;
  assign n23013 = ~n9092 & n20883 ;
  assign n23011 = n9081 & n23010 ;
  assign n23006 = n10131 & ~n20876 ;
  assign n23005 = n9085 & n20882 ;
  assign n23007 = n23006 ^ n23005 ;
  assign n23008 = n23007 ^ x5 ;
  assign n23012 = n23011 ^ n23008 ;
  assign n23014 = n23013 ^ n23012 ;
  assign n22695 = n22315 ^ n22303 ;
  assign n22690 = n9085 & n20883 ;
  assign n22689 = n10131 & n20882 ;
  assign n22691 = n22690 ^ n22689 ;
  assign n22692 = n22691 ^ x5 ;
  assign n22688 = n9081 & ~n22672 ;
  assign n22693 = n22692 ^ n22688 ;
  assign n22687 = ~n9092 & ~n21025 ;
  assign n22694 = n22693 ^ n22687 ;
  assign n22696 = n22695 ^ n22694 ;
  assign n22704 = n9081 & ~n22546 ;
  assign n22702 = n9085 & ~n21025 ;
  assign n22700 = n10131 & n20883 ;
  assign n22698 = n22208 ^ n21957 ;
  assign n22699 = n22698 ^ x5 ;
  assign n22701 = n22700 ^ n22699 ;
  assign n22703 = n22702 ^ n22701 ;
  assign n22705 = n22704 ^ n22703 ;
  assign n22697 = ~n9092 & ~n20887 ;
  assign n22706 = n22705 ^ n22697 ;
  assign n22714 = n9081 & n22415 ;
  assign n22710 = n22205 ^ n21969 ;
  assign n22711 = n22710 ^ x5 ;
  assign n22709 = n10131 & ~n21025 ;
  assign n22712 = n22711 ^ n22709 ;
  assign n22708 = n9085 & ~n20887 ;
  assign n22713 = n22712 ^ n22708 ;
  assign n22715 = n22714 ^ n22713 ;
  assign n22707 = ~n9092 & ~n20894 ;
  assign n22716 = n22715 ^ n22707 ;
  assign n22724 = n9081 & n22307 ;
  assign n22720 = n22202 ^ n21984 ;
  assign n22721 = n22720 ^ x5 ;
  assign n22719 = n10131 & ~n20887 ;
  assign n22722 = n22721 ^ n22719 ;
  assign n22718 = n9085 & ~n20894 ;
  assign n22723 = n22722 ^ n22718 ;
  assign n22725 = n22724 ^ n22723 ;
  assign n22717 = ~n9092 & n20897 ;
  assign n22726 = n22725 ^ n22717 ;
  assign n22734 = n9081 & n21954 ;
  assign n22730 = n22199 ^ n21994 ;
  assign n22731 = n22730 ^ x5 ;
  assign n22729 = n10131 & ~n20894 ;
  assign n22732 = n22731 ^ n22729 ;
  assign n22728 = n9085 & n20897 ;
  assign n22733 = n22732 ^ n22728 ;
  assign n22735 = n22734 ^ n22733 ;
  assign n22727 = ~n9092 & n20898 ;
  assign n22736 = n22735 ^ n22727 ;
  assign n22977 = n22197 ^ n22186 ;
  assign n22745 = n22183 ^ n22004 ;
  assign n22743 = ~n9092 & n20902 ;
  assign n22741 = n9081 & ~n21972 ;
  assign n22738 = n9085 & ~n21012 ;
  assign n22737 = n10131 & n20898 ;
  assign n22739 = n22738 ^ n22737 ;
  assign n22740 = n22739 ^ x5 ;
  assign n22742 = n22741 ^ n22740 ;
  assign n22744 = n22743 ^ n22742 ;
  assign n22746 = n22745 ^ n22744 ;
  assign n22755 = n22180 ^ n22014 ;
  assign n22753 = ~n9092 & n20903 ;
  assign n22751 = n9081 & n21735 ;
  assign n22748 = n9085 & n20902 ;
  assign n22747 = n10131 & ~n21012 ;
  assign n22749 = n22748 ^ n22747 ;
  assign n22750 = n22749 ^ x5 ;
  assign n22752 = n22751 ^ n22750 ;
  assign n22754 = n22753 ^ n22752 ;
  assign n22756 = n22755 ^ n22754 ;
  assign n22765 = n22177 ^ n22024 ;
  assign n22763 = ~n9092 & n20910 ;
  assign n22761 = n9081 & ~n21744 ;
  assign n22758 = n9085 & n20903 ;
  assign n22757 = n10131 & n20902 ;
  assign n22759 = n22758 ^ n22757 ;
  assign n22760 = n22759 ^ x5 ;
  assign n22762 = n22761 ^ n22760 ;
  assign n22764 = n22763 ^ n22762 ;
  assign n22766 = n22765 ^ n22764 ;
  assign n22775 = n22175 ^ n22025 ;
  assign n22776 = n22775 ^ x5 ;
  assign n22774 = ~n9092 & n20913 ;
  assign n22777 = n22776 ^ n22774 ;
  assign n22773 = n9085 & n20910 ;
  assign n22778 = n22777 ^ n22773 ;
  assign n22768 = n20903 ^ n9089 ;
  assign n22769 = n22768 ^ n20903 ;
  assign n22770 = ~n21755 & n22769 ;
  assign n22771 = n22770 ^ n20903 ;
  assign n22772 = n9077 & n22771 ;
  assign n22779 = n22778 ^ n22772 ;
  assign n22949 = n22162 ^ n22154 ;
  assign n22788 = n22149 ^ n22141 ;
  assign n22786 = ~n9092 & n20994 ;
  assign n22784 = n9081 & ~n21087 ;
  assign n22781 = n10131 & n20913 ;
  assign n22780 = n9085 & ~n20922 ;
  assign n22782 = n22781 ^ n22780 ;
  assign n22783 = n22782 ^ x5 ;
  assign n22785 = n22784 ^ n22783 ;
  assign n22787 = n22786 ^ n22785 ;
  assign n22789 = n22788 ^ n22787 ;
  assign n22797 = ~n9092 & n20962 ;
  assign n22795 = n9081 & ~n21920 ;
  assign n22792 = n9085 & n20994 ;
  assign n22791 = n10131 & ~n20922 ;
  assign n22793 = n22792 ^ n22791 ;
  assign n22794 = n22793 ^ x5 ;
  assign n22796 = n22795 ^ n22794 ;
  assign n22798 = n22797 ^ n22796 ;
  assign n22790 = n22136 ^ n22035 ;
  assign n22799 = n22798 ^ n22790 ;
  assign n22930 = n22134 ^ n22123 ;
  assign n22807 = n9081 & n21109 ;
  assign n22803 = n22120 ^ n22045 ;
  assign n22804 = n22803 ^ x5 ;
  assign n22802 = n10131 & n20962 ;
  assign n22805 = n22804 ^ n22802 ;
  assign n22801 = n9085 & ~n20969 ;
  assign n22806 = n22805 ^ n22801 ;
  assign n22808 = n22807 ^ n22806 ;
  assign n22800 = ~n9092 & ~n20963 ;
  assign n22809 = n22808 ^ n22800 ;
  assign n22817 = n9081 & n21114 ;
  assign n22813 = n22118 ^ n22108 ;
  assign n22814 = n22813 ^ x5 ;
  assign n22812 = n10131 & ~n20969 ;
  assign n22815 = n22814 ^ n22812 ;
  assign n22811 = n9085 & ~n20963 ;
  assign n22816 = n22815 ^ n22811 ;
  assign n22818 = n22817 ^ n22816 ;
  assign n22810 = ~n9092 & n20970 ;
  assign n22819 = n22818 ^ n22810 ;
  assign n22828 = n22103 ^ n22095 ;
  assign n22823 = n9085 & n20970 ;
  assign n22822 = n10131 & ~n20963 ;
  assign n22824 = n22823 ^ n22822 ;
  assign n22825 = n22824 ^ x5 ;
  assign n22821 = n9081 & n21240 ;
  assign n22826 = n22825 ^ n22821 ;
  assign n22820 = ~n9092 & ~n20924 ;
  assign n22827 = n22826 ^ n22820 ;
  assign n22829 = n22828 ^ n22827 ;
  assign n22838 = n22082 ^ n22074 ;
  assign n22833 = n9085 & ~n20924 ;
  assign n22832 = n10131 & n20970 ;
  assign n22834 = n22833 ^ n22832 ;
  assign n22835 = n22834 ^ x5 ;
  assign n22831 = n9081 & ~n21251 ;
  assign n22836 = n22835 ^ n22831 ;
  assign n22830 = ~n9092 & n20499 ;
  assign n22837 = n22836 ^ n22830 ;
  assign n22839 = n22838 ^ n22837 ;
  assign n22848 = n22059 ^ n22046 ;
  assign n22849 = n22848 ^ n22068 ;
  assign n22843 = n9085 & n20499 ;
  assign n22842 = n10131 & ~n20924 ;
  assign n22844 = n22843 ^ n22842 ;
  assign n22845 = n22844 ^ x5 ;
  assign n22841 = n9081 & n21211 ;
  assign n22846 = n22845 ^ n22841 ;
  assign n22840 = ~n9092 & ~n20925 ;
  assign n22847 = n22846 ^ n22840 ;
  assign n22850 = n22849 ^ n22847 ;
  assign n22855 = n9085 & n20941 ;
  assign n22854 = n10131 & ~n20925 ;
  assign n22856 = n22855 ^ n22854 ;
  assign n22852 = ~n9092 & n20939 ;
  assign n22851 = n9081 & ~n21188 ;
  assign n22853 = n22852 ^ n22851 ;
  assign n22857 = n22856 ^ n22853 ;
  assign n22858 = n22857 ^ x5 ;
  assign n22865 = n9085 & ~n20925 ;
  assign n22864 = n10131 & n20499 ;
  assign n22866 = n22865 ^ n22864 ;
  assign n22862 = ~n9092 & n20941 ;
  assign n22861 = n9081 & ~n21124 ;
  assign n22863 = n22862 ^ n22861 ;
  assign n22867 = n22866 ^ n22863 ;
  assign n22859 = n22058 ^ n22050 ;
  assign n22860 = n22859 ^ n22857 ;
  assign n22868 = n22867 ^ n22860 ;
  assign n22869 = n22858 & ~n22868 ;
  assign n22870 = n7128 & ~n20927 ;
  assign n22871 = n9077 & n20926 ;
  assign n22872 = x5 & ~n22871 ;
  assign n22873 = ~n20927 & n22872 ;
  assign n22874 = ~n18627 & n22873 ;
  assign n22875 = n22874 ^ n22872 ;
  assign n22884 = n9089 & n22871 ;
  assign n22885 = n22884 ^ n9092 ;
  assign n22886 = n20927 & ~n22885 ;
  assign n22887 = n22886 ^ n9092 ;
  assign n22879 = n9077 & n20939 ;
  assign n22888 = n22887 ^ n22879 ;
  assign n22878 = n9085 & n20926 ;
  assign n22889 = n22888 ^ n22878 ;
  assign n22890 = n22875 & n22889 ;
  assign n22891 = ~n22870 & ~n22890 ;
  assign n22898 = n10131 & n20941 ;
  assign n22896 = n9085 & n20939 ;
  assign n22893 = ~n9092 & n20926 ;
  assign n22892 = n9081 & n21172 ;
  assign n22894 = n22893 ^ n22892 ;
  assign n22895 = n22894 ^ x5 ;
  assign n22897 = n22896 ^ n22895 ;
  assign n22899 = n22898 ^ n22897 ;
  assign n22900 = n22891 & n22899 ;
  assign n22901 = n22900 ^ n22899 ;
  assign n22902 = n7140 & ~n20927 ;
  assign n22903 = n22902 ^ n22047 ;
  assign n22905 = n22901 & n22903 ;
  assign n22904 = n22903 ^ n22901 ;
  assign n22906 = n22905 ^ n22904 ;
  assign n22907 = n22905 ^ n22859 ;
  assign n22908 = n22867 ^ x5 ;
  assign n22909 = n22908 ^ n22905 ;
  assign n22910 = n22907 & ~n22909 ;
  assign n22911 = n22910 ^ n22859 ;
  assign n22912 = n22906 & ~n22911 ;
  assign n22913 = n22869 & n22912 ;
  assign n22914 = n22913 ^ n22911 ;
  assign n22915 = n22914 ^ n22847 ;
  assign n22916 = n22850 & n22915 ;
  assign n22917 = n22916 ^ n22847 ;
  assign n22918 = n22917 ^ n22837 ;
  assign n22919 = n22839 & n22918 ;
  assign n22920 = n22919 ^ n22837 ;
  assign n22921 = n22920 ^ n22827 ;
  assign n22922 = n22829 & n22921 ;
  assign n22923 = n22922 ^ n22827 ;
  assign n22924 = n22923 ^ n22813 ;
  assign n22925 = n22819 & n22924 ;
  assign n22926 = n22925 ^ n22813 ;
  assign n22927 = n22926 ^ n22803 ;
  assign n22928 = n22809 & n22927 ;
  assign n22929 = n22928 ^ n22803 ;
  assign n22931 = n22930 ^ n22929 ;
  assign n22938 = ~n9092 & ~n20969 ;
  assign n22936 = n9081 & n21630 ;
  assign n22933 = n9085 & n20962 ;
  assign n22932 = n10131 & n20994 ;
  assign n22934 = n22933 ^ n22932 ;
  assign n22935 = n22934 ^ x5 ;
  assign n22937 = n22936 ^ n22935 ;
  assign n22939 = n22938 ^ n22937 ;
  assign n22940 = n22939 ^ n22929 ;
  assign n22941 = ~n22931 & ~n22940 ;
  assign n22942 = n22941 ^ n22930 ;
  assign n22943 = n22942 ^ n22790 ;
  assign n22944 = n22799 & n22943 ;
  assign n22945 = n22944 ^ n22798 ;
  assign n22946 = n22945 ^ n22787 ;
  assign n22947 = ~n22789 & n22946 ;
  assign n22948 = n22947 ^ n22787 ;
  assign n22950 = n22949 ^ n22948 ;
  assign n22960 = n9085 & n20913 ;
  assign n22958 = ~n9092 & ~n20922 ;
  assign n22957 = n22949 ^ x5 ;
  assign n22959 = n22958 ^ n22957 ;
  assign n22961 = n22960 ^ n22959 ;
  assign n22952 = n20910 ^ n9089 ;
  assign n22953 = n22952 ^ n20910 ;
  assign n22954 = n22951 & n22953 ;
  assign n22955 = n22954 ^ n20910 ;
  assign n22956 = n9077 & n22955 ;
  assign n22962 = n22961 ^ n22956 ;
  assign n22963 = n22950 & n22962 ;
  assign n22964 = n22963 ^ n22949 ;
  assign n22965 = n22964 ^ n22775 ;
  assign n22966 = n22779 & n22965 ;
  assign n22967 = n22966 ^ n22775 ;
  assign n22968 = n22967 ^ n22764 ;
  assign n22969 = ~n22766 & n22968 ;
  assign n22970 = n22969 ^ n22764 ;
  assign n22971 = n22970 ^ n22754 ;
  assign n22972 = n22756 & n22971 ;
  assign n22973 = n22972 ^ n22754 ;
  assign n22974 = n22973 ^ n22744 ;
  assign n22975 = n22746 & n22974 ;
  assign n22976 = n22975 ^ n22744 ;
  assign n22978 = n22977 ^ n22976 ;
  assign n22985 = n9081 & ~n21966 ;
  assign n22983 = n9085 & n20898 ;
  assign n22981 = n10131 & n20897 ;
  assign n22980 = n22977 ^ x5 ;
  assign n22982 = n22981 ^ n22980 ;
  assign n22984 = n22983 ^ n22982 ;
  assign n22986 = n22985 ^ n22984 ;
  assign n22979 = ~n9092 & ~n21012 ;
  assign n22987 = n22986 ^ n22979 ;
  assign n22988 = ~n22978 & ~n22987 ;
  assign n22989 = n22988 ^ n22977 ;
  assign n22990 = n22989 ^ n22730 ;
  assign n22991 = n22736 & ~n22990 ;
  assign n22992 = n22991 ^ n22730 ;
  assign n22993 = n22992 ^ n22720 ;
  assign n22994 = n22726 & n22993 ;
  assign n22995 = n22994 ^ n22720 ;
  assign n22996 = n22995 ^ n22710 ;
  assign n22997 = n22716 & n22996 ;
  assign n22998 = n22997 ^ n22710 ;
  assign n22999 = n22998 ^ n22698 ;
  assign n23000 = ~n22706 & ~n22999 ;
  assign n23001 = n23000 ^ n22698 ;
  assign n23002 = n23001 ^ n22694 ;
  assign n23003 = n22696 & ~n23002 ;
  assign n23004 = n23003 ^ n22694 ;
  assign n23015 = n23014 ^ n23004 ;
  assign n23019 = n22315 ^ n22211 ;
  assign n23020 = ~n22303 & n23019 ;
  assign n23016 = n22422 ^ n22412 ;
  assign n23017 = n23016 ^ n22314 ;
  assign n23018 = n23017 ^ n23014 ;
  assign n23021 = n23020 ^ n23018 ;
  assign n23022 = n23015 & n23021 ;
  assign n23023 = n23022 ^ n23014 ;
  assign n23025 = n23024 ^ n23023 ;
  assign n23034 = n9081 & n23033 ;
  assign n23030 = n9085 & ~n20876 ;
  assign n23028 = n10131 & ~n20872 ;
  assign n23027 = n23024 ^ x5 ;
  assign n23029 = n23028 ^ n23027 ;
  assign n23031 = n23030 ^ n23029 ;
  assign n23035 = n23034 ^ n23031 ;
  assign n23026 = ~n9092 & n20882 ;
  assign n23036 = n23035 ^ n23026 ;
  assign n23037 = ~n23025 & ~n23036 ;
  assign n23038 = n23037 ^ n23024 ;
  assign n23636 = n23038 ^ n22676 ;
  assign n23637 = n22686 & ~n23636 ;
  assign n23638 = n23637 ^ n22676 ;
  assign n23831 = n23809 ^ n23638 ;
  assign n23832 = n23814 & n23831 ;
  assign n23828 = ~n9092 & n20865 ;
  assign n23059 = n21051 ^ n21032 ;
  assign n23825 = n23059 ^ n20852 ;
  assign n23826 = n9081 & ~n23825 ;
  assign n23822 = n10131 & n20852 ;
  assign n23821 = n9085 & n20861 ;
  assign n23823 = n23822 ^ n23821 ;
  assign n23824 = n23823 ^ x5 ;
  assign n23827 = n23826 ^ n23824 ;
  assign n23829 = n23828 ^ n23827 ;
  assign n23830 = n23829 ^ n23809 ;
  assign n23833 = n23832 ^ n23830 ;
  assign n23998 = n23997 ^ n23989 ;
  assign n24098 = n23998 ^ n23829 ;
  assign n24099 = ~n23833 & n24098 ;
  assign n24100 = n24099 ^ n23998 ;
  assign n24927 = n24926 ^ n24100 ;
  assign n24928 = n24927 ^ n24925 ;
  assign n24929 = n24925 ^ n24440 ;
  assign n24930 = n24929 ^ n24443 ;
  assign n24931 = n24930 ^ n24925 ;
  assign n24932 = ~n24928 & n24931 ;
  assign n24933 = n24932 ^ n24925 ;
  assign n24934 = n24430 & n24933 ;
  assign n24945 = n24944 ^ n24934 ;
  assign n24922 = n7141 & n20861 ;
  assign n24920 = n7135 & ~n23825 ;
  assign n24917 = n7146 & n20865 ;
  assign n24916 = n8054 & n20852 ;
  assign n24918 = n24917 ^ n24916 ;
  assign n24919 = n24918 ^ x8 ;
  assign n24921 = n24920 ^ n24919 ;
  assign n24923 = n24922 ^ n24921 ;
  assign n24904 = n5703 & n21954 ;
  assign n24902 = n5700 & n20897 ;
  assign n24900 = n5702 & ~n20894 ;
  assign n24895 = n4916 & n20902 ;
  assign n24888 = n4504 & ~n20922 ;
  assign n24887 = n4491 & n20910 ;
  assign n24889 = n24888 ^ n24887 ;
  assign n24885 = ~n4496 & n20913 ;
  assign n24884 = n4492 & n21667 ;
  assign n24886 = n24885 ^ n24884 ;
  assign n24890 = n24889 ^ n24886 ;
  assign n24891 = n24890 ^ x23 ;
  assign n24851 = n446 & n20962 ;
  assign n24849 = n12861 & ~n20969 ;
  assign n24847 = ~n487 & n20994 ;
  assign n24835 = n5218 ^ n1906 ;
  assign n24834 = n13874 ^ n733 ;
  assign n24836 = n24835 ^ n24834 ;
  assign n24837 = n24836 ^ n13152 ;
  assign n24838 = n24837 ^ n4771 ;
  assign n24830 = n743 ^ n612 ;
  assign n24831 = n24830 ^ n4790 ;
  assign n24828 = n2460 ^ n774 ;
  assign n24829 = n24828 ^ n935 ;
  assign n24832 = n24831 ^ n24829 ;
  assign n24833 = n24832 ^ n3702 ;
  assign n24839 = n24838 ^ n24833 ;
  assign n24840 = n24839 ^ n4355 ;
  assign n24841 = ~n13227 & ~n24840 ;
  assign n24825 = ~n3733 & ~n20925 ;
  assign n24824 = n3726 & n20499 ;
  assign n24826 = n24825 ^ n24824 ;
  assign n24821 = n3520 & n21124 ;
  assign n24820 = n24383 ^ n3520 ;
  assign n24822 = n24821 ^ n24820 ;
  assign n24823 = x31 & n24822 ;
  assign n24827 = n24826 ^ n24823 ;
  assign n24842 = n24841 ^ n24827 ;
  assign n24817 = n24391 ^ n24375 ;
  assign n24818 = n24388 & ~n24817 ;
  assign n24819 = n24818 ^ n24391 ;
  assign n24843 = n24842 ^ n24819 ;
  assign n24814 = n3484 & n20970 ;
  assign n24807 = n20963 ^ x29 ;
  assign n24808 = n24807 ^ x28 ;
  assign n24809 = n24808 ^ n20963 ;
  assign n24810 = ~n21686 & n24809 ;
  assign n24811 = n24810 ^ n20963 ;
  assign n24812 = n650 & ~n24811 ;
  assign n24813 = n24812 ^ x29 ;
  assign n24815 = n24814 ^ n24813 ;
  assign n24806 = n831 & ~n20924 ;
  assign n24816 = n24815 ^ n24806 ;
  assign n24844 = n24843 ^ n24816 ;
  assign n24803 = n24357 ^ n24346 ;
  assign n24804 = ~n24393 & n24803 ;
  assign n24805 = n24804 ^ n24357 ;
  assign n24845 = n24844 ^ n24805 ;
  assign n24846 = n24845 ^ x26 ;
  assign n24848 = n24847 ^ n24846 ;
  assign n24850 = n24849 ^ n24848 ;
  assign n24852 = n24851 ^ n24850 ;
  assign n24802 = ~n3501 & n21630 ;
  assign n24853 = n24852 ^ n24802 ;
  assign n24799 = n24339 & ~n24394 ;
  assign n24798 = n24394 ^ n24339 ;
  assign n24800 = n24799 ^ n24798 ;
  assign n24854 = n24853 ^ n24800 ;
  assign n24879 = n24395 & ~n24854 ;
  assign n24871 = ~n24331 & ~n24399 ;
  assign n24795 = n24394 ^ n24342 ;
  assign n24796 = ~n24343 & ~n24795 ;
  assign n24797 = n24796 ^ n24394 ;
  assign n24872 = n24799 ^ n24797 ;
  assign n24875 = n24853 & n24872 ;
  assign n24876 = n24875 ^ n24799 ;
  assign n24877 = n24871 & ~n24876 ;
  assign n24860 = n24399 ^ n24331 ;
  assign n24880 = n24877 ^ n24860 ;
  assign n24881 = n24879 & n24880 ;
  assign n24878 = n24877 ^ n24871 ;
  assign n24882 = n24881 ^ n24878 ;
  assign n24794 = n24331 & n24399 ;
  assign n24801 = n24800 ^ n24797 ;
  assign n24856 = ~n24801 & n24853 ;
  assign n24857 = n24856 ^ n24800 ;
  assign n24858 = n24794 & ~n24857 ;
  assign n24861 = n24860 ^ n24858 ;
  assign n24862 = n24853 ^ n24342 ;
  assign n24863 = n24862 ^ n24853 ;
  assign n24864 = n24853 ^ n24394 ;
  assign n24865 = n24864 ^ n24853 ;
  assign n24866 = n24863 & ~n24865 ;
  assign n24867 = n24866 ^ n24853 ;
  assign n24868 = ~n24395 & ~n24867 ;
  assign n24869 = n24861 & n24868 ;
  assign n24859 = n24858 ^ n24794 ;
  assign n24870 = n24869 ^ n24859 ;
  assign n24883 = n24882 ^ n24870 ;
  assign n24892 = n24891 ^ n24883 ;
  assign n24893 = n24892 ^ x20 ;
  assign n24789 = n21735 ^ n4685 ;
  assign n24790 = n24789 ^ n21735 ;
  assign n24791 = ~n21734 & ~n24790 ;
  assign n24792 = n24791 ^ n21735 ;
  assign n24793 = n4678 & n24792 ;
  assign n24894 = n24893 ^ n24793 ;
  assign n24896 = n24895 ^ n24894 ;
  assign n24788 = n14027 & n20903 ;
  assign n24897 = n24896 ^ n24788 ;
  assign n24785 = n24320 ^ n24308 ;
  assign n24786 = ~n24401 & n24785 ;
  assign n24787 = n24786 ^ n24320 ;
  assign n24898 = n24897 ^ n24787 ;
  assign n24899 = n24898 ^ x17 ;
  assign n24901 = n24900 ^ n24899 ;
  assign n24903 = n24902 ^ n24901 ;
  assign n24905 = n24904 ^ n24903 ;
  assign n24784 = n20731 & n20898 ;
  assign n24906 = n24905 ^ n24784 ;
  assign n24781 = n24402 ^ n24300 ;
  assign n24782 = ~n24409 & ~n24781 ;
  assign n24783 = n24782 ^ n24402 ;
  assign n24907 = n24906 ^ n24783 ;
  assign n24759 = x13 & ~x14 ;
  assign n24760 = ~n4898 & ~n20887 ;
  assign n24761 = n24759 & n24760 ;
  assign n24762 = n24761 ^ n4898 ;
  assign n24756 = n4896 & n15433 ;
  assign n24757 = ~n20887 & n24756 ;
  assign n24758 = n24757 ^ n4896 ;
  assign n24763 = n24762 ^ n24758 ;
  assign n24766 = n24758 ^ x13 ;
  assign n24767 = n21025 & ~n24766 ;
  assign n24768 = n24767 ^ x13 ;
  assign n24769 = ~n24763 & ~n24768 ;
  assign n24770 = n24769 ^ n24762 ;
  assign n24771 = n24770 ^ x14 ;
  assign n24775 = n24771 ^ n6060 ;
  assign n24776 = x13 & ~n22545 ;
  assign n24777 = n24775 & n24776 ;
  assign n24773 = n6060 & n22546 ;
  assign n24772 = n20883 & n24771 ;
  assign n24774 = n24773 ^ n24772 ;
  assign n24778 = n24777 ^ n24774 ;
  assign n24779 = n24770 ^ n6062 ;
  assign n24780 = ~n24778 & ~n24779 ;
  assign n24908 = n24907 ^ n24780 ;
  assign n24753 = n24410 ^ n24293 ;
  assign n24754 = ~n24418 & ~n24753 ;
  assign n24755 = n24754 ^ n24410 ;
  assign n24909 = n24908 ^ n24755 ;
  assign n24743 = n6655 & n20882 ;
  assign n24742 = n6658 & ~n20872 ;
  assign n24744 = n24743 ^ n24742 ;
  assign n24745 = n24744 ^ x11 ;
  assign n24741 = n15413 & n23033 ;
  assign n24746 = n24745 ^ n24741 ;
  assign n24740 = n6650 & ~n20876 ;
  assign n24747 = n24746 ^ n24740 ;
  assign n24749 = n24747 ^ n24285 ;
  assign n24748 = n24747 ^ n24419 ;
  assign n24750 = n24749 ^ n24748 ;
  assign n24751 = ~n24290 & ~n24750 ;
  assign n24752 = n24751 ^ n24749 ;
  assign n24910 = n24909 ^ n24752 ;
  assign n24912 = n24910 ^ n24269 ;
  assign n24911 = n24910 ^ n24420 ;
  assign n24913 = n24912 ^ n24911 ;
  assign n24914 = n24277 & n24913 ;
  assign n24915 = n24914 ^ n24912 ;
  assign n24924 = n24923 ^ n24915 ;
  assign n24946 = n24945 ^ n24924 ;
  assign n24993 = n24992 ^ n24946 ;
  assign n24706 = n24079 ^ n20834 ;
  assign n24707 = n24706 ^ n24079 ;
  assign n24463 = n24462 ^ n24461 ;
  assign n24701 = n24700 ^ x1 ;
  assign n24703 = n24702 ^ n24701 ;
  assign n24704 = n24463 & n24703 ;
  assign n24705 = n24704 ^ n24701 ;
  assign n24081 = n24079 ^ x2 ;
  assign n24708 = n24705 ^ n24081 ;
  assign n24709 = n24708 ^ n24705 ;
  assign n24710 = n24709 ^ n24079 ;
  assign n24711 = n24707 & n24710 ;
  assign n24712 = n24711 ^ n24079 ;
  assign n24713 = ~x1 & n24712 ;
  assign n24714 = n24713 ^ n24708 ;
  assign n24715 = ~x0 & ~n24714 ;
  assign n24716 = n24715 ^ n24705 ;
  assign n24451 = n24443 ^ n24440 ;
  assign n24452 = n24451 ^ n24100 ;
  assign n24431 = n24430 ^ n24100 ;
  assign n24453 = n24431 ^ n24430 ;
  assign n24732 = ~n24440 & ~n24453 ;
  assign n24733 = n24732 ^ n24430 ;
  assign n24734 = ~n24452 & n24733 ;
  assign n23047 = n20861 ^ n20852 ;
  assign n23048 = n23047 ^ n20852 ;
  assign n23049 = n20852 ^ x2 ;
  assign n23052 = n23049 ^ n20852 ;
  assign n23053 = n23048 & n23052 ;
  assign n23054 = n23053 ^ n20852 ;
  assign n23055 = ~x1 & n23054 ;
  assign n23042 = n20836 ^ x1 ;
  assign n21068 = n20836 ^ x2 ;
  assign n23043 = n23042 ^ n21068 ;
  assign n23044 = n23041 & n23043 ;
  assign n23045 = n23044 ^ n23042 ;
  assign n23050 = n23049 ^ n23045 ;
  assign n23056 = n23055 ^ n23050 ;
  assign n23057 = ~x0 & n23056 ;
  assign n23039 = n23038 ^ n22686 ;
  assign n23046 = n23045 ^ n23039 ;
  assign n23058 = n23057 ^ n23046 ;
  assign n23613 = n20872 ^ n20865 ;
  assign n23614 = n23613 ^ n20865 ;
  assign n23609 = n20861 ^ x1 ;
  assign n23066 = n20861 ^ x2 ;
  assign n23610 = n23609 ^ n23066 ;
  assign n23611 = n23608 & n23610 ;
  assign n23612 = n23611 ^ n23609 ;
  assign n23078 = n20865 ^ x2 ;
  assign n23615 = n23612 ^ n23078 ;
  assign n23616 = n23615 ^ n23612 ;
  assign n23617 = n23616 ^ n20865 ;
  assign n23618 = ~n23614 & n23617 ;
  assign n23619 = n23618 ^ n20865 ;
  assign n23620 = ~x1 & n23619 ;
  assign n23621 = n23620 ^ n23615 ;
  assign n23622 = ~x0 & n23621 ;
  assign n23623 = n23622 ^ n23612 ;
  assign n23086 = n20872 ^ x2 ;
  assign n23089 = n23086 ^ n20872 ;
  assign n23090 = ~n20876 & n23089 ;
  assign n23091 = n23090 ^ n20872 ;
  assign n23092 = ~x1 & ~n23091 ;
  assign n23077 = n20865 ^ x1 ;
  assign n23079 = n23078 ^ n23077 ;
  assign n23080 = n22682 & n23079 ;
  assign n23081 = n23080 ^ n23077 ;
  assign n23087 = n23086 ^ n23081 ;
  assign n23093 = n23092 ^ n23087 ;
  assign n23094 = ~x0 & ~n23093 ;
  assign n23082 = n23001 ^ n22696 ;
  assign n23083 = n23082 ^ n23081 ;
  assign n23095 = n23094 ^ n23083 ;
  assign n23120 = n20882 ^ x2 ;
  assign n23123 = n23120 ^ n20882 ;
  assign n23124 = n20883 & n23123 ;
  assign n23125 = n23124 ^ n20882 ;
  assign n23126 = ~x1 & n23125 ;
  assign n23112 = n20876 ^ x1 ;
  assign n23102 = n20876 ^ x2 ;
  assign n23113 = n23112 ^ n23102 ;
  assign n23114 = n23009 & n23113 ;
  assign n23115 = n23114 ^ n23112 ;
  assign n23121 = n23120 ^ n23115 ;
  assign n23127 = n23126 ^ n23121 ;
  assign n23128 = ~x0 & ~n23127 ;
  assign n23116 = n22995 ^ n22716 ;
  assign n23117 = n23116 ^ n23115 ;
  assign n23129 = n23128 ^ n23117 ;
  assign n23152 = n21025 ^ n20887 ;
  assign n23153 = n23152 ^ n21025 ;
  assign n23154 = n21025 ^ x2 ;
  assign n23157 = n23154 ^ n23152 ;
  assign n23158 = ~n23153 & ~n23157 ;
  assign n23159 = n23158 ^ n23152 ;
  assign n23160 = ~x1 & n23159 ;
  assign n23146 = n20883 ^ x1 ;
  assign n23136 = n20883 ^ x2 ;
  assign n23147 = n23146 ^ n23136 ;
  assign n23148 = n22545 & n23147 ;
  assign n23149 = n23148 ^ n23146 ;
  assign n23155 = n23154 ^ n23149 ;
  assign n23161 = n23160 ^ n23155 ;
  assign n23162 = ~x0 & ~n23161 ;
  assign n23150 = n22989 ^ n22736 ;
  assign n23151 = n23150 ^ n23149 ;
  assign n23163 = n23162 ^ n23151 ;
  assign n23169 = n22987 ^ n22976 ;
  assign n23588 = n23169 ^ n23150 ;
  assign n23173 = n20887 ^ x2 ;
  assign n23176 = n23173 ^ n20887 ;
  assign n23177 = ~n20894 & n23176 ;
  assign n23178 = n23177 ^ n20887 ;
  assign n23179 = ~x1 & ~n23178 ;
  assign n23164 = n21025 ^ x1 ;
  assign n23165 = n23164 ^ x2 ;
  assign n23166 = n23165 ^ n21025 ;
  assign n23167 = n22414 & n23166 ;
  assign n23168 = n23167 ^ n23164 ;
  assign n23174 = n23173 ^ n23168 ;
  assign n23180 = n23179 ^ n23174 ;
  assign n23181 = ~x0 & n23180 ;
  assign n23170 = n23169 ^ n23168 ;
  assign n23182 = n23181 ^ n23170 ;
  assign n23187 = n22973 ^ n22746 ;
  assign n23585 = n23187 ^ n23169 ;
  assign n23191 = n20894 ^ x2 ;
  assign n23194 = n23191 ^ n20894 ;
  assign n23195 = n20897 & n23194 ;
  assign n23196 = n23195 ^ n20894 ;
  assign n23197 = ~x1 & ~n23196 ;
  assign n23183 = n20887 ^ x1 ;
  assign n23184 = n23183 ^ n23173 ;
  assign n23185 = n22306 & n23184 ;
  assign n23186 = n23185 ^ n23183 ;
  assign n23192 = n23191 ^ n23186 ;
  assign n23198 = n23197 ^ n23192 ;
  assign n23199 = ~x0 & n23198 ;
  assign n23188 = n23187 ^ n23186 ;
  assign n23200 = n23199 ^ n23188 ;
  assign n23208 = n20897 ^ x2 ;
  assign n23211 = n23208 ^ n20897 ;
  assign n23212 = n20898 & n23211 ;
  assign n23213 = n23212 ^ n20897 ;
  assign n23214 = ~x1 & n23213 ;
  assign n23202 = n20894 ^ x1 ;
  assign n23203 = n23202 ^ n23191 ;
  assign n23204 = n21953 & n23203 ;
  assign n23205 = n23204 ^ n23202 ;
  assign n23209 = n23208 ^ n23205 ;
  assign n23215 = n23214 ^ n23209 ;
  assign n23216 = ~x0 & ~n23215 ;
  assign n23217 = n23216 ^ n23205 ;
  assign n23582 = n23217 ^ n23187 ;
  assign n23226 = n20898 ^ x2 ;
  assign n23229 = n23226 ^ n20898 ;
  assign n23230 = ~n21012 & n23229 ;
  assign n23231 = n23230 ^ n20898 ;
  assign n23232 = ~x1 & n23231 ;
  assign n23219 = n20897 ^ x1 ;
  assign n23220 = n23219 ^ n23208 ;
  assign n23221 = n21965 & n23220 ;
  assign n23222 = n23221 ^ n23219 ;
  assign n23227 = n23226 ^ n23222 ;
  assign n23233 = n23232 ^ n23227 ;
  assign n23234 = ~x0 & n23233 ;
  assign n23201 = n22967 ^ n22766 ;
  assign n23223 = n23222 ^ n23201 ;
  assign n23235 = n23234 ^ n23223 ;
  assign n23261 = n20898 ^ x1 ;
  assign n23253 = n21012 ^ x2 ;
  assign n23254 = n23253 ^ n21012 ;
  assign n23255 = n21012 ^ n20902 ;
  assign n23256 = n23255 ^ n23253 ;
  assign n23257 = n23254 & n23256 ;
  assign n23258 = n23257 ^ n23253 ;
  assign n23259 = ~x1 & ~n23258 ;
  assign n23260 = n23259 ^ n23253 ;
  assign n23262 = n23261 ^ n23260 ;
  assign n23263 = n23262 ^ x2 ;
  assign n23264 = n23263 ^ x1 ;
  assign n23265 = n23264 ^ n23262 ;
  assign n23266 = n23262 ^ n21971 ;
  assign n23267 = n23266 ^ n23262 ;
  assign n23268 = n23265 & n23267 ;
  assign n23269 = n23268 ^ n23262 ;
  assign n23270 = x0 & ~n23269 ;
  assign n23271 = n23270 ^ n23260 ;
  assign n23575 = n23271 ^ n23201 ;
  assign n23252 = n22962 ^ n22948 ;
  assign n23272 = n23271 ^ n23252 ;
  assign n23273 = n23272 ^ n23271 ;
  assign n23238 = n21012 ^ x1 ;
  assign n23239 = n23238 ^ x2 ;
  assign n23240 = n23239 ^ n21012 ;
  assign n23241 = n21734 & n23240 ;
  assign n23242 = n23241 ^ n23238 ;
  assign n23274 = n23273 ^ n23242 ;
  assign n23243 = n20902 ^ x2 ;
  assign n23246 = n23243 ^ n20902 ;
  assign n23247 = n20903 & n23246 ;
  assign n23248 = n23247 ^ n20902 ;
  assign n23249 = ~x1 & n23248 ;
  assign n23244 = n23243 ^ n23242 ;
  assign n23250 = n23249 ^ n23244 ;
  assign n23251 = ~x0 & ~n23250 ;
  assign n23275 = n23274 ^ n23251 ;
  assign n23282 = n20903 ^ x1 ;
  assign n23281 = n20903 ^ x2 ;
  assign n23283 = n23282 ^ n23281 ;
  assign n23284 = n21755 & n23283 ;
  assign n23285 = n23284 ^ n23282 ;
  assign n23279 = n22942 ^ n22799 ;
  assign n23295 = n23285 ^ n23279 ;
  assign n23286 = n20910 ^ x2 ;
  assign n23289 = n23286 ^ n20910 ;
  assign n23290 = n20913 & n23289 ;
  assign n23291 = n23290 ^ n20910 ;
  assign n23292 = ~x1 & n23291 ;
  assign n23287 = n23286 ^ n23285 ;
  assign n23293 = n23292 ^ n23287 ;
  assign n23294 = ~x0 & n23293 ;
  assign n23296 = n23295 ^ n23294 ;
  assign n23303 = n20913 ^ x2 ;
  assign n23306 = n23303 ^ n20913 ;
  assign n23307 = ~n20922 & n23306 ;
  assign n23308 = n23307 ^ n20913 ;
  assign n23309 = ~x1 & n23308 ;
  assign n23298 = n20910 ^ x1 ;
  assign n23299 = n23298 ^ n23286 ;
  assign n23300 = ~n21000 & n23299 ;
  assign n23301 = n23300 ^ n23298 ;
  assign n23304 = n23303 ^ n23301 ;
  assign n23310 = n23309 ^ n23304 ;
  assign n23311 = ~x0 & n23310 ;
  assign n23312 = n23311 ^ n23301 ;
  assign n23297 = n22939 ^ n22931 ;
  assign n23313 = n23312 ^ n23297 ;
  assign n23546 = n23312 ^ n23279 ;
  assign n23315 = n22926 ^ n22809 ;
  assign n23544 = n23315 ^ n23279 ;
  assign n23319 = n20922 ^ x2 ;
  assign n23318 = n20922 ^ x1 ;
  assign n23320 = n23319 ^ n23318 ;
  assign n23321 = ~n21395 & n23320 ;
  assign n23322 = n23321 ^ n23318 ;
  assign n23314 = n22923 ^ n22819 ;
  assign n23332 = n23322 ^ n23314 ;
  assign n23317 = n21394 ^ n20994 ;
  assign n23327 = x2 & n23317 ;
  assign n23328 = n23327 ^ n20994 ;
  assign n23329 = ~x1 & n23328 ;
  assign n23323 = n20994 ^ x2 ;
  assign n23324 = n23323 ^ n23322 ;
  assign n23330 = n23329 ^ n23324 ;
  assign n23331 = ~x0 & ~n23330 ;
  assign n23333 = n23332 ^ n23331 ;
  assign n23338 = n21630 ^ x2 ;
  assign n23337 = n20994 ^ x1 ;
  assign n23339 = n23338 ^ n23337 ;
  assign n23340 = ~n20991 & n23339 ;
  assign n23341 = n23340 ^ n23337 ;
  assign n23336 = n20962 ^ x2 ;
  assign n23342 = n23341 ^ n23336 ;
  assign n23343 = n23342 ^ n23341 ;
  assign n23344 = n23343 ^ n20962 ;
  assign n23345 = ~n20969 & n23344 ;
  assign n23346 = n23345 ^ n20962 ;
  assign n23347 = ~x1 & n23346 ;
  assign n23348 = n23347 ^ n23342 ;
  assign n23349 = ~x0 & n23348 ;
  assign n23350 = n23349 ^ n23341 ;
  assign n23334 = n22920 ^ n22829 ;
  assign n23351 = n23350 ^ n23334 ;
  assign n23519 = n23350 ^ n23314 ;
  assign n23353 = n22917 ^ n22839 ;
  assign n23517 = n23353 ^ n23314 ;
  assign n23376 = n22903 ^ n22858 ;
  assign n23377 = ~n22904 & n23376 ;
  assign n23356 = n20970 ^ n20924 ;
  assign n23357 = n23356 ^ n20970 ;
  assign n23358 = n20970 ^ x2 ;
  assign n23359 = n23358 ^ n20970 ;
  assign n23360 = ~n23357 & n23359 ;
  assign n23361 = n23360 ^ n20970 ;
  assign n23362 = ~x1 & n23361 ;
  assign n23363 = n23362 ^ n23358 ;
  assign n23355 = n20963 ^ x1 ;
  assign n23364 = n23363 ^ n23355 ;
  assign n23365 = n23364 ^ x2 ;
  assign n23366 = n23365 ^ x1 ;
  assign n23367 = n23366 ^ n23364 ;
  assign n23368 = n23364 ^ n21239 ;
  assign n23369 = n23368 ^ n23364 ;
  assign n23370 = n23367 & n23369 ;
  assign n23371 = n23370 ^ n23364 ;
  assign n23372 = x0 & ~n23371 ;
  assign n23373 = n23372 ^ n23363 ;
  assign n23375 = n23373 ^ n22868 ;
  assign n23378 = n23377 ^ n23375 ;
  assign n23450 = n22899 ^ n22890 ;
  assign n23451 = n23450 ^ n22870 ;
  assign n23441 = x2 & ~n20939 ;
  assign n23429 = n20941 ^ n10828 ;
  assign n23430 = n23429 ^ n20941 ;
  assign n23431 = n21170 & n23430 ;
  assign n23432 = n23431 ^ n20941 ;
  assign n23433 = x0 & n23432 ;
  assign n23442 = n21142 & ~n23433 ;
  assign n23443 = n23441 & n23442 ;
  assign n23437 = n10854 & n20926 ;
  assign n23435 = n10850 & n20939 ;
  assign n23434 = n23433 ^ x3 ;
  assign n23436 = n23435 ^ n23434 ;
  assign n23438 = n23437 ^ n23436 ;
  assign n23439 = n9077 & ~n23438 ;
  assign n23440 = ~n20927 & n23439 ;
  assign n23444 = n23443 ^ n23440 ;
  assign n22876 = n22875 ^ x5 ;
  assign n23407 = n22889 ^ n22876 ;
  assign n23403 = n10854 & n20941 ;
  assign n23402 = n10850 & ~n20925 ;
  assign n23404 = n23403 ^ n23402 ;
  assign n23397 = n20499 ^ n10828 ;
  assign n23398 = n23397 ^ n20499 ;
  assign n23399 = ~n21123 & n23398 ;
  assign n23400 = n23399 ^ n20499 ;
  assign n23401 = x0 & n23400 ;
  assign n23405 = n23404 ^ n23401 ;
  assign n23406 = n23405 ^ x2 ;
  assign n23408 = n23407 ^ n23406 ;
  assign n23417 = n10854 & n20939 ;
  assign n23416 = n10850 & n20941 ;
  assign n23418 = n23417 ^ n23416 ;
  assign n23411 = n20925 ^ n10828 ;
  assign n23412 = n23411 ^ n20925 ;
  assign n23413 = n21187 & n23412 ;
  assign n23414 = n23413 ^ n20925 ;
  assign n23415 = x0 & ~n23414 ;
  assign n23419 = n23418 ^ n23415 ;
  assign n23445 = n23419 ^ x2 ;
  assign n23422 = n11206 & ~n20927 ;
  assign n23423 = n23422 ^ n22871 ;
  assign n23446 = n23445 ^ n23423 ;
  assign n23447 = ~n23408 & n23446 ;
  assign n23448 = n23444 & n23447 ;
  assign n23449 = n23448 ^ n23407 ;
  assign n23452 = n23451 ^ n23449 ;
  assign n23420 = n23419 ^ n23405 ;
  assign n23421 = n23420 ^ n23407 ;
  assign n23424 = n23423 ^ n23407 ;
  assign n23425 = n23424 ^ n23407 ;
  assign n23426 = n23421 & n23425 ;
  assign n23427 = n23426 ^ n23407 ;
  assign n23428 = ~n23408 & ~n23427 ;
  assign n23453 = n23452 ^ n23428 ;
  assign n23458 = n10828 & n21210 ;
  assign n23456 = n20924 ^ x1 ;
  assign n23459 = n23458 ^ n23456 ;
  assign n23469 = n23459 ^ n23451 ;
  assign n23460 = n20499 ^ x2 ;
  assign n23463 = n23460 ^ n20499 ;
  assign n23464 = ~n20925 & n23463 ;
  assign n23465 = n23464 ^ n20499 ;
  assign n23466 = ~x1 & n23465 ;
  assign n23461 = n23460 ^ n23459 ;
  assign n23467 = n23466 ^ n23461 ;
  assign n23468 = ~x0 & ~n23467 ;
  assign n23470 = n23469 ^ n23468 ;
  assign n23471 = ~n23453 & ~n23470 ;
  assign n23472 = n23471 ^ n23451 ;
  assign n23477 = n23472 ^ n23373 ;
  assign n23383 = n20924 ^ n20499 ;
  assign n23384 = n23383 ^ n20924 ;
  assign n23389 = x2 & n23384 ;
  assign n23390 = n23389 ^ n20924 ;
  assign n23391 = ~x1 & ~n23390 ;
  assign n23385 = n20924 ^ x2 ;
  assign n23379 = n20970 ^ x1 ;
  assign n23380 = n23379 ^ n23358 ;
  assign n23381 = n20954 & n23380 ;
  assign n23382 = n23381 ^ n23379 ;
  assign n23386 = n23385 ^ n23382 ;
  assign n23392 = n23391 ^ n23386 ;
  assign n23393 = ~x0 & ~n23392 ;
  assign n23394 = n23393 ^ n23382 ;
  assign n23473 = n23472 ^ n23394 ;
  assign n23474 = n22904 ^ n22858 ;
  assign n23475 = n23474 ^ n23394 ;
  assign n23476 = n23473 & ~n23475 ;
  assign n23478 = n23477 ^ n23476 ;
  assign n23479 = n23378 & n23478 ;
  assign n23352 = n22914 ^ n22850 ;
  assign n23374 = n23373 ^ n23352 ;
  assign n23480 = n23479 ^ n23374 ;
  assign n23484 = n20969 ^ x1 ;
  assign n23483 = n20969 ^ x2 ;
  assign n23485 = n23484 ^ n23483 ;
  assign n23486 = n21106 & n23485 ;
  assign n23487 = n23486 ^ n23484 ;
  assign n23497 = n23487 ^ n23352 ;
  assign n23488 = n20963 ^ x2 ;
  assign n23491 = n23488 ^ n20963 ;
  assign n23492 = n20970 & n23491 ;
  assign n23493 = n23492 ^ n20963 ;
  assign n23494 = ~x1 & ~n23493 ;
  assign n23489 = n23488 ^ n23487 ;
  assign n23495 = n23494 ^ n23489 ;
  assign n23496 = ~x0 & n23495 ;
  assign n23498 = n23497 ^ n23496 ;
  assign n23499 = n23480 & ~n23498 ;
  assign n23354 = n23353 ^ n23352 ;
  assign n23500 = n23499 ^ n23354 ;
  assign n23502 = n20962 ^ x1 ;
  assign n23503 = n23502 ^ n23336 ;
  assign n23504 = ~n21108 & n23503 ;
  assign n23505 = n23504 ^ n23502 ;
  assign n23514 = n23505 ^ n23353 ;
  assign n23501 = n20974 ^ n20969 ;
  assign n23506 = n23505 ^ n23483 ;
  assign n23507 = n23506 ^ n23505 ;
  assign n23508 = n23507 ^ n20969 ;
  assign n23509 = ~n23501 & n23508 ;
  assign n23510 = n23509 ^ n20969 ;
  assign n23511 = ~x1 & ~n23510 ;
  assign n23512 = n23511 ^ n23506 ;
  assign n23513 = ~x0 & ~n23512 ;
  assign n23515 = n23514 ^ n23513 ;
  assign n23516 = n23500 & n23515 ;
  assign n23518 = n23517 ^ n23516 ;
  assign n23520 = n23519 ^ n23518 ;
  assign n23521 = ~n23351 & n23520 ;
  assign n23522 = n23521 ^ n23518 ;
  assign n23523 = ~n23333 & n23522 ;
  assign n23316 = n23315 ^ n23314 ;
  assign n23524 = n23523 ^ n23316 ;
  assign n23525 = n20995 ^ n20922 ;
  assign n23526 = n23319 ^ n20922 ;
  assign n23527 = n23525 & n23526 ;
  assign n23528 = n23527 ^ n20922 ;
  assign n23529 = ~x1 & ~n23528 ;
  assign n23530 = n23529 ^ n23319 ;
  assign n23541 = n23530 ^ n23315 ;
  assign n23531 = n20913 ^ x1 ;
  assign n23532 = n23531 ^ n23530 ;
  assign n23533 = n23532 ^ x2 ;
  assign n23534 = n23533 ^ x1 ;
  assign n23535 = n23534 ^ n23532 ;
  assign n23536 = n23532 ^ n20999 ;
  assign n23537 = n23536 ^ n23532 ;
  assign n23538 = n23535 & n23537 ;
  assign n23539 = n23538 ^ n23532 ;
  assign n23540 = x0 & ~n23539 ;
  assign n23542 = n23541 ^ n23540 ;
  assign n23543 = n23524 & ~n23542 ;
  assign n23545 = n23544 ^ n23543 ;
  assign n23547 = n23546 ^ n23545 ;
  assign n23548 = n23313 & n23547 ;
  assign n23549 = n23548 ^ n23545 ;
  assign n23550 = ~n23296 & ~n23549 ;
  assign n23276 = n22945 ^ n22789 ;
  assign n23280 = n23279 ^ n23276 ;
  assign n23551 = n23550 ^ n23280 ;
  assign n23554 = n20902 ^ x1 ;
  assign n23555 = n23554 ^ n23243 ;
  assign n23556 = n21743 & n23555 ;
  assign n23557 = n23556 ^ n23554 ;
  assign n23566 = n23557 ^ n23276 ;
  assign n23552 = n20910 ^ n20903 ;
  assign n23553 = n23552 ^ n20903 ;
  assign n23558 = n23557 ^ n23281 ;
  assign n23559 = n23558 ^ n23557 ;
  assign n23560 = n23559 ^ n20903 ;
  assign n23561 = n23553 & n23560 ;
  assign n23562 = n23561 ^ n20903 ;
  assign n23563 = ~x1 & n23562 ;
  assign n23564 = n23563 ^ n23558 ;
  assign n23565 = ~x0 & n23564 ;
  assign n23567 = n23566 ^ n23565 ;
  assign n23568 = n23551 & ~n23567 ;
  assign n23277 = n23276 ^ n23271 ;
  assign n23278 = n23277 ^ n23272 ;
  assign n23569 = n23568 ^ n23278 ;
  assign n23570 = ~n23275 & ~n23569 ;
  assign n23571 = n23570 ^ n23272 ;
  assign n23572 = n23271 ^ n22964 ;
  assign n23573 = n23572 ^ n22779 ;
  assign n23574 = ~n23571 & ~n23573 ;
  assign n23576 = n23575 ^ n23574 ;
  assign n23577 = ~n23235 & n23576 ;
  assign n23218 = n23217 ^ n23201 ;
  assign n23578 = n23577 ^ n23218 ;
  assign n23579 = n23217 ^ n22970 ;
  assign n23580 = n23579 ^ n22756 ;
  assign n23581 = n23578 & ~n23580 ;
  assign n23583 = n23582 ^ n23581 ;
  assign n23584 = ~n23200 & ~n23583 ;
  assign n23586 = n23585 ^ n23584 ;
  assign n23587 = n23182 & ~n23586 ;
  assign n23589 = n23588 ^ n23587 ;
  assign n23590 = ~n23163 & n23589 ;
  assign n23591 = n23590 ^ n23150 ;
  assign n23596 = n23591 ^ n23116 ;
  assign n23139 = n23136 ^ n20883 ;
  assign n23140 = ~n21025 & n23139 ;
  assign n23141 = n23140 ^ n20883 ;
  assign n23142 = ~x1 & n23141 ;
  assign n23130 = n20882 ^ x1 ;
  assign n23131 = n23130 ^ n23120 ;
  assign n23132 = n22671 & n23131 ;
  assign n23133 = n23132 ^ n23130 ;
  assign n23137 = n23136 ^ n23133 ;
  assign n23143 = n23142 ^ n23137 ;
  assign n23144 = ~x0 & n23143 ;
  assign n23145 = n23144 ^ n23133 ;
  assign n23592 = n23591 ^ n23145 ;
  assign n23593 = n22992 ^ n22726 ;
  assign n23594 = n23593 ^ n23145 ;
  assign n23595 = ~n23592 & ~n23594 ;
  assign n23597 = n23596 ^ n23595 ;
  assign n23598 = ~n23129 & ~n23597 ;
  assign n23599 = n23598 ^ n23116 ;
  assign n23604 = n23599 ^ n23082 ;
  assign n23105 = n23102 ^ n20876 ;
  assign n23106 = n20882 & n23105 ;
  assign n23107 = n23106 ^ n20876 ;
  assign n23108 = ~x1 & ~n23107 ;
  assign n23096 = n20872 ^ x1 ;
  assign n23097 = n23096 ^ n23086 ;
  assign n23098 = n23032 & n23097 ;
  assign n23099 = n23098 ^ n23096 ;
  assign n23103 = n23102 ^ n23099 ;
  assign n23109 = n23108 ^ n23103 ;
  assign n23110 = ~x0 & n23109 ;
  assign n23111 = n23110 ^ n23099 ;
  assign n23600 = n23599 ^ n23111 ;
  assign n23601 = n22998 ^ n22706 ;
  assign n23602 = n23601 ^ n23111 ;
  assign n23603 = ~n23600 & ~n23602 ;
  assign n23605 = n23604 ^ n23603 ;
  assign n23606 = ~n23095 & ~n23605 ;
  assign n23607 = n23606 ^ n23082 ;
  assign n23624 = n23623 ^ n23607 ;
  assign n23625 = n23021 ^ n23004 ;
  assign n23626 = n23625 ^ n23607 ;
  assign n23627 = ~n23624 & n23626 ;
  assign n23628 = n23627 ^ n23623 ;
  assign n23069 = n23066 ^ n20861 ;
  assign n23070 = n20865 & n23069 ;
  assign n23071 = n23070 ^ n20861 ;
  assign n23072 = ~x1 & n23071 ;
  assign n23060 = n20852 ^ x1 ;
  assign n23061 = n23060 ^ n23049 ;
  assign n23062 = n23059 & n23061 ;
  assign n23063 = n23062 ^ n23060 ;
  assign n23067 = n23066 ^ n23063 ;
  assign n23073 = n23072 ^ n23067 ;
  assign n23074 = ~x0 & n23073 ;
  assign n23075 = n23074 ^ n23063 ;
  assign n23629 = n23628 ^ n23075 ;
  assign n23630 = n23036 ^ n23023 ;
  assign n23631 = n23630 ^ n23628 ;
  assign n23632 = n23629 & n23631 ;
  assign n23076 = n23075 ^ n23039 ;
  assign n23633 = n23632 ^ n23076 ;
  assign n23634 = ~n23058 & ~n23633 ;
  assign n21062 = n20837 ^ x1 ;
  assign n20840 = n20837 ^ x2 ;
  assign n21063 = n21062 ^ n20840 ;
  assign n21064 = n21061 & n21063 ;
  assign n21065 = n21064 ^ n21062 ;
  assign n21069 = n21068 ^ n21065 ;
  assign n21070 = n21069 ^ n21065 ;
  assign n21071 = n21070 ^ n20836 ;
  assign n21072 = n20852 & n21071 ;
  assign n21073 = n21072 ^ n20836 ;
  assign n21074 = ~x1 & n21073 ;
  assign n21075 = n21074 ^ n21069 ;
  assign n21076 = ~x0 & n21075 ;
  assign n21077 = n21076 ^ n21065 ;
  assign n23040 = n23039 ^ n21077 ;
  assign n23635 = n23634 ^ n23040 ;
  assign n23815 = n23814 ^ n21077 ;
  assign n23816 = n23815 ^ n23638 ;
  assign n23817 = ~n23635 & n23816 ;
  assign n23818 = n23817 ^ n21077 ;
  assign n20838 = n20837 ^ n20836 ;
  assign n20839 = n20838 ^ n20837 ;
  assign n20841 = n20840 ^ n20837 ;
  assign n20842 = n20839 & n20841 ;
  assign n20843 = n20842 ^ n20837 ;
  assign n20844 = ~x1 & n20843 ;
  assign n20845 = n20844 ^ n20840 ;
  assign n23819 = n23818 ^ n20845 ;
  assign n20835 = n20834 ^ x1 ;
  assign n20846 = n20845 ^ n20835 ;
  assign n20847 = n20846 ^ x2 ;
  assign n20848 = n20847 ^ x1 ;
  assign n20849 = n20848 ^ n20846 ;
  assign n21058 = n20849 & n21055 ;
  assign n21059 = n21058 ^ n20846 ;
  assign n21060 = x0 & n21059 ;
  assign n23820 = n23819 ^ n21060 ;
  assign n23834 = n23833 ^ n23818 ;
  assign n23999 = n23998 ^ n23834 ;
  assign n24000 = n23820 & n23999 ;
  assign n24001 = n24000 ^ n23818 ;
  assign n24087 = n20834 ^ x2 ;
  assign n24004 = n24003 ^ n24002 ;
  assign n24080 = n24079 ^ x1 ;
  assign n24082 = n24081 ^ n24080 ;
  assign n24083 = n24004 & n24082 ;
  assign n24084 = n24083 ^ n24080 ;
  assign n24088 = n24087 ^ n24084 ;
  assign n24089 = n24088 ^ n24084 ;
  assign n24090 = n24089 ^ n20834 ;
  assign n24091 = n20837 & n24090 ;
  assign n24092 = n24091 ^ n20834 ;
  assign n24093 = ~x1 & n24092 ;
  assign n24094 = n24093 ^ n24088 ;
  assign n24095 = ~x0 & n24094 ;
  assign n24096 = n24095 ^ n24084 ;
  assign n24720 = ~n24001 & ~n24096 ;
  assign n24441 = n24440 ^ n24430 ;
  assign n24721 = n24451 ^ n24441 ;
  assign n24722 = n24721 ^ n24441 ;
  assign n24723 = n24443 ^ n24441 ;
  assign n24724 = ~n24100 & n24723 ;
  assign n24725 = n24724 ^ n24441 ;
  assign n24726 = n24722 & ~n24725 ;
  assign n24727 = n24726 ^ n24441 ;
  assign n24728 = n24720 & ~n24727 ;
  assign n24729 = n24728 ^ n24720 ;
  assign n24449 = n24096 ^ n24001 ;
  assign n24735 = n24729 ^ n24449 ;
  assign n24736 = n24734 & n24735 ;
  assign n24737 = n24736 ^ n24728 ;
  assign n24738 = n24716 & n24737 ;
  assign n24097 = n24001 & n24096 ;
  assign n24442 = n24441 ^ n24431 ;
  assign n24444 = n24443 ^ n24430 ;
  assign n24445 = n24444 ^ n24441 ;
  assign n24446 = n24442 & n24445 ;
  assign n24447 = n24446 ^ n24441 ;
  assign n24448 = n24097 & ~n24447 ;
  assign n24459 = n24448 ^ n24097 ;
  assign n24450 = n24449 ^ n24448 ;
  assign n24454 = n24444 ^ n24430 ;
  assign n24455 = n24453 & n24454 ;
  assign n24456 = n24455 ^ n24430 ;
  assign n24457 = n24452 & n24456 ;
  assign n24458 = n24450 & n24457 ;
  assign n24460 = n24459 ^ n24458 ;
  assign n24718 = ~n24460 & n24716 ;
  assign n24717 = n24716 ^ n24460 ;
  assign n24719 = n24718 ^ n24717 ;
  assign n24739 = n24738 ^ n24719 ;
  assign n24994 = n24993 ^ n24739 ;
  assign n25251 = n24980 ^ n24700 ;
  assign n25252 = n25251 ^ n24980 ;
  assign n25007 = ~n24948 & ~n24980 ;
  assign n25006 = ~n24947 & n24980 ;
  assign n25008 = n25007 ^ n25006 ;
  assign n25040 = n3942 ^ n476 ;
  assign n25035 = ~n24965 & n24970 ;
  assign n25038 = ~n24967 & n25035 ;
  assign n25034 = n24970 ^ n24965 ;
  assign n25036 = n25035 ^ n25034 ;
  assign n25037 = n24967 & n25036 ;
  assign n25039 = n25038 ^ n25037 ;
  assign n25041 = n25040 ^ n25039 ;
  assign n25027 = ~n12755 & n24214 ;
  assign n25028 = n25027 ^ n33 ;
  assign n25029 = x31 & ~n20645 ;
  assign n25030 = ~n25028 & n25029 ;
  assign n25031 = n25030 ^ n25028 ;
  assign n25032 = n25031 ^ n24952 ;
  assign n25024 = n24972 ^ n24952 ;
  assign n25025 = n24957 & n25024 ;
  assign n25026 = n25025 ^ n24952 ;
  assign n25033 = n25032 ^ n25026 ;
  assign n25042 = n25041 ^ n25033 ;
  assign n25018 = n24976 ^ n24668 ;
  assign n25009 = n24608 & n24611 ;
  assign n25010 = n24973 ^ n24696 ;
  assign n25011 = n24973 ^ n24668 ;
  assign n25012 = n24974 ^ n24973 ;
  assign n25013 = n25011 & n25012 ;
  assign n25014 = n25010 & n25013 ;
  assign n25015 = n25014 ^ n25010 ;
  assign n25016 = n25015 ^ n24696 ;
  assign n25017 = ~n25009 & ~n25016 ;
  assign n25019 = n25009 ^ n24973 ;
  assign n25020 = n25019 ^ n24978 ;
  assign n25021 = ~n25017 & n25020 ;
  assign n25022 = ~n25018 & n25021 ;
  assign n25023 = n25022 ^ n25017 ;
  assign n25043 = n25042 ^ n25023 ;
  assign n25044 = n25043 ^ x1 ;
  assign n25045 = n25044 ^ x2 ;
  assign n25046 = n25045 ^ n25043 ;
  assign n25047 = n25008 & n25046 ;
  assign n25048 = n25047 ^ n25044 ;
  assign n25253 = n25048 ^ n24981 ;
  assign n25254 = n25253 ^ n25048 ;
  assign n25255 = n25254 ^ n24980 ;
  assign n25256 = ~n25252 & n25255 ;
  assign n25257 = n25256 ^ n24980 ;
  assign n25258 = ~x1 & ~n25257 ;
  assign n25259 = n25258 ^ n25253 ;
  assign n25260 = ~x0 & ~n25259 ;
  assign n25245 = n24079 ^ n24004 ;
  assign n25053 = ~x4 & ~n24004 ;
  assign n25246 = n25245 ^ n25053 ;
  assign n25247 = n19158 & ~n25246 ;
  assign n25235 = n7146 & n20861 ;
  assign n25234 = n8054 & n20836 ;
  assign n25236 = n25235 ^ n25234 ;
  assign n25237 = n25236 ^ x8 ;
  assign n25233 = n7135 & ~n24433 ;
  assign n25238 = n25237 ^ n25233 ;
  assign n25232 = n7141 & n20852 ;
  assign n25239 = n25238 ^ n25232 ;
  assign n25213 = n6655 & ~n20876 ;
  assign n25212 = n6650 & ~n20872 ;
  assign n25214 = n25213 ^ n25212 ;
  assign n25215 = n25214 ^ n6656 ;
  assign n25216 = n25215 ^ x11 ;
  assign n25217 = n25214 ^ x11 ;
  assign n25221 = n25217 ^ n6657 ;
  assign n25222 = ~x10 & ~n22682 ;
  assign n25223 = n25221 & n25222 ;
  assign n25219 = n6657 & ~n22683 ;
  assign n25218 = ~n20865 & n25217 ;
  assign n25220 = n25219 ^ n25218 ;
  assign n25224 = n25223 ^ n25220 ;
  assign n25225 = ~n25216 & ~n25224 ;
  assign n25062 = ~n6072 & ~n21025 ;
  assign n25061 = ~n6074 & n20883 ;
  assign n25063 = n25062 ^ n25061 ;
  assign n25195 = n5703 & n22307 ;
  assign n25188 = n4916 & ~n21012 ;
  assign n25182 = ~n24870 & ~n24890 ;
  assign n25183 = n25182 ^ x23 ;
  assign n25184 = ~n24883 & n25183 ;
  assign n25177 = n4504 & n20913 ;
  assign n25176 = n4491 & n20903 ;
  assign n25178 = n25177 ^ n25176 ;
  assign n25174 = ~n4496 & n20910 ;
  assign n25173 = n4492 & ~n21756 ;
  assign n25175 = n25174 ^ n25173 ;
  assign n25179 = n25178 ^ n25175 ;
  assign n25172 = n24882 ^ x23 ;
  assign n25180 = n25179 ^ n25172 ;
  assign n25160 = n12861 & n20962 ;
  assign n25159 = n446 & n20994 ;
  assign n25161 = n25160 ^ n25159 ;
  assign n25164 = n25161 ^ x26 ;
  assign n25165 = n25164 ^ n20922 ;
  assign n25162 = n67 ^ x25 ;
  assign n25163 = n21395 & ~n25162 ;
  assign n25166 = n25165 ^ n25163 ;
  assign n25167 = ~n25161 & n25166 ;
  assign n25168 = n25167 ^ n25164 ;
  assign n25169 = n64 & ~n25168 ;
  assign n25170 = n25169 ^ n25164 ;
  assign n25154 = n3484 & ~n20963 ;
  assign n25147 = n20969 ^ x29 ;
  assign n25148 = n25147 ^ x28 ;
  assign n25149 = n25148 ^ n20969 ;
  assign n25150 = ~n21106 & n25149 ;
  assign n25151 = n25150 ^ n20969 ;
  assign n25152 = n650 & ~n25151 ;
  assign n25153 = n25152 ^ x29 ;
  assign n25155 = n25154 ^ n25153 ;
  assign n25146 = n831 & n20970 ;
  assign n25156 = n25155 ^ n25146 ;
  assign n25122 = n3732 ^ x31 ;
  assign n25121 = ~n35 & n20499 ;
  assign n25132 = n25121 ^ n20925 ;
  assign n25133 = n25132 ^ n25121 ;
  assign n25135 = ~n25122 & ~n25133 ;
  assign n25136 = n25135 ^ n25121 ;
  assign n25137 = n13181 & ~n25136 ;
  assign n25128 = x31 & ~n20945 ;
  assign n25129 = n25128 ^ n20924 ;
  assign n25130 = n3520 & ~n25129 ;
  assign n25123 = n25122 ^ n25121 ;
  assign n25124 = n25123 ^ x31 ;
  assign n25131 = n25130 ^ n25124 ;
  assign n25138 = n25137 ^ n25131 ;
  assign n25115 = n24821 ^ n3720 ;
  assign n25116 = ~n13181 & ~n25115 ;
  assign n25117 = n25116 ^ n3720 ;
  assign n25118 = ~n20499 & ~n25117 ;
  assign n25139 = n25138 ^ n25118 ;
  assign n25097 = n13911 ^ n876 ;
  assign n25107 = n13883 ^ n2171 ;
  assign n25106 = n2076 ^ n1290 ;
  assign n25108 = n25107 ^ n25106 ;
  assign n25104 = n197 ^ n155 ;
  assign n25103 = n4780 ^ n296 ;
  assign n25105 = n25104 ^ n25103 ;
  assign n25109 = n25108 ^ n25105 ;
  assign n25110 = n25109 ^ n6490 ;
  assign n25100 = n2209 ^ n791 ;
  assign n25098 = n3539 ^ n1906 ;
  assign n25099 = n25098 ^ n1094 ;
  assign n25101 = n25100 ^ n25099 ;
  assign n25102 = n25101 ^ n6304 ;
  assign n25111 = n25110 ^ n25102 ;
  assign n25112 = n25111 ^ n3148 ;
  assign n25113 = ~n25097 & ~n25112 ;
  assign n25094 = n24827 ^ n24819 ;
  assign n25095 = ~n24842 & n25094 ;
  assign n25096 = n25095 ^ n24827 ;
  assign n25114 = n25113 ^ n25096 ;
  assign n25140 = n25139 ^ n25114 ;
  assign n25141 = n25140 ^ n24816 ;
  assign n25142 = n25141 ^ n25140 ;
  assign n25143 = n25142 ^ n24805 ;
  assign n25144 = ~n24844 & n25143 ;
  assign n25145 = n25144 ^ n25141 ;
  assign n25157 = n25156 ^ n25145 ;
  assign n25091 = n24845 ^ n24797 ;
  assign n25092 = ~n24853 & n25091 ;
  assign n25093 = n25092 ^ n24845 ;
  assign n25158 = n25157 ^ n25093 ;
  assign n25171 = n25170 ^ n25158 ;
  assign n25181 = n25180 ^ n25171 ;
  assign n25185 = n25184 ^ n25181 ;
  assign n25186 = n25185 ^ x20 ;
  assign n25086 = n20898 ^ n4685 ;
  assign n25087 = n25086 ^ n20898 ;
  assign n25088 = ~n21971 & n25087 ;
  assign n25089 = n25088 ^ n20898 ;
  assign n25090 = n4678 & n25089 ;
  assign n25187 = n25186 ^ n25090 ;
  assign n25189 = n25188 ^ n25187 ;
  assign n25085 = n14027 & n20902 ;
  assign n25190 = n25189 ^ n25085 ;
  assign n25082 = n24892 ^ n24787 ;
  assign n25083 = ~n24897 & ~n25082 ;
  assign n25084 = n25083 ^ n24892 ;
  assign n25191 = n25190 ^ n25084 ;
  assign n25192 = n25191 ^ x17 ;
  assign n25081 = n5702 & ~n20887 ;
  assign n25193 = n25192 ^ n25081 ;
  assign n25080 = n5700 & ~n20894 ;
  assign n25194 = n25193 ^ n25080 ;
  assign n25196 = n25195 ^ n25194 ;
  assign n25079 = n20731 & n20897 ;
  assign n25197 = n25196 ^ n25079 ;
  assign n25076 = n24898 ^ n24783 ;
  assign n25077 = ~n24906 & n25076 ;
  assign n25078 = n25077 ^ n24898 ;
  assign n25198 = n25197 ^ n25078 ;
  assign n25199 = n25198 ^ x14 ;
  assign n25064 = n20882 ^ x13 ;
  assign n25065 = n25064 ^ n20882 ;
  assign n25069 = ~n22671 & n25065 ;
  assign n25070 = n25069 ^ n20882 ;
  assign n25071 = n6063 & n25070 ;
  assign n25200 = n25199 ^ n25071 ;
  assign n25201 = n25200 ^ n25198 ;
  assign n25072 = ~n22671 & ~n25065 ;
  assign n25073 = n25072 ^ n20882 ;
  assign n25074 = n6060 & ~n25073 ;
  assign n25075 = n25074 ^ n16242 ;
  assign n25202 = n25201 ^ n25075 ;
  assign n25203 = n25202 ^ n25071 ;
  assign n25204 = ~n25063 & ~n25203 ;
  assign n25205 = n25204 ^ n25200 ;
  assign n25058 = n24907 ^ n24755 ;
  assign n25059 = ~n24908 & ~n25058 ;
  assign n25060 = n25059 ^ n24907 ;
  assign n25206 = n25205 ^ n25060 ;
  assign n25208 = n25206 ^ n24747 ;
  assign n25207 = n25206 ^ n24909 ;
  assign n25209 = n25208 ^ n25207 ;
  assign n25210 = n24752 & n25209 ;
  assign n25211 = n25210 ^ n25208 ;
  assign n25226 = n25225 ^ n25211 ;
  assign n25228 = n25226 ^ n24910 ;
  assign n25227 = n25226 ^ n24923 ;
  assign n25229 = n25228 ^ n25227 ;
  assign n25230 = n24915 & n25229 ;
  assign n25231 = n25230 ^ n25228 ;
  assign n25240 = n25239 ^ n25231 ;
  assign n25241 = n25240 ^ x5 ;
  assign n25057 = ~n9092 & n20837 ;
  assign n25242 = n25241 ^ n25057 ;
  assign n25056 = n9085 & n20834 ;
  assign n25243 = n25242 ^ n25056 ;
  assign n25054 = n25053 ^ n24079 ;
  assign n25055 = n25052 & n25054 ;
  assign n25244 = n25243 ^ n25055 ;
  assign n25248 = n25247 ^ n25244 ;
  assign n25049 = n24943 ^ n24924 ;
  assign n25050 = n24945 & n25049 ;
  assign n25051 = n25050 ^ n24943 ;
  assign n25249 = n25248 ^ n25051 ;
  assign n25250 = n25249 ^ n25048 ;
  assign n25261 = n25260 ^ n25250 ;
  assign n24995 = n24737 ^ n24718 ;
  assign n24996 = n24995 ^ n24738 ;
  assign n25003 = n24996 ^ n24946 ;
  assign n25004 = n24993 & n25003 ;
  assign n25005 = n25004 ^ n24992 ;
  assign n25262 = n25261 ^ n25005 ;
  assign n24997 = n24996 ^ n24719 ;
  assign n25000 = n24993 & n24997 ;
  assign n25001 = n25000 ^ n24719 ;
  assign n25002 = ~n24738 & n25001 ;
  assign n25263 = n25262 ^ n25002 ;
  assign n25514 = n25002 & ~n25262 ;
  assign n25507 = n7135 & ~n24427 ;
  assign n25505 = n7146 & n20852 ;
  assign n25503 = n8054 & n20837 ;
  assign n25495 = n5703 & n22415 ;
  assign n25488 = n4916 & n20898 ;
  assign n25471 = n25171 & ~n25179 ;
  assign n25474 = n25471 ^ n25179 ;
  assign n25475 = n25474 ^ n25171 ;
  assign n25479 = n25475 ^ n25179 ;
  assign n25480 = ~x23 & ~n25479 ;
  assign n25481 = ~n24882 & n25474 ;
  assign n25482 = ~n25182 & n25481 ;
  assign n25483 = n25480 & ~n25482 ;
  assign n25472 = x23 & ~n25471 ;
  assign n25473 = n25182 ^ n24870 ;
  assign n25476 = ~n24882 & ~n25475 ;
  assign n25477 = n25473 & n25476 ;
  assign n25478 = n25472 & ~n25477 ;
  assign n25484 = n25483 ^ n25478 ;
  assign n25468 = n4492 & ~n21744 ;
  assign n25466 = n4504 & n20910 ;
  assign n25464 = n4491 & n20902 ;
  assign n25451 = n3213 ^ n409 ;
  assign n25452 = n25451 ^ n1272 ;
  assign n25449 = n1198 ^ n141 ;
  assign n25450 = n25449 ^ n871 ;
  assign n25453 = n25452 ^ n25450 ;
  assign n25454 = n25453 ^ n3647 ;
  assign n25445 = n3884 ^ n1150 ;
  assign n25444 = n1059 ^ n91 ;
  assign n25446 = n25445 ^ n25444 ;
  assign n25442 = n14544 ^ n2465 ;
  assign n25443 = n25442 ^ n1028 ;
  assign n25447 = n25446 ^ n25443 ;
  assign n25441 = n13242 ^ n2370 ;
  assign n25448 = n25447 ^ n25441 ;
  assign n25455 = n25454 ^ n25448 ;
  assign n25456 = n25455 ^ n3682 ;
  assign n25457 = ~n2556 & ~n25456 ;
  assign n25438 = x31 & n25121 ;
  assign n25437 = ~n3733 & ~n20924 ;
  assign n25439 = n25438 ^ n25437 ;
  assign n25432 = n20970 ^ x31 ;
  assign n25433 = n25432 ^ n20970 ;
  assign n25434 = ~n21456 & n25433 ;
  assign n25435 = n25434 ^ n20970 ;
  assign n25436 = n3520 & n25435 ;
  assign n25440 = n25439 ^ n25436 ;
  assign n25458 = n25457 ^ n25440 ;
  assign n25427 = n25139 ^ n25096 ;
  assign n25428 = n25114 & n25427 ;
  assign n25429 = n25428 ^ n25139 ;
  assign n25459 = n25458 ^ n25429 ;
  assign n25425 = n831 & ~n20963 ;
  assign n25419 = n25156 ^ n25140 ;
  assign n25420 = ~n25145 & ~n25419 ;
  assign n25421 = n25420 ^ n25140 ;
  assign n25422 = n25421 ^ x29 ;
  assign n25414 = n20962 ^ n4536 ;
  assign n25415 = n25414 ^ n20962 ;
  assign n25416 = n21596 & n25415 ;
  assign n25417 = n25416 ^ n20962 ;
  assign n25418 = n650 & n25417 ;
  assign n25423 = n25422 ^ n25418 ;
  assign n25411 = n3484 & ~n20969 ;
  assign n25424 = n25423 ^ n25411 ;
  assign n25426 = n25425 ^ n25424 ;
  assign n25460 = n25459 ^ n25426 ;
  assign n25390 = n12861 & n20994 ;
  assign n25389 = n446 & ~n20922 ;
  assign n25391 = n25390 ^ n25389 ;
  assign n25392 = n25391 ^ n65 ;
  assign n25393 = n25391 ^ x26 ;
  assign n25394 = n25393 ^ n67 ;
  assign n25395 = n25394 ^ x25 ;
  assign n25396 = n25395 ^ n20913 ;
  assign n25397 = n25396 ^ n25393 ;
  assign n25398 = n25397 ^ n20999 ;
  assign n25399 = n25398 ^ n25397 ;
  assign n25400 = n25393 & ~n25399 ;
  assign n25401 = n25400 ^ n25394 ;
  assign n25402 = n25397 ^ n20913 ;
  assign n25403 = ~n25399 & ~n25402 ;
  assign n25404 = n25403 ^ n20913 ;
  assign n25405 = ~n25394 & ~n25404 ;
  assign n25406 = ~n25401 & n25405 ;
  assign n25407 = n25406 ^ n25403 ;
  assign n25408 = n25407 ^ n67 ;
  assign n25409 = n25408 ^ n20913 ;
  assign n25410 = ~n25392 & n25409 ;
  assign n25461 = n25460 ^ n25410 ;
  assign n25386 = n25170 ^ n25093 ;
  assign n25387 = ~n25158 & ~n25386 ;
  assign n25388 = n25387 ^ n25170 ;
  assign n25462 = n25461 ^ n25388 ;
  assign n25463 = n25462 ^ x23 ;
  assign n25465 = n25464 ^ n25463 ;
  assign n25467 = n25466 ^ n25465 ;
  assign n25469 = n25468 ^ n25467 ;
  assign n25385 = ~n4496 & n20903 ;
  assign n25470 = n25469 ^ n25385 ;
  assign n25485 = n25484 ^ n25470 ;
  assign n25486 = n25485 ^ x20 ;
  assign n25380 = n20897 ^ n4685 ;
  assign n25381 = n25380 ^ n20897 ;
  assign n25382 = ~n23665 & n25381 ;
  assign n25383 = n25382 ^ n20897 ;
  assign n25384 = n4678 & n25383 ;
  assign n25487 = n25486 ^ n25384 ;
  assign n25489 = n25488 ^ n25487 ;
  assign n25379 = n14027 & ~n21012 ;
  assign n25490 = n25489 ^ n25379 ;
  assign n25376 = n25185 ^ n25084 ;
  assign n25377 = ~n25190 & n25376 ;
  assign n25378 = n25377 ^ n25185 ;
  assign n25491 = n25490 ^ n25378 ;
  assign n25492 = n25491 ^ x17 ;
  assign n25375 = n5702 & ~n21025 ;
  assign n25493 = n25492 ^ n25375 ;
  assign n25374 = n5700 & ~n20887 ;
  assign n25494 = n25493 ^ n25374 ;
  assign n25496 = n25495 ^ n25494 ;
  assign n25373 = n20731 & ~n20894 ;
  assign n25497 = n25496 ^ n25373 ;
  assign n25370 = n25191 ^ n25078 ;
  assign n25371 = n25197 & ~n25370 ;
  assign n25372 = n25371 ^ n25191 ;
  assign n25498 = n25497 ^ n25372 ;
  assign n25354 = ~n6072 & n20883 ;
  assign n25353 = ~n6074 & n20882 ;
  assign n25355 = n25354 ^ n25353 ;
  assign n25356 = n25355 ^ n6060 ;
  assign n25357 = n25356 ^ x14 ;
  assign n25367 = n6063 & n23009 ;
  assign n25358 = n25355 ^ n6062 ;
  assign n25359 = n23010 ^ n20876 ;
  assign n25362 = n20876 ^ x13 ;
  assign n25363 = n25362 ^ n20876 ;
  assign n25364 = ~n25359 & ~n25363 ;
  assign n25365 = n25364 ^ n20876 ;
  assign n25366 = n25358 & n25365 ;
  assign n25368 = n25367 ^ n25366 ;
  assign n25369 = ~n25357 & ~n25368 ;
  assign n25499 = n25498 ^ n25369 ;
  assign n25350 = n25198 ^ n25060 ;
  assign n25351 = n25205 & ~n25350 ;
  assign n25352 = n25351 ^ n25198 ;
  assign n25500 = n25499 ^ n25352 ;
  assign n25340 = n6655 & ~n20872 ;
  assign n25339 = n6658 & n20861 ;
  assign n25341 = n25340 ^ n25339 ;
  assign n25342 = n25341 ^ x11 ;
  assign n25338 = n15413 & ~n23640 ;
  assign n25343 = n25342 ^ n25338 ;
  assign n25337 = n6650 & n20865 ;
  assign n25344 = n25343 ^ n25337 ;
  assign n25346 = n25344 ^ n25206 ;
  assign n25345 = n25344 ^ n25225 ;
  assign n25347 = n25346 ^ n25345 ;
  assign n25348 = n25211 & ~n25347 ;
  assign n25349 = n25348 ^ n25346 ;
  assign n25501 = n25500 ^ n25349 ;
  assign n25502 = n25501 ^ x8 ;
  assign n25504 = n25503 ^ n25502 ;
  assign n25506 = n25505 ^ n25504 ;
  assign n25508 = n25507 ^ n25506 ;
  assign n25336 = n7141 & n20836 ;
  assign n25509 = n25508 ^ n25336 ;
  assign n25333 = n25239 ^ n25226 ;
  assign n25334 = ~n25231 & ~n25333 ;
  assign n25335 = n25334 ^ n25226 ;
  assign n25510 = n25509 ^ n25335 ;
  assign n25315 = ~n9092 & n20834 ;
  assign n25314 = n9085 & n24079 ;
  assign n25316 = n25315 ^ n25314 ;
  assign n25317 = n25316 ^ n9079 ;
  assign n25318 = n25316 ^ x5 ;
  assign n25323 = n25318 ^ n19158 ;
  assign n25324 = ~x4 & ~n24463 ;
  assign n25325 = n25323 & n25324 ;
  assign n25320 = n24700 ^ n24463 ;
  assign n25321 = n19158 & n25320 ;
  assign n25319 = n24700 & n25318 ;
  assign n25322 = n25321 ^ n25319 ;
  assign n25326 = n25325 ^ n25322 ;
  assign n25327 = ~n25317 & ~n25326 ;
  assign n25328 = n25327 ^ n25240 ;
  assign n25329 = n25328 ^ n25327 ;
  assign n25330 = n25329 ^ n25051 ;
  assign n25331 = ~n25248 & ~n25330 ;
  assign n25332 = n25331 ^ n25328 ;
  assign n25511 = n25510 ^ n25332 ;
  assign n25311 = n25249 ^ n25005 ;
  assign n25312 = ~n25261 & ~n25311 ;
  assign n25313 = n25312 ^ n25249 ;
  assign n25512 = n25511 ^ n25313 ;
  assign n25289 = n25043 ^ x2 ;
  assign n25290 = n25289 ^ n25043 ;
  assign n25291 = n25043 ^ n24980 ;
  assign n25292 = n25291 ^ n25043 ;
  assign n25293 = n25290 & ~n25292 ;
  assign n25294 = n25293 ^ n25043 ;
  assign n25295 = ~x1 & n25294 ;
  assign n25296 = n25295 ^ n25289 ;
  assign n25286 = n25037 & n25041 ;
  assign n25282 = n25040 ^ n482 ;
  assign n25283 = ~n25038 & n25282 ;
  assign n25266 = ~n25026 & n25031 ;
  assign n25280 = n25023 & n25266 ;
  assign n25277 = n25041 ^ n3513 ;
  assign n25264 = n25026 ^ n25023 ;
  assign n25265 = n25264 ^ n25031 ;
  assign n25267 = n25033 ^ n24952 ;
  assign n25268 = n25267 ^ n25266 ;
  assign n25269 = n25265 & ~n25268 ;
  assign n25278 = n25277 ^ n25269 ;
  assign n25276 = n482 & n25035 ;
  assign n25279 = n25278 ^ n25276 ;
  assign n25281 = n25280 ^ n25279 ;
  assign n25284 = n25283 ^ n25281 ;
  assign n25270 = n25269 ^ n25265 ;
  assign n25271 = n25041 ^ n24952 ;
  assign n25272 = n25265 ^ n25041 ;
  assign n25273 = n25271 & ~n25272 ;
  assign n25274 = ~n25270 & n25273 ;
  assign n25285 = n25284 ^ n25274 ;
  assign n25287 = n25286 ^ n25285 ;
  assign n25288 = n25287 ^ x1 ;
  assign n25297 = n25296 ^ n25288 ;
  assign n25298 = n25297 ^ x2 ;
  assign n25299 = n25298 ^ x1 ;
  assign n25300 = n25299 ^ n25297 ;
  assign n25303 = n25006 & n25043 ;
  assign n25301 = ~n25007 & ~n25043 ;
  assign n25302 = n25301 ^ n25043 ;
  assign n25304 = n25303 ^ n25302 ;
  assign n25307 = n25300 & n25304 ;
  assign n25308 = n25307 ^ n25297 ;
  assign n25309 = x0 & ~n25308 ;
  assign n25310 = n25309 ^ n25296 ;
  assign n25513 = n25512 ^ n25310 ;
  assign n25515 = n25514 ^ n25513 ;
  assign n25692 = ~n25287 & ~n25301 ;
  assign n25693 = ~n25303 & ~n25692 ;
  assign n25711 = x0 & ~x2 ;
  assign n25712 = n25693 & n25711 ;
  assign n25695 = ~x0 & n25287 ;
  assign n25707 = n25695 ^ n10713 ;
  assign n25703 = ~n25043 & n25287 ;
  assign n25705 = n25703 ^ n25693 ;
  assign n25706 = ~x1 & n25705 ;
  assign n25708 = n25707 ^ n25706 ;
  assign n25704 = n10702 & n25703 ;
  assign n25709 = n25708 ^ n25704 ;
  assign n25694 = n25693 ^ x2 ;
  assign n25696 = n25695 ^ n25694 ;
  assign n25697 = n25696 ^ n25693 ;
  assign n25698 = n25693 ^ n25043 ;
  assign n25699 = n25698 ^ n25693 ;
  assign n25700 = n25697 & n25699 ;
  assign n25701 = n25700 ^ n25693 ;
  assign n25702 = n11240 & ~n25701 ;
  assign n25710 = n25709 ^ n25702 ;
  assign n25713 = n25712 ^ n25710 ;
  assign n25691 = ~n25513 & n25514 ;
  assign n25714 = n25713 ^ n25691 ;
  assign n25682 = n25510 ^ n25327 ;
  assign n25683 = n25332 & ~n25682 ;
  assign n25684 = n25683 ^ n25327 ;
  assign n25679 = n9085 & ~n24700 ;
  assign n25672 = n7146 & n20836 ;
  assign n25671 = n8054 & n20834 ;
  assign n25673 = n25672 ^ n25671 ;
  assign n25669 = n7141 & n20837 ;
  assign n25668 = n7135 & ~n24936 ;
  assign n25670 = n25669 ^ n25668 ;
  assign n25674 = n25673 ^ n25670 ;
  assign n25675 = n25674 ^ x8 ;
  assign n25664 = n6650 & n20861 ;
  assign n25662 = n15413 & ~n23825 ;
  assign n25659 = n6655 & n20865 ;
  assign n25658 = n6658 & n20852 ;
  assign n25660 = n25659 ^ n25658 ;
  assign n25661 = n25660 ^ x11 ;
  assign n25663 = n25662 ^ n25661 ;
  assign n25665 = n25664 ^ n25663 ;
  assign n25649 = n25498 ^ n25352 ;
  assign n25650 = n25499 & n25649 ;
  assign n25651 = n25650 ^ n25498 ;
  assign n25646 = ~n6072 & n20882 ;
  assign n25644 = ~n6074 & ~n20876 ;
  assign n25639 = n5703 & ~n22546 ;
  assign n25637 = n5700 & ~n21025 ;
  assign n25635 = n5702 & n20883 ;
  assign n25630 = n4916 & n20897 ;
  assign n25624 = n4492 & n21735 ;
  assign n25622 = n4504 & n20903 ;
  assign n25620 = n4491 & ~n21012 ;
  assign n25615 = n25410 ^ n25388 ;
  assign n25616 = ~n25461 & ~n25615 ;
  assign n25617 = n25616 ^ n25410 ;
  assign n25601 = n3699 ^ n490 ;
  assign n25602 = n25601 ^ n11888 ;
  assign n25600 = n2392 ^ n568 ;
  assign n25603 = n25602 ^ n25600 ;
  assign n25598 = n658 ^ n371 ;
  assign n25599 = n25598 ^ n837 ;
  assign n25604 = n25603 ^ n25599 ;
  assign n25595 = n4779 ^ n2856 ;
  assign n25596 = n25595 ^ n4362 ;
  assign n25597 = n25596 ^ n14857 ;
  assign n25605 = n25604 ^ n25597 ;
  assign n25606 = n25605 ^ n2658 ;
  assign n25607 = n25606 ^ n6474 ;
  assign n25608 = ~n6418 & ~n25607 ;
  assign n25585 = n21240 ^ n20970 ;
  assign n25584 = n21240 ^ n20924 ;
  assign n25586 = n25585 ^ n25584 ;
  assign n25589 = x30 & ~n25586 ;
  assign n25590 = n25589 ^ n25585 ;
  assign n25591 = ~n3520 & n25590 ;
  assign n25592 = n25591 ^ n21240 ;
  assign n25593 = x31 & n25592 ;
  assign n25581 = ~n35 & n20963 ;
  assign n25579 = ~n35 & ~n20970 ;
  assign n25580 = n25579 ^ n20963 ;
  assign n25582 = n25581 ^ n25580 ;
  assign n25583 = ~n3514 & ~n25582 ;
  assign n25594 = n25593 ^ n25583 ;
  assign n25609 = n25608 ^ n25594 ;
  assign n25576 = n25440 ^ n25429 ;
  assign n25577 = ~n25458 & n25576 ;
  assign n25578 = n25577 ^ n25440 ;
  assign n25610 = n25609 ^ n25578 ;
  assign n25573 = n25459 ^ n25421 ;
  assign n25574 = n25426 & n25573 ;
  assign n25575 = n25574 ^ n25459 ;
  assign n25611 = n25610 ^ n25575 ;
  assign n25570 = n3484 & n20962 ;
  assign n25563 = n20994 ^ x29 ;
  assign n25564 = n25563 ^ x28 ;
  assign n25565 = n25564 ^ n20994 ;
  assign n25566 = n21631 & n25565 ;
  assign n25567 = n25566 ^ n20994 ;
  assign n25568 = n650 & n25567 ;
  assign n25569 = n25568 ^ x29 ;
  assign n25571 = n25570 ^ n25569 ;
  assign n25562 = n831 & ~n20969 ;
  assign n25572 = n25571 ^ n25562 ;
  assign n25612 = n25611 ^ n25572 ;
  assign n25551 = n446 & n20913 ;
  assign n25550 = n12861 & ~n20922 ;
  assign n25552 = n25551 ^ n25550 ;
  assign n25561 = n25552 ^ x26 ;
  assign n25613 = n25612 ^ n25561 ;
  assign n25554 = n20910 ^ n467 ;
  assign n25553 = n25552 ^ n20910 ;
  assign n25555 = n25554 ^ n25553 ;
  assign n25556 = n25554 ^ n21000 ;
  assign n25557 = n25556 ^ n25554 ;
  assign n25558 = n25555 & ~n25557 ;
  assign n25559 = n25558 ^ n25554 ;
  assign n25560 = n64 & n25559 ;
  assign n25614 = n25613 ^ n25560 ;
  assign n25618 = n25617 ^ n25614 ;
  assign n25619 = n25618 ^ x23 ;
  assign n25621 = n25620 ^ n25619 ;
  assign n25623 = n25622 ^ n25621 ;
  assign n25625 = n25624 ^ n25623 ;
  assign n25549 = ~n4496 & n20902 ;
  assign n25626 = n25625 ^ n25549 ;
  assign n25546 = n25484 ^ n25462 ;
  assign n25547 = n25470 & n25546 ;
  assign n25548 = n25547 ^ n25484 ;
  assign n25627 = n25626 ^ n25548 ;
  assign n25628 = n25627 ^ x20 ;
  assign n23953 = n21954 ^ n20894 ;
  assign n25541 = n20894 ^ n4685 ;
  assign n25542 = n25541 ^ n20894 ;
  assign n25543 = ~n23953 & n25542 ;
  assign n25544 = n25543 ^ n20894 ;
  assign n25545 = n4678 & ~n25544 ;
  assign n25629 = n25628 ^ n25545 ;
  assign n25631 = n25630 ^ n25629 ;
  assign n25540 = n14027 & n20898 ;
  assign n25632 = n25631 ^ n25540 ;
  assign n25537 = n25485 ^ n25378 ;
  assign n25538 = n25490 & ~n25537 ;
  assign n25539 = n25538 ^ n25485 ;
  assign n25633 = n25632 ^ n25539 ;
  assign n25634 = n25633 ^ x17 ;
  assign n25636 = n25635 ^ n25634 ;
  assign n25638 = n25637 ^ n25636 ;
  assign n25640 = n25639 ^ n25638 ;
  assign n25536 = n20731 & ~n20887 ;
  assign n25641 = n25640 ^ n25536 ;
  assign n25533 = n25491 ^ n25372 ;
  assign n25534 = ~n25497 & ~n25533 ;
  assign n25535 = n25534 ^ n25491 ;
  assign n25642 = n25641 ^ n25535 ;
  assign n25643 = n25642 ^ x14 ;
  assign n25645 = n25644 ^ n25643 ;
  assign n25647 = n25646 ^ n25645 ;
  assign n25528 = n20872 ^ n4899 ;
  assign n25529 = n25528 ^ n20872 ;
  assign n25530 = ~n23032 & n25529 ;
  assign n25531 = n25530 ^ n20872 ;
  assign n25532 = n4897 & ~n25531 ;
  assign n25648 = n25647 ^ n25532 ;
  assign n25652 = n25651 ^ n25648 ;
  assign n25654 = n25652 ^ n25344 ;
  assign n25653 = n25652 ^ n25500 ;
  assign n25655 = n25654 ^ n25653 ;
  assign n25656 = n25349 & ~n25655 ;
  assign n25657 = n25656 ^ n25654 ;
  assign n25666 = n25665 ^ n25657 ;
  assign n25524 = n25501 ^ n25335 ;
  assign n25525 = ~n25509 & n25524 ;
  assign n25526 = n25525 ^ n25501 ;
  assign n25667 = n25666 ^ n25526 ;
  assign n25676 = n25675 ^ n25667 ;
  assign n25677 = n25676 ^ x5 ;
  assign n25517 = n24980 ^ n24949 ;
  assign n25518 = n25517 ^ n24980 ;
  assign n25519 = n24980 ^ n9089 ;
  assign n25520 = n25519 ^ n24980 ;
  assign n25521 = ~n25518 & n25520 ;
  assign n25522 = n25521 ^ n24980 ;
  assign n25523 = n9077 & ~n25522 ;
  assign n25678 = n25677 ^ n25523 ;
  assign n25680 = n25679 ^ n25678 ;
  assign n25516 = ~n9092 & n24079 ;
  assign n25681 = n25680 ^ n25516 ;
  assign n25685 = n25684 ^ n25681 ;
  assign n25686 = n25685 ^ n25313 ;
  assign n25687 = n25686 ^ n25310 ;
  assign n25688 = n25687 ^ n25685 ;
  assign n25689 = ~n25512 & ~n25688 ;
  assign n25690 = n25689 ^ n25686 ;
  assign n25715 = n25714 ^ n25690 ;
  assign n25896 = n25043 ^ n25008 ;
  assign n25897 = n9081 & ~n25896 ;
  assign n25894 = n9085 & ~n24980 ;
  assign n25892 = n10131 & n25043 ;
  assign n25886 = n7146 & n20837 ;
  assign n25885 = n8054 & n24079 ;
  assign n25887 = n25886 ^ n25885 ;
  assign n25883 = n7141 & n20834 ;
  assign n25882 = n7135 & ~n25245 ;
  assign n25884 = n25883 ^ n25882 ;
  assign n25888 = n25887 ^ n25884 ;
  assign n25875 = n25651 ^ n25642 ;
  assign n25876 = ~n25648 & n25875 ;
  assign n25877 = n25876 ^ n25642 ;
  assign n25872 = ~n6074 & ~n20872 ;
  assign n25870 = ~n6072 & ~n20876 ;
  assign n25865 = n5703 & ~n22672 ;
  assign n25858 = n4916 & ~n20894 ;
  assign n25851 = n20887 ^ x20 ;
  assign n25852 = n25851 ^ x19 ;
  assign n25853 = n25852 ^ n20887 ;
  assign n25854 = ~n22306 & n25853 ;
  assign n25855 = n25854 ^ n20887 ;
  assign n25856 = n4678 & ~n25855 ;
  assign n25857 = n25856 ^ x20 ;
  assign n25859 = n25858 ^ n25857 ;
  assign n25850 = n14027 & n20897 ;
  assign n25860 = n25859 ^ n25850 ;
  assign n25841 = n4492 & ~n21972 ;
  assign n25839 = n4504 & n20902 ;
  assign n25837 = n4491 & n20898 ;
  assign n25830 = n3484 & n20994 ;
  assign n25825 = n25575 ^ n25572 ;
  assign n25826 = ~n25611 & ~n25825 ;
  assign n25827 = n25826 ^ n25572 ;
  assign n25828 = n25827 ^ x29 ;
  assign n25820 = n20922 ^ n4536 ;
  assign n25821 = n25820 ^ n20922 ;
  assign n25822 = n21395 & n25821 ;
  assign n25823 = n25822 ^ n20922 ;
  assign n25824 = n650 & ~n25823 ;
  assign n25829 = n25828 ^ n25824 ;
  assign n25831 = n25830 ^ n25829 ;
  assign n25817 = n831 & n20962 ;
  assign n25832 = n25831 ^ n25817 ;
  assign n25809 = x31 & ~n25579 ;
  assign n25810 = n33 & n20963 ;
  assign n25811 = n25809 & ~n25810 ;
  assign n25812 = n3520 & ~n21114 ;
  assign n25813 = n25811 & ~n25812 ;
  assign n25806 = ~n35 & n20974 ;
  assign n25807 = n25806 ^ n20969 ;
  assign n25808 = ~n3514 & ~n25807 ;
  assign n25814 = n25813 ^ n25808 ;
  assign n25796 = n313 ^ n153 ;
  assign n25794 = n1069 ^ n141 ;
  assign n25795 = n25794 ^ n104 ;
  assign n25797 = n25796 ^ n25795 ;
  assign n25793 = n15090 ^ n3650 ;
  assign n25798 = n25797 ^ n25793 ;
  assign n25799 = n25798 ^ n25100 ;
  assign n25789 = n5635 ^ n577 ;
  assign n25788 = n378 ^ n118 ;
  assign n25790 = n25789 ^ n25788 ;
  assign n25787 = n11921 ^ n1890 ;
  assign n25791 = n25790 ^ n25787 ;
  assign n25783 = n1739 ^ n1135 ;
  assign n25782 = n2358 ^ n710 ;
  assign n25784 = n25783 ^ n25782 ;
  assign n25780 = n4941 ^ n304 ;
  assign n25781 = n25780 ^ n1600 ;
  assign n25785 = n25784 ^ n25781 ;
  assign n25786 = n25785 ^ n2566 ;
  assign n25792 = n25791 ^ n25786 ;
  assign n25800 = n25799 ^ n25792 ;
  assign n25801 = n25800 ^ n3634 ;
  assign n25802 = ~n4259 & ~n25801 ;
  assign n25815 = n25814 ^ n25802 ;
  assign n25777 = n25594 ^ n25578 ;
  assign n25778 = ~n25609 & n25777 ;
  assign n25779 = n25778 ^ n25594 ;
  assign n25816 = n25815 ^ n25779 ;
  assign n25833 = n25832 ^ n25816 ;
  assign n25772 = n12861 & n20913 ;
  assign n25771 = n446 & n20910 ;
  assign n25773 = n25772 ^ n25771 ;
  assign n25774 = n25773 ^ x26 ;
  assign n25770 = ~n487 & n20903 ;
  assign n25775 = n25774 ^ n25770 ;
  assign n25769 = ~n3501 & ~n21756 ;
  assign n25776 = n25775 ^ n25769 ;
  assign n25834 = n25833 ^ n25776 ;
  assign n25766 = n25617 ^ n25612 ;
  assign n25767 = ~n25614 & ~n25766 ;
  assign n25768 = n25767 ^ n25617 ;
  assign n25835 = n25834 ^ n25768 ;
  assign n25836 = n25835 ^ x23 ;
  assign n25838 = n25837 ^ n25836 ;
  assign n25840 = n25839 ^ n25838 ;
  assign n25842 = n25841 ^ n25840 ;
  assign n25765 = ~n4496 & ~n21012 ;
  assign n25843 = n25842 ^ n25765 ;
  assign n25762 = n25618 ^ n25548 ;
  assign n25763 = ~n25626 & n25762 ;
  assign n25764 = n25763 ^ n25618 ;
  assign n25844 = n25843 ^ n25764 ;
  assign n25845 = n25844 ^ n25627 ;
  assign n25846 = n25845 ^ n25844 ;
  assign n25847 = n25846 ^ n25539 ;
  assign n25848 = n25632 & n25847 ;
  assign n25849 = n25848 ^ n25845 ;
  assign n25861 = n25860 ^ n25849 ;
  assign n25862 = n25861 ^ x17 ;
  assign n25761 = n5702 & n20882 ;
  assign n25863 = n25862 ^ n25761 ;
  assign n25760 = n5700 & n20883 ;
  assign n25864 = n25863 ^ n25760 ;
  assign n25866 = n25865 ^ n25864 ;
  assign n25759 = n20731 & ~n21025 ;
  assign n25867 = n25866 ^ n25759 ;
  assign n25756 = n25633 ^ n25535 ;
  assign n25757 = n25641 & ~n25756 ;
  assign n25758 = n25757 ^ n25633 ;
  assign n25868 = n25867 ^ n25758 ;
  assign n25869 = n25868 ^ x14 ;
  assign n25871 = n25870 ^ n25869 ;
  assign n25873 = n25872 ^ n25871 ;
  assign n25750 = n20865 ^ n4899 ;
  assign n25751 = n25750 ^ n20865 ;
  assign n25753 = ~n22682 & n25751 ;
  assign n25754 = n25753 ^ n20865 ;
  assign n25755 = n4897 & n25754 ;
  assign n25874 = n25873 ^ n25755 ;
  assign n25878 = n25877 ^ n25874 ;
  assign n25747 = n25665 ^ n25652 ;
  assign n25748 = n25657 & n25747 ;
  assign n25749 = n25748 ^ n25652 ;
  assign n25879 = n25878 ^ n25749 ;
  assign n25742 = n6655 & n20861 ;
  assign n25741 = n6658 & n20836 ;
  assign n25743 = n25742 ^ n25741 ;
  assign n25744 = n25743 ^ x11 ;
  assign n25740 = n15413 & ~n24433 ;
  assign n25745 = n25744 ^ n25740 ;
  assign n25739 = n6650 & n20852 ;
  assign n25746 = n25745 ^ n25739 ;
  assign n25880 = n25879 ^ n25746 ;
  assign n25881 = n25880 ^ n25674 ;
  assign n25889 = n25888 ^ n25881 ;
  assign n25737 = n25675 ^ n25666 ;
  assign n25738 = n25667 & n25737 ;
  assign n25890 = n25889 ^ n25738 ;
  assign n25891 = n25890 ^ x5 ;
  assign n25893 = n25892 ^ n25891 ;
  assign n25895 = n25894 ^ n25893 ;
  assign n25898 = n25897 ^ n25895 ;
  assign n25736 = ~n9092 & ~n24700 ;
  assign n25899 = n25898 ^ n25736 ;
  assign n25733 = n25684 ^ n25676 ;
  assign n25734 = n25681 & n25733 ;
  assign n25735 = n25734 ^ n25684 ;
  assign n25900 = n25899 ^ n25735 ;
  assign n25720 = n25703 ^ n25695 ;
  assign n25721 = x1 & ~n25720 ;
  assign n25722 = n25721 ^ n25695 ;
  assign n25723 = n25722 ^ x2 ;
  assign n25724 = n10728 ^ n10702 ;
  assign n25725 = n25703 ^ n25692 ;
  assign n25726 = n25724 & n25725 ;
  assign n25727 = n25726 ^ n10702 ;
  assign n25728 = ~n25723 & ~n25727 ;
  assign n25729 = ~n25721 & n25728 ;
  assign n25730 = ~x2 & n25729 ;
  assign n25731 = n25730 ^ n25728 ;
  assign n25732 = n25731 ^ n25727 ;
  assign n25901 = n25900 ^ n25732 ;
  assign n25718 = ~n25685 & n25690 ;
  assign n25716 = n25691 ^ n25690 ;
  assign n25717 = n25714 & ~n25716 ;
  assign n25719 = n25718 ^ n25717 ;
  assign n25902 = n25901 ^ n25719 ;
  assign n26093 = n7135 & n25320 ;
  assign n26091 = n7146 & n20834 ;
  assign n26089 = n8054 & ~n24700 ;
  assign n26081 = n20865 ^ x14 ;
  assign n25974 = n20861 ^ x13 ;
  assign n25973 = n20861 ^ x14 ;
  assign n25975 = n25974 ^ n25973 ;
  assign n25976 = n23608 & n25975 ;
  assign n25977 = n25976 ^ n25974 ;
  assign n26082 = n26081 ^ n25977 ;
  assign n26078 = ~n23614 & n25751 ;
  assign n26079 = n26078 ^ n20865 ;
  assign n26080 = ~n6066 & n26079 ;
  assign n26083 = n26082 ^ n26080 ;
  assign n26084 = ~n4897 & n26083 ;
  assign n26073 = n5703 & n23010 ;
  assign n26071 = n5702 & ~n20876 ;
  assign n26069 = n5700 & n20882 ;
  assign n26063 = n14027 & ~n20894 ;
  assign n26062 = n4916 & ~n20887 ;
  assign n26064 = n26063 ^ n26062 ;
  assign n26060 = n4678 & n22415 ;
  assign n26059 = n4683 & ~n22414 ;
  assign n26061 = n26060 ^ n26059 ;
  assign n26065 = n26064 ^ n26061 ;
  assign n26066 = n26065 ^ x20 ;
  assign n26054 = n4492 & ~n21966 ;
  assign n26052 = n4504 & ~n21012 ;
  assign n26050 = n4491 & n20897 ;
  assign n26037 = x31 & ~n25581 ;
  assign n26038 = n33 & n20969 ;
  assign n26039 = n26037 & ~n26038 ;
  assign n26040 = n3520 & ~n21109 ;
  assign n26041 = n26039 & ~n26040 ;
  assign n26032 = n20962 ^ n35 ;
  assign n26033 = n26032 ^ n20962 ;
  assign n26034 = ~n20973 & ~n26033 ;
  assign n26035 = n26034 ^ n20962 ;
  assign n26036 = ~n3514 & n26035 ;
  assign n26042 = n26041 ^ n26036 ;
  assign n26024 = n1243 ^ n265 ;
  assign n26023 = n675 ^ n197 ;
  assign n26025 = n26024 ^ n26023 ;
  assign n26021 = n819 ^ n693 ;
  assign n26022 = n26021 ^ n238 ;
  assign n26026 = n26025 ^ n26022 ;
  assign n26018 = n5332 ^ n1543 ;
  assign n26019 = n26018 ^ n2234 ;
  assign n26020 = n26019 ^ n756 ;
  assign n26027 = n26026 ^ n26020 ;
  assign n26017 = n4033 ^ n3879 ;
  assign n26028 = n26027 ^ n26017 ;
  assign n26029 = n26028 ^ n15124 ;
  assign n26030 = ~n5089 & ~n26029 ;
  assign n26043 = n26042 ^ n26030 ;
  assign n26014 = n25814 ^ n25779 ;
  assign n26015 = ~n25815 & n26014 ;
  assign n26016 = n26015 ^ n25814 ;
  assign n26044 = n26043 ^ n26016 ;
  assign n26011 = n3484 & ~n20922 ;
  assign n26004 = n20913 ^ x29 ;
  assign n26005 = n26004 ^ x28 ;
  assign n26006 = n26005 ^ n20913 ;
  assign n26007 = ~n21088 & n26006 ;
  assign n26008 = n26007 ^ n20913 ;
  assign n26009 = n650 & n26008 ;
  assign n26010 = n26009 ^ x29 ;
  assign n26012 = n26011 ^ n26010 ;
  assign n26003 = n831 & n20994 ;
  assign n26013 = n26012 ^ n26003 ;
  assign n26045 = n26044 ^ n26013 ;
  assign n26000 = n25827 ^ n25816 ;
  assign n26001 = n25832 & ~n26000 ;
  assign n26002 = n26001 ^ n25827 ;
  assign n26046 = n26045 ^ n26002 ;
  assign n25995 = n446 & n20903 ;
  assign n25994 = n12861 & n20910 ;
  assign n25996 = n25995 ^ n25994 ;
  assign n25997 = n25996 ^ x26 ;
  assign n25993 = ~n487 & n20902 ;
  assign n25998 = n25997 ^ n25993 ;
  assign n25992 = ~n3501 & ~n21744 ;
  assign n25999 = n25998 ^ n25992 ;
  assign n26047 = n26046 ^ n25999 ;
  assign n25989 = n25776 ^ n25768 ;
  assign n25990 = ~n25834 & ~n25989 ;
  assign n25991 = n25990 ^ n25776 ;
  assign n26048 = n26047 ^ n25991 ;
  assign n26049 = n26048 ^ x23 ;
  assign n26051 = n26050 ^ n26049 ;
  assign n26053 = n26052 ^ n26051 ;
  assign n26055 = n26054 ^ n26053 ;
  assign n25988 = ~n4496 & n20898 ;
  assign n26056 = n26055 ^ n25988 ;
  assign n25985 = n25835 ^ n25764 ;
  assign n25986 = n25843 & ~n25985 ;
  assign n25987 = n25986 ^ n25835 ;
  assign n26057 = n26056 ^ n25987 ;
  assign n25982 = n25860 ^ n25844 ;
  assign n25983 = ~n25849 & ~n25982 ;
  assign n25984 = n25983 ^ n25844 ;
  assign n26058 = n26057 ^ n25984 ;
  assign n26067 = n26066 ^ n26058 ;
  assign n26068 = n26067 ^ x17 ;
  assign n26070 = n26069 ^ n26068 ;
  assign n26072 = n26071 ^ n26070 ;
  assign n26074 = n26073 ^ n26072 ;
  assign n25981 = n20731 & n20883 ;
  assign n26075 = n26074 ^ n25981 ;
  assign n25978 = n25861 ^ n25758 ;
  assign n25979 = ~n25867 & ~n25978 ;
  assign n25980 = n25979 ^ n25861 ;
  assign n26076 = n26075 ^ n25980 ;
  assign n26077 = n26076 ^ n25977 ;
  assign n26085 = n26084 ^ n26077 ;
  assign n25970 = n25877 ^ n25868 ;
  assign n25971 = ~n25874 & n25970 ;
  assign n25972 = n25971 ^ n25868 ;
  assign n26086 = n26085 ^ n25972 ;
  assign n25962 = n6650 & n20836 ;
  assign n25955 = n20837 ^ x11 ;
  assign n25956 = n25955 ^ x10 ;
  assign n25957 = n25956 ^ n20837 ;
  assign n25958 = ~n21061 & n25957 ;
  assign n25959 = n25958 ^ n20837 ;
  assign n25960 = n6648 & n25959 ;
  assign n25961 = n25960 ^ x11 ;
  assign n25963 = n25962 ^ n25961 ;
  assign n25953 = n6655 & n20852 ;
  assign n25964 = n25963 ^ n25953 ;
  assign n25965 = n25964 ^ n25749 ;
  assign n25966 = n25965 ^ n25746 ;
  assign n25967 = n25966 ^ n25964 ;
  assign n25968 = n25879 & n25967 ;
  assign n25969 = n25968 ^ n25965 ;
  assign n26087 = n26086 ^ n25969 ;
  assign n26088 = n26087 ^ x8 ;
  assign n26090 = n26089 ^ n26088 ;
  assign n26092 = n26091 ^ n26090 ;
  assign n26094 = n26093 ^ n26092 ;
  assign n25952 = n7141 & n24079 ;
  assign n26095 = n26094 ^ n25952 ;
  assign n25941 = n25675 & ~n25889 ;
  assign n25942 = ~n25526 & n25666 ;
  assign n25943 = n25942 ^ n25667 ;
  assign n25944 = n25942 ^ n25880 ;
  assign n25945 = n25888 ^ x8 ;
  assign n25946 = n25945 ^ n25942 ;
  assign n25947 = n25944 & ~n25946 ;
  assign n25948 = n25947 ^ n25880 ;
  assign n25949 = ~n25943 & ~n25948 ;
  assign n25950 = n25941 & n25949 ;
  assign n25951 = n25950 ^ n25948 ;
  assign n26096 = n26095 ^ n25951 ;
  assign n25937 = n25304 ^ n25287 ;
  assign n25938 = n9081 & n25937 ;
  assign n25935 = ~n9092 & ~n24980 ;
  assign n25933 = n9085 & n25043 ;
  assign n25934 = n25933 ^ x5 ;
  assign n25936 = n25935 ^ n25934 ;
  assign n25939 = n25938 ^ n25936 ;
  assign n25932 = n10131 & ~n25287 ;
  assign n25940 = n25939 ^ n25932 ;
  assign n26097 = n26096 ^ n25940 ;
  assign n25929 = n25890 ^ n25735 ;
  assign n25930 = n25899 & ~n25929 ;
  assign n25931 = n25930 ^ n25890 ;
  assign n26098 = n26097 ^ n25931 ;
  assign n25925 = x2 & n11240 ;
  assign n25926 = n25703 & n25925 ;
  assign n25927 = n25926 ^ x2 ;
  assign n25903 = n25690 & n25713 ;
  assign n25920 = n25903 ^ n25713 ;
  assign n25908 = n25685 & n25690 ;
  assign n25909 = n25908 ^ n25690 ;
  assign n25921 = n25920 ^ n25909 ;
  assign n25922 = n25921 ^ n25732 ;
  assign n25923 = ~n25901 & n25922 ;
  assign n25924 = n25923 ^ n25900 ;
  assign n25928 = n25927 ^ n25924 ;
  assign n26099 = n26098 ^ n25928 ;
  assign n25904 = n25691 & ~n25903 ;
  assign n25915 = n25908 ^ n25901 ;
  assign n25905 = n25901 ^ n25690 ;
  assign n25906 = n25905 ^ n25713 ;
  assign n25907 = n25901 ^ n25685 ;
  assign n25910 = n25909 ^ n25901 ;
  assign n25911 = n25910 ^ n25901 ;
  assign n25912 = ~n25907 & n25911 ;
  assign n25913 = n25912 ^ n25901 ;
  assign n25914 = ~n25906 & ~n25913 ;
  assign n25916 = n25915 ^ n25914 ;
  assign n25917 = n25916 ^ n25713 ;
  assign n25918 = n25917 ^ n25713 ;
  assign n25919 = n25904 & ~n25918 ;
  assign n26100 = n26099 ^ n25919 ;
  assign n26101 = ~n25924 & n25927 ;
  assign n26102 = n26098 & ~n26101 ;
  assign n26103 = n26102 ^ n25928 ;
  assign n26282 = n7141 & ~n24700 ;
  assign n26280 = n7135 & n25517 ;
  assign n26277 = n7146 & n24079 ;
  assign n26276 = n8054 & ~n24980 ;
  assign n26278 = n26277 ^ n26276 ;
  assign n26279 = n26278 ^ x8 ;
  assign n26281 = n26280 ^ n26279 ;
  assign n26283 = n26282 ^ n26281 ;
  assign n26267 = n26086 ^ n25964 ;
  assign n26268 = n25969 & n26267 ;
  assign n26269 = n26268 ^ n25964 ;
  assign n26264 = n15413 & ~n24936 ;
  assign n26254 = n5703 & n23033 ;
  assign n26252 = n5700 & ~n20876 ;
  assign n26250 = n5702 & ~n20872 ;
  assign n26244 = ~n4496 & n20897 ;
  assign n26241 = n4490 & ~n21953 ;
  assign n26240 = n14007 & n21954 ;
  assign n26242 = n26241 ^ n26240 ;
  assign n26217 = ~n35 & n20962 ;
  assign n26215 = ~n3520 & ~n20994 ;
  assign n26214 = n20994 ^ n3520 ;
  assign n26216 = n26215 ^ n26214 ;
  assign n26218 = n26217 ^ n26216 ;
  assign n26228 = n26218 ^ n21630 ;
  assign n26221 = n21630 ^ n20962 ;
  assign n26220 = n21630 ^ n20969 ;
  assign n26222 = n26221 ^ n26220 ;
  assign n26225 = x30 & ~n26222 ;
  assign n26226 = n26225 ^ n26221 ;
  assign n26227 = ~n3520 & n26226 ;
  assign n26229 = n26228 ^ n26227 ;
  assign n26230 = x31 & ~n26229 ;
  assign n26207 = n24830 ^ n4142 ;
  assign n26205 = n1414 ^ n178 ;
  assign n26204 = n1553 ^ n255 ;
  assign n26206 = n26205 ^ n26204 ;
  assign n26208 = n26207 ^ n26206 ;
  assign n26201 = n5107 ^ n360 ;
  assign n26202 = n26201 ^ n490 ;
  assign n26199 = n3251 ^ n1366 ;
  assign n26200 = n26199 ^ n2161 ;
  assign n26203 = n26202 ^ n26200 ;
  assign n26209 = n26208 ^ n26203 ;
  assign n26195 = n2045 ^ n982 ;
  assign n26194 = n14531 ^ n2583 ;
  assign n26196 = n26195 ^ n26194 ;
  assign n26197 = n26196 ^ n13882 ;
  assign n26198 = n26197 ^ n25599 ;
  assign n26210 = n26209 ^ n26198 ;
  assign n26211 = n14328 ^ n5125 ;
  assign n26212 = n26211 ^ n3148 ;
  assign n26213 = ~n26210 & ~n26212 ;
  assign n26219 = n26218 ^ n26213 ;
  assign n26231 = n26230 ^ n26219 ;
  assign n26191 = n26042 ^ n26016 ;
  assign n26192 = ~n26043 & n26191 ;
  assign n26193 = n26192 ^ n26042 ;
  assign n26232 = n26231 ^ n26193 ;
  assign n26188 = n831 & ~n20922 ;
  assign n26181 = n20910 ^ x29 ;
  assign n26182 = n26181 ^ x28 ;
  assign n26183 = n26182 ^ n20910 ;
  assign n26184 = n22951 & n26183 ;
  assign n26185 = n26184 ^ n20910 ;
  assign n26186 = n650 & n26185 ;
  assign n26187 = n26186 ^ x29 ;
  assign n26189 = n26188 ^ n26187 ;
  assign n26180 = n3484 & n20913 ;
  assign n26190 = n26189 ^ n26180 ;
  assign n26233 = n26232 ^ n26190 ;
  assign n26177 = n26013 ^ n26002 ;
  assign n26178 = ~n26045 & n26177 ;
  assign n26179 = n26178 ^ n26013 ;
  assign n26234 = n26233 ^ n26179 ;
  assign n26172 = n12861 & n20903 ;
  assign n26171 = n446 & n20902 ;
  assign n26173 = n26172 ^ n26171 ;
  assign n26174 = n26173 ^ x26 ;
  assign n26170 = ~n487 & ~n21012 ;
  assign n26175 = n26174 ^ n26170 ;
  assign n26169 = ~n3501 & n21735 ;
  assign n26176 = n26175 ^ n26169 ;
  assign n26235 = n26234 ^ n26176 ;
  assign n26166 = n25999 ^ n25991 ;
  assign n26167 = ~n26047 & n26166 ;
  assign n26168 = n26167 ^ n25999 ;
  assign n26236 = n26235 ^ n26168 ;
  assign n26237 = n26236 ^ x23 ;
  assign n26165 = n4504 & n20898 ;
  assign n26238 = n26237 ^ n26165 ;
  assign n26164 = n14008 & ~n20894 ;
  assign n26239 = n26238 ^ n26164 ;
  assign n26243 = n26242 ^ n26239 ;
  assign n26245 = n26244 ^ n26243 ;
  assign n26161 = n26048 ^ n25987 ;
  assign n26162 = ~n26056 & ~n26161 ;
  assign n26163 = n26162 ^ n26048 ;
  assign n26246 = n26245 ^ n26163 ;
  assign n26158 = n4916 & ~n21025 ;
  assign n26156 = n4683 & n20883 ;
  assign n26154 = n14027 & ~n20887 ;
  assign n26153 = n4684 & ~n22546 ;
  assign n26155 = n26154 ^ n26153 ;
  assign n26157 = n26156 ^ n26155 ;
  assign n26159 = n26158 ^ n26157 ;
  assign n26160 = n26159 ^ n26065 ;
  assign n26247 = n26246 ^ n26160 ;
  assign n26151 = n26066 ^ n26057 ;
  assign n26152 = ~n26058 & ~n26151 ;
  assign n26248 = n26247 ^ n26152 ;
  assign n26249 = n26248 ^ x17 ;
  assign n26251 = n26250 ^ n26249 ;
  assign n26253 = n26252 ^ n26251 ;
  assign n26255 = n26254 ^ n26253 ;
  assign n26150 = n20731 & n20882 ;
  assign n26256 = n26255 ^ n26150 ;
  assign n26147 = n26067 ^ n25980 ;
  assign n26148 = n26075 & ~n26147 ;
  assign n26149 = n26148 ^ n26067 ;
  assign n26257 = n26256 ^ n26149 ;
  assign n26126 = n20861 ^ n4899 ;
  assign n26127 = n26126 ^ n20861 ;
  assign n26128 = n20865 & n26127 ;
  assign n26129 = n26128 ^ n20861 ;
  assign n26130 = n4899 ^ x12 ;
  assign n26131 = n26130 ^ n20861 ;
  assign n26132 = n26131 ^ x13 ;
  assign n26133 = n26132 ^ n4899 ;
  assign n26134 = n26133 ^ n20861 ;
  assign n26135 = ~n26129 & ~n26134 ;
  assign n26136 = n26135 ^ n26131 ;
  assign n26258 = n26257 ^ n26136 ;
  assign n26137 = n20852 ^ x13 ;
  assign n26138 = n26137 ^ n26136 ;
  assign n26139 = n26138 ^ x13 ;
  assign n26140 = n26139 ^ x14 ;
  assign n26141 = n26140 ^ n26138 ;
  assign n26142 = n26138 ^ n23059 ;
  assign n26143 = n26142 ^ n26138 ;
  assign n26144 = n26141 & n26143 ;
  assign n26145 = n26144 ^ n26138 ;
  assign n26146 = n4897 & ~n26145 ;
  assign n26259 = n26258 ^ n26146 ;
  assign n26123 = n26076 ^ n25972 ;
  assign n26124 = ~n26085 & n26123 ;
  assign n26125 = n26124 ^ n26076 ;
  assign n26260 = n26259 ^ n26125 ;
  assign n26261 = n26260 ^ x11 ;
  assign n26122 = n6658 & n20834 ;
  assign n26262 = n26261 ^ n26122 ;
  assign n26121 = n6655 & n20836 ;
  assign n26263 = n26262 ^ n26121 ;
  assign n26265 = n26264 ^ n26263 ;
  assign n26120 = n6650 & n20837 ;
  assign n26266 = n26265 ^ n26120 ;
  assign n26270 = n26269 ^ n26266 ;
  assign n26271 = n26270 ^ n26087 ;
  assign n26272 = n26271 ^ n25951 ;
  assign n26273 = n26272 ^ n26270 ;
  assign n26274 = n26095 & n26273 ;
  assign n26275 = n26274 ^ n26271 ;
  assign n26284 = n26283 ^ n26275 ;
  assign n26115 = ~n9092 & n25043 ;
  assign n26114 = n9081 & n25693 ;
  assign n26116 = n26115 ^ n26114 ;
  assign n26117 = n26116 ^ n9085 ;
  assign n26111 = n10131 & ~n25043 ;
  assign n26112 = n26111 ^ n9085 ;
  assign n26113 = n25287 & n26112 ;
  assign n26118 = n26117 ^ n26113 ;
  assign n26119 = n26118 ^ n5328 ;
  assign n26285 = n26284 ^ n26119 ;
  assign n26104 = n25940 ^ n25931 ;
  assign n26105 = n26097 & ~n26104 ;
  assign n26106 = n26105 ^ n26096 ;
  assign n26286 = n26285 ^ n26106 ;
  assign n26287 = n26286 ^ n25919 ;
  assign n26288 = n26287 ^ n26101 ;
  assign n26289 = n26288 ^ n26102 ;
  assign n26290 = n26289 ^ n26286 ;
  assign n26291 = n26103 & n26290 ;
  assign n26292 = n26291 ^ n26287 ;
  assign n26504 = n26098 ^ n25927 ;
  assign n26505 = n26504 ^ n25924 ;
  assign n26506 = n26286 ^ n26101 ;
  assign n26507 = ~n26505 & ~n26506 ;
  assign n26508 = n25919 & n26507 ;
  assign n26488 = n26285 ^ n26101 ;
  assign n26489 = n26106 ^ n26101 ;
  assign n26490 = ~n26488 & ~n26489 ;
  assign n26501 = n26490 ^ n26285 ;
  assign n26491 = n26488 ^ n25928 ;
  assign n26492 = n26491 ^ n26490 ;
  assign n26493 = n26285 ^ n25931 ;
  assign n26494 = n26493 ^ n26285 ;
  assign n26495 = n26285 ^ n26096 ;
  assign n26496 = n26495 ^ n26285 ;
  assign n26497 = n26494 & n26496 ;
  assign n26498 = n26497 ^ n26285 ;
  assign n26499 = n26102 & ~n26498 ;
  assign n26500 = n26492 & n26499 ;
  assign n26502 = n26501 ^ n26500 ;
  assign n26476 = n9092 ^ x5 ;
  assign n26473 = n9091 ^ n9077 ;
  assign n26474 = n26473 ^ n25933 ;
  assign n26475 = n25287 & ~n26474 ;
  assign n26477 = n26476 ^ n26475 ;
  assign n26472 = n9081 & n25725 ;
  assign n26478 = n26477 ^ n26472 ;
  assign n26479 = n26283 ^ n26270 ;
  assign n26480 = ~n26275 & ~n26479 ;
  assign n26481 = n26480 ^ n26270 ;
  assign n26483 = ~n26478 & ~n26481 ;
  assign n26452 = n4916 & n20883 ;
  assign n26443 = n3484 & n20910 ;
  assign n26436 = n20903 ^ x29 ;
  assign n26437 = n26436 ^ x28 ;
  assign n26438 = n26437 ^ n20903 ;
  assign n26439 = ~n21755 & n26438 ;
  assign n26440 = n26439 ^ n20903 ;
  assign n26441 = n650 & n26440 ;
  assign n26442 = n26441 ^ x29 ;
  assign n26444 = n26443 ^ n26442 ;
  assign n26435 = n831 & n20913 ;
  assign n26445 = n26444 ^ n26435 ;
  assign n26421 = n6422 ^ n5071 ;
  assign n26422 = n26421 ^ n13780 ;
  assign n26423 = n26422 ^ n12472 ;
  assign n26424 = n26423 ^ n2457 ;
  assign n26415 = n797 ^ n678 ;
  assign n26413 = n418 ^ n400 ;
  assign n26414 = n26413 ^ n1074 ;
  assign n26416 = n26415 ^ n26414 ;
  assign n26411 = n13014 ^ n794 ;
  assign n26412 = n26411 ^ n4793 ;
  assign n26417 = n26416 ^ n26412 ;
  assign n26418 = n13130 ^ n2864 ;
  assign n26419 = n26418 ^ n349 ;
  assign n26420 = ~n26417 & n26419 ;
  assign n26425 = n26424 ^ n26420 ;
  assign n26426 = ~n2855 & n26425 ;
  assign n26427 = ~n596 & n26426 ;
  assign n26428 = n26427 ^ x2 ;
  assign n26408 = n12533 & ~n26215 ;
  assign n26406 = ~n35 & n20994 ;
  assign n26403 = x31 & n21395 ;
  assign n26404 = n26403 ^ n20922 ;
  assign n26405 = n3520 & n26404 ;
  assign n26407 = n26406 ^ n26405 ;
  assign n26409 = n26408 ^ n26407 ;
  assign n26400 = x31 & n26217 ;
  assign n26410 = n26409 ^ n26400 ;
  assign n26429 = n26428 ^ n26410 ;
  assign n26430 = n26429 ^ n26213 ;
  assign n26431 = n26430 ^ n26429 ;
  assign n26432 = n26431 ^ n26193 ;
  assign n26433 = n26231 & ~n26432 ;
  assign n26434 = n26433 ^ n26430 ;
  assign n26446 = n26445 ^ n26434 ;
  assign n26397 = n26190 ^ n26179 ;
  assign n26398 = n26233 & n26397 ;
  assign n26399 = n26398 ^ n26190 ;
  assign n26447 = n26446 ^ n26399 ;
  assign n26392 = n12861 & n20902 ;
  assign n26391 = n446 & ~n21012 ;
  assign n26393 = n26392 ^ n26391 ;
  assign n26394 = n26393 ^ x26 ;
  assign n26390 = ~n487 & n20898 ;
  assign n26395 = n26394 ^ n26390 ;
  assign n26389 = ~n3501 & ~n21972 ;
  assign n26396 = n26395 ^ n26389 ;
  assign n26448 = n26447 ^ n26396 ;
  assign n26379 = x23 & n22306 ;
  assign n26378 = n4490 & n22307 ;
  assign n26380 = n26379 ^ n26378 ;
  assign n26376 = n4504 & n20897 ;
  assign n26374 = n4490 ^ n4488 ;
  assign n26375 = ~n20887 & n26374 ;
  assign n26377 = n26376 ^ n26375 ;
  assign n26381 = n26380 ^ n26377 ;
  assign n26373 = ~n4496 & ~n20894 ;
  assign n26382 = n26381 ^ n26373 ;
  assign n26372 = n14005 & ~n22306 ;
  assign n26383 = n26382 ^ n26372 ;
  assign n26384 = n26383 ^ n26176 ;
  assign n26385 = n26384 ^ n26383 ;
  assign n26386 = n26385 ^ n26168 ;
  assign n26387 = n26235 & n26386 ;
  assign n26388 = n26387 ^ n26384 ;
  assign n26449 = n26448 ^ n26388 ;
  assign n26450 = n26449 ^ x20 ;
  assign n26367 = n20882 ^ n4685 ;
  assign n26368 = n26367 ^ n20882 ;
  assign n26369 = ~n22671 & n26368 ;
  assign n26370 = n26369 ^ n20882 ;
  assign n26371 = n4678 & n26370 ;
  assign n26451 = n26450 ^ n26371 ;
  assign n26453 = n26452 ^ n26451 ;
  assign n26366 = n14027 & ~n21025 ;
  assign n26454 = n26453 ^ n26366 ;
  assign n26363 = n26236 ^ n26163 ;
  assign n26364 = n26245 & ~n26363 ;
  assign n26365 = n26364 ^ n26236 ;
  assign n26455 = n26454 ^ n26365 ;
  assign n26352 = n26066 & n26247 ;
  assign n26353 = ~n25984 & ~n26057 ;
  assign n26354 = n26353 ^ n26058 ;
  assign n26355 = n26353 ^ n26246 ;
  assign n26356 = n26159 ^ x20 ;
  assign n26357 = n26356 ^ n26353 ;
  assign n26358 = ~n26355 & ~n26357 ;
  assign n26359 = n26358 ^ n26246 ;
  assign n26360 = n26354 & n26359 ;
  assign n26361 = n26352 & n26360 ;
  assign n26362 = n26361 ^ n26359 ;
  assign n26456 = n26455 ^ n26362 ;
  assign n26350 = n20731 & ~n20876 ;
  assign n26348 = n5703 & ~n22683 ;
  assign n26345 = n5700 & ~n20872 ;
  assign n26344 = n5702 & n20865 ;
  assign n26346 = n26345 ^ n26344 ;
  assign n26347 = n26346 ^ x17 ;
  assign n26349 = n26348 ^ n26347 ;
  assign n26351 = n26350 ^ n26349 ;
  assign n26457 = n26456 ^ n26351 ;
  assign n26319 = ~n6074 & n20852 ;
  assign n26318 = ~n6072 & n20861 ;
  assign n26320 = n26319 ^ n26318 ;
  assign n26321 = n26320 ^ n6060 ;
  assign n26322 = n26321 ^ x14 ;
  assign n26340 = n20836 ^ n6063 ;
  assign n26326 = n26320 ^ n6062 ;
  assign n26327 = n24433 ^ n20836 ;
  assign n26328 = n26327 ^ n20836 ;
  assign n26329 = n26328 ^ n20836 ;
  assign n26330 = n20836 ^ n17542 ;
  assign n26331 = n26330 ^ n20836 ;
  assign n26332 = ~n26329 & ~n26331 ;
  assign n26333 = n26332 ^ n20836 ;
  assign n26334 = ~n26326 & ~n26333 ;
  assign n26341 = n26340 ^ n26334 ;
  assign n26339 = ~n17542 & ~n23041 ;
  assign n26342 = n26341 ^ n26339 ;
  assign n26343 = ~n26322 & n26342 ;
  assign n26458 = n26457 ^ n26343 ;
  assign n26315 = n26248 ^ n26149 ;
  assign n26316 = ~n26256 & ~n26315 ;
  assign n26317 = n26316 ^ n26248 ;
  assign n26459 = n26458 ^ n26317 ;
  assign n26310 = n6655 & n20837 ;
  assign n26309 = n6658 & n24079 ;
  assign n26311 = n26310 ^ n26309 ;
  assign n26312 = n26311 ^ x11 ;
  assign n26308 = n15413 & ~n25245 ;
  assign n26313 = n26312 ^ n26308 ;
  assign n26307 = n6650 & n20834 ;
  assign n26314 = n26313 ^ n26307 ;
  assign n26460 = n26459 ^ n26314 ;
  assign n26304 = n26257 ^ n26125 ;
  assign n26305 = n26259 & n26304 ;
  assign n26306 = n26305 ^ n26257 ;
  assign n26461 = n26460 ^ n26306 ;
  assign n26301 = n26269 ^ n26260 ;
  assign n26302 = n26266 & ~n26301 ;
  assign n26303 = n26302 ^ n26269 ;
  assign n26462 = n26461 ^ n26303 ;
  assign n26299 = n7141 & ~n24980 ;
  assign n26297 = n7135 & ~n25896 ;
  assign n26294 = n7146 & ~n24700 ;
  assign n26293 = n8054 & n25043 ;
  assign n26295 = n26294 ^ n26293 ;
  assign n26296 = n26295 ^ x8 ;
  assign n26298 = n26297 ^ n26296 ;
  assign n26300 = n26299 ^ n26298 ;
  assign n26463 = n26462 ^ n26300 ;
  assign n26464 = n26284 ^ x2 ;
  assign n26465 = n26284 ^ x5 ;
  assign n26466 = n26465 ^ n26118 ;
  assign n26467 = ~n26464 & n26466 ;
  assign n26468 = n26467 ^ x2 ;
  assign n26470 = ~n26463 & ~n26468 ;
  assign n26486 = n26483 ^ n26470 ;
  assign n26482 = n26481 ^ n26478 ;
  assign n26484 = n26483 ^ n26482 ;
  assign n26469 = n26468 ^ n26463 ;
  assign n26471 = n26470 ^ n26469 ;
  assign n26485 = n26484 ^ n26471 ;
  assign n26487 = n26486 ^ n26485 ;
  assign n26503 = n26502 ^ n26487 ;
  assign n26509 = n26508 ^ n26503 ;
  assign n26705 = ~n26503 & n26508 ;
  assign n26702 = n26502 ^ n26482 ;
  assign n26703 = n26487 & n26702 ;
  assign n26696 = n6650 & n24079 ;
  assign n26694 = n15413 & n25320 ;
  assign n26691 = n6655 & n20834 ;
  assign n26690 = n6658 & ~n24700 ;
  assign n26692 = n26691 ^ n26690 ;
  assign n26693 = n26692 ^ x11 ;
  assign n26695 = n26694 ^ n26693 ;
  assign n26697 = n26696 ^ n26695 ;
  assign n26678 = n26449 ^ n26365 ;
  assign n26679 = n26454 & n26678 ;
  assign n26680 = n26679 ^ n26449 ;
  assign n26672 = n14027 & n20883 ;
  assign n26671 = n4684 & n23010 ;
  assign n26673 = n26672 ^ n26671 ;
  assign n26674 = n26673 ^ x20 ;
  assign n26670 = n4683 & ~n20876 ;
  assign n26675 = n26674 ^ n26670 ;
  assign n26669 = n4916 & n20882 ;
  assign n26676 = n26675 ^ n26669 ;
  assign n26659 = n26399 ^ n26396 ;
  assign n26660 = ~n26447 & n26659 ;
  assign n26661 = n26660 ^ n26396 ;
  assign n26637 = n12861 & ~n21012 ;
  assign n26636 = n446 & n20898 ;
  assign n26638 = n26637 ^ n26636 ;
  assign n26639 = n26638 ^ n65 ;
  assign n26640 = n26638 ^ x26 ;
  assign n26641 = n26640 ^ n67 ;
  assign n26642 = n26641 ^ x25 ;
  assign n26643 = n26642 ^ n20897 ;
  assign n26644 = n26643 ^ n26640 ;
  assign n26645 = n26644 ^ n21965 ;
  assign n26646 = n26645 ^ n26644 ;
  assign n26647 = n26640 & ~n26646 ;
  assign n26648 = n26647 ^ n26641 ;
  assign n26649 = n26644 ^ n20897 ;
  assign n26650 = ~n26646 & ~n26649 ;
  assign n26651 = n26650 ^ n20897 ;
  assign n26652 = ~n26641 & ~n26651 ;
  assign n26653 = ~n26648 & n26652 ;
  assign n26654 = n26653 ^ n26650 ;
  assign n26655 = n26654 ^ n67 ;
  assign n26656 = n26655 ^ n20897 ;
  assign n26657 = ~n26639 & n26656 ;
  assign n26633 = n831 & n20910 ;
  assign n26608 = n12815 ^ n782 ;
  assign n26609 = n26608 ^ n266 ;
  assign n26607 = n4777 ^ n589 ;
  assign n26610 = n26609 ^ n26607 ;
  assign n26611 = n26610 ^ n1946 ;
  assign n26620 = n4242 ^ n272 ;
  assign n26621 = n26620 ^ n260 ;
  assign n26619 = n1208 ^ n697 ;
  assign n26622 = n26621 ^ n26619 ;
  assign n26623 = n26622 ^ n2398 ;
  assign n26616 = n1396 ^ n1149 ;
  assign n26615 = n1742 ^ n1113 ;
  assign n26617 = n26616 ^ n26615 ;
  assign n26613 = n3987 ^ n1549 ;
  assign n26612 = n3673 ^ n2856 ;
  assign n26614 = n26613 ^ n26612 ;
  assign n26618 = n26617 ^ n26614 ;
  assign n26624 = n26623 ^ n26618 ;
  assign n26625 = n26624 ^ n3190 ;
  assign n26626 = ~n15201 & ~n26625 ;
  assign n26627 = ~n26611 & n26626 ;
  assign n26604 = n26427 ^ n26410 ;
  assign n26605 = ~n26428 & n26604 ;
  assign n26606 = n26605 ^ x2 ;
  assign n26628 = n26627 ^ n26606 ;
  assign n26629 = n26628 ^ x2 ;
  assign n26595 = n21087 ^ n20922 ;
  assign n26596 = ~n23912 & n26595 ;
  assign n26593 = ~n35 & ~n20922 ;
  assign n26591 = n21087 ^ n3726 ;
  assign n26592 = n26591 ^ n26406 ;
  assign n26594 = n26593 ^ n26592 ;
  assign n26597 = n26596 ^ n26594 ;
  assign n26583 = n26406 ^ n20922 ;
  assign n26584 = n26583 ^ n3726 ;
  assign n26585 = n26584 ^ n26583 ;
  assign n26586 = n26583 ^ n20913 ;
  assign n26587 = n26586 ^ n26583 ;
  assign n26588 = n26585 & ~n26587 ;
  assign n26589 = n26588 ^ n26583 ;
  assign n26590 = ~x31 & ~n26589 ;
  assign n26598 = n26597 ^ n26590 ;
  assign n26600 = n26598 ^ n26429 ;
  assign n26599 = n26598 ^ n26445 ;
  assign n26601 = n26600 ^ n26599 ;
  assign n26602 = n26434 & ~n26601 ;
  assign n26603 = n26602 ^ n26600 ;
  assign n26630 = n26629 ^ n26603 ;
  assign n26631 = n26630 ^ x29 ;
  assign n26577 = n21744 ^ n20902 ;
  assign n26578 = n20902 ^ n4536 ;
  assign n26579 = n26578 ^ n20902 ;
  assign n26580 = ~n26577 & n26579 ;
  assign n26581 = n26580 ^ n20902 ;
  assign n26582 = n650 & n26581 ;
  assign n26632 = n26631 ^ n26582 ;
  assign n26634 = n26633 ^ n26632 ;
  assign n26575 = n3484 & n20903 ;
  assign n26635 = n26634 ^ n26575 ;
  assign n26658 = n26657 ^ n26635 ;
  assign n26662 = n26661 ^ n26658 ;
  assign n26570 = n4504 & ~n20894 ;
  assign n26569 = n4491 & ~n21025 ;
  assign n26571 = n26570 ^ n26569 ;
  assign n26572 = n26571 ^ x23 ;
  assign n26568 = n4492 & n22415 ;
  assign n26573 = n26572 ^ n26568 ;
  assign n26567 = ~n4496 & ~n20887 ;
  assign n26574 = n26573 ^ n26567 ;
  assign n26663 = n26662 ^ n26574 ;
  assign n26665 = n26663 ^ n26383 ;
  assign n26664 = n26663 ^ n26448 ;
  assign n26666 = n26665 ^ n26664 ;
  assign n26667 = n26388 & n26666 ;
  assign n26668 = n26667 ^ n26665 ;
  assign n26677 = n26676 ^ n26668 ;
  assign n26681 = n26680 ^ n26677 ;
  assign n26562 = n5700 & n20865 ;
  assign n26561 = n5702 & n20861 ;
  assign n26563 = n26562 ^ n26561 ;
  assign n26564 = n26563 ^ x17 ;
  assign n26560 = n5703 & ~n23640 ;
  assign n26565 = n26564 ^ n26560 ;
  assign n26559 = n20731 & ~n20872 ;
  assign n26566 = n26565 ^ n26559 ;
  assign n26682 = n26681 ^ n26566 ;
  assign n26556 = n26362 ^ n26351 ;
  assign n26557 = ~n26456 & ~n26556 ;
  assign n26558 = n26557 ^ n26362 ;
  assign n26683 = n26682 ^ n26558 ;
  assign n26539 = ~x13 & ~n21061 ;
  assign n26538 = ~x14 & n21061 ;
  assign n26540 = n26539 ^ n26538 ;
  assign n26541 = n6062 & n20837 ;
  assign n26543 = ~n6072 & n20852 ;
  assign n26542 = ~n6074 & n20836 ;
  assign n26544 = n26543 ^ n26542 ;
  assign n26545 = x14 & n26544 ;
  assign n26546 = n26541 & ~n26545 ;
  assign n26547 = n26540 & n26546 ;
  assign n26548 = n26544 ^ n6060 ;
  assign n26549 = n26548 ^ x14 ;
  assign n26550 = n26541 ^ n6062 ;
  assign n26551 = n26545 ^ n26538 ;
  assign n26552 = ~n26539 & ~n26551 ;
  assign n26553 = n26550 & n26552 ;
  assign n26554 = ~n26549 & ~n26553 ;
  assign n26555 = ~n26547 & n26554 ;
  assign n26684 = n26683 ^ n26555 ;
  assign n26685 = n26684 ^ n26343 ;
  assign n26686 = n26685 ^ n26317 ;
  assign n26687 = n26686 ^ n26684 ;
  assign n26688 = n26458 & n26687 ;
  assign n26689 = n26688 ^ n26685 ;
  assign n26698 = n26697 ^ n26689 ;
  assign n26518 = n7146 & ~n24980 ;
  assign n26517 = n7141 & n25043 ;
  assign n26519 = n26518 ^ n26517 ;
  assign n26520 = n26519 ^ n7129 ;
  assign n26521 = n26520 ^ x8 ;
  assign n26522 = n26519 ^ x8 ;
  assign n26523 = n26522 ^ n7130 ;
  assign n26530 = n25287 & n26523 ;
  assign n26526 = ~x7 & ~n26523 ;
  assign n26527 = n26526 ^ n7131 ;
  assign n26528 = ~n25304 & ~n26527 ;
  assign n26529 = n26528 ^ n7130 ;
  assign n26531 = n26530 ^ n26529 ;
  assign n26532 = ~n26521 & ~n26531 ;
  assign n26533 = n26532 ^ n26314 ;
  assign n26534 = n26533 ^ n26306 ;
  assign n26535 = n26534 ^ n26532 ;
  assign n26536 = ~n26460 & ~n26535 ;
  assign n26537 = n26536 ^ n26533 ;
  assign n26699 = n26698 ^ n26537 ;
  assign n26510 = ~n9092 & n25703 ;
  assign n26511 = n26510 ^ x5 ;
  assign n26512 = n26511 ^ n26300 ;
  assign n26513 = n26512 ^ n26511 ;
  assign n26514 = n26513 ^ n26303 ;
  assign n26515 = ~n26462 & n26514 ;
  assign n26516 = n26515 ^ n26512 ;
  assign n26700 = n26699 ^ n26516 ;
  assign n26701 = n26700 ^ n26486 ;
  assign n26704 = n26703 ^ n26701 ;
  assign n26706 = n26705 ^ n26704 ;
  assign n26917 = ~n26704 & n26705 ;
  assign n26911 = n26698 ^ n26532 ;
  assign n26912 = ~n26537 & n26911 ;
  assign n26913 = n26912 ^ n26532 ;
  assign n26906 = n7141 & ~n25287 ;
  assign n26905 = n7135 & n25693 ;
  assign n26907 = n26906 ^ n26905 ;
  assign n26903 = n7146 ^ x8 ;
  assign n26900 = n8054 & n25287 ;
  assign n26901 = n26900 ^ n7146 ;
  assign n26902 = ~n25043 & n26901 ;
  assign n26904 = n26903 ^ n26902 ;
  assign n26908 = n26907 ^ n26904 ;
  assign n26863 = ~n6072 & n20836 ;
  assign n26862 = ~n6074 & n20837 ;
  assign n26864 = n26863 ^ n26862 ;
  assign n26865 = n26864 ^ n6060 ;
  assign n26866 = n26865 ^ x14 ;
  assign n26884 = n20834 ^ n6063 ;
  assign n26870 = n26864 ^ n6062 ;
  assign n26874 = n20834 ^ n17542 ;
  assign n26875 = n26874 ^ n20834 ;
  assign n26876 = ~n21055 & ~n26875 ;
  assign n26877 = n26876 ^ n20834 ;
  assign n26878 = ~n26870 & ~n26877 ;
  assign n26885 = n26884 ^ n26878 ;
  assign n26867 = n26864 ^ n17542 ;
  assign n26868 = n26867 ^ x14 ;
  assign n26869 = n26868 ^ n17542 ;
  assign n26881 = n26869 & n26878 ;
  assign n26882 = n26881 ^ n17542 ;
  assign n26883 = ~n21055 & ~n26882 ;
  assign n26886 = n26885 ^ n26883 ;
  assign n26887 = ~n26866 & n26886 ;
  assign n26852 = n14027 & n20882 ;
  assign n26845 = n20872 ^ x20 ;
  assign n26846 = n26845 ^ x19 ;
  assign n26847 = n26846 ^ n20872 ;
  assign n26848 = ~n23032 & n26847 ;
  assign n26849 = n26848 ^ n20872 ;
  assign n26850 = n4678 & ~n26849 ;
  assign n26851 = n26850 ^ x20 ;
  assign n26853 = n26852 ^ n26851 ;
  assign n26844 = n4916 & ~n20876 ;
  assign n26854 = n26853 ^ n26844 ;
  assign n26836 = ~n4496 & ~n21025 ;
  assign n26834 = n4492 & ~n22546 ;
  assign n26831 = n4504 & ~n20887 ;
  assign n26830 = n4491 & n20883 ;
  assign n26832 = n26831 ^ n26830 ;
  assign n26833 = n26832 ^ x23 ;
  assign n26835 = n26834 ^ n26833 ;
  assign n26837 = n26836 ^ n26835 ;
  assign n26814 = n3128 ^ n3003 ;
  assign n26812 = n589 ^ n557 ;
  assign n26810 = n1903 ^ n836 ;
  assign n26811 = n26810 ^ n642 ;
  assign n26813 = n26812 ^ n26811 ;
  assign n26815 = n26814 ^ n26813 ;
  assign n26816 = n26815 ^ n4978 ;
  assign n26807 = n1819 ^ n100 ;
  assign n26806 = n3850 ^ n1785 ;
  assign n26808 = n26807 ^ n26806 ;
  assign n26809 = n26808 ^ n14526 ;
  assign n26817 = n26816 ^ n26809 ;
  assign n26818 = n26817 ^ n1498 ;
  assign n26819 = n26818 ^ n2624 ;
  assign n26820 = ~n1277 & ~n26819 ;
  assign n26804 = n26627 ^ n26427 ;
  assign n26805 = n26605 & ~n26804 ;
  assign n26821 = n26820 ^ n26805 ;
  assign n26777 = n21001 ^ n20910 ;
  assign n26800 = ~n33 & n26777 ;
  assign n26794 = n26629 ^ n26598 ;
  assign n26795 = n26603 & n26794 ;
  assign n26796 = n26795 ^ n26598 ;
  assign n21649 = n20913 ^ n20910 ;
  assign n26789 = n20910 ^ n35 ;
  assign n26790 = n26789 ^ n20910 ;
  assign n26791 = n21649 & ~n26790 ;
  assign n26792 = n26791 ^ n20910 ;
  assign n26793 = ~n3514 & n26792 ;
  assign n26797 = n26796 ^ n26793 ;
  assign n26787 = n3722 & n20913 ;
  assign n26798 = n26797 ^ n26787 ;
  assign n26801 = n26798 ^ n26797 ;
  assign n26802 = n26800 & n26801 ;
  assign n26775 = n26593 ^ n20913 ;
  assign n26776 = n26775 ^ n26593 ;
  assign n26782 = n3520 & n26777 ;
  assign n26783 = ~n26776 & n26782 ;
  assign n26784 = n26783 ^ n26776 ;
  assign n26785 = n26784 ^ n26775 ;
  assign n26786 = x31 & n26785 ;
  assign n26799 = n26798 ^ n26786 ;
  assign n26803 = n26802 ^ n26799 ;
  assign n26822 = n26821 ^ n26803 ;
  assign n26770 = n12861 & n20898 ;
  assign n26769 = n446 & n20897 ;
  assign n26771 = n26770 ^ n26769 ;
  assign n26772 = n26771 ^ x26 ;
  assign n26768 = ~n487 & ~n20894 ;
  assign n26773 = n26772 ^ n26768 ;
  assign n26767 = ~n3501 & n21954 ;
  assign n26774 = n26773 ^ n26767 ;
  assign n26823 = n26822 ^ n26774 ;
  assign n26764 = n3484 & n20902 ;
  assign n26757 = n21735 ^ x29 ;
  assign n26758 = n26757 ^ x28 ;
  assign n26759 = n26758 ^ n21735 ;
  assign n26760 = ~n21734 & ~n26759 ;
  assign n26761 = n26760 ^ n21735 ;
  assign n26762 = n650 & n26761 ;
  assign n26763 = n26762 ^ x29 ;
  assign n26765 = n26764 ^ n26763 ;
  assign n26756 = n831 & n20903 ;
  assign n26766 = n26765 ^ n26756 ;
  assign n26824 = n26823 ^ n26766 ;
  assign n26825 = n26824 ^ n26657 ;
  assign n26826 = n26825 ^ n26630 ;
  assign n26827 = n26826 ^ n26824 ;
  assign n26828 = n26635 & n26827 ;
  assign n26829 = n26828 ^ n26825 ;
  assign n26838 = n26837 ^ n26829 ;
  assign n26839 = n26838 ^ n26661 ;
  assign n26840 = n26839 ^ n26574 ;
  assign n26841 = n26840 ^ n26838 ;
  assign n26842 = n26662 & n26841 ;
  assign n26843 = n26842 ^ n26839 ;
  assign n26855 = n26854 ^ n26843 ;
  assign n26743 = n20731 & n20865 ;
  assign n26742 = n5700 & n20861 ;
  assign n26744 = n26743 ^ n26742 ;
  assign n26745 = n26744 ^ n5694 ;
  assign n26746 = n26744 ^ x17 ;
  assign n26750 = n26746 ^ n5696 ;
  assign n26751 = ~x16 & ~n23059 ;
  assign n26752 = n26750 & n26751 ;
  assign n26748 = n5696 & ~n23825 ;
  assign n26747 = ~n20852 & n26746 ;
  assign n26749 = n26748 ^ n26747 ;
  assign n26753 = n26752 ^ n26749 ;
  assign n26754 = ~n26745 & ~n26753 ;
  assign n26739 = n26676 ^ n26663 ;
  assign n26740 = n26668 & n26739 ;
  assign n26741 = n26740 ^ n26663 ;
  assign n26755 = n26754 ^ n26741 ;
  assign n26856 = n26855 ^ n26755 ;
  assign n26857 = n26856 ^ n26680 ;
  assign n26858 = n26857 ^ n26566 ;
  assign n26859 = n26858 ^ n26856 ;
  assign n26860 = n26681 & n26859 ;
  assign n26861 = n26860 ^ n26857 ;
  assign n26888 = n26887 ^ n26861 ;
  assign n26736 = n26558 ^ n26555 ;
  assign n26737 = n26683 & n26736 ;
  assign n26738 = n26737 ^ n26555 ;
  assign n26889 = n26888 ^ n26738 ;
  assign n26734 = n6650 & ~n24700 ;
  assign n26732 = n15413 & n25517 ;
  assign n26729 = n6655 & n24079 ;
  assign n26728 = n6658 & ~n24980 ;
  assign n26730 = n26729 ^ n26728 ;
  assign n26731 = n26730 ^ x11 ;
  assign n26733 = n26732 ^ n26731 ;
  assign n26735 = n26734 ^ n26733 ;
  assign n26890 = n26889 ^ n26735 ;
  assign n26892 = n26890 ^ n26684 ;
  assign n26891 = n26890 ^ n26697 ;
  assign n26893 = n26892 ^ n26891 ;
  assign n26894 = ~n26689 & n26893 ;
  assign n26895 = n26894 ^ n26892 ;
  assign n26909 = n26908 ^ n26895 ;
  assign n26910 = n26909 ^ x5 ;
  assign n26914 = n26913 ^ n26910 ;
  assign n26725 = n26699 ^ n26511 ;
  assign n26726 = n26516 & n26725 ;
  assign n26727 = n26726 ^ n26511 ;
  assign n26915 = n26914 ^ n26727 ;
  assign n26707 = n26700 ^ n26471 ;
  assign n26709 = n26502 ^ n26481 ;
  assign n26708 = n26700 ^ n26478 ;
  assign n26710 = n26709 ^ n26708 ;
  assign n26711 = n26710 ^ n26708 ;
  assign n26712 = n26708 ^ n26482 ;
  assign n26713 = n26712 ^ n26708 ;
  assign n26714 = ~n26711 & n26713 ;
  assign n26715 = n26714 ^ n26708 ;
  assign n26716 = ~n26707 & n26715 ;
  assign n26717 = n26716 ^ n26471 ;
  assign n26718 = ~n26470 & n26717 ;
  assign n26719 = ~n26708 & ~n26709 ;
  assign n26720 = n26700 ^ n26481 ;
  assign n26721 = n26719 & ~n26720 ;
  assign n26722 = n26721 ^ n26700 ;
  assign n26723 = n26718 & n26722 ;
  assign n26724 = n26723 ^ n26717 ;
  assign n26916 = n26915 ^ n26724 ;
  assign n26918 = n26917 ^ n26916 ;
  assign n27093 = n26913 ^ n26909 ;
  assign n27094 = n26910 & n27093 ;
  assign n27081 = n4916 & ~n20872 ;
  assign n27080 = n4681 & ~n22683 ;
  assign n27082 = n27081 ^ n27080 ;
  assign n27077 = n4682 & n20865 ;
  assign n27076 = ~n4679 & ~n22682 ;
  assign n27078 = n27077 ^ n27076 ;
  assign n27074 = n14027 & ~n20876 ;
  assign n27073 = ~x20 & n22682 ;
  assign n27075 = n27074 ^ n27073 ;
  assign n27079 = n27078 ^ n27075 ;
  assign n27083 = n27082 ^ n27079 ;
  assign n27069 = ~n4496 & n20883 ;
  assign n27062 = n26837 ^ n26824 ;
  assign n27063 = ~n26829 & n27062 ;
  assign n27064 = n27063 ^ n26824 ;
  assign n27065 = n27064 ^ x23 ;
  assign n27061 = n4504 & ~n21025 ;
  assign n27066 = n27065 ^ n27061 ;
  assign n27060 = n4491 & n20882 ;
  assign n27067 = n27066 ^ n27060 ;
  assign n27059 = n4492 & ~n22672 ;
  assign n27068 = n27067 ^ n27059 ;
  assign n27070 = n27069 ^ n27068 ;
  assign n27052 = n26606 & ~n26627 ;
  assign n27053 = ~n26820 & n27052 ;
  assign n27037 = n26627 & n26820 ;
  assign n27038 = ~n26606 & n27037 ;
  assign n27054 = n27053 ^ n27038 ;
  assign n27055 = ~x2 & n27054 ;
  assign n27048 = n3484 & ~n21012 ;
  assign n27041 = n20898 ^ x29 ;
  assign n27042 = n27041 ^ x28 ;
  assign n27043 = n27042 ^ n20898 ;
  assign n27044 = ~n21971 & n27043 ;
  assign n27045 = n27044 ^ n20898 ;
  assign n27046 = n650 & n27045 ;
  assign n27047 = n27046 ^ x29 ;
  assign n27049 = n27048 ^ n27047 ;
  assign n27040 = n831 & n20902 ;
  assign n27050 = n27049 ^ n27040 ;
  assign n27028 = n4793 ^ n710 ;
  assign n27029 = n27028 ^ n2849 ;
  assign n27030 = n27029 ^ n13241 ;
  assign n27026 = n5120 ^ n4806 ;
  assign n27023 = n567 ^ n226 ;
  assign n27024 = n27023 ^ n153 ;
  assign n27021 = n615 ^ n219 ;
  assign n27022 = n27021 ^ n506 ;
  assign n27025 = n27024 ^ n27022 ;
  assign n27027 = n27026 ^ n27025 ;
  assign n27031 = n27030 ^ n27027 ;
  assign n27032 = n27031 ^ n23753 ;
  assign n27033 = n27032 ^ n3572 ;
  assign n27034 = ~n2396 & ~n27033 ;
  assign n27035 = n27034 ^ x5 ;
  assign n27011 = n20903 ^ x30 ;
  assign n27012 = n27011 ^ n20903 ;
  assign n27013 = n23553 & n27012 ;
  assign n27014 = n27013 ^ n20903 ;
  assign n27015 = ~n3520 & n27014 ;
  assign n27016 = n27015 ^ n20903 ;
  assign n27017 = n27016 ^ n21756 ;
  assign n27004 = n21756 ^ n20910 ;
  assign n27003 = n21756 ^ n20913 ;
  assign n27005 = n27004 ^ n27003 ;
  assign n27006 = n27004 ^ x30 ;
  assign n27007 = n27006 ^ n27004 ;
  assign n27008 = n27005 & n27007 ;
  assign n27009 = n27008 ^ n27004 ;
  assign n27010 = ~n3520 & ~n27009 ;
  assign n27018 = n27017 ^ n27010 ;
  assign n27019 = x31 & ~n27018 ;
  assign n27020 = n27019 ^ n27016 ;
  assign n27036 = n27035 ^ n27020 ;
  assign n27039 = n27038 ^ n27036 ;
  assign n27051 = n27050 ^ n27039 ;
  assign n27056 = n27055 ^ n27051 ;
  assign n27000 = n26821 ^ n26796 ;
  assign n27001 = n26803 & n27000 ;
  assign n27002 = n27001 ^ n26821 ;
  assign n27057 = n27056 ^ n27002 ;
  assign n26974 = n12861 & n20897 ;
  assign n26973 = n446 & ~n20894 ;
  assign n26975 = n26974 ^ n26973 ;
  assign n26976 = n26975 ^ n65 ;
  assign n26977 = n26975 ^ x26 ;
  assign n26978 = n26977 ^ n67 ;
  assign n26979 = n26978 ^ x25 ;
  assign n26980 = n26979 ^ n20887 ;
  assign n26981 = n26980 ^ n26977 ;
  assign n26982 = n26981 ^ n22306 ;
  assign n26983 = n26982 ^ n26981 ;
  assign n26984 = n26977 & ~n26983 ;
  assign n26985 = n26984 ^ n26978 ;
  assign n26986 = n26981 ^ n20887 ;
  assign n26987 = ~n26983 & ~n26986 ;
  assign n26988 = n26987 ^ n20887 ;
  assign n26989 = ~n26978 & n26988 ;
  assign n26990 = ~n26985 & n26989 ;
  assign n26991 = n26990 ^ n26987 ;
  assign n26992 = n26991 ^ n67 ;
  assign n26993 = n26992 ^ n20887 ;
  assign n26994 = ~n26976 & ~n26993 ;
  assign n26995 = n26994 ^ n26774 ;
  assign n26996 = n26995 ^ n26766 ;
  assign n26997 = n26996 ^ n26994 ;
  assign n26998 = n26823 & n26997 ;
  assign n26999 = n26998 ^ n26995 ;
  assign n27058 = n27057 ^ n26999 ;
  assign n27071 = n27070 ^ n27058 ;
  assign n26970 = n26854 ^ n26838 ;
  assign n26971 = ~n26843 & ~n26970 ;
  assign n26972 = n26971 ^ n26838 ;
  assign n27072 = n27071 ^ n26972 ;
  assign n27084 = n27083 ^ n27072 ;
  assign n26965 = n5700 & n20852 ;
  assign n26964 = n5702 & n20836 ;
  assign n26966 = n26965 ^ n26964 ;
  assign n26967 = n26966 ^ x17 ;
  assign n26963 = n5703 & ~n24433 ;
  assign n26968 = n26967 ^ n26963 ;
  assign n26962 = n20731 & n20861 ;
  assign n26969 = n26968 ^ n26962 ;
  assign n27085 = n27084 ^ n26969 ;
  assign n26959 = n26855 ^ n26741 ;
  assign n26960 = n26755 & ~n26959 ;
  assign n26961 = n26960 ^ n26855 ;
  assign n27086 = n27085 ^ n26961 ;
  assign n26943 = ~x13 & ~n24004 ;
  assign n26944 = n26943 ^ n24079 ;
  assign n26951 = n6060 & n26944 ;
  assign n26948 = ~n6072 & n20837 ;
  assign n26947 = ~n6074 & n20834 ;
  assign n26949 = n26948 ^ n26947 ;
  assign n26950 = n26949 ^ x14 ;
  assign n26952 = n26951 ^ n26950 ;
  assign n26945 = n26944 ^ n24004 ;
  assign n26946 = n6063 & ~n26945 ;
  assign n26953 = n26952 ^ n26946 ;
  assign n26955 = n26953 ^ n26856 ;
  assign n26954 = n26953 ^ n26887 ;
  assign n26956 = n26955 ^ n26954 ;
  assign n26957 = n26861 & ~n26956 ;
  assign n26958 = n26957 ^ n26955 ;
  assign n27087 = n27086 ^ n26958 ;
  assign n26941 = n6650 & ~n24980 ;
  assign n26939 = n15413 & ~n25896 ;
  assign n26936 = n6655 & ~n24700 ;
  assign n26935 = n6658 & n25043 ;
  assign n26937 = n26936 ^ n26935 ;
  assign n26938 = n26937 ^ x11 ;
  assign n26940 = n26939 ^ n26938 ;
  assign n26942 = n26941 ^ n26940 ;
  assign n27088 = n27087 ^ n26942 ;
  assign n26932 = n26738 ^ n26735 ;
  assign n26933 = n26889 & ~n26932 ;
  assign n26934 = n26933 ^ n26738 ;
  assign n27089 = n27088 ^ n26934 ;
  assign n26927 = n7146 ^ n7141 ;
  assign n26928 = n26927 ^ n26517 ;
  assign n26929 = n25287 & n26928 ;
  assign n26930 = n26929 ^ n26903 ;
  assign n26926 = n7135 & n25725 ;
  assign n26931 = n26930 ^ n26926 ;
  assign n27090 = n27089 ^ n26931 ;
  assign n26923 = n26908 ^ n26890 ;
  assign n26924 = n26895 & n26923 ;
  assign n26925 = n26924 ^ n26890 ;
  assign n27091 = n27090 ^ n26925 ;
  assign n27092 = n27091 ^ x5 ;
  assign n27095 = n27094 ^ n27092 ;
  assign n26920 = n26727 ^ n26724 ;
  assign n26921 = n26915 & n26920 ;
  assign n26919 = n26916 & ~n26917 ;
  assign n26922 = n26921 ^ n26919 ;
  assign n27096 = n27095 ^ n26922 ;
  assign n27301 = n27095 ^ n26915 ;
  assign n27302 = n26916 & ~n27301 ;
  assign n27303 = n26917 & n27302 ;
  assign n27298 = n26931 ^ n26925 ;
  assign n27299 = ~n27090 & n27298 ;
  assign n27300 = n27299 ^ n26931 ;
  assign n27304 = n27303 ^ n27300 ;
  assign n27271 = n26909 & ~n26913 ;
  assign n27272 = n27271 ^ n27093 ;
  assign n27280 = n27271 ^ n27091 ;
  assign n27273 = n27091 & ~n27271 ;
  assign n27281 = n27280 ^ n27273 ;
  assign n27274 = n26727 ^ x5 ;
  assign n27277 = ~n26920 & n27274 ;
  assign n27278 = n27277 ^ n26727 ;
  assign n27279 = ~n27273 & n27278 ;
  assign n27282 = n27281 ^ n27279 ;
  assign n27283 = n27091 ^ n26724 ;
  assign n27284 = n27283 ^ n26724 ;
  assign n27285 = n27284 ^ n26727 ;
  assign n27288 = n27284 ^ n27092 ;
  assign n27289 = n27288 ^ n27284 ;
  assign n27290 = n27283 & ~n27289 ;
  assign n27291 = ~n27285 & n27290 ;
  assign n27292 = n27291 ^ n27285 ;
  assign n27293 = n27292 ^ n26727 ;
  assign n27294 = ~n27282 & ~n27293 ;
  assign n27295 = ~n27272 & n27294 ;
  assign n27296 = n27295 ^ n27282 ;
  assign n27267 = n7146 & n25703 ;
  assign n27268 = n27267 ^ x8 ;
  assign n27264 = n26942 ^ n26934 ;
  assign n27265 = n27088 & n27264 ;
  assign n27266 = n27265 ^ n27087 ;
  assign n27269 = n27268 ^ n27266 ;
  assign n27259 = n27086 ^ n26953 ;
  assign n27260 = n26958 & n27259 ;
  assign n27261 = n27260 ^ n26953 ;
  assign n27248 = n27057 ^ n26994 ;
  assign n27249 = ~n26999 & ~n27248 ;
  assign n27250 = n27249 ^ n26994 ;
  assign n27242 = n12861 & ~n20894 ;
  assign n27241 = n446 & ~n20887 ;
  assign n27243 = n27242 ^ n27241 ;
  assign n27244 = n27243 ^ x26 ;
  assign n27240 = ~n487 & ~n21025 ;
  assign n27245 = n27244 ^ n27240 ;
  assign n27239 = ~n3501 & n22415 ;
  assign n27246 = n27245 ^ n27239 ;
  assign n27224 = n3484 & n20898 ;
  assign n27217 = n20897 ^ x29 ;
  assign n27218 = n27217 ^ x28 ;
  assign n27219 = n27218 ^ n20897 ;
  assign n27220 = ~n23665 & n27219 ;
  assign n27221 = n27220 ^ n20897 ;
  assign n27222 = n650 & n27221 ;
  assign n27223 = n27222 ^ x29 ;
  assign n27225 = n27224 ^ n27223 ;
  assign n27216 = n831 & ~n21012 ;
  assign n27226 = n27225 ^ n27216 ;
  assign n27227 = n27226 ^ n27020 ;
  assign n27209 = n27053 ^ n27035 ;
  assign n27208 = n27038 ^ n27020 ;
  assign n27210 = n27209 ^ n27208 ;
  assign n27211 = ~n27054 & ~n27210 ;
  assign n27212 = n27211 ^ n27208 ;
  assign n27213 = n27035 ^ x2 ;
  assign n27214 = n27213 ^ n27020 ;
  assign n27215 = ~n27212 & ~n27214 ;
  assign n27228 = n27227 ^ n27215 ;
  assign n27201 = n3539 ^ n868 ;
  assign n27197 = n245 ^ n90 ;
  assign n27198 = n27197 ^ n6484 ;
  assign n27199 = n27198 ^ n12491 ;
  assign n27200 = n27199 ^ n1369 ;
  assign n27202 = n27201 ^ n27200 ;
  assign n27194 = n5302 ^ n3846 ;
  assign n27192 = n862 ^ n558 ;
  assign n27191 = n3022 ^ n589 ;
  assign n27193 = n27192 ^ n27191 ;
  assign n27195 = n27194 ^ n27193 ;
  assign n27196 = n27195 ^ n2053 ;
  assign n27203 = n27202 ^ n27196 ;
  assign n27186 = n1099 ^ n109 ;
  assign n27185 = n12406 ^ n206 ;
  assign n27187 = n27186 ^ n27185 ;
  assign n27188 = n27187 ^ n12394 ;
  assign n27189 = n27188 ^ n997 ;
  assign n27182 = n2516 ^ n1927 ;
  assign n27183 = n27182 ^ n6434 ;
  assign n27180 = n5614 ^ n1339 ;
  assign n27181 = n27180 ^ n1896 ;
  assign n27184 = n27183 ^ n27181 ;
  assign n27190 = n27189 ^ n27184 ;
  assign n27204 = n27203 ^ n27190 ;
  assign n27205 = ~n1470 & ~n27204 ;
  assign n27178 = n5328 & ~n27035 ;
  assign n27179 = n27178 ^ x2 ;
  assign n27206 = n27205 ^ n27179 ;
  assign n27172 = x30 & n20903 ;
  assign n27158 = n21744 ^ n20903 ;
  assign n27157 = n21744 ^ n20910 ;
  assign n27159 = n27158 ^ n27157 ;
  assign n27162 = x30 & n27159 ;
  assign n27163 = n27162 ^ n27158 ;
  assign n27164 = ~n3520 & ~n27163 ;
  assign n27165 = n27164 ^ n21744 ;
  assign n27166 = n27165 ^ n20902 ;
  assign n27167 = n27166 ^ n27165 ;
  assign n27173 = n27172 ^ n27167 ;
  assign n27174 = ~n3520 & n27173 ;
  assign n27175 = n27174 ^ n27166 ;
  assign n27176 = ~x31 & ~n27175 ;
  assign n27177 = n27176 ^ n27165 ;
  assign n27207 = n27206 ^ n27177 ;
  assign n27233 = n27228 ^ n27207 ;
  assign n27234 = n27233 ^ n27050 ;
  assign n27235 = n27234 ^ n27233 ;
  assign n27236 = n27235 ^ n27002 ;
  assign n27237 = ~n27056 & ~n27236 ;
  assign n27238 = n27237 ^ n27234 ;
  assign n27247 = n27246 ^ n27238 ;
  assign n27251 = n27250 ^ n27247 ;
  assign n27155 = ~n4496 & n20882 ;
  assign n27153 = n4492 & n23010 ;
  assign n27150 = n4504 & n20883 ;
  assign n27149 = n4491 & ~n20876 ;
  assign n27151 = n27150 ^ n27149 ;
  assign n27152 = n27151 ^ x23 ;
  assign n27154 = n27153 ^ n27152 ;
  assign n27156 = n27155 ^ n27154 ;
  assign n27252 = n27251 ^ n27156 ;
  assign n27146 = n27064 ^ n27058 ;
  assign n27147 = n27070 & ~n27146 ;
  assign n27148 = n27147 ^ n27064 ;
  assign n27253 = n27252 ^ n27148 ;
  assign n27143 = n4916 & n20865 ;
  assign n27136 = n20861 ^ x20 ;
  assign n27137 = n27136 ^ x19 ;
  assign n27138 = n27137 ^ n20861 ;
  assign n27139 = ~n23608 & n27138 ;
  assign n27140 = n27139 ^ n20861 ;
  assign n27141 = n4678 & n27140 ;
  assign n27142 = n27141 ^ x20 ;
  assign n27144 = n27143 ^ n27142 ;
  assign n27135 = n14027 & ~n20872 ;
  assign n27145 = n27144 ^ n27135 ;
  assign n27254 = n27253 ^ n27145 ;
  assign n27132 = n27083 ^ n26972 ;
  assign n27133 = ~n27072 & n27132 ;
  assign n27134 = n27133 ^ n27083 ;
  assign n27255 = n27254 ^ n27134 ;
  assign n27130 = n20731 & n20852 ;
  assign n27128 = n5703 & ~n24427 ;
  assign n27125 = n5700 & n20836 ;
  assign n27124 = n5702 & n20837 ;
  assign n27126 = n27125 ^ n27124 ;
  assign n27127 = n27126 ^ x17 ;
  assign n27129 = n27128 ^ n27127 ;
  assign n27131 = n27130 ^ n27129 ;
  assign n27256 = n27255 ^ n27131 ;
  assign n27121 = n26969 ^ n26961 ;
  assign n27122 = ~n27085 & ~n27121 ;
  assign n27123 = n27122 ^ n26969 ;
  assign n27257 = n27256 ^ n27123 ;
  assign n27116 = n24079 ^ x14 ;
  assign n27107 = n24700 ^ x13 ;
  assign n27106 = n24700 ^ x14 ;
  assign n27108 = n27107 ^ n27106 ;
  assign n27109 = n24463 & n27108 ;
  assign n27110 = n27109 ^ n27107 ;
  assign n27117 = n27116 ^ n27110 ;
  assign n27111 = n24079 ^ n4899 ;
  assign n27112 = n27111 ^ n24079 ;
  assign n27113 = n24707 & n27112 ;
  assign n27114 = n27113 ^ n24079 ;
  assign n27115 = ~n6066 & n27114 ;
  assign n27118 = n27117 ^ n27115 ;
  assign n27119 = ~n4897 & ~n27118 ;
  assign n27120 = n27119 ^ n27110 ;
  assign n27258 = n27257 ^ n27120 ;
  assign n27262 = n27261 ^ n27258 ;
  assign n27101 = n6650 & n25043 ;
  assign n27099 = n6658 & n25287 ;
  assign n27100 = n27099 ^ n6658 ;
  assign n27102 = n27101 ^ n27100 ;
  assign n27103 = n27102 ^ x11 ;
  assign n27098 = n6655 & ~n24980 ;
  assign n27104 = n27103 ^ n27098 ;
  assign n27097 = n15413 & n25937 ;
  assign n27105 = n27104 ^ n27097 ;
  assign n27263 = n27262 ^ n27105 ;
  assign n27270 = n27269 ^ n27263 ;
  assign n27297 = n27296 ^ n27270 ;
  assign n27305 = n27304 ^ n27297 ;
  assign n27306 = n27300 ^ n27270 ;
  assign n27307 = n27306 ^ n27296 ;
  assign n27310 = n27266 ^ n27263 ;
  assign n27478 = n6650 & ~n25287 ;
  assign n27477 = n15413 & n25693 ;
  assign n27479 = n27478 ^ n27477 ;
  assign n27476 = n6655 ^ x11 ;
  assign n27480 = n27479 ^ n27476 ;
  assign n27474 = n27099 ^ n6655 ;
  assign n27475 = ~n25043 & n27474 ;
  assign n27481 = n27480 ^ n27475 ;
  assign n27448 = ~n6074 & ~n24700 ;
  assign n27447 = ~n6072 & n24079 ;
  assign n27449 = n27448 ^ n27447 ;
  assign n27450 = n27449 ^ n6060 ;
  assign n27451 = n27450 ^ x14 ;
  assign n27468 = n24980 ^ n6063 ;
  assign n27455 = n27449 ^ n6062 ;
  assign n27458 = n24980 ^ n17542 ;
  assign n27459 = n27458 ^ n24980 ;
  assign n27460 = ~n25518 & ~n27459 ;
  assign n27461 = n27460 ^ n24980 ;
  assign n27462 = ~n27455 & n27461 ;
  assign n27469 = n27468 ^ n27462 ;
  assign n27452 = n27449 ^ n17542 ;
  assign n27453 = n27452 ^ x14 ;
  assign n27454 = n27453 ^ n17542 ;
  assign n27463 = n27462 ^ n17542 ;
  assign n27464 = n27463 ^ n17542 ;
  assign n27465 = n27454 & n27464 ;
  assign n27466 = n27465 ^ n17542 ;
  assign n27467 = ~n24949 & ~n27466 ;
  assign n27470 = n27469 ^ n27467 ;
  assign n27471 = ~n27451 & ~n27470 ;
  assign n27436 = n5700 & n20837 ;
  assign n27435 = n5702 & n20834 ;
  assign n27437 = n27436 ^ n27435 ;
  assign n27438 = n27437 ^ x17 ;
  assign n27434 = n5703 & ~n24936 ;
  assign n27439 = n27438 ^ n27434 ;
  assign n27433 = n20731 & n20836 ;
  assign n27440 = n27439 ^ n27433 ;
  assign n27424 = n4678 & ~n23059 ;
  assign n27425 = x20 & n27424 ;
  assign n27419 = n4682 & n20852 ;
  assign n27418 = n4916 & n20861 ;
  assign n27420 = n27419 ^ n27418 ;
  assign n27416 = n14027 & n20865 ;
  assign n27415 = n4681 & ~n23825 ;
  assign n27417 = n27416 ^ n27415 ;
  assign n27421 = n27420 ^ n27417 ;
  assign n27422 = n27421 ^ x20 ;
  assign n27426 = n27425 ^ n27422 ;
  assign n27404 = n4504 & n20882 ;
  assign n27403 = n4491 & ~n20872 ;
  assign n27405 = n27404 ^ n27403 ;
  assign n27406 = n27405 ^ x23 ;
  assign n27402 = n4492 & n23033 ;
  assign n27407 = n27406 ^ n27402 ;
  assign n27401 = ~n4496 & ~n20876 ;
  assign n27408 = n27407 ^ n27401 ;
  assign n27392 = n3484 & n20897 ;
  assign n27379 = n21735 ^ n20902 ;
  assign n27378 = n21735 ^ n20903 ;
  assign n27380 = n27379 ^ n27378 ;
  assign n27383 = x30 & n27380 ;
  assign n27384 = n27383 ^ n27379 ;
  assign n27385 = ~n3520 & n27384 ;
  assign n27386 = n27385 ^ n21735 ;
  assign n27387 = x31 & n27386 ;
  assign n27371 = n13647 ^ n4352 ;
  assign n27368 = n11823 ^ n490 ;
  assign n27369 = n27368 ^ n3103 ;
  assign n27367 = n2354 ^ n952 ;
  assign n27370 = n27369 ^ n27367 ;
  assign n27372 = n27371 ^ n27370 ;
  assign n27363 = n1842 ^ n999 ;
  assign n27364 = n27363 ^ n1654 ;
  assign n27365 = n27364 ^ n4181 ;
  assign n27366 = n27365 ^ n2862 ;
  assign n27373 = n27372 ^ n27366 ;
  assign n27356 = n1677 ^ n379 ;
  assign n27357 = n27356 ^ n697 ;
  assign n27355 = n726 ^ n202 ;
  assign n27358 = n27357 ^ n27355 ;
  assign n27359 = n27358 ^ n842 ;
  assign n27360 = n27359 ^ n3552 ;
  assign n27352 = n1286 ^ n1198 ;
  assign n27351 = n1492 ^ n1171 ;
  assign n27353 = n27352 ^ n27351 ;
  assign n27349 = n797 ^ n143 ;
  assign n27346 = n2621 ^ n122 ;
  assign n27347 = n27346 ^ n848 ;
  assign n27348 = n27347 ^ n520 ;
  assign n27350 = n27349 ^ n27348 ;
  assign n27354 = n27353 ^ n27350 ;
  assign n27361 = n27360 ^ n27354 ;
  assign n27362 = n27361 ^ n3993 ;
  assign n27374 = n27373 ^ n27362 ;
  assign n27375 = ~n13252 & ~n27374 ;
  assign n27344 = n27179 ^ n27177 ;
  assign n27345 = ~n27206 & ~n27344 ;
  assign n27376 = n27375 ^ n27345 ;
  assign n27341 = n35 & ~n23255 ;
  assign n27342 = n27341 ^ n20902 ;
  assign n27343 = ~n3514 & n27342 ;
  assign n27377 = n27376 ^ n27343 ;
  assign n27388 = n27387 ^ n27377 ;
  assign n27336 = n27226 ^ n27207 ;
  assign n27337 = n27228 & n27336 ;
  assign n27338 = n27337 ^ n27226 ;
  assign n27389 = n27388 ^ n27338 ;
  assign n27390 = n27389 ^ x29 ;
  assign n27331 = n20894 ^ n4536 ;
  assign n27332 = n27331 ^ n20894 ;
  assign n27333 = ~n23953 & n27332 ;
  assign n27334 = n27333 ^ n20894 ;
  assign n27335 = n650 & ~n27334 ;
  assign n27391 = n27390 ^ n27335 ;
  assign n27393 = n27392 ^ n27391 ;
  assign n27330 = n831 & n20898 ;
  assign n27394 = n27393 ^ n27330 ;
  assign n27318 = n12861 & ~n20887 ;
  assign n27317 = n446 & ~n21025 ;
  assign n27319 = n27318 ^ n27317 ;
  assign n27320 = n27319 ^ n65 ;
  assign n27321 = n27319 ^ x26 ;
  assign n27325 = n27321 ^ n67 ;
  assign n27326 = ~x25 & ~n22545 ;
  assign n27327 = n27325 & n27326 ;
  assign n27323 = n67 & ~n22546 ;
  assign n27322 = ~n20883 & n27321 ;
  assign n27324 = n27323 ^ n27322 ;
  assign n27328 = n27327 ^ n27324 ;
  assign n27329 = ~n27320 & ~n27328 ;
  assign n27395 = n27394 ^ n27329 ;
  assign n27397 = n27395 ^ n27233 ;
  assign n27396 = n27395 ^ n27246 ;
  assign n27398 = n27397 ^ n27396 ;
  assign n27399 = n27238 & n27398 ;
  assign n27400 = n27399 ^ n27397 ;
  assign n27409 = n27408 ^ n27400 ;
  assign n27410 = n27409 ^ n27250 ;
  assign n27411 = n27410 ^ n27156 ;
  assign n27412 = n27411 ^ n27409 ;
  assign n27413 = ~n27251 & ~n27412 ;
  assign n27414 = n27413 ^ n27410 ;
  assign n27427 = n27426 ^ n27414 ;
  assign n27428 = n27427 ^ n27145 ;
  assign n27429 = n27428 ^ n27427 ;
  assign n27430 = n27429 ^ n27148 ;
  assign n27431 = n27253 & n27430 ;
  assign n27432 = n27431 ^ n27428 ;
  assign n27441 = n27440 ^ n27432 ;
  assign n27442 = n27441 ^ n27131 ;
  assign n27443 = n27442 ^ n27441 ;
  assign n27444 = n27443 ^ n27134 ;
  assign n27445 = ~n27255 & ~n27444 ;
  assign n27446 = n27445 ^ n27442 ;
  assign n27472 = n27471 ^ n27446 ;
  assign n27314 = n27123 ^ n27120 ;
  assign n27315 = n27257 & ~n27314 ;
  assign n27316 = n27315 ^ n27123 ;
  assign n27473 = n27472 ^ n27316 ;
  assign n27482 = n27481 ^ n27473 ;
  assign n27483 = n27482 ^ x8 ;
  assign n27311 = n27261 ^ n27105 ;
  assign n27312 = ~n27262 & n27311 ;
  assign n27313 = n27312 ^ n27261 ;
  assign n27484 = n27483 ^ n27313 ;
  assign n27485 = n27484 ^ n27268 ;
  assign n27486 = n27485 ^ n27484 ;
  assign n27487 = n27486 ^ n27266 ;
  assign n27488 = n27310 & n27487 ;
  assign n27489 = n27488 ^ n27485 ;
  assign n27308 = ~n27270 & n27296 ;
  assign n27309 = n27308 ^ n27303 ;
  assign n27490 = n27489 ^ n27309 ;
  assign n27491 = n27490 ^ n27297 ;
  assign n27492 = n27491 ^ n27308 ;
  assign n27493 = n27492 ^ n27489 ;
  assign n27494 = n27307 & ~n27493 ;
  assign n27495 = n27494 ^ n27490 ;
  assign n27671 = n27489 ^ n27308 ;
  assign n27672 = ~n27307 & n27671 ;
  assign n27673 = n27303 & n27672 ;
  assign n27664 = n27440 ^ n27427 ;
  assign n27665 = ~n27432 & ~n27664 ;
  assign n27666 = n27665 ^ n27427 ;
  assign n27661 = n5703 & ~n25245 ;
  assign n27659 = n5700 & n20834 ;
  assign n27657 = n5702 & n24079 ;
  assign n27646 = n27376 ^ n27338 ;
  assign n27647 = ~n27388 & ~n27646 ;
  assign n27648 = n27647 ^ n27376 ;
  assign n27635 = n1195 ^ n985 ;
  assign n27634 = n14549 ^ n2863 ;
  assign n27636 = n27635 ^ n27634 ;
  assign n27631 = n3453 ^ n2627 ;
  assign n27632 = n27631 ^ n2043 ;
  assign n27630 = n13211 ^ n12789 ;
  assign n27633 = n27632 ^ n27630 ;
  assign n27637 = n27636 ^ n27633 ;
  assign n27638 = n27637 ^ n2978 ;
  assign n27639 = n5347 ^ n2590 ;
  assign n27640 = n27639 ^ n903 ;
  assign n27641 = ~n27638 & ~n27640 ;
  assign n27642 = n27641 ^ n27205 ;
  assign n27643 = n27642 ^ x8 ;
  assign n27612 = ~n35 & n21012 ;
  assign n27613 = n27612 ^ x29 ;
  assign n27604 = n21972 ^ n20902 ;
  assign n27603 = n21972 ^ n21012 ;
  assign n27605 = n27604 ^ n27603 ;
  assign n27608 = ~x30 & ~n27605 ;
  assign n27609 = n27608 ^ n27604 ;
  assign n27610 = ~n3520 & ~n27609 ;
  assign n27611 = n27610 ^ n21972 ;
  assign n27614 = n27613 ^ n27611 ;
  assign n27615 = n27614 ^ n20898 ;
  assign n27616 = n27615 ^ x30 ;
  assign n27617 = n27616 ^ n27614 ;
  assign n27618 = n27614 ^ x29 ;
  assign n27619 = n27618 ^ n20898 ;
  assign n27620 = n27619 ^ n27614 ;
  assign n27621 = ~n27617 & n27620 ;
  assign n27622 = n27621 ^ n27614 ;
  assign n27623 = ~x31 & ~n27622 ;
  assign n27624 = n27623 ^ n27611 ;
  assign n27625 = n27624 ^ n27205 ;
  assign n27626 = n27625 ^ n27375 ;
  assign n27627 = n27626 ^ n27624 ;
  assign n27628 = n27345 & ~n27627 ;
  assign n27629 = n27628 ^ n27625 ;
  assign n27644 = n27643 ^ n27629 ;
  assign n27601 = n831 & n20897 ;
  assign n27599 = n3484 & ~n20894 ;
  assign n27592 = n20887 ^ x29 ;
  assign n27593 = n27592 ^ x28 ;
  assign n27594 = n27593 ^ n20887 ;
  assign n27595 = ~n22306 & n27594 ;
  assign n27596 = n27595 ^ n20887 ;
  assign n27597 = n650 & ~n27596 ;
  assign n27598 = n27597 ^ x29 ;
  assign n27600 = n27599 ^ n27598 ;
  assign n27602 = n27601 ^ n27600 ;
  assign n27645 = n27644 ^ n27602 ;
  assign n27649 = n27648 ^ n27645 ;
  assign n27587 = n12861 & ~n21025 ;
  assign n27586 = n446 & n20883 ;
  assign n27588 = n27587 ^ n27586 ;
  assign n27589 = n27588 ^ x26 ;
  assign n27585 = ~n487 & n20882 ;
  assign n27590 = n27589 ^ n27585 ;
  assign n27584 = ~n3501 & ~n22672 ;
  assign n27591 = n27590 ^ n27584 ;
  assign n27650 = n27649 ^ n27591 ;
  assign n27581 = n27389 ^ n27329 ;
  assign n27582 = ~n27394 & n27581 ;
  assign n27583 = n27582 ^ n27389 ;
  assign n27651 = n27650 ^ n27583 ;
  assign n27578 = n27408 ^ n27395 ;
  assign n27579 = n27400 & n27578 ;
  assign n27580 = n27579 ^ n27395 ;
  assign n27652 = n27651 ^ n27580 ;
  assign n27576 = ~n4496 & ~n20872 ;
  assign n27574 = n4492 & ~n22683 ;
  assign n27571 = n4504 & ~n20876 ;
  assign n27570 = n4491 & n20865 ;
  assign n27572 = n27571 ^ n27570 ;
  assign n27573 = n27572 ^ x23 ;
  assign n27575 = n27574 ^ n27573 ;
  assign n27577 = n27576 ^ n27575 ;
  assign n27653 = n27652 ^ n27577 ;
  assign n27567 = n14027 & n20861 ;
  assign n27560 = n20836 ^ x20 ;
  assign n27561 = n27560 ^ x19 ;
  assign n27562 = n27561 ^ n20836 ;
  assign n27563 = ~n26327 & n27562 ;
  assign n27564 = n27563 ^ n20836 ;
  assign n27565 = n4678 & n27564 ;
  assign n27566 = n27565 ^ x20 ;
  assign n27568 = n27567 ^ n27566 ;
  assign n27559 = n4916 & n20852 ;
  assign n27569 = n27568 ^ n27559 ;
  assign n27654 = n27653 ^ n27569 ;
  assign n27556 = n27426 ^ n27409 ;
  assign n27557 = ~n27414 & n27556 ;
  assign n27558 = n27557 ^ n27409 ;
  assign n27655 = n27654 ^ n27558 ;
  assign n27656 = n27655 ^ x17 ;
  assign n27658 = n27657 ^ n27656 ;
  assign n27660 = n27659 ^ n27658 ;
  assign n27662 = n27661 ^ n27660 ;
  assign n27555 = n20731 & n20837 ;
  assign n27663 = n27662 ^ n27555 ;
  assign n27667 = n27666 ^ n27663 ;
  assign n27534 = ~n6072 & ~n24700 ;
  assign n27533 = ~n6074 & ~n24980 ;
  assign n27535 = n27534 ^ n27533 ;
  assign n27536 = n27535 ^ n6060 ;
  assign n27537 = n27536 ^ x14 ;
  assign n27547 = n6063 & n25008 ;
  assign n27538 = n27535 ^ n6062 ;
  assign n27539 = n25896 ^ n25043 ;
  assign n27542 = n25043 ^ x13 ;
  assign n27543 = n27542 ^ n25043 ;
  assign n27544 = ~n27539 & ~n27543 ;
  assign n27545 = n27544 ^ n25043 ;
  assign n27546 = n27538 & ~n27545 ;
  assign n27548 = n27547 ^ n27546 ;
  assign n27549 = ~n27537 & ~n27548 ;
  assign n27551 = n27549 ^ n27441 ;
  assign n27550 = n27549 ^ n27471 ;
  assign n27552 = n27551 ^ n27550 ;
  assign n27553 = ~n27446 & n27552 ;
  assign n27554 = n27553 ^ n27551 ;
  assign n27668 = n27667 ^ n27554 ;
  assign n27529 = n27482 ^ n27313 ;
  assign n27530 = n27483 & ~n27529 ;
  assign n27531 = n27530 ^ x8 ;
  assign n27526 = n27481 ^ n27316 ;
  assign n27527 = ~n27473 & n27526 ;
  assign n27528 = n27527 ^ n27481 ;
  assign n27532 = n27531 ^ n27528 ;
  assign n27669 = n27668 ^ n27532 ;
  assign n27503 = n27266 & n27300 ;
  assign n27502 = n27300 ^ n27266 ;
  assign n27504 = n27503 ^ n27502 ;
  assign n27505 = n27504 ^ n27484 ;
  assign n27507 = n27268 ^ n27263 ;
  assign n27510 = n27507 ^ n27266 ;
  assign n27511 = ~n27502 & n27510 ;
  assign n27506 = ~n27263 & n27268 ;
  assign n27512 = n27511 ^ n27506 ;
  assign n27513 = n27505 & n27512 ;
  assign n27514 = n27513 ^ n27484 ;
  assign n27518 = n27502 ^ n27484 ;
  assign n27519 = ~n27506 & ~n27518 ;
  assign n27515 = n27506 ^ n27484 ;
  assign n27508 = n27507 ^ n27506 ;
  assign n27516 = n27515 ^ n27508 ;
  assign n27517 = ~n27503 & n27516 ;
  assign n27520 = n27519 ^ n27517 ;
  assign n27521 = ~n27281 & n27520 ;
  assign n27522 = ~n27279 & n27521 ;
  assign n27523 = ~n27296 & n27522 ;
  assign n27524 = n27514 & ~n27523 ;
  assign n27497 = n6655 ^ n6650 ;
  assign n27498 = n27497 ^ n27101 ;
  assign n27499 = n25287 & n27498 ;
  assign n27500 = n27499 ^ n27476 ;
  assign n27496 = n15413 & n25725 ;
  assign n27501 = n27500 ^ n27496 ;
  assign n27525 = n27524 ^ n27501 ;
  assign n27670 = n27669 ^ n27525 ;
  assign n27674 = n27673 ^ n27670 ;
  assign n27819 = n27669 ^ n27524 ;
  assign n27820 = ~n27525 & ~n27819 ;
  assign n27813 = n27667 ^ n27549 ;
  assign n27814 = n27554 & n27813 ;
  assign n27815 = n27814 ^ n27549 ;
  assign n27816 = n27815 ^ x11 ;
  assign n27812 = n6655 & n25703 ;
  assign n27817 = n27816 ^ n27812 ;
  assign n27804 = n4916 & n20836 ;
  assign n27797 = n20837 ^ x20 ;
  assign n27798 = n27797 ^ x19 ;
  assign n27799 = n27798 ^ n20837 ;
  assign n27800 = ~n21061 & n27799 ;
  assign n27801 = n27800 ^ n20837 ;
  assign n27802 = n4678 & n27801 ;
  assign n27803 = n27802 ^ x20 ;
  assign n27805 = n27804 ^ n27803 ;
  assign n27796 = n14027 & n20852 ;
  assign n27806 = n27805 ^ n27796 ;
  assign n27786 = n27591 ^ n27583 ;
  assign n27787 = ~n27650 & ~n27786 ;
  assign n27788 = n27787 ^ n27591 ;
  assign n27779 = n27643 ^ n27624 ;
  assign n27780 = ~n27629 & n27779 ;
  assign n27781 = n27780 ^ n27624 ;
  assign n27772 = x31 & ~n27612 ;
  assign n27773 = n33 & ~n20898 ;
  assign n27774 = n27772 & ~n27773 ;
  assign n27775 = n3520 & n21966 ;
  assign n27776 = n27774 & ~n27775 ;
  assign n23206 = n20898 ^ n20897 ;
  assign n27769 = ~n35 & n23206 ;
  assign n27770 = n27769 ^ n20897 ;
  assign n27771 = ~n3514 & n27770 ;
  assign n27777 = n27776 ^ n27771 ;
  assign n27760 = n13759 ^ n4740 ;
  assign n27757 = n13885 ^ n1272 ;
  assign n27756 = n27197 ^ n1399 ;
  assign n27758 = n27757 ^ n27756 ;
  assign n27754 = n945 ^ n239 ;
  assign n27752 = n4786 ^ n244 ;
  assign n27753 = n27752 ^ n841 ;
  assign n27755 = n27754 ^ n27753 ;
  assign n27759 = n27758 ^ n27755 ;
  assign n27761 = n27760 ^ n27759 ;
  assign n27762 = n27761 ^ n4202 ;
  assign n27763 = n27762 ^ n822 ;
  assign n27764 = ~n2363 & ~n27763 ;
  assign n27749 = n27205 ^ x8 ;
  assign n27750 = ~n27642 & n27749 ;
  assign n27751 = n27750 ^ x8 ;
  assign n27765 = n27764 ^ n27751 ;
  assign n27778 = n27777 ^ n27765 ;
  assign n27782 = n27781 ^ n27778 ;
  assign n27746 = n3484 & ~n20887 ;
  assign n27739 = n22415 ^ x29 ;
  assign n27740 = n27739 ^ x28 ;
  assign n27741 = n27740 ^ n22415 ;
  assign n27742 = ~n23652 & ~n27741 ;
  assign n27743 = n27742 ^ n22415 ;
  assign n27744 = n650 & n27743 ;
  assign n27745 = n27744 ^ x29 ;
  assign n27747 = n27746 ^ n27745 ;
  assign n27738 = n831 & ~n20894 ;
  assign n27748 = n27747 ^ n27738 ;
  assign n27783 = n27782 ^ n27748 ;
  assign n27735 = n27648 ^ n27602 ;
  assign n27736 = ~n27645 & ~n27735 ;
  assign n27737 = n27736 ^ n27648 ;
  assign n27784 = n27783 ^ n27737 ;
  assign n27723 = n12861 & n20883 ;
  assign n27722 = n446 & n20882 ;
  assign n27724 = n27723 ^ n27722 ;
  assign n27725 = n27724 ^ n65 ;
  assign n27726 = n27724 ^ x26 ;
  assign n27730 = n27726 ^ n67 ;
  assign n27731 = ~x25 & ~n23009 ;
  assign n27732 = n27730 & n27731 ;
  assign n27728 = n67 & n23010 ;
  assign n27727 = n20876 & n27726 ;
  assign n27729 = n27728 ^ n27727 ;
  assign n27733 = n27732 ^ n27729 ;
  assign n27734 = ~n27725 & ~n27733 ;
  assign n27785 = n27784 ^ n27734 ;
  assign n27789 = n27788 ^ n27785 ;
  assign n27717 = n4504 & ~n20872 ;
  assign n27716 = n4491 & n20861 ;
  assign n27718 = n27717 ^ n27716 ;
  assign n27719 = n27718 ^ x23 ;
  assign n27715 = n4492 & ~n23640 ;
  assign n27720 = n27719 ^ n27715 ;
  assign n27714 = ~n4496 & n20865 ;
  assign n27721 = n27720 ^ n27714 ;
  assign n27790 = n27789 ^ n27721 ;
  assign n27791 = n27790 ^ n27580 ;
  assign n27792 = n27791 ^ n27577 ;
  assign n27793 = n27792 ^ n27790 ;
  assign n27794 = n27652 & n27793 ;
  assign n27795 = n27794 ^ n27791 ;
  assign n27807 = n27806 ^ n27795 ;
  assign n27711 = n27569 ^ n27558 ;
  assign n27712 = n27654 & n27711 ;
  assign n27713 = n27712 ^ n27569 ;
  assign n27808 = n27807 ^ n27713 ;
  assign n27709 = n20731 & n20834 ;
  assign n27707 = n5703 & n25320 ;
  assign n27704 = n5702 & ~n24700 ;
  assign n27703 = n5700 & n24079 ;
  assign n27705 = n27704 ^ n27703 ;
  assign n27706 = n27705 ^ x17 ;
  assign n27708 = n27707 ^ n27706 ;
  assign n27710 = n27709 ^ n27708 ;
  assign n27809 = n27808 ^ n27710 ;
  assign n27700 = n27666 ^ n27655 ;
  assign n27701 = ~n27663 & ~n27700 ;
  assign n27702 = n27701 ^ n27666 ;
  assign n27810 = n27809 ^ n27702 ;
  assign n27679 = ~n6072 & ~n24980 ;
  assign n27678 = ~n6074 & n25043 ;
  assign n27680 = n27679 ^ n27678 ;
  assign n27681 = n27680 ^ n6060 ;
  assign n27682 = n27681 ^ x14 ;
  assign n27685 = n25287 ^ n6063 ;
  assign n27686 = n27685 ^ x13 ;
  assign n27687 = n27686 ^ n25287 ;
  assign n27692 = ~n25304 & ~n27687 ;
  assign n27693 = ~x13 & n27692 ;
  assign n27696 = n27693 ^ n27692 ;
  assign n27683 = n27680 ^ x14 ;
  assign n27684 = n27683 ^ n6063 ;
  assign n27688 = n27687 ^ n27684 ;
  assign n27690 = n27688 ^ n27687 ;
  assign n27694 = n27693 ^ n25287 ;
  assign n27695 = n27690 & n27694 ;
  assign n27697 = n27696 ^ n27695 ;
  assign n27698 = n27697 ^ n6063 ;
  assign n27699 = ~n27682 & ~n27698 ;
  assign n27811 = n27810 ^ n27699 ;
  assign n27818 = n27817 ^ n27811 ;
  assign n27821 = n27820 ^ n27818 ;
  assign n27676 = n27668 ^ n27531 ;
  assign n27677 = ~n27532 & n27676 ;
  assign n27822 = n27821 ^ n27677 ;
  assign n27675 = ~n27670 & n27673 ;
  assign n27823 = n27822 ^ n27675 ;
  assign n27992 = n27675 & n27822 ;
  assign n27985 = n16242 & n25693 ;
  assign n27983 = ~n6072 & ~n25043 ;
  assign n27980 = n8464 ^ n4898 ;
  assign n27979 = ~n6074 & n25287 ;
  assign n27981 = n27980 ^ n27979 ;
  assign n27977 = n4897 & ~n4899 ;
  assign n27978 = n25703 & n27977 ;
  assign n27982 = n27981 ^ n27978 ;
  assign n27984 = n27983 ^ n27982 ;
  assign n27986 = n27985 ^ n27984 ;
  assign n27974 = n25693 ^ n8434 ;
  assign n27975 = n8434 ^ x14 ;
  assign n27976 = ~n27974 & n27975 ;
  assign n27987 = n27986 ^ n27976 ;
  assign n27965 = n5700 & ~n24700 ;
  assign n27958 = n24980 ^ x17 ;
  assign n27959 = n27958 ^ x16 ;
  assign n27960 = n27959 ^ n24980 ;
  assign n27961 = ~n25518 & n27960 ;
  assign n27962 = n27961 ^ n24980 ;
  assign n27963 = n5693 & ~n27962 ;
  assign n27964 = n27963 ^ x17 ;
  assign n27966 = n27965 ^ n27964 ;
  assign n27957 = n20731 & n24079 ;
  assign n27967 = n27966 ^ n27957 ;
  assign n27948 = n4916 & n20837 ;
  assign n27941 = n20834 ^ x20 ;
  assign n27942 = n27941 ^ x19 ;
  assign n27943 = n27942 ^ n20834 ;
  assign n27944 = ~n21055 & n27943 ;
  assign n27945 = n27944 ^ n20834 ;
  assign n27946 = n4678 & n27945 ;
  assign n27947 = n27946 ^ x20 ;
  assign n27949 = n27948 ^ n27947 ;
  assign n27940 = n14027 & n20836 ;
  assign n27950 = n27949 ^ n27940 ;
  assign n27932 = ~n4496 & n20861 ;
  assign n27930 = n4492 & ~n23825 ;
  assign n27927 = n4504 & n20865 ;
  assign n27926 = n4491 & n20852 ;
  assign n27928 = n27927 ^ n27926 ;
  assign n27929 = n27928 ^ x23 ;
  assign n27931 = n27930 ^ n27929 ;
  assign n27933 = n27932 ^ n27931 ;
  assign n27915 = n446 & ~n20876 ;
  assign n27914 = n12861 & n20882 ;
  assign n27916 = n27915 ^ n27914 ;
  assign n27917 = n27916 ^ x26 ;
  assign n27913 = ~n487 & ~n20872 ;
  assign n27918 = n27917 ^ n27913 ;
  assign n27912 = ~n3501 & n23033 ;
  assign n27919 = n27918 ^ n27912 ;
  assign n27891 = ~n35 & n20897 ;
  assign n27889 = ~n3520 & n20894 ;
  assign n27888 = n20894 ^ n3520 ;
  assign n27890 = n27889 ^ n27888 ;
  assign n27892 = n27891 ^ n27890 ;
  assign n27902 = n27892 ^ n21954 ;
  assign n27895 = n21954 ^ n20897 ;
  assign n27894 = n21954 ^ n20898 ;
  assign n27896 = n27895 ^ n27894 ;
  assign n27899 = x30 & n27896 ;
  assign n27900 = n27899 ^ n27895 ;
  assign n27901 = ~n3520 & n27900 ;
  assign n27903 = n27902 ^ n27901 ;
  assign n27904 = x31 & n27903 ;
  assign n27883 = n14561 ^ n13223 ;
  assign n27880 = n4130 ^ n2618 ;
  assign n27879 = n4751 ^ n1968 ;
  assign n27881 = n27880 ^ n27879 ;
  assign n27877 = n13846 ^ n1060 ;
  assign n27874 = n1899 ^ n918 ;
  assign n27875 = n27874 ^ n1652 ;
  assign n27872 = n1254 ^ n192 ;
  assign n27873 = n27872 ^ n202 ;
  assign n27876 = n27875 ^ n27873 ;
  assign n27878 = n27877 ^ n27876 ;
  assign n27882 = n27881 ^ n27878 ;
  assign n27884 = n27883 ^ n27882 ;
  assign n27885 = ~n27190 & ~n27884 ;
  assign n27886 = ~n5089 & n27885 ;
  assign n27870 = n27777 ^ n27751 ;
  assign n27871 = ~n27765 & n27870 ;
  assign n27887 = n27886 ^ n27871 ;
  assign n27893 = n27892 ^ n27887 ;
  assign n27905 = n27904 ^ n27893 ;
  assign n27867 = n3484 & ~n21025 ;
  assign n27860 = n20883 ^ x29 ;
  assign n27861 = n27860 ^ x28 ;
  assign n27862 = n27861 ^ n20883 ;
  assign n27863 = ~n22545 & n27862 ;
  assign n27864 = n27863 ^ n20883 ;
  assign n27865 = n650 & n27864 ;
  assign n27866 = n27865 ^ x29 ;
  assign n27868 = n27867 ^ n27866 ;
  assign n27858 = n831 & ~n20887 ;
  assign n27869 = n27868 ^ n27858 ;
  assign n27906 = n27905 ^ n27869 ;
  assign n27907 = n27906 ^ n27781 ;
  assign n27908 = n27907 ^ n27748 ;
  assign n27909 = n27908 ^ n27906 ;
  assign n27910 = n27782 & ~n27909 ;
  assign n27911 = n27910 ^ n27907 ;
  assign n27920 = n27919 ^ n27911 ;
  assign n27921 = n27920 ^ n27734 ;
  assign n27922 = n27921 ^ n27920 ;
  assign n27923 = n27922 ^ n27737 ;
  assign n27924 = n27784 & n27923 ;
  assign n27925 = n27924 ^ n27921 ;
  assign n27934 = n27933 ^ n27925 ;
  assign n27935 = n27934 ^ n27788 ;
  assign n27936 = n27935 ^ n27721 ;
  assign n27937 = n27936 ^ n27934 ;
  assign n27938 = n27789 & n27937 ;
  assign n27939 = n27938 ^ n27935 ;
  assign n27951 = n27950 ^ n27939 ;
  assign n27953 = n27951 ^ n27790 ;
  assign n27952 = n27951 ^ n27806 ;
  assign n27954 = n27953 ^ n27952 ;
  assign n27955 = n27795 & n27954 ;
  assign n27956 = n27955 ^ n27953 ;
  assign n27968 = n27967 ^ n27956 ;
  assign n27969 = n27968 ^ n27710 ;
  assign n27970 = n27969 ^ n27968 ;
  assign n27971 = n27970 ^ n27713 ;
  assign n27972 = ~n27808 & n27971 ;
  assign n27973 = n27972 ^ n27969 ;
  assign n27988 = n27987 ^ n27973 ;
  assign n27989 = n27988 ^ x11 ;
  assign n27854 = n27702 ^ n27699 ;
  assign n27855 = n27810 & n27854 ;
  assign n27856 = n27855 ^ n27699 ;
  assign n27851 = n27815 ^ n27811 ;
  assign n27852 = ~n27817 & ~n27851 ;
  assign n27853 = n27852 ^ n27815 ;
  assign n27857 = n27856 ^ n27853 ;
  assign n27990 = n27989 ^ n27857 ;
  assign n27832 = n27818 ^ n27676 ;
  assign n27824 = n27676 ^ n27528 ;
  assign n27825 = n27676 ^ n27524 ;
  assign n27826 = n27825 ^ n27676 ;
  assign n27827 = n27676 ^ n27501 ;
  assign n27828 = n27827 ^ n27676 ;
  assign n27829 = ~n27826 & ~n27828 ;
  assign n27830 = n27829 ^ n27676 ;
  assign n27831 = ~n27824 & n27830 ;
  assign n27833 = n27832 ^ n27831 ;
  assign n27834 = n27831 ^ n27531 ;
  assign n27835 = n27834 ^ n27831 ;
  assign n27838 = n27676 & ~n27835 ;
  assign n27839 = n27838 ^ n27831 ;
  assign n27840 = n27833 & n27839 ;
  assign n27841 = n27840 ^ n27818 ;
  assign n27842 = n27501 & n27841 ;
  assign n27843 = n27524 & n27818 ;
  assign n27844 = n27668 ^ n27528 ;
  assign n27845 = n27532 & ~n27844 ;
  assign n27846 = n27845 ^ n27528 ;
  assign n27847 = n27843 & ~n27846 ;
  assign n27848 = n27847 ^ n27524 ;
  assign n27849 = n27842 & n27848 ;
  assign n27850 = n27849 ^ n27841 ;
  assign n27991 = n27990 ^ n27850 ;
  assign n27993 = n27992 ^ n27991 ;
  assign n28135 = ~n27991 & n27992 ;
  assign n28126 = n14027 & n20837 ;
  assign n28124 = n4916 & n20834 ;
  assign n28119 = n27950 ^ n27934 ;
  assign n28120 = ~n27939 & ~n28119 ;
  assign n28121 = n28120 ^ n27934 ;
  assign n28122 = n28121 ^ x20 ;
  assign n28113 = n25245 ^ n24079 ;
  assign n28114 = n24079 ^ n4685 ;
  assign n28115 = n28114 ^ n24079 ;
  assign n28116 = ~n28113 & n28115 ;
  assign n28117 = n28116 ^ n24079 ;
  assign n28118 = n4678 & n28117 ;
  assign n28123 = n28122 ^ n28118 ;
  assign n28125 = n28124 ^ n28123 ;
  assign n28127 = n28126 ^ n28125 ;
  assign n28107 = n27919 ^ n27906 ;
  assign n28108 = n27911 & ~n28107 ;
  assign n28109 = n28108 ^ n27906 ;
  assign n28104 = ~n487 & n20865 ;
  assign n28102 = n12861 & ~n20876 ;
  assign n28100 = n446 & ~n20872 ;
  assign n28088 = n27751 & ~n27777 ;
  assign n28093 = n28088 ^ n27870 ;
  assign n28094 = ~n27886 & n28093 ;
  assign n28089 = n27886 & n28088 ;
  assign n28095 = n28094 ^ n28089 ;
  assign n28096 = ~n27764 & n28095 ;
  assign n28078 = n5110 ^ n2642 ;
  assign n28076 = n2432 ^ n1191 ;
  assign n28074 = n12551 ^ n499 ;
  assign n28073 = n27346 ^ n621 ;
  assign n28075 = n28074 ^ n28073 ;
  assign n28077 = n28076 ^ n28075 ;
  assign n28079 = n28078 ^ n28077 ;
  assign n28080 = n28079 ^ n2027 ;
  assign n28081 = n28080 ^ n2094 ;
  assign n28083 = n12321 ^ n193 ;
  assign n28082 = n5129 ^ n987 ;
  assign n28084 = n28083 ^ n28082 ;
  assign n28085 = n28084 ^ n1092 ;
  assign n28086 = ~n28081 & ~n28085 ;
  assign n28087 = n28086 ^ x11 ;
  assign n28090 = n28089 ^ n28087 ;
  assign n28071 = x31 & n27891 ;
  assign n28069 = ~n35 & ~n20894 ;
  assign n28067 = n12533 & ~n27889 ;
  assign n28064 = x31 & ~n22306 ;
  assign n28065 = n28064 ^ n20887 ;
  assign n28066 = n3520 & n28065 ;
  assign n28068 = n28067 ^ n28066 ;
  assign n28070 = n28069 ^ n28068 ;
  assign n28072 = n28071 ^ n28070 ;
  assign n28091 = n28090 ^ n28072 ;
  assign n28057 = n27887 ^ n27869 ;
  assign n28058 = ~n27905 & ~n28057 ;
  assign n28059 = n28058 ^ n27887 ;
  assign n28092 = n28091 ^ n28059 ;
  assign n28097 = n28096 ^ n28092 ;
  assign n28055 = n3484 & n20883 ;
  assign n28051 = n831 & ~n21025 ;
  assign n28050 = n653 & ~n22671 ;
  assign n28052 = n28051 ^ n28050 ;
  assign n28053 = n28052 ^ x29 ;
  assign n28047 = ~x28 & ~n22671 ;
  assign n28048 = n28047 ^ n20882 ;
  assign n28049 = n650 & n28048 ;
  assign n28054 = n28053 ^ n28049 ;
  assign n28056 = n28055 ^ n28054 ;
  assign n28098 = n28097 ^ n28056 ;
  assign n28099 = n28098 ^ x26 ;
  assign n28101 = n28100 ^ n28099 ;
  assign n28103 = n28102 ^ n28101 ;
  assign n28105 = n28104 ^ n28103 ;
  assign n28044 = ~n3501 & ~n22683 ;
  assign n28106 = n28105 ^ n28044 ;
  assign n28110 = n28109 ^ n28106 ;
  assign n28039 = n4504 & n20861 ;
  assign n28038 = n4491 & n20836 ;
  assign n28040 = n28039 ^ n28038 ;
  assign n28041 = n28040 ^ x23 ;
  assign n28037 = n4492 & ~n24433 ;
  assign n28042 = n28041 ^ n28037 ;
  assign n28036 = ~n4496 & n20852 ;
  assign n28043 = n28042 ^ n28036 ;
  assign n28111 = n28110 ^ n28043 ;
  assign n28033 = n27933 ^ n27920 ;
  assign n28034 = ~n27925 & n28033 ;
  assign n28035 = n28034 ^ n27920 ;
  assign n28112 = n28111 ^ n28035 ;
  assign n28128 = n28127 ^ n28112 ;
  assign n28031 = n20731 & ~n24700 ;
  assign n28029 = n5703 & ~n25896 ;
  assign n28026 = n5700 & ~n24980 ;
  assign n28025 = n5702 & n25043 ;
  assign n28027 = n28026 ^ n28025 ;
  assign n28028 = n28027 ^ x17 ;
  assign n28030 = n28029 ^ n28028 ;
  assign n28032 = n28031 ^ n28030 ;
  assign n28129 = n28128 ^ n28032 ;
  assign n28022 = n27967 ^ n27951 ;
  assign n28023 = ~n27956 & ~n28022 ;
  assign n28024 = n28023 ^ n27951 ;
  assign n28130 = n28129 ^ n28024 ;
  assign n28004 = n25287 ^ x13 ;
  assign n28013 = ~n4898 & n28004 ;
  assign n28006 = n25043 ^ x14 ;
  assign n28014 = n25287 & n28006 ;
  assign n28015 = n28014 ^ x14 ;
  assign n28016 = n28013 & ~n28015 ;
  assign n28005 = n4896 & ~n28004 ;
  assign n28009 = ~n25287 & ~n28006 ;
  assign n28010 = n28009 ^ n25043 ;
  assign n28011 = n28005 & ~n28010 ;
  assign n28012 = n28011 ^ x14 ;
  assign n28017 = n28016 ^ n28012 ;
  assign n28018 = n28017 ^ x13 ;
  assign n28019 = n4897 & n25725 ;
  assign n28020 = n28018 & n28019 ;
  assign n28021 = n28020 ^ n28017 ;
  assign n28131 = n28130 ^ n28021 ;
  assign n28001 = n27987 ^ n27968 ;
  assign n28002 = ~n27973 & n28001 ;
  assign n28003 = n28002 ^ n27968 ;
  assign n28132 = n28131 ^ n28003 ;
  assign n27997 = n27856 ^ x11 ;
  assign n27998 = n27988 ^ n27856 ;
  assign n27994 = n27853 ^ n27850 ;
  assign n27999 = n27998 ^ n27994 ;
  assign n28000 = n27997 & ~n27999 ;
  assign n28133 = n28132 ^ n28000 ;
  assign n27995 = n27988 ^ n27850 ;
  assign n27996 = ~n27994 & n27995 ;
  assign n28134 = n28133 ^ n27996 ;
  assign n28136 = n28135 ^ n28134 ;
  assign n28281 = ~n6072 & n25703 ;
  assign n28273 = ~n4496 & n20836 ;
  assign n28271 = n4492 & ~n24427 ;
  assign n28268 = n4504 & n20852 ;
  assign n28267 = n4491 & n20837 ;
  assign n28269 = n28268 ^ n28267 ;
  assign n28270 = n28269 ^ x23 ;
  assign n28272 = n28271 ^ n28270 ;
  assign n28274 = n28273 ^ n28272 ;
  assign n28257 = n28059 ^ n28056 ;
  assign n28258 = ~n28097 & ~n28257 ;
  assign n28259 = n28258 ^ n28056 ;
  assign n28246 = n28094 ^ n28072 ;
  assign n28244 = n28087 ^ n28072 ;
  assign n28245 = ~n28095 & n28244 ;
  assign n28247 = n28246 ^ n28245 ;
  assign n28248 = n28087 ^ n27764 ;
  assign n28249 = n28248 ^ n28072 ;
  assign n28250 = n28247 & ~n28249 ;
  assign n28251 = n28250 ^ n28072 ;
  assign n28238 = n28086 ^ n27764 ;
  assign n28239 = n27764 ^ x11 ;
  assign n28240 = ~n28238 & n28239 ;
  assign n28241 = n28240 ^ x11 ;
  assign n28226 = n3116 ^ n765 ;
  assign n28225 = n4311 ^ n1311 ;
  assign n28227 = n28226 ^ n28225 ;
  assign n28228 = n28227 ^ n13039 ;
  assign n28229 = n28228 ^ n14574 ;
  assign n28231 = n2069 ^ n819 ;
  assign n28232 = n28231 ^ n736 ;
  assign n28230 = n2132 ^ n332 ;
  assign n28233 = n28232 ^ n28230 ;
  assign n28234 = n28233 ^ n26203 ;
  assign n28235 = n28234 ^ n25799 ;
  assign n28236 = n28235 ^ n12420 ;
  assign n28237 = ~n28229 & ~n28236 ;
  assign n28242 = n28241 ^ n28237 ;
  assign n28222 = ~n3724 & ~n20887 ;
  assign n28221 = n3726 & ~n21025 ;
  assign n28223 = n28222 ^ n28221 ;
  assign n28212 = n22415 ^ n20887 ;
  assign n28211 = n22415 ^ n20894 ;
  assign n28213 = n28212 ^ n28211 ;
  assign n28216 = x30 & n28213 ;
  assign n28217 = n28216 ^ n28212 ;
  assign n28218 = ~n3520 & ~n28217 ;
  assign n28219 = n28218 ^ n22415 ;
  assign n28220 = x31 & n28219 ;
  assign n28224 = n28223 ^ n28220 ;
  assign n28243 = n28242 ^ n28224 ;
  assign n28255 = n28251 ^ n28243 ;
  assign n28208 = n3484 & n20882 ;
  assign n28201 = n20876 ^ x29 ;
  assign n28202 = n28201 ^ x28 ;
  assign n28203 = n28202 ^ n20876 ;
  assign n28204 = ~n25359 & n28203 ;
  assign n28205 = n28204 ^ n20876 ;
  assign n28206 = n650 & ~n28205 ;
  assign n28207 = n28206 ^ x29 ;
  assign n28209 = n28208 ^ n28207 ;
  assign n28200 = n831 & n20883 ;
  assign n28210 = n28209 ^ n28200 ;
  assign n28256 = n28255 ^ n28210 ;
  assign n28260 = n28259 ^ n28256 ;
  assign n28195 = n12861 & ~n20872 ;
  assign n28194 = n446 & n20865 ;
  assign n28196 = n28195 ^ n28194 ;
  assign n28197 = n28196 ^ x26 ;
  assign n28193 = ~n487 & n20861 ;
  assign n28198 = n28197 ^ n28193 ;
  assign n28192 = ~n3501 & ~n23640 ;
  assign n28199 = n28198 ^ n28192 ;
  assign n28261 = n28260 ^ n28199 ;
  assign n28262 = n28261 ^ n28109 ;
  assign n28263 = n28262 ^ n28098 ;
  assign n28264 = n28263 ^ n28261 ;
  assign n28265 = ~n28106 & ~n28264 ;
  assign n28266 = n28265 ^ n28262 ;
  assign n28275 = n28274 ^ n28266 ;
  assign n28189 = n28043 ^ n28035 ;
  assign n28190 = ~n28111 & n28189 ;
  assign n28191 = n28190 ^ n28043 ;
  assign n28276 = n28275 ^ n28191 ;
  assign n28186 = n4916 & n24079 ;
  assign n28178 = n25320 ^ n24700 ;
  assign n28179 = n24700 ^ x20 ;
  assign n28180 = n28179 ^ x19 ;
  assign n28181 = n28180 ^ n24700 ;
  assign n28182 = ~n28178 & n28181 ;
  assign n28183 = n28182 ^ n24700 ;
  assign n28184 = n4678 & ~n28183 ;
  assign n28185 = n28184 ^ x20 ;
  assign n28187 = n28186 ^ n28185 ;
  assign n28177 = n14027 & n20834 ;
  assign n28188 = n28187 ^ n28177 ;
  assign n28277 = n28276 ^ n28188 ;
  assign n28174 = n28121 ^ n28112 ;
  assign n28175 = ~n28127 & n28174 ;
  assign n28176 = n28175 ^ n28121 ;
  assign n28278 = n28277 ^ n28176 ;
  assign n28171 = n5703 & n25937 ;
  assign n28169 = n20731 & ~n24980 ;
  assign n28167 = n5700 & n25043 ;
  assign n28168 = n28167 ^ x17 ;
  assign n28170 = n28169 ^ n28168 ;
  assign n28172 = n28171 ^ n28170 ;
  assign n28166 = n5702 & ~n25287 ;
  assign n28173 = n28172 ^ n28166 ;
  assign n28279 = n28278 ^ n28173 ;
  assign n28280 = n28279 ^ x14 ;
  assign n28282 = n28281 ^ n28280 ;
  assign n28163 = n28032 ^ n28024 ;
  assign n28164 = n28129 & ~n28163 ;
  assign n28165 = n28164 ^ n28032 ;
  assign n28283 = n28282 ^ n28165 ;
  assign n28160 = n28021 ^ n28003 ;
  assign n28161 = ~n28131 & ~n28160 ;
  assign n28162 = n28161 ^ n28021 ;
  assign n28284 = n28283 ^ n28162 ;
  assign n28138 = n27850 & ~n27988 ;
  assign n28139 = n28138 ^ n27995 ;
  assign n28140 = n28138 ^ n28132 ;
  assign n28142 = n28138 ^ x11 ;
  assign n28141 = n28138 ^ n27853 ;
  assign n28143 = n28142 ^ n28141 ;
  assign n28144 = n28142 ^ n27857 ;
  assign n28145 = n28144 ^ n28142 ;
  assign n28146 = ~n28143 & ~n28145 ;
  assign n28147 = n28146 ^ n28142 ;
  assign n28148 = ~n28140 & n28147 ;
  assign n28149 = n28148 ^ n28132 ;
  assign n28150 = n28132 ^ n27856 ;
  assign n28151 = n28132 ^ n27853 ;
  assign n28152 = n28132 ^ x11 ;
  assign n28153 = ~n28151 & n28152 ;
  assign n28154 = ~n28150 & n28153 ;
  assign n28155 = n28154 ^ n28150 ;
  assign n28156 = n28155 ^ n27856 ;
  assign n28157 = n28149 & ~n28156 ;
  assign n28158 = ~n28139 & n28157 ;
  assign n28159 = n28158 ^ n28149 ;
  assign n28285 = n28284 ^ n28159 ;
  assign n28137 = ~n28134 & n28135 ;
  assign n28286 = n28285 ^ n28137 ;
  assign n28414 = n28162 ^ n28159 ;
  assign n28415 = n28284 & n28414 ;
  assign n28416 = n28415 ^ n28159 ;
  assign n28409 = n28176 ^ n28173 ;
  assign n28410 = n28278 & ~n28409 ;
  assign n28411 = n28410 ^ n28173 ;
  assign n28404 = n5703 & n25693 ;
  assign n28403 = n5700 ^ x17 ;
  assign n28405 = n28404 ^ n28403 ;
  assign n28402 = n20731 & n25043 ;
  assign n28406 = n28405 ^ n28402 ;
  assign n28395 = n5702 ^ n5700 ;
  assign n28396 = n28395 ^ n5700 ;
  assign n28399 = ~n25043 & n28396 ;
  assign n28400 = n28399 ^ n5700 ;
  assign n28401 = n25287 & n28400 ;
  assign n28407 = n28406 ^ n28401 ;
  assign n28386 = n4916 & ~n24700 ;
  assign n28379 = n24980 ^ x20 ;
  assign n28380 = n28379 ^ x19 ;
  assign n28381 = n28380 ^ n24980 ;
  assign n28382 = ~n25518 & n28381 ;
  assign n28383 = n28382 ^ n24980 ;
  assign n28384 = n4678 & ~n28383 ;
  assign n28385 = n28384 ^ x20 ;
  assign n28387 = n28386 ^ n28385 ;
  assign n28378 = n14027 & n24079 ;
  assign n28388 = n28387 ^ n28378 ;
  assign n28369 = ~n4496 & n20837 ;
  assign n28362 = n20834 ^ x23 ;
  assign n28363 = n28362 ^ x22 ;
  assign n28364 = n28363 ^ n20834 ;
  assign n28365 = ~n21055 & n28364 ;
  assign n28366 = n28365 ^ n20834 ;
  assign n28367 = n4488 & n28366 ;
  assign n28368 = n28367 ^ x23 ;
  assign n28370 = n28369 ^ n28368 ;
  assign n28361 = n4504 & n20836 ;
  assign n28371 = n28370 ^ n28361 ;
  assign n28342 = n11833 ^ n2639 ;
  assign n28340 = n12053 ^ n1250 ;
  assign n28338 = n1012 ^ n615 ;
  assign n28337 = n3063 ^ n1876 ;
  assign n28339 = n28338 ^ n28337 ;
  assign n28341 = n28340 ^ n28339 ;
  assign n28343 = n28342 ^ n28341 ;
  assign n28344 = n28343 ^ n2922 ;
  assign n28335 = n12561 ^ n3446 ;
  assign n28336 = n28335 ^ n4967 ;
  assign n28345 = n28344 ^ n28336 ;
  assign n28346 = ~n13141 & ~n28345 ;
  assign n28347 = n28346 ^ n28237 ;
  assign n28316 = n3520 & n22546 ;
  assign n28319 = x30 & ~n21025 ;
  assign n28320 = n28319 ^ n20883 ;
  assign n28321 = ~n3520 & n28320 ;
  assign n28322 = n28321 ^ n20883 ;
  assign n28323 = ~x31 & n28322 ;
  assign n28330 = n28323 ^ x31 ;
  assign n28327 = ~x29 & n23152 ;
  assign n28328 = n28327 ^ n20887 ;
  assign n28329 = n12015 & n28328 ;
  assign n28331 = n28330 ^ n28329 ;
  assign n28332 = n28331 ^ n28323 ;
  assign n28333 = n28316 & n28332 ;
  assign n28334 = n28333 ^ n28331 ;
  assign n28348 = n28347 ^ n28334 ;
  assign n28313 = n28237 & ~n28241 ;
  assign n28314 = n28313 ^ n28242 ;
  assign n28312 = n28210 & n28251 ;
  assign n28315 = n28314 ^ n28312 ;
  assign n28349 = n28348 ^ n28315 ;
  assign n28309 = n28251 ^ n28210 ;
  assign n28310 = n28309 ^ n28224 ;
  assign n28311 = ~n28243 & ~n28310 ;
  assign n28350 = n28349 ^ n28311 ;
  assign n28351 = n28350 ^ x29 ;
  assign n28304 = n20872 ^ n4536 ;
  assign n28305 = n28304 ^ n20872 ;
  assign n28306 = ~n23032 & n28305 ;
  assign n28307 = n28306 ^ n20872 ;
  assign n28308 = n650 & ~n28307 ;
  assign n28352 = n28351 ^ n28308 ;
  assign n28301 = n831 & n20882 ;
  assign n28353 = n28352 ^ n28301 ;
  assign n28300 = n3484 & ~n20876 ;
  assign n28354 = n28353 ^ n28300 ;
  assign n28295 = n12861 & n20865 ;
  assign n28294 = ~n487 & n20852 ;
  assign n28296 = n28295 ^ n28294 ;
  assign n28297 = n28296 ^ x26 ;
  assign n28293 = n446 & n20861 ;
  assign n28298 = n28297 ^ n28293 ;
  assign n28292 = ~n3501 & ~n23825 ;
  assign n28299 = n28298 ^ n28292 ;
  assign n28355 = n28354 ^ n28299 ;
  assign n28356 = n28355 ^ n28259 ;
  assign n28357 = n28356 ^ n28199 ;
  assign n28358 = n28357 ^ n28355 ;
  assign n28359 = ~n28260 & n28358 ;
  assign n28360 = n28359 ^ n28356 ;
  assign n28372 = n28371 ^ n28360 ;
  assign n28374 = n28372 ^ n28261 ;
  assign n28373 = n28372 ^ n28274 ;
  assign n28375 = n28374 ^ n28373 ;
  assign n28376 = n28266 & ~n28375 ;
  assign n28377 = n28376 ^ n28374 ;
  assign n28389 = n28388 ^ n28377 ;
  assign n28390 = n28389 ^ n28188 ;
  assign n28391 = n28390 ^ n28389 ;
  assign n28392 = n28391 ^ n28191 ;
  assign n28393 = ~n28276 & n28392 ;
  assign n28394 = n28393 ^ n28390 ;
  assign n28408 = n28407 ^ n28394 ;
  assign n28412 = n28411 ^ n28408 ;
  assign n28413 = n28412 ^ x14 ;
  assign n28417 = n28416 ^ n28413 ;
  assign n28288 = n28279 ^ n28165 ;
  assign n28289 = ~n28282 & ~n28288 ;
  assign n28290 = n28289 ^ n28279 ;
  assign n28287 = n28137 & ~n28285 ;
  assign n28291 = n28290 ^ n28287 ;
  assign n28418 = n28417 ^ n28291 ;
  assign n28573 = n28413 ^ n28290 ;
  assign n28576 = n28291 & ~n28573 ;
  assign n28574 = n28573 ^ n28287 ;
  assign n28575 = ~n28416 & n28574 ;
  assign n28577 = n28576 ^ n28575 ;
  assign n28559 = n446 & n20852 ;
  assign n28558 = n12861 & n20861 ;
  assign n28560 = n28559 ^ n28558 ;
  assign n28561 = n28560 ^ x26 ;
  assign n28557 = ~n487 & n20836 ;
  assign n28562 = n28561 ^ n28557 ;
  assign n28556 = ~n3501 & ~n24433 ;
  assign n28563 = n28562 ^ n28556 ;
  assign n28547 = n3484 & ~n20872 ;
  assign n28540 = n20865 ^ x29 ;
  assign n28541 = n28540 ^ x28 ;
  assign n28542 = n28541 ^ n20865 ;
  assign n28543 = ~n22682 & n28542 ;
  assign n28544 = n28543 ^ n20865 ;
  assign n28545 = n650 & n28544 ;
  assign n28546 = n28545 ^ x29 ;
  assign n28548 = n28547 ^ n28546 ;
  assign n28539 = n831 & ~n20876 ;
  assign n28549 = n28548 ^ n28539 ;
  assign n28529 = n13839 ^ n2953 ;
  assign n28526 = n3561 ^ n116 ;
  assign n28527 = n28526 ^ n1739 ;
  assign n28524 = n2240 ^ n90 ;
  assign n28525 = n28524 ^ n273 ;
  assign n28528 = n28527 ^ n28525 ;
  assign n28530 = n28529 ^ n28528 ;
  assign n28523 = n4802 ^ n1620 ;
  assign n28531 = n28530 ^ n28523 ;
  assign n28532 = n28531 ^ n6417 ;
  assign n28533 = n28532 ^ n13639 ;
  assign n28534 = ~n1993 & ~n28533 ;
  assign n28535 = n28534 ^ x14 ;
  assign n28520 = ~n3724 & n20883 ;
  assign n28519 = n3726 & n20882 ;
  assign n28521 = n28520 ^ n28519 ;
  assign n28510 = n22672 ^ n20883 ;
  assign n28509 = n22672 ^ n21025 ;
  assign n28511 = n28510 ^ n28509 ;
  assign n28514 = x30 & ~n28511 ;
  assign n28515 = n28514 ^ n28510 ;
  assign n28516 = ~n3520 & ~n28515 ;
  assign n28517 = n28516 ^ n22672 ;
  assign n28518 = x31 & ~n28517 ;
  assign n28522 = n28521 ^ n28518 ;
  assign n28536 = n28535 ^ n28522 ;
  assign n28480 = n28313 ^ n28210 ;
  assign n28458 = n28237 ^ n28224 ;
  assign n28459 = n28348 ^ n28241 ;
  assign n28460 = n28459 ^ n28224 ;
  assign n28461 = n28460 ^ n28348 ;
  assign n28462 = ~n28458 & ~n28461 ;
  assign n28463 = n28462 ^ n28459 ;
  assign n28465 = n28463 ^ n28312 ;
  assign n28468 = n28465 ^ n28310 ;
  assign n28481 = n28480 ^ n28468 ;
  assign n28482 = n28481 ^ n28251 ;
  assign n28487 = n28482 ^ n28468 ;
  assign n28475 = n28224 ^ n28210 ;
  assign n28476 = n28475 ^ n28224 ;
  assign n28477 = n28463 & n28476 ;
  assign n28478 = n28477 ^ n28224 ;
  assign n28479 = ~n28309 & ~n28478 ;
  assign n28484 = n28482 ^ n28463 ;
  assign n28488 = ~n28479 & n28484 ;
  assign n28489 = n28487 & n28488 ;
  assign n28483 = n28482 ^ n28313 ;
  assign n28485 = n28484 ^ n28483 ;
  assign n28486 = n28485 ^ n28479 ;
  assign n28490 = n28489 ^ n28486 ;
  assign n28470 = n28465 ^ n28309 ;
  assign n28464 = n28313 ^ n28309 ;
  assign n28466 = n28465 ^ n28464 ;
  assign n28467 = n28466 ^ n28465 ;
  assign n28469 = n28468 ^ n28467 ;
  assign n28471 = n28470 ^ n28469 ;
  assign n28472 = n28471 ^ n28463 ;
  assign n28491 = n28490 ^ n28472 ;
  assign n28492 = n28312 ^ n28242 ;
  assign n28493 = n28492 ^ n28309 ;
  assign n28494 = ~n28243 & ~n28493 ;
  assign n28495 = n28494 ^ n28242 ;
  assign n28496 = ~n28348 & n28495 ;
  assign n28497 = n28496 ^ n28348 ;
  assign n28500 = n28497 ^ n28494 ;
  assign n28501 = n28500 ^ n28497 ;
  assign n28504 = n28496 & ~n28501 ;
  assign n28505 = n28237 & n28504 ;
  assign n28506 = n28505 ^ n28237 ;
  assign n28498 = n28497 ^ n28237 ;
  assign n28507 = n28506 ^ n28498 ;
  assign n28508 = n28491 & n28507 ;
  assign n28537 = n28536 ^ n28508 ;
  assign n28456 = n28346 ^ n28334 ;
  assign n28457 = ~n28347 & n28456 ;
  assign n28538 = n28537 ^ n28457 ;
  assign n28550 = n28549 ^ n28538 ;
  assign n28551 = n28550 ^ n28350 ;
  assign n28552 = n28551 ^ n28299 ;
  assign n28553 = n28552 ^ n28550 ;
  assign n28554 = n28354 & n28553 ;
  assign n28555 = n28554 ^ n28551 ;
  assign n28564 = n28563 ^ n28555 ;
  assign n28453 = n28371 ^ n28355 ;
  assign n28454 = n28360 & n28453 ;
  assign n28455 = n28454 ^ n28355 ;
  assign n28565 = n28564 ^ n28455 ;
  assign n28448 = n4504 & n20837 ;
  assign n28447 = n4491 & n24079 ;
  assign n28449 = n28448 ^ n28447 ;
  assign n28450 = n28449 ^ x23 ;
  assign n28446 = n4492 & ~n25245 ;
  assign n28451 = n28450 ^ n28446 ;
  assign n28445 = ~n4496 & n20834 ;
  assign n28452 = n28451 ^ n28445 ;
  assign n28566 = n28565 ^ n28452 ;
  assign n28442 = n4916 & ~n24980 ;
  assign n28435 = n25043 ^ x20 ;
  assign n28436 = n28435 ^ x19 ;
  assign n28437 = n28436 ^ n25043 ;
  assign n28438 = ~n27539 & n28437 ;
  assign n28439 = n28438 ^ n25043 ;
  assign n28440 = n4678 & n28439 ;
  assign n28441 = n28440 ^ x20 ;
  assign n28443 = n28442 ^ n28441 ;
  assign n28434 = n14027 & ~n24700 ;
  assign n28444 = n28443 ^ n28434 ;
  assign n28567 = n28566 ^ n28444 ;
  assign n28431 = n28388 ^ n28372 ;
  assign n28432 = ~n28377 & n28431 ;
  assign n28433 = n28432 ^ n28372 ;
  assign n28568 = n28567 ^ n28433 ;
  assign n28428 = n20731 ^ x17 ;
  assign n28425 = n20731 ^ n5700 ;
  assign n28426 = n28425 ^ n28167 ;
  assign n28427 = n25287 & n28426 ;
  assign n28429 = n28428 ^ n28427 ;
  assign n28424 = n5703 & n25725 ;
  assign n28430 = n28429 ^ n28424 ;
  assign n28569 = n28568 ^ n28430 ;
  assign n28421 = n28407 ^ n28389 ;
  assign n28422 = ~n28394 & ~n28421 ;
  assign n28423 = n28422 ^ n28389 ;
  assign n28570 = n28569 ^ n28423 ;
  assign n28571 = n28570 ^ x14 ;
  assign n28419 = n28411 ^ x14 ;
  assign n28420 = n28412 & n28419 ;
  assign n28572 = n28571 ^ n28420 ;
  assign n28578 = n28577 ^ n28572 ;
  assign n28707 = n28573 ^ n28416 ;
  assign n28708 = n28573 ^ n28572 ;
  assign n28709 = n28707 & n28708 ;
  assign n28710 = n28287 & n28709 ;
  assign n28702 = n20731 & n25703 ;
  assign n28691 = n12861 & n20852 ;
  assign n28690 = n446 & n20836 ;
  assign n28692 = n28691 ^ n28690 ;
  assign n28693 = n28692 ^ x26 ;
  assign n28689 = ~n487 & n20837 ;
  assign n28694 = n28693 ^ n28689 ;
  assign n28688 = ~n3501 & ~n24427 ;
  assign n28695 = n28694 ^ n28688 ;
  assign n28677 = n20883 & n24214 ;
  assign n28676 = ~n3733 & n20882 ;
  assign n28678 = n28677 ^ n28676 ;
  assign n28674 = n3726 & ~n23009 ;
  assign n28673 = n3520 & n23010 ;
  assign n28675 = n28674 ^ n28673 ;
  assign n28679 = n28678 ^ n28675 ;
  assign n28655 = n28534 ^ n28237 ;
  assign n28660 = n15192 ^ n1480 ;
  assign n28661 = n28660 ^ n14344 ;
  assign n28662 = n28661 ^ n3437 ;
  assign n28657 = n1597 ^ n219 ;
  assign n28656 = n2050 ^ n1054 ;
  assign n28658 = n28657 ^ n28656 ;
  assign n28659 = n28658 ^ n24196 ;
  assign n28663 = n28662 ^ n28659 ;
  assign n28664 = n28663 ^ n5345 ;
  assign n28665 = n28664 ^ n13921 ;
  assign n28666 = n28665 ^ n5112 ;
  assign n28667 = ~n2980 & ~n28666 ;
  assign n28668 = n28667 ^ x14 ;
  assign n28669 = n28668 ^ n28534 ;
  assign n28670 = n28669 ^ n28667 ;
  assign n28671 = ~n28655 & n28670 ;
  assign n28672 = n28671 ^ n28668 ;
  assign n28680 = n28679 ^ n28672 ;
  assign n28645 = n28535 ^ n28237 ;
  assign n28646 = n28645 ^ n28522 ;
  assign n28649 = n28522 ^ n28334 ;
  assign n28650 = n28649 ^ n28535 ;
  assign n28651 = n28456 & n28650 ;
  assign n28652 = n28651 ^ n28535 ;
  assign n28653 = ~n28646 & n28652 ;
  assign n28654 = n28653 ^ n28522 ;
  assign n28681 = n28680 ^ n28654 ;
  assign n28633 = ~x28 & ~n23608 ;
  assign n28642 = n28633 ^ n23640 ;
  assign n28643 = n653 & ~n28642 ;
  assign n28638 = n831 & ~n20872 ;
  assign n28637 = n3484 & n20865 ;
  assign n28639 = n28638 ^ n28637 ;
  assign n28640 = n28639 ^ n651 ;
  assign n28634 = n28633 ^ n20861 ;
  assign n28636 = ~n28634 & n28635 ;
  assign n28641 = n28640 ^ n28636 ;
  assign n28644 = n28643 ^ n28641 ;
  assign n28682 = n28681 ^ n28644 ;
  assign n28683 = n28682 ^ n28549 ;
  assign n28684 = n28683 ^ n28682 ;
  assign n28685 = n28684 ^ n28508 ;
  assign n28686 = ~n28538 & ~n28685 ;
  assign n28687 = n28686 ^ n28683 ;
  assign n28696 = n28695 ^ n28687 ;
  assign n28630 = n28563 ^ n28550 ;
  assign n28631 = n28555 & n28630 ;
  assign n28632 = n28631 ^ n28550 ;
  assign n28697 = n28696 ^ n28632 ;
  assign n28628 = ~n4496 & n24079 ;
  assign n28626 = n4492 & n25320 ;
  assign n28623 = n4504 & n20834 ;
  assign n28622 = n4491 & ~n24700 ;
  assign n28624 = n28623 ^ n28622 ;
  assign n28625 = n28624 ^ x23 ;
  assign n28627 = n28626 ^ n28625 ;
  assign n28629 = n28628 ^ n28627 ;
  assign n28698 = n28697 ^ n28629 ;
  assign n28619 = n28455 ^ n28452 ;
  assign n28620 = n28565 & n28619 ;
  assign n28621 = n28620 ^ n28455 ;
  assign n28699 = n28698 ^ n28621 ;
  assign n28617 = n14027 & ~n24980 ;
  assign n28613 = n4683 & ~n25304 ;
  assign n28612 = n4678 & n25937 ;
  assign n28614 = n28613 ^ n28612 ;
  assign n28611 = n4916 & n25043 ;
  assign n28615 = n28614 ^ n28611 ;
  assign n28616 = n28615 ^ x20 ;
  assign n28618 = n28617 ^ n28616 ;
  assign n28700 = n28699 ^ n28618 ;
  assign n28701 = n28700 ^ x17 ;
  assign n28703 = n28702 ^ n28701 ;
  assign n28608 = n28444 ^ n28433 ;
  assign n28609 = n28567 & n28608 ;
  assign n28610 = n28609 ^ n28444 ;
  assign n28704 = n28703 ^ n28610 ;
  assign n28582 = n28408 ^ n28290 ;
  assign n28583 = n28408 ^ x14 ;
  assign n28584 = ~n28582 & ~n28583 ;
  assign n28585 = n28584 ^ x14 ;
  assign n28586 = n28570 & ~n28585 ;
  assign n28587 = n28585 ^ n28570 ;
  assign n28588 = n28587 ^ n28586 ;
  assign n28589 = ~n28411 & ~n28588 ;
  assign n28590 = n28589 ^ n28416 ;
  assign n28592 = n28416 ^ n28290 ;
  assign n28591 = n28570 ^ n28416 ;
  assign n28593 = n28592 ^ n28591 ;
  assign n28594 = n28593 ^ n28592 ;
  assign n28595 = n28594 ^ n28571 ;
  assign n28596 = n28595 ^ n28594 ;
  assign n28597 = n28594 ^ n28593 ;
  assign n28598 = n28597 ^ n28594 ;
  assign n28599 = n28594 ^ n28582 ;
  assign n28600 = n28599 ^ n28594 ;
  assign n28601 = n28598 & ~n28600 ;
  assign n28602 = ~n28596 & n28601 ;
  assign n28603 = n28602 ^ n28596 ;
  assign n28604 = n28603 ^ n28595 ;
  assign n28605 = ~n28590 & ~n28604 ;
  assign n28606 = n28605 ^ n28416 ;
  assign n28607 = ~n28586 & n28606 ;
  assign n28705 = n28704 ^ n28607 ;
  assign n28579 = n28430 ^ n28423 ;
  assign n28580 = n28569 & ~n28579 ;
  assign n28581 = n28580 ^ n28430 ;
  assign n28706 = n28705 ^ n28581 ;
  assign n28711 = n28710 ^ n28706 ;
  assign n28815 = n28700 ^ n28610 ;
  assign n28816 = ~n28703 & ~n28815 ;
  assign n28817 = n28816 ^ n28700 ;
  assign n28811 = n28621 ^ n28618 ;
  assign n28812 = n28699 & n28811 ;
  assign n28813 = n28812 ^ n28618 ;
  assign n28806 = n4916 & ~n25287 ;
  assign n28799 = n25693 ^ x20 ;
  assign n28800 = n28799 ^ x19 ;
  assign n28801 = n28800 ^ n25693 ;
  assign n28802 = n25705 & ~n28801 ;
  assign n28803 = n28802 ^ n25693 ;
  assign n28804 = n4678 & n28803 ;
  assign n28805 = n28804 ^ x20 ;
  assign n28807 = n28806 ^ n28805 ;
  assign n28798 = n14027 & n25043 ;
  assign n28808 = n28807 ^ n28798 ;
  assign n28789 = ~n4496 & ~n24700 ;
  assign n28782 = n24980 ^ x23 ;
  assign n28783 = n28782 ^ x22 ;
  assign n28784 = n28783 ^ n24980 ;
  assign n28785 = ~n25518 & n28784 ;
  assign n28786 = n28785 ^ n24980 ;
  assign n28787 = n4488 & ~n28786 ;
  assign n28788 = n28787 ^ x23 ;
  assign n28790 = n28789 ^ n28788 ;
  assign n28781 = n4504 & n24079 ;
  assign n28791 = n28790 ^ n28781 ;
  assign n28766 = n13789 ^ n564 ;
  assign n28763 = n4267 ^ n2069 ;
  assign n28764 = n28763 ^ n2690 ;
  assign n28761 = n15103 ^ n12563 ;
  assign n28762 = n28761 ^ n5332 ;
  assign n28765 = n28764 ^ n28762 ;
  assign n28767 = n28766 ^ n28765 ;
  assign n28760 = n12028 ^ n2905 ;
  assign n28768 = n28767 ^ n28760 ;
  assign n28769 = n5001 ^ n1867 ;
  assign n28770 = ~n28768 & ~n28769 ;
  assign n28758 = n28679 ^ n28667 ;
  assign n28759 = ~n28672 & n28758 ;
  assign n28771 = n28770 ^ n28759 ;
  assign n28746 = n3520 ^ x31 ;
  assign n28747 = n28746 ^ n20872 ;
  assign n28748 = n28747 ^ n20872 ;
  assign n28749 = n28748 ^ x31 ;
  assign n28752 = ~x31 & ~n20872 ;
  assign n28750 = n20876 ^ x31 ;
  assign n28751 = n5281 & ~n28750 ;
  assign n28753 = n28752 ^ n28751 ;
  assign n28754 = ~n28749 & n28753 ;
  assign n28755 = n28754 ^ n28752 ;
  assign n28756 = n28755 ^ x31 ;
  assign n28740 = n23033 ^ n20882 ;
  assign n28743 = n35 & n28740 ;
  assign n28744 = n28743 ^ n20882 ;
  assign n28745 = n4851 & ~n28744 ;
  assign n28757 = n28756 ^ n28745 ;
  assign n28772 = n28771 ^ n28757 ;
  assign n28737 = n3484 & n20861 ;
  assign n28730 = n20852 ^ x29 ;
  assign n28731 = n28730 ^ x28 ;
  assign n28732 = n28731 ^ n20852 ;
  assign n28733 = ~n23059 & n28732 ;
  assign n28734 = n28733 ^ n20852 ;
  assign n28735 = n650 & n28734 ;
  assign n28736 = n28735 ^ x29 ;
  assign n28738 = n28737 ^ n28736 ;
  assign n28728 = n831 & n20865 ;
  assign n28739 = n28738 ^ n28728 ;
  assign n28773 = n28772 ^ n28739 ;
  assign n28725 = n28654 ^ n28644 ;
  assign n28726 = ~n28681 & n28725 ;
  assign n28727 = n28726 ^ n28654 ;
  assign n28774 = n28773 ^ n28727 ;
  assign n28720 = n446 & n20837 ;
  assign n28719 = ~n487 & n20834 ;
  assign n28721 = n28720 ^ n28719 ;
  assign n28722 = n28721 ^ x26 ;
  assign n28718 = n12861 & n20836 ;
  assign n28723 = n28722 ^ n28718 ;
  assign n28717 = ~n3501 & ~n24936 ;
  assign n28724 = n28723 ^ n28717 ;
  assign n28775 = n28774 ^ n28724 ;
  assign n28777 = n28775 ^ n28682 ;
  assign n28776 = n28775 ^ n28695 ;
  assign n28778 = n28777 ^ n28776 ;
  assign n28779 = ~n28687 & ~n28778 ;
  assign n28780 = n28779 ^ n28777 ;
  assign n28792 = n28791 ^ n28780 ;
  assign n28793 = n28792 ^ n28632 ;
  assign n28794 = n28793 ^ n28629 ;
  assign n28795 = n28794 ^ n28792 ;
  assign n28796 = ~n28697 & n28795 ;
  assign n28797 = n28796 ^ n28793 ;
  assign n28809 = n28808 ^ n28797 ;
  assign n28810 = n28809 ^ x17 ;
  assign n28814 = n28813 ^ n28810 ;
  assign n28818 = n28817 ^ n28814 ;
  assign n28715 = ~n28706 & n28710 ;
  assign n28712 = n28607 ^ n28581 ;
  assign n28713 = ~n28705 & n28712 ;
  assign n28714 = n28713 ^ n28607 ;
  assign n28716 = n28715 ^ n28714 ;
  assign n28819 = n28818 ^ n28716 ;
  assign n28913 = n28814 ^ n28715 ;
  assign n28916 = ~n28716 & ~n28913 ;
  assign n28914 = n28913 ^ n28714 ;
  assign n28915 = n28817 & n28914 ;
  assign n28917 = n28916 ^ n28915 ;
  assign n28904 = ~n3501 & ~n25245 ;
  assign n28901 = n446 & n20834 ;
  assign n28899 = n12861 & n20837 ;
  assign n28895 = n28727 ^ n28724 ;
  assign n28896 = n28774 & n28895 ;
  assign n28897 = n28896 ^ n28724 ;
  assign n28898 = n28897 ^ x26 ;
  assign n28900 = n28899 ^ n28898 ;
  assign n28902 = n28901 ^ n28900 ;
  assign n28894 = ~n487 & n24079 ;
  assign n28903 = n28902 ^ n28894 ;
  assign n28905 = n28904 ^ n28903 ;
  assign n28890 = n831 & n20861 ;
  assign n28883 = n28770 ^ n28679 ;
  assign n28884 = ~n28759 & n28883 ;
  assign n28885 = n28884 ^ n28679 ;
  assign n28881 = n28770 ^ x17 ;
  assign n28875 = n12032 ^ n382 ;
  assign n28873 = n882 ^ n250 ;
  assign n28872 = n12406 ^ n88 ;
  assign n28874 = n28873 ^ n28872 ;
  assign n28876 = n28875 ^ n28874 ;
  assign n28868 = n2397 ^ n297 ;
  assign n28867 = n24205 ^ n743 ;
  assign n28869 = n28868 ^ n28867 ;
  assign n28870 = n28869 ^ n1646 ;
  assign n28871 = n28870 ^ n12433 ;
  assign n28877 = n28876 ^ n28871 ;
  assign n28878 = n28877 ^ n1469 ;
  assign n28879 = n28878 ^ n4783 ;
  assign n28880 = ~n3767 & ~n28879 ;
  assign n28882 = n28881 ^ n28880 ;
  assign n28886 = n28885 ^ n28882 ;
  assign n28861 = x31 & ~n20876 ;
  assign n28862 = n28861 ^ n20872 ;
  assign n28863 = ~n5281 & ~n28862 ;
  assign n28853 = x31 & ~n22682 ;
  assign n28854 = n28853 ^ n20865 ;
  assign n28855 = n28854 ^ n20872 ;
  assign n28864 = n28863 ^ n28855 ;
  assign n28865 = ~n3520 & ~n28864 ;
  assign n28866 = n28865 ^ n28854 ;
  assign n28887 = n28886 ^ n28866 ;
  assign n28888 = n28887 ^ x29 ;
  assign n28848 = n20836 ^ n4536 ;
  assign n28849 = n28848 ^ n20836 ;
  assign n28850 = ~n26327 & n28849 ;
  assign n28851 = n28850 ^ n20836 ;
  assign n28852 = n650 & n28851 ;
  assign n28889 = n28888 ^ n28852 ;
  assign n28891 = n28890 ^ n28889 ;
  assign n28847 = n3484 & n20852 ;
  assign n28892 = n28891 ^ n28847 ;
  assign n28844 = n28757 ^ n28739 ;
  assign n28845 = ~n28772 & n28844 ;
  assign n28846 = n28845 ^ n28757 ;
  assign n28893 = n28892 ^ n28846 ;
  assign n28906 = n28905 ^ n28893 ;
  assign n28842 = ~n4496 & ~n24980 ;
  assign n28840 = n4492 & ~n25896 ;
  assign n28837 = n4504 & ~n24700 ;
  assign n28836 = n4491 & n25043 ;
  assign n28838 = n28837 ^ n28836 ;
  assign n28839 = n28838 ^ x23 ;
  assign n28841 = n28840 ^ n28839 ;
  assign n28843 = n28842 ^ n28841 ;
  assign n28907 = n28906 ^ n28843 ;
  assign n28833 = n28791 ^ n28775 ;
  assign n28834 = n28780 & ~n28833 ;
  assign n28835 = n28834 ^ n28775 ;
  assign n28908 = n28907 ^ n28835 ;
  assign n28827 = n14027 ^ n4916 ;
  assign n28828 = n28827 ^ n28611 ;
  assign n28829 = n25287 & n28828 ;
  assign n28831 = n28829 ^ n14026 ;
  assign n28826 = n4684 & n25725 ;
  assign n28832 = n28831 ^ n28826 ;
  assign n28909 = n28908 ^ n28832 ;
  assign n28823 = n28808 ^ n28792 ;
  assign n28824 = n28797 & n28823 ;
  assign n28825 = n28824 ^ n28792 ;
  assign n28910 = n28909 ^ n28825 ;
  assign n28911 = n28910 ^ x17 ;
  assign n28820 = n28813 ^ n28809 ;
  assign n28821 = n28813 ^ x17 ;
  assign n28822 = ~n28820 & n28821 ;
  assign n28912 = n28911 ^ n28822 ;
  assign n28918 = n28917 ^ n28912 ;
  assign n29021 = n28818 ^ n28714 ;
  assign n29022 = n28912 ^ n28714 ;
  assign n29023 = ~n29021 & n29022 ;
  assign n29024 = n28715 & n29023 ;
  assign n29016 = n14027 & n25703 ;
  assign n29007 = n12861 & n20834 ;
  assign n29006 = n446 & n24079 ;
  assign n29008 = n29007 ^ n29006 ;
  assign n29009 = n29008 ^ x26 ;
  assign n29005 = ~n487 & ~n24700 ;
  assign n29010 = n29009 ^ n29005 ;
  assign n29004 = ~n3501 & n25320 ;
  assign n29011 = n29010 ^ n29004 ;
  assign n28994 = n28880 ^ n28770 ;
  assign n28995 = n28881 & ~n28994 ;
  assign n28996 = n28995 ^ x17 ;
  assign n28985 = n12493 ^ n4132 ;
  assign n28986 = n28985 ^ n6491 ;
  assign n28983 = n2785 ^ n1451 ;
  assign n28981 = n1358 ^ n567 ;
  assign n28979 = n15120 ^ n426 ;
  assign n28980 = n28979 ^ n641 ;
  assign n28982 = n28981 ^ n28980 ;
  assign n28984 = n28983 ^ n28982 ;
  assign n28987 = n28986 ^ n28984 ;
  assign n28988 = n28987 ^ n1072 ;
  assign n28989 = n28988 ^ n2954 ;
  assign n28990 = n27373 ^ n6233 ;
  assign n28991 = ~n28989 & ~n28990 ;
  assign n28971 = x30 & n20865 ;
  assign n28972 = n28971 ^ n20861 ;
  assign n28973 = ~n3520 & n28972 ;
  assign n28974 = n28973 ^ n20861 ;
  assign n28975 = n28974 ^ n23640 ;
  assign n28962 = n23640 ^ n20865 ;
  assign n28961 = n23640 ^ n20872 ;
  assign n28963 = n28962 ^ n28961 ;
  assign n28966 = x30 & ~n28963 ;
  assign n28967 = n28966 ^ n28962 ;
  assign n28968 = ~n3520 & ~n28967 ;
  assign n28976 = n28975 ^ n28968 ;
  assign n28977 = x31 & ~n28976 ;
  assign n28978 = n28977 ^ n28974 ;
  assign n28992 = n28991 ^ n28978 ;
  assign n28958 = n28885 ^ n28866 ;
  assign n28959 = ~n28886 & n28958 ;
  assign n28960 = n28959 ^ n28885 ;
  assign n28993 = n28992 ^ n28960 ;
  assign n28997 = n28996 ^ n28993 ;
  assign n28955 = n3484 & n20836 ;
  assign n28948 = n20837 ^ x29 ;
  assign n28949 = n28948 ^ x28 ;
  assign n28950 = n28949 ^ n20837 ;
  assign n28951 = ~n21061 & n28950 ;
  assign n28952 = n28951 ^ n20837 ;
  assign n28953 = n650 & n28952 ;
  assign n28954 = n28953 ^ x29 ;
  assign n28956 = n28955 ^ n28954 ;
  assign n28947 = n831 & n20852 ;
  assign n28957 = n28956 ^ n28947 ;
  assign n28998 = n28997 ^ n28957 ;
  assign n28999 = n28998 ^ n28887 ;
  assign n29000 = n28999 ^ n28998 ;
  assign n29001 = n29000 ^ n28846 ;
  assign n29002 = ~n28892 & ~n29001 ;
  assign n29003 = n29002 ^ n28999 ;
  assign n29012 = n29011 ^ n29003 ;
  assign n28944 = n28897 ^ n28893 ;
  assign n28945 = n28905 & ~n28944 ;
  assign n28946 = n28945 ^ n28897 ;
  assign n29013 = n29012 ^ n28946 ;
  assign n28938 = ~n4496 & n25043 ;
  assign n28937 = n4491 & n25287 ;
  assign n28939 = n28938 ^ n28937 ;
  assign n28940 = n28939 ^ n4491 ;
  assign n28941 = n28940 ^ x23 ;
  assign n28936 = n4504 & ~n24980 ;
  assign n28942 = n28941 ^ n28936 ;
  assign n28935 = n4492 & n25937 ;
  assign n28943 = n28942 ^ n28935 ;
  assign n29014 = n29013 ^ n28943 ;
  assign n29015 = n29014 ^ x20 ;
  assign n29017 = n29016 ^ n29015 ;
  assign n28932 = n28843 ^ n28835 ;
  assign n28933 = ~n28907 & ~n28932 ;
  assign n28934 = n28933 ^ n28843 ;
  assign n29018 = n29017 ^ n28934 ;
  assign n28929 = n28832 ^ n28825 ;
  assign n28930 = n28909 & n28929 ;
  assign n28931 = n28930 ^ n28832 ;
  assign n29019 = n29018 ^ n28931 ;
  assign n28919 = n28817 ^ n28714 ;
  assign n28920 = n28912 & n28919 ;
  assign n28921 = n28910 ^ n28813 ;
  assign n28922 = n28910 ^ n28809 ;
  assign n28923 = n28911 & n28922 ;
  assign n28924 = n28921 & n28923 ;
  assign n28925 = n28924 ^ n28910 ;
  assign n28926 = n28925 ^ n28817 ;
  assign n28927 = n28920 & ~n28926 ;
  assign n28928 = n28927 ^ n28925 ;
  assign n29020 = n29019 ^ n28928 ;
  assign n29025 = n29024 ^ n29020 ;
  assign n29122 = n29014 ^ n28934 ;
  assign n29123 = n29017 & n29122 ;
  assign n29124 = n29123 ^ n29014 ;
  assign n29118 = n28946 ^ n28943 ;
  assign n29119 = ~n29013 & n29118 ;
  assign n29120 = n29119 ^ n28943 ;
  assign n29112 = ~n4496 & ~n25287 ;
  assign n29111 = n4492 & n25693 ;
  assign n29113 = n29112 ^ n29111 ;
  assign n29110 = n4504 ^ x23 ;
  assign n29114 = n29113 ^ n29110 ;
  assign n29108 = n28937 ^ n4504 ;
  assign n29109 = ~n25043 & n29108 ;
  assign n29115 = n29114 ^ n29109 ;
  assign n29099 = n3484 & n20837 ;
  assign n29062 = n28978 ^ n28960 ;
  assign n29094 = n28960 ^ n28957 ;
  assign n29095 = ~n29062 & ~n29094 ;
  assign n29088 = n6259 ^ n4285 ;
  assign n29084 = n14330 ^ n732 ;
  assign n29082 = n15103 ^ n667 ;
  assign n29083 = n29082 ^ n284 ;
  assign n29085 = n29084 ^ n29083 ;
  assign n29079 = n1998 ^ n760 ;
  assign n29077 = n13253 ^ n280 ;
  assign n29078 = n29077 ^ n2969 ;
  assign n29080 = n29079 ^ n29078 ;
  assign n29081 = n29080 ^ n26610 ;
  assign n29086 = n29085 ^ n29081 ;
  assign n29087 = n29086 ^ n3753 ;
  assign n29089 = n29088 ^ n29087 ;
  assign n29090 = ~n1470 & ~n29089 ;
  assign n29091 = n29090 ^ n28991 ;
  assign n29075 = ~n23825 & n23912 ;
  assign n29073 = ~n3733 & ~n20861 ;
  assign n29067 = x30 & ~n20865 ;
  assign n29068 = n29067 ^ n20852 ;
  assign n29069 = ~n3520 & n29068 ;
  assign n29070 = n29069 ^ n20852 ;
  assign n29071 = n28746 & ~n29070 ;
  assign n29072 = n29071 ^ n3514 ;
  assign n29074 = n29073 ^ n29072 ;
  assign n29076 = n29075 ^ n29074 ;
  assign n29092 = n29091 ^ n29076 ;
  assign n29060 = n28996 ^ n28991 ;
  assign n29061 = n28991 ^ n28957 ;
  assign n29063 = n29062 ^ n29061 ;
  assign n29064 = n29060 & n29063 ;
  assign n29093 = n29092 ^ n29064 ;
  assign n29096 = n29095 ^ n29093 ;
  assign n29097 = n29096 ^ x29 ;
  assign n29055 = n20834 ^ n4536 ;
  assign n29056 = n29055 ^ n20834 ;
  assign n29057 = ~n21055 & n29056 ;
  assign n29058 = n29057 ^ n20834 ;
  assign n29059 = n650 & n29058 ;
  assign n29098 = n29097 ^ n29059 ;
  assign n29100 = n29099 ^ n29098 ;
  assign n29054 = n831 & n20836 ;
  assign n29101 = n29100 ^ n29054 ;
  assign n29033 = n446 & ~n24700 ;
  assign n29032 = n12861 & n24079 ;
  assign n29034 = n29033 ^ n29032 ;
  assign n29035 = n29034 ^ n65 ;
  assign n29036 = n29034 ^ x26 ;
  assign n29037 = n29036 ^ n67 ;
  assign n29038 = n29037 ^ x25 ;
  assign n29039 = n29038 ^ n24980 ;
  assign n29040 = n29039 ^ n29036 ;
  assign n29041 = n29040 ^ n24949 ;
  assign n29042 = n29041 ^ n29040 ;
  assign n29043 = n29036 & ~n29042 ;
  assign n29044 = n29043 ^ n29037 ;
  assign n29045 = n29040 ^ n24980 ;
  assign n29046 = ~n29042 & ~n29045 ;
  assign n29047 = n29046 ^ n24980 ;
  assign n29048 = ~n29037 & n29047 ;
  assign n29049 = ~n29044 & n29048 ;
  assign n29050 = n29049 ^ n29046 ;
  assign n29051 = n29050 ^ n67 ;
  assign n29052 = n29051 ^ n24980 ;
  assign n29053 = ~n29035 & ~n29052 ;
  assign n29102 = n29101 ^ n29053 ;
  assign n29104 = n29102 ^ n28998 ;
  assign n29103 = n29102 ^ n29011 ;
  assign n29105 = n29104 ^ n29103 ;
  assign n29106 = n29003 & ~n29105 ;
  assign n29107 = n29106 ^ n29104 ;
  assign n29116 = n29115 ^ n29107 ;
  assign n29117 = n29116 ^ x20 ;
  assign n29121 = n29120 ^ n29117 ;
  assign n29125 = n29124 ^ n29121 ;
  assign n29026 = n29018 ^ n28928 ;
  assign n29029 = n28931 ^ n28928 ;
  assign n29030 = ~n29026 & ~n29029 ;
  assign n29027 = n29026 ^ n28931 ;
  assign n29028 = ~n29024 & n29027 ;
  assign n29031 = n29030 ^ n29028 ;
  assign n29126 = n29125 ^ n29031 ;
  assign n29244 = n29115 ^ n29102 ;
  assign n29245 = ~n29107 & n29244 ;
  assign n29246 = n29245 ^ n29102 ;
  assign n29216 = ~n28957 & ~n28960 ;
  assign n29217 = n29216 ^ n29094 ;
  assign n29218 = n29216 ^ n29092 ;
  assign n29220 = n29216 ^ n28996 ;
  assign n29219 = n29216 ^ n28978 ;
  assign n29221 = n29220 ^ n29219 ;
  assign n29222 = n29219 ^ n28992 ;
  assign n29223 = n29222 ^ n29219 ;
  assign n29224 = ~n29221 & n29223 ;
  assign n29225 = n29224 ^ n29219 ;
  assign n29226 = ~n29218 & n29225 ;
  assign n29227 = n29226 ^ n29092 ;
  assign n29228 = n29092 ^ n28978 ;
  assign n29229 = n29092 ^ n28996 ;
  assign n29230 = n29092 ^ n28991 ;
  assign n29231 = ~n29229 & n29230 ;
  assign n29232 = n29228 & n29231 ;
  assign n29233 = n29232 ^ n29228 ;
  assign n29234 = n29233 ^ n28978 ;
  assign n29235 = n29227 & ~n29234 ;
  assign n29236 = n29217 & n29235 ;
  assign n29237 = n29236 ^ n29227 ;
  assign n29205 = n356 ^ n283 ;
  assign n29204 = n1809 ^ n273 ;
  assign n29206 = n29205 ^ n29204 ;
  assign n29202 = n794 ^ n542 ;
  assign n29201 = n13143 ^ n3408 ;
  assign n29203 = n29202 ^ n29201 ;
  assign n29207 = n29206 ^ n29203 ;
  assign n29208 = n29207 ^ n2904 ;
  assign n29209 = n29208 ^ n15116 ;
  assign n29198 = n5058 ^ n1528 ;
  assign n29199 = n29198 ^ n1297 ;
  assign n29200 = n29199 ^ n14332 ;
  assign n29210 = n29209 ^ n29200 ;
  assign n29211 = n29210 ^ n1568 ;
  assign n29212 = ~n4335 & ~n29211 ;
  assign n29213 = n29212 ^ x20 ;
  assign n29196 = n29076 ^ n28991 ;
  assign n29197 = ~n29091 & ~n29196 ;
  assign n29214 = n29213 ^ n29197 ;
  assign n29192 = n33 & ~n20852 ;
  assign n29186 = x30 & n20852 ;
  assign n29187 = n29186 ^ n20836 ;
  assign n29188 = ~n3520 & n29187 ;
  assign n29189 = n29188 ^ n20836 ;
  assign n29190 = ~x31 & n29189 ;
  assign n29179 = x30 & ~n20861 ;
  assign n29180 = n29179 ^ n24433 ;
  assign n29181 = ~n3520 & n29180 ;
  assign n29182 = n29181 ^ n24433 ;
  assign n29183 = x31 & ~n29182 ;
  assign n29191 = n29190 ^ n29183 ;
  assign n29193 = n29191 ^ n29190 ;
  assign n29194 = n29192 & n29193 ;
  assign n29195 = n29194 ^ n29191 ;
  assign n29215 = n29214 ^ n29195 ;
  assign n29238 = n29237 ^ n29215 ;
  assign n29172 = n831 & n20837 ;
  assign n29171 = n3484 & n20834 ;
  assign n29173 = n29172 ^ n29171 ;
  assign n29174 = n29173 ^ n651 ;
  assign n29166 = ~x28 & ~n24004 ;
  assign n29169 = n29166 ^ n24079 ;
  assign n29170 = n28635 & ~n29169 ;
  assign n29175 = n29174 ^ n29170 ;
  assign n29167 = n29166 ^ n25245 ;
  assign n29168 = n653 & ~n29167 ;
  assign n29176 = n29175 ^ n29168 ;
  assign n29239 = n29238 ^ n29176 ;
  assign n29149 = n12861 & ~n24700 ;
  assign n29148 = n446 & ~n24980 ;
  assign n29150 = n29149 ^ n29148 ;
  assign n29151 = n29150 ^ n65 ;
  assign n29153 = n29150 ^ x26 ;
  assign n29156 = n29153 ^ n67 ;
  assign n29157 = ~x25 & ~n25008 ;
  assign n29158 = n29156 & n29157 ;
  assign n29154 = ~n25043 & n29153 ;
  assign n29152 = n67 & ~n25896 ;
  assign n29155 = n29154 ^ n29152 ;
  assign n29159 = n29158 ^ n29155 ;
  assign n29160 = ~n29151 & ~n29159 ;
  assign n29161 = n29160 ^ n29096 ;
  assign n29162 = n29161 ^ n29053 ;
  assign n29163 = n29162 ^ n29160 ;
  assign n29164 = ~n29101 & n29163 ;
  assign n29165 = n29164 ^ n29161 ;
  assign n29240 = n29239 ^ n29165 ;
  assign n29241 = n29240 ^ n29110 ;
  assign n29145 = n4504 ^ n4496 ;
  assign n29146 = n29145 ^ n28938 ;
  assign n29147 = n25287 & ~n29146 ;
  assign n29242 = n29241 ^ n29147 ;
  assign n29144 = n4492 & n25725 ;
  assign n29243 = n29242 ^ n29144 ;
  assign n29247 = n29246 ^ n29243 ;
  assign n29140 = n29120 ^ n29116 ;
  assign n29141 = n29120 ^ x20 ;
  assign n29142 = n29140 & n29141 ;
  assign n29143 = n29142 ^ x20 ;
  assign n29248 = n29247 ^ n29143 ;
  assign n29131 = n29124 ^ n29018 ;
  assign n29132 = n29131 ^ n29029 ;
  assign n29133 = n29132 ^ n29131 ;
  assign n29134 = n29124 ^ n28931 ;
  assign n29135 = n29134 ^ n29131 ;
  assign n29136 = ~n29133 & n29135 ;
  assign n29137 = n29136 ^ n29131 ;
  assign n29138 = ~n29125 & n29137 ;
  assign n29139 = n29138 ^ n29124 ;
  assign n29249 = n29248 ^ n29139 ;
  assign n29127 = n29020 & n29024 ;
  assign n29128 = n28928 & n28931 ;
  assign n29129 = n29128 ^ n29125 ;
  assign n29130 = n29127 & ~n29129 ;
  assign n29250 = n29249 ^ n29130 ;
  assign n29331 = n29130 & ~n29249 ;
  assign n29328 = n29246 ^ n29240 ;
  assign n29329 = n29243 & ~n29328 ;
  assign n29330 = n29329 ^ n29246 ;
  assign n29332 = n29331 ^ n29330 ;
  assign n29323 = n29239 ^ n29160 ;
  assign n29324 = n29165 & n29323 ;
  assign n29325 = n29324 ^ n29160 ;
  assign n29320 = n4504 & n25703 ;
  assign n29321 = n29320 ^ x23 ;
  assign n29315 = n831 & n20834 ;
  assign n29313 = n3484 & n24079 ;
  assign n29307 = n29213 ^ n28991 ;
  assign n29308 = n29307 ^ n29195 ;
  assign n29309 = n29214 & ~n29308 ;
  assign n29310 = n29309 ^ n29195 ;
  assign n29311 = n29310 ^ x29 ;
  assign n29302 = n24700 ^ n4536 ;
  assign n29303 = n29302 ^ n24700 ;
  assign n29304 = ~n28178 & n29303 ;
  assign n29305 = n29304 ^ n24700 ;
  assign n29306 = n650 & ~n29305 ;
  assign n29312 = n29311 ^ n29306 ;
  assign n29314 = n29313 ^ n29312 ;
  assign n29316 = n29315 ^ n29314 ;
  assign n29296 = n29212 ^ n28991 ;
  assign n29297 = n28991 ^ x20 ;
  assign n29298 = ~n29296 & n29297 ;
  assign n29299 = n29298 ^ x20 ;
  assign n29286 = n1039 ^ n433 ;
  assign n29287 = n29286 ^ n506 ;
  assign n29285 = n673 ^ n635 ;
  assign n29288 = n29287 ^ n29285 ;
  assign n29283 = n2243 ^ n1982 ;
  assign n29282 = n3995 ^ n1500 ;
  assign n29284 = n29283 ^ n29282 ;
  assign n29289 = n29288 ^ n29284 ;
  assign n29290 = n29289 ^ n2204 ;
  assign n29291 = n29290 ^ n3571 ;
  assign n29292 = n29291 ^ n13930 ;
  assign n29293 = n15196 ^ n3767 ;
  assign n29294 = n29293 ^ n2352 ;
  assign n29295 = ~n29292 & ~n29294 ;
  assign n29300 = n29299 ^ n29295 ;
  assign n29276 = ~n35 & n20836 ;
  assign n29274 = ~n3520 & ~n20837 ;
  assign n29273 = n20837 ^ n3520 ;
  assign n29275 = n29274 ^ n29273 ;
  assign n29277 = n29276 ^ n29275 ;
  assign n29278 = n29277 ^ n24427 ;
  assign n29266 = n24427 ^ n20852 ;
  assign n29265 = n24427 ^ n20836 ;
  assign n29267 = n29266 ^ n29265 ;
  assign n29270 = ~x30 & n29267 ;
  assign n29271 = n29270 ^ n29266 ;
  assign n29272 = ~n3520 & ~n29271 ;
  assign n29279 = n29278 ^ n29272 ;
  assign n29280 = x31 & n29279 ;
  assign n29281 = n29280 ^ n29277 ;
  assign n29301 = n29300 ^ n29281 ;
  assign n29317 = n29316 ^ n29301 ;
  assign n29262 = n29237 ^ n29176 ;
  assign n29263 = ~n29238 & n29262 ;
  assign n29264 = n29263 ^ n29237 ;
  assign n29318 = n29317 ^ n29264 ;
  assign n29257 = n12861 & ~n24980 ;
  assign n29256 = n446 & n25043 ;
  assign n29258 = n29257 ^ n29256 ;
  assign n29259 = n29258 ^ x26 ;
  assign n29255 = ~n487 & ~n25287 ;
  assign n29260 = n29259 ^ n29255 ;
  assign n29254 = ~n3501 & n25937 ;
  assign n29261 = n29260 ^ n29254 ;
  assign n29319 = n29318 ^ n29261 ;
  assign n29322 = n29321 ^ n29319 ;
  assign n29326 = n29325 ^ n29322 ;
  assign n29251 = n29143 ^ n29139 ;
  assign n29252 = n29248 & n29251 ;
  assign n29253 = n29252 ^ n29139 ;
  assign n29327 = n29326 ^ n29253 ;
  assign n29333 = n29332 ^ n29327 ;
  assign n29398 = n29264 ^ n29261 ;
  assign n29399 = ~n29318 & n29398 ;
  assign n29400 = n29399 ^ n29261 ;
  assign n29393 = ~n3501 & n25693 ;
  assign n29392 = n446 ^ x26 ;
  assign n29394 = n29393 ^ n29392 ;
  assign n29391 = n12861 & n25043 ;
  assign n29395 = n29394 ^ n29391 ;
  assign n29388 = ~n487 & ~n25043 ;
  assign n29389 = n29388 ^ n446 ;
  assign n29390 = n25287 & n29389 ;
  assign n29396 = n29395 ^ n29390 ;
  assign n29376 = n12533 & ~n29274 ;
  assign n29373 = ~n35 & n20837 ;
  assign n29365 = n1036 ^ n811 ;
  assign n29364 = n1982 ^ n1283 ;
  assign n29366 = n29365 ^ n29364 ;
  assign n29362 = n15001 ^ n2852 ;
  assign n29360 = n375 ^ n266 ;
  assign n29359 = n1185 ^ n106 ;
  assign n29361 = n29360 ^ n29359 ;
  assign n29363 = n29362 ^ n29361 ;
  assign n29367 = n29366 ^ n29363 ;
  assign n29368 = n29367 ^ n27359 ;
  assign n29369 = n29368 ^ n12909 ;
  assign n29370 = n29369 ^ n23734 ;
  assign n29371 = ~n4197 & ~n29370 ;
  assign n29357 = n29299 ^ n29281 ;
  assign n29358 = ~n29300 & ~n29357 ;
  assign n29372 = n29371 ^ n29358 ;
  assign n29374 = n29373 ^ n29372 ;
  assign n29354 = x31 & ~n21055 ;
  assign n29355 = n29354 ^ n20834 ;
  assign n29356 = n3520 & ~n29355 ;
  assign n29375 = n29374 ^ n29356 ;
  assign n29377 = n29376 ^ n29375 ;
  assign n29351 = x31 & n29276 ;
  assign n29378 = n29377 ^ n29351 ;
  assign n29348 = n29310 ^ n29301 ;
  assign n29349 = n29316 & n29348 ;
  assign n29350 = n29349 ^ n29310 ;
  assign n29379 = n29378 ^ n29350 ;
  assign n29380 = n29379 ^ x29 ;
  assign n29347 = n3484 & ~n24700 ;
  assign n29381 = n29380 ^ n29347 ;
  assign n29346 = n831 & n24079 ;
  assign n29382 = n29381 ^ n29346 ;
  assign n29341 = n24980 ^ n4536 ;
  assign n29342 = n29341 ^ n24980 ;
  assign n29343 = ~n25518 & n29342 ;
  assign n29344 = n29343 ^ n24980 ;
  assign n29345 = n650 & ~n29344 ;
  assign n29383 = n29382 ^ n29345 ;
  assign n29397 = n29396 ^ n29383 ;
  assign n29401 = n29400 ^ n29397 ;
  assign n29402 = n29401 ^ x23 ;
  assign n29338 = n29319 ^ n29253 ;
  assign n29339 = ~n29322 & ~n29338 ;
  assign n29336 = n29322 ^ n29253 ;
  assign n29337 = ~n29325 & ~n29336 ;
  assign n29340 = n29339 ^ n29337 ;
  assign n29403 = n29402 ^ n29340 ;
  assign n29334 = n29330 ^ n29327 ;
  assign n29335 = ~n29332 & ~n29334 ;
  assign n29404 = n29403 ^ n29335 ;
  assign n29480 = n29372 ^ n29350 ;
  assign n29481 = ~n29378 & ~n29480 ;
  assign n29482 = n29481 ^ n29372 ;
  assign n29475 = n29371 ^ x23 ;
  assign n29469 = n1999 ^ n448 ;
  assign n29468 = n5097 ^ n683 ;
  assign n29470 = n29469 ^ n29468 ;
  assign n29466 = n1834 ^ n259 ;
  assign n29467 = n29466 ^ n857 ;
  assign n29471 = n29470 ^ n29467 ;
  assign n29465 = n4808 ^ n1781 ;
  assign n29472 = n29471 ^ n29465 ;
  assign n29473 = n29472 ^ n387 ;
  assign n29474 = n29473 ^ n12646 ;
  assign n29476 = n29475 ^ n29474 ;
  assign n29462 = n29371 ^ n29295 ;
  assign n29463 = ~n29358 & ~n29462 ;
  assign n29464 = n29463 ^ n29295 ;
  assign n29477 = n29476 ^ n29464 ;
  assign n29459 = x31 & n29373 ;
  assign n29458 = ~n3733 & n20834 ;
  assign n29460 = n29459 ^ n29458 ;
  assign n29455 = x31 & ~n28113 ;
  assign n29456 = n29455 ^ n24079 ;
  assign n29457 = n3520 & n29456 ;
  assign n29461 = n29460 ^ n29457 ;
  assign n29478 = n29477 ^ n29461 ;
  assign n29448 = n3484 & ~n24980 ;
  assign n29441 = n25043 ^ x29 ;
  assign n29442 = n29441 ^ x28 ;
  assign n29443 = n29442 ^ n25043 ;
  assign n29444 = ~n27539 & n29443 ;
  assign n29445 = n29444 ^ n25043 ;
  assign n29446 = n650 & n29445 ;
  assign n29447 = n29446 ^ x29 ;
  assign n29449 = n29448 ^ n29447 ;
  assign n29440 = n831 & ~n24700 ;
  assign n29450 = n29449 ^ n29440 ;
  assign n29479 = n29478 ^ n29450 ;
  assign n29483 = n29482 ^ n29479 ;
  assign n29438 = n446 & n25703 ;
  assign n29435 = n12861 & ~n25287 ;
  assign n29434 = ~n3501 & n25725 ;
  assign n29436 = n29435 ^ n29434 ;
  assign n29437 = n29436 ^ x26 ;
  assign n29439 = n29438 ^ n29437 ;
  assign n29484 = n29483 ^ n29439 ;
  assign n29430 = n29400 ^ x23 ;
  assign n29431 = n29401 & n29430 ;
  assign n29432 = n29431 ^ x23 ;
  assign n29427 = n29396 ^ n29379 ;
  assign n29428 = ~n29383 & ~n29427 ;
  assign n29429 = n29428 ^ n29379 ;
  assign n29433 = n29432 ^ n29429 ;
  assign n29485 = n29484 ^ n29433 ;
  assign n29408 = n29402 ^ n29325 ;
  assign n29409 = n29325 ^ n29319 ;
  assign n29410 = n29408 & n29409 ;
  assign n29411 = n29330 ^ n29325 ;
  assign n29412 = n29410 & n29411 ;
  assign n29413 = n29412 ^ n29402 ;
  assign n29414 = ~n29321 & n29413 ;
  assign n29415 = n29330 ^ n29319 ;
  assign n29416 = ~n29409 & ~n29415 ;
  assign n29417 = n29416 ^ n29325 ;
  assign n29418 = n29402 & n29417 ;
  assign n29419 = ~n29414 & ~n29418 ;
  assign n29420 = n29413 ^ n29321 ;
  assign n29421 = n29420 ^ n29414 ;
  assign n29422 = n29417 ^ n29402 ;
  assign n29423 = n29422 ^ n29418 ;
  assign n29424 = ~n29421 & n29423 ;
  assign n29425 = ~n29253 & n29424 ;
  assign n29426 = n29419 & ~n29425 ;
  assign n29486 = n29485 ^ n29426 ;
  assign n29405 = n29403 ^ n29330 ;
  assign n29406 = n29331 & ~n29334 ;
  assign n29407 = ~n29405 & n29406 ;
  assign n29487 = n29486 ^ n29407 ;
  assign n29567 = n29407 & n29486 ;
  assign n29564 = n29433 ^ n29426 ;
  assign n29565 = n29485 & n29564 ;
  assign n29544 = n24675 ^ n14523 ;
  assign n29550 = ~n386 & ~n2112 ;
  assign n29547 = n4267 ^ n2303 ;
  assign n29546 = n5631 ^ n5134 ;
  assign n29548 = n29547 ^ n29546 ;
  assign n29545 = n357 ^ n223 ;
  assign n29549 = n29548 ^ n29545 ;
  assign n29551 = n29550 ^ n29549 ;
  assign n29552 = ~n29544 & n29551 ;
  assign n29553 = n14284 ^ n2345 ;
  assign n29554 = n29553 ^ n12795 ;
  assign n29555 = n29554 ^ n315 ;
  assign n29556 = n29552 & ~n29555 ;
  assign n29557 = ~n14999 & n29556 ;
  assign n29541 = n29474 ^ n29371 ;
  assign n29542 = n29475 & ~n29541 ;
  assign n29543 = n29542 ^ x23 ;
  assign n29558 = n29557 ^ n29543 ;
  assign n29533 = n24700 ^ n24079 ;
  assign n29534 = n29533 ^ n24700 ;
  assign n29535 = x30 & n29534 ;
  assign n29536 = n29535 ^ n24700 ;
  assign n29537 = ~n3520 & ~n29536 ;
  assign n29521 = n25320 ^ n20834 ;
  assign n29520 = n25320 ^ n24079 ;
  assign n29522 = n29521 ^ n29520 ;
  assign n29525 = ~x30 & n29522 ;
  assign n29526 = n29525 ^ n29521 ;
  assign n29527 = ~n3520 & n29526 ;
  assign n29528 = n29527 ^ n25320 ;
  assign n29529 = n29528 ^ n24700 ;
  assign n29538 = n29537 ^ n29529 ;
  assign n29539 = ~x31 & ~n29538 ;
  assign n29540 = n29539 ^ n29528 ;
  assign n29559 = n29558 ^ n29540 ;
  assign n29517 = n29464 ^ n29461 ;
  assign n29518 = n29477 & ~n29517 ;
  assign n29519 = n29518 ^ n29464 ;
  assign n29560 = n29559 ^ n29519 ;
  assign n29498 = n831 & ~n24980 ;
  assign n29497 = n3484 & n25043 ;
  assign n29499 = n29498 ^ n29497 ;
  assign n29500 = n29499 ^ n651 ;
  assign n29503 = n25287 ^ n653 ;
  assign n29504 = n29503 ^ x28 ;
  assign n29505 = n29504 ^ n25287 ;
  assign n29501 = n29499 ^ x29 ;
  assign n29502 = n29501 ^ n653 ;
  assign n29506 = n29505 ^ n29502 ;
  assign n29507 = n29506 ^ n29502 ;
  assign n29509 = ~n25304 & ~n29507 ;
  assign n29510 = ~x28 & n29509 ;
  assign n29513 = n29510 ^ n29509 ;
  assign n29508 = n29507 ^ n29506 ;
  assign n29511 = n29510 ^ n25287 ;
  assign n29512 = n29508 & n29511 ;
  assign n29514 = n29513 ^ n29512 ;
  assign n29515 = n29514 ^ n653 ;
  assign n29516 = ~n29500 & ~n29515 ;
  assign n29561 = n29560 ^ n29516 ;
  assign n29495 = n12861 & n25703 ;
  assign n29491 = n29482 ^ n29450 ;
  assign n29492 = ~n29479 & ~n29491 ;
  assign n29493 = n29492 ^ n29482 ;
  assign n29494 = n29493 ^ x26 ;
  assign n29496 = n29495 ^ n29494 ;
  assign n29562 = n29561 ^ n29496 ;
  assign n29489 = ~n29439 & n29483 ;
  assign n29488 = ~n29429 & n29432 ;
  assign n29490 = n29489 ^ n29488 ;
  assign n29563 = n29562 ^ n29490 ;
  assign n29566 = n29565 ^ n29563 ;
  assign n29568 = n29567 ^ n29566 ;
  assign n29644 = ~n29566 & n29567 ;
  assign n29639 = n29519 ^ n29516 ;
  assign n29640 = ~n29560 & n29639 ;
  assign n29641 = n29640 ^ n29516 ;
  assign n29626 = n482 ^ n372 ;
  assign n29625 = n351 ^ n349 ;
  assign n29627 = n29626 ^ n29625 ;
  assign n29628 = n24675 ^ n473 ;
  assign n29629 = n29628 ^ n717 ;
  assign n29630 = n29627 & ~n29629 ;
  assign n29631 = ~n12697 & n29630 ;
  assign n29623 = n29543 ^ n29540 ;
  assign n29624 = ~n29558 & n29623 ;
  assign n29632 = n29631 ^ n29624 ;
  assign n29604 = n24700 ^ x31 ;
  assign n29605 = n29604 ^ n33 ;
  assign n29606 = n29605 ^ n3724 ;
  assign n29633 = n29632 ^ n29606 ;
  assign n29610 = n29606 ^ n24980 ;
  assign n29611 = n29610 ^ n29606 ;
  assign n29612 = ~n33 & ~n29611 ;
  assign n29613 = n29612 ^ n29606 ;
  assign n29614 = ~x31 & n29613 ;
  assign n29634 = n29633 ^ n29614 ;
  assign n29617 = n25517 ^ n24079 ;
  assign n29620 = n35 & n29617 ;
  assign n29621 = n29620 ^ n24079 ;
  assign n29622 = n4851 & ~n29621 ;
  assign n29635 = n29634 ^ n29622 ;
  assign n29607 = n29606 ^ x31 ;
  assign n29615 = n29604 & ~n29614 ;
  assign n29616 = n29607 & n29615 ;
  assign n29636 = n29635 ^ n29616 ;
  assign n29637 = n29636 ^ x26 ;
  assign n29601 = n3484 & ~n25287 ;
  assign n29594 = n25693 ^ x29 ;
  assign n29595 = n29594 ^ x28 ;
  assign n29596 = n29595 ^ n25693 ;
  assign n29597 = n25705 & ~n29596 ;
  assign n29598 = n29597 ^ n25693 ;
  assign n29599 = n650 & n29598 ;
  assign n29600 = n29599 ^ x29 ;
  assign n29602 = n29601 ^ n29600 ;
  assign n29593 = n831 & n25043 ;
  assign n29603 = n29602 ^ n29593 ;
  assign n29638 = n29637 ^ n29603 ;
  assign n29642 = n29641 ^ n29638 ;
  assign n29569 = n29488 ^ n29433 ;
  assign n29571 = ~n29483 & ~n29569 ;
  assign n29573 = ~n29488 & n29489 ;
  assign n29574 = ~n29426 & n29573 ;
  assign n29572 = ~n29488 & ~n29562 ;
  assign n29575 = n29574 ^ n29572 ;
  assign n29576 = n29575 ^ n29574 ;
  assign n29577 = n29571 & n29576 ;
  assign n29578 = n29577 ^ n29575 ;
  assign n29579 = n29439 ^ n29426 ;
  assign n29580 = n29572 ^ n29483 ;
  assign n29581 = n29580 ^ n29439 ;
  assign n29582 = n29579 & ~n29581 ;
  assign n29583 = n29582 ^ n29439 ;
  assign n29584 = ~n29578 & ~n29583 ;
  assign n29586 = n29584 ^ n29578 ;
  assign n29570 = n29562 & ~n29569 ;
  assign n29585 = n29570 & n29584 ;
  assign n29587 = n29586 ^ n29585 ;
  assign n29589 = n29587 ^ n29561 ;
  assign n29588 = n29587 ^ n29493 ;
  assign n29590 = n29589 ^ n29588 ;
  assign n29591 = n29496 & n29590 ;
  assign n29592 = n29591 ^ n29589 ;
  assign n29643 = n29642 ^ n29592 ;
  assign n29645 = n29644 ^ n29643 ;
  assign n29683 = n831 & ~n25287 ;
  assign n29682 = n3481 & n25725 ;
  assign n29684 = n29683 ^ n29682 ;
  assign n29679 = n29631 ^ n29557 ;
  assign n29680 = ~n29624 & ~n29679 ;
  assign n29673 = x29 ^ x26 ;
  assign n29672 = n3940 ^ n477 ;
  assign n29674 = n29673 ^ n29672 ;
  assign n29675 = n29674 ^ n29557 ;
  assign n29676 = n29675 ^ n29631 ;
  assign n29660 = x30 & ~n25251 ;
  assign n29661 = n29660 ^ n24980 ;
  assign n29662 = n28746 & ~n29661 ;
  assign n29663 = n29662 ^ x30 ;
  assign n29677 = n29676 ^ n29663 ;
  assign n29664 = n29663 ^ n25043 ;
  assign n29667 = n29664 ^ n25008 ;
  assign n29668 = n29667 ^ n29664 ;
  assign n29669 = x31 & ~n29668 ;
  assign n29670 = n29669 ^ n29664 ;
  assign n29671 = n3520 & n29670 ;
  assign n29678 = n29677 ^ n29671 ;
  assign n29681 = n29680 ^ n29678 ;
  assign n29685 = n29684 ^ n29681 ;
  assign n29654 = n29603 ^ x26 ;
  assign n29653 = n29641 ^ n29632 ;
  assign n29655 = n29654 ^ n29653 ;
  assign n29656 = n29636 & n29655 ;
  assign n29686 = n29685 ^ n29656 ;
  assign n29650 = n29641 ^ n29603 ;
  assign n29651 = n29641 ^ x26 ;
  assign n29652 = n29650 & n29651 ;
  assign n29687 = n29686 ^ n29652 ;
  assign n29647 = n29642 ^ n29587 ;
  assign n29648 = ~n29592 & n29647 ;
  assign n29646 = n29643 & ~n29644 ;
  assign n29649 = n29648 ^ n29646 ;
  assign n29688 = n29687 ^ n29649 ;
  assign y0 = ~n24994 ;
  assign y1 = ~n25263 ;
  assign y2 = ~n25515 ;
  assign y3 = n25715 ;
  assign y4 = n25902 ;
  assign y5 = ~n26100 ;
  assign y6 = ~n26292 ;
  assign y7 = ~n26509 ;
  assign y8 = ~n26706 ;
  assign y9 = n26918 ;
  assign y10 = n27096 ;
  assign y11 = ~n27305 ;
  assign y12 = n27495 ;
  assign y13 = ~n27674 ;
  assign y14 = n27823 ;
  assign y15 = ~n27993 ;
  assign y16 = ~n28136 ;
  assign y17 = ~n28286 ;
  assign y18 = n28418 ;
  assign y19 = n28578 ;
  assign y20 = ~n28711 ;
  assign y21 = ~n28819 ;
  assign y22 = ~n28918 ;
  assign y23 = n29025 ;
  assign y24 = n29126 ;
  assign y25 = ~n29250 ;
  assign y26 = ~n29333 ;
  assign y27 = n29404 ;
  assign y28 = n29487 ;
  assign y29 = ~n29568 ;
  assign y30 = n29645 ;
  assign y31 = ~n29688 ;
endmodule
