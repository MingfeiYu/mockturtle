module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n137 , n139 , n140 , n141 , n142 , n143 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n159 , n160 , n163 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n176 , n177 , n178 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n191 , n192 , n193 , n195 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n208 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n257 , n258 , n259 , n262 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n275 , n276 , n277 , n278 , n279 , n281 , n282 , n283 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n316 , n317 , n318 , n319 , n320 , n322 , n323 , n324 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n362 , n363 , n364 , n366 , n367 , n368 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n430 , n431 , n432 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n485 , n486 , n487 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n545 , n546 , n547 , n548 , n549 , n550 , n552 , n553 , n554 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n591 , n592 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n620 , n621 , n622 , n623 , n624 , n626 , n627 , n628 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n689 , n690 , n691 , n692 , n693 , n695 , n696 , n697 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n730 , n731 , n732 , n733 , n734 , n735 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n762 , n763 , n764 , n765 , n766 , n768 , n769 , n770 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n846 , n847 , n848 , n850 , n851 , n852 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n927 , n928 , n929 , n930 , n931 , n933 , n934 , n935 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n969 , n971 , n972 , n973 , n974 , n975 , n976 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1019 , n1020 , n1021 , n1023 , n1024 , n1025 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1109 , n1110 , n1111 , n1113 , n1114 , n1115 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1200 , n1201 , n1202 , n1204 , n1205 , n1206 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1244 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1296 , n1297 , n1298 , n1300 , n1301 , n1302 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1553 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1898 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3217 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3732 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4298 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4888 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6208 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6953 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7686 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8395 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8497 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8918 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8969 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9284 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9383 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9860 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16657 , n16658 , n16659 , n16660 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16823 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16850 , n16852 , n16853 , n16854 , n16855 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18034 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18838 , n18839 , n18840 , n18841 , n18842 , n18844 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18870 , n18871 , n18872 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18885 , n18886 , n18887 , n18889 , n18890 , n18891 , n18892 , n18893 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19275 , n19276 , n19277 , n19278 , n19279 , n19282 , n19283 , n19284 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19299 , n19300 , n19301 , n19302 , n19303 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19409 , n19410 , n19411 , n19413 , n19415 , n19417 , n19419 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19445 , n19446 , n19447 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19460 , n19461 , n19462 , n19464 , n19465 , n19466 , n19467 , n19468 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19780 , n19781 , n19782 , n19783 , n19784 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19843 , n19847 , n19848 , n19849 , n19850 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19868 , n19869 , n19870 , n19871 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19884 , n19885 , n19886 , n19887 , n19888 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19993 , n19994 , n19995 , n20001 , n20002 , n20003 , n20004 , n20005 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20084 , n20085 , n20086 , n20087 , n20089 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20319 , n20321 , n20322 , n20323 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20347 , n20348 , n20349 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20402 , n20403 , n20404 , n20406 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20416 , n20417 , n20418 , n20420 , n20422 , n20424 , n20426 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20452 , n20453 , n20454 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20467 , n20468 , n20469 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20600 , n20602 , n20603 , n20604 , n20606 , n20607 , n20609 , n20610 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20651 , n20652 , n20653 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20833 , n20834 , n20835 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 ;
  assign n129 = x0 & x64 ;
  assign n131 = x0 & x65 ;
  assign n130 = x1 & x64 ;
  assign n132 = n131 ^ n130 ;
  assign n142 = x1 & x65 ;
  assign n145 = n142 ^ x66 ;
  assign n146 = x64 & ~n145 ;
  assign n147 = n146 ^ x66 ;
  assign n148 = x0 & n147 ;
  assign n139 = x0 & ~x66 ;
  assign n140 = n139 ^ x2 ;
  assign n141 = x64 & n140 ;
  assign n143 = n142 ^ n141 ;
  assign n149 = n148 ^ n143 ;
  assign n151 = ~x64 & ~x65 ;
  assign n176 = ~x66 & n151 ;
  assign n177 = n176 ^ x64 ;
  assign n178 = x2 & ~n177 ;
  assign n181 = ~x0 & ~n142 ;
  assign n182 = n178 & n181 ;
  assign n172 = x3 & x64 ;
  assign n173 = n172 ^ x2 ;
  assign n180 = n178 ^ n173 ;
  assign n183 = n182 ^ n180 ;
  assign n166 = x2 & x65 ;
  assign n167 = n166 ^ x66 ;
  assign n168 = ~x1 & n167 ;
  assign n152 = n151 ^ x64 ;
  assign n153 = n152 ^ x65 ;
  assign n154 = ~x66 & n153 ;
  assign n150 = x65 & x66 ;
  assign n155 = n154 ^ n150 ;
  assign n10145 = x2 ^ x1 ;
  assign n159 = n155 & n10145 ;
  assign n157 = x67 ^ x1 ;
  assign n160 = n159 ^ n157 ;
  assign n137 = x66 ^ x2 ;
  assign n163 = n160 ^ n137 ;
  assign n169 = n168 ^ n163 ;
  assign n170 = ~x0 & n169 ;
  assign n171 = n170 ^ n160 ;
  assign n184 = n183 ^ n171 ;
  assign n217 = n171 & n183 ;
  assign n211 = x2 & x66 ;
  assign n212 = n211 ^ x67 ;
  assign n213 = ~x1 & n212 ;
  assign n186 = x67 & ~n154 ;
  assign n185 = ~x67 & ~n150 ;
  assign n187 = n186 ^ n185 ;
  assign n191 = n187 & n10145 ;
  assign n189 = x68 ^ x1 ;
  assign n192 = n191 ^ n189 ;
  assign n156 = x67 ^ x2 ;
  assign n208 = n192 ^ n156 ;
  assign n214 = n213 ^ n208 ;
  assign n215 = ~x0 & n214 ;
  assign n201 = x65 ^ x3 ;
  assign n202 = x3 ^ x2 ;
  assign n203 = ~n201 & n202 ;
  assign n197 = x2 & x3 ;
  assign n198 = n197 ^ x4 ;
  assign n199 = ~x64 & n198 ;
  assign n193 = x4 ^ x2 ;
  assign n200 = n199 ^ n193 ;
  assign n204 = n203 ^ n200 ;
  assign n205 = n204 ^ n192 ;
  assign n216 = n215 ^ n205 ;
  assign n218 = n217 ^ n216 ;
  assign n259 = x1 ^ x0 ;
  assign n265 = x2 & x67 ;
  assign n266 = n265 ^ x68 ;
  assign n267 = ~n259 & n266 ;
  assign n252 = ~x68 & ~n186 ;
  assign n251 = x68 & ~n185 ;
  assign n253 = n252 ^ n251 ;
  assign n257 = n253 & n10145 ;
  assign n255 = x69 ^ x1 ;
  assign n258 = n257 ^ n255 ;
  assign n188 = x68 ^ x2 ;
  assign n262 = n258 ^ n188 ;
  assign n268 = n267 ^ n262 ;
  assign n269 = ~x0 & n268 ;
  assign n270 = n269 ^ n258 ;
  assign n247 = x66 & n202 ;
  assign n233 = x5 ^ x4 ;
  assign n234 = n202 & ~n233 ;
  assign n235 = n234 ^ n202 ;
  assign n243 = x65 & n235 ;
  assign n236 = x5 ^ x3 ;
  assign n237 = ~n202 & n236 ;
  assign n238 = n233 & n237 ;
  assign n244 = n243 ^ n238 ;
  assign n245 = ~x64 & n244 ;
  assign n246 = n245 ^ n238 ;
  assign n248 = n247 ^ n246 ;
  assign n195 = x4 ^ x3 ;
  assign n231 = n195 & ~n202 ;
  assign n232 = x65 & n231 ;
  assign n249 = n248 ^ n232 ;
  assign n222 = n193 ^ x65 ;
  assign n223 = ~x64 & ~n222 ;
  assign n224 = n223 ^ n193 ;
  assign n225 = n202 ^ x64 ;
  assign n226 = n225 ^ x5 ;
  assign n227 = ~n224 & ~n226 ;
  assign n228 = n227 ^ x64 ;
  assign n229 = x5 & ~n228 ;
  assign n230 = n229 ^ x5 ;
  assign n250 = n249 ^ n230 ;
  assign n271 = n270 ^ n250 ;
  assign n219 = n217 ^ n204 ;
  assign n220 = n216 & n219 ;
  assign n221 = n220 ^ n204 ;
  assign n272 = n271 ^ n221 ;
  assign n307 = n270 ^ n221 ;
  assign n308 = n271 & n307 ;
  assign n309 = n308 ^ n270 ;
  assign n298 = x65 & n238 ;
  assign n297 = x67 & n234 ;
  assign n299 = n298 ^ n297 ;
  assign n300 = n299 ^ x5 ;
  assign n295 = n155 ^ x67 ;
  assign n296 = n235 & ~n295 ;
  assign n301 = n300 ^ n296 ;
  assign n294 = x66 & n231 ;
  assign n302 = n301 ^ n294 ;
  assign n293 = n229 & ~n249 ;
  assign n303 = n302 ^ n293 ;
  assign n291 = x6 ^ x5 ;
  assign n292 = x64 & n291 ;
  assign n304 = n303 ^ n292 ;
  assign n276 = x69 & ~n252 ;
  assign n275 = ~x69 & ~n251 ;
  assign n277 = n276 ^ n275 ;
  assign n281 = n277 & n10145 ;
  assign n279 = x70 ^ x1 ;
  assign n282 = n281 ^ n279 ;
  assign n305 = n304 ^ n282 ;
  assign n286 = x2 & x68 ;
  assign n287 = n286 ^ x69 ;
  assign n288 = ~x1 & n287 ;
  assign n254 = x69 ^ x2 ;
  assign n283 = n282 ^ n254 ;
  assign n289 = n288 ^ n283 ;
  assign n290 = ~x0 & n289 ;
  assign n306 = n305 ^ n290 ;
  assign n310 = n309 ^ n306 ;
  assign n354 = x67 & n231 ;
  assign n351 = n187 ^ x68 ;
  assign n352 = n235 & ~n351 ;
  assign n347 = x66 & n238 ;
  assign n346 = x68 & n234 ;
  assign n348 = n347 ^ n346 ;
  assign n349 = n348 ^ x5 ;
  assign n344 = ~x7 & x64 ;
  assign n335 = ~x5 & ~x6 ;
  assign n336 = n335 ^ n291 ;
  assign n341 = x65 & ~n335 ;
  assign n342 = n341 ^ x64 ;
  assign n343 = n336 & n342 ;
  assign n345 = n344 ^ n343 ;
  assign n350 = n349 ^ n345 ;
  assign n353 = n352 ^ n350 ;
  assign n355 = n354 ^ n353 ;
  assign n332 = ~n293 & n302 ;
  assign n333 = ~n292 & n332 ;
  assign n334 = n333 ^ n302 ;
  assign n356 = n355 ^ n334 ;
  assign n317 = ~x70 & ~n276 ;
  assign n316 = x70 & ~n275 ;
  assign n318 = n317 ^ n316 ;
  assign n322 = n318 & n10145 ;
  assign n320 = x71 ^ x1 ;
  assign n323 = n322 ^ n320 ;
  assign n357 = n356 ^ n323 ;
  assign n327 = x2 & x69 ;
  assign n328 = n327 ^ x70 ;
  assign n329 = ~x1 & n328 ;
  assign n278 = x70 ^ x2 ;
  assign n324 = n323 ^ n278 ;
  assign n330 = n329 ^ n324 ;
  assign n331 = ~x0 & n330 ;
  assign n358 = n357 ^ n331 ;
  assign n311 = n309 ^ n304 ;
  assign n312 = ~n306 & n311 ;
  assign n313 = n312 ^ n309 ;
  assign n359 = n358 ^ n313 ;
  assign n413 = n356 ^ n313 ;
  assign n414 = n358 & n413 ;
  assign n415 = n414 ^ n356 ;
  assign n407 = n345 ^ n334 ;
  assign n408 = n355 & n407 ;
  assign n409 = n408 ^ n345 ;
  assign n405 = x68 & n231 ;
  assign n395 = ~n292 & ~n345 ;
  assign n390 = x7 ^ x6 ;
  assign n391 = ~n291 & n390 ;
  assign n392 = x65 & n391 ;
  assign n383 = x8 ^ x7 ;
  assign n384 = n291 & ~n383 ;
  assign n385 = n384 ^ n291 ;
  assign n388 = ~n152 & n385 ;
  assign n387 = x66 & n291 ;
  assign n389 = n388 ^ n387 ;
  assign n393 = n392 ^ n389 ;
  assign n382 = n335 & n344 ;
  assign n394 = n393 ^ n382 ;
  assign n396 = n395 ^ n394 ;
  assign n397 = n396 ^ n393 ;
  assign n380 = n344 ^ x64 ;
  assign n381 = ~n336 & n380 ;
  assign n398 = n397 ^ n381 ;
  assign n399 = ~x8 & ~n398 ;
  assign n400 = n399 ^ n396 ;
  assign n401 = n400 ^ x5 ;
  assign n379 = x67 & n238 ;
  assign n402 = n401 ^ n379 ;
  assign n378 = x69 & n234 ;
  assign n403 = n402 ^ n378 ;
  assign n376 = n253 ^ x69 ;
  assign n377 = n235 & ~n376 ;
  assign n404 = n403 ^ n377 ;
  assign n406 = n405 ^ n404 ;
  assign n410 = n409 ^ n406 ;
  assign n360 = x71 ^ x70 ;
  assign n362 = n318 & n360 ;
  assign n366 = ~n362 & n10145 ;
  assign n364 = x72 ^ x1 ;
  assign n367 = n366 ^ n364 ;
  assign n411 = n410 ^ n367 ;
  assign n371 = x2 & x70 ;
  assign n372 = n371 ^ x71 ;
  assign n373 = ~x1 & n372 ;
  assign n319 = x71 ^ x2 ;
  assign n368 = n367 ^ n319 ;
  assign n374 = n373 ^ n368 ;
  assign n375 = ~x0 & n374 ;
  assign n412 = n411 ^ n375 ;
  assign n416 = n415 ^ n412 ;
  assign n468 = x69 & n231 ;
  assign n454 = x8 ^ x6 ;
  assign n455 = ~n291 & n454 ;
  assign n456 = n383 & n455 ;
  assign n457 = x65 & n456 ;
  assign n453 = x67 & n384 ;
  assign n458 = n457 ^ n453 ;
  assign n459 = n458 ^ x8 ;
  assign n452 = ~n295 & n385 ;
  assign n460 = n459 ^ n452 ;
  assign n451 = x66 & n391 ;
  assign n461 = n460 ^ n451 ;
  assign n449 = x9 ^ x8 ;
  assign n450 = x64 & n449 ;
  assign n462 = n461 ^ n450 ;
  assign n447 = x8 & n396 ;
  assign n448 = ~n394 & n447 ;
  assign n463 = n462 ^ n448 ;
  assign n464 = n463 ^ x5 ;
  assign n446 = x68 & n238 ;
  assign n465 = n464 ^ n446 ;
  assign n445 = x70 & n234 ;
  assign n466 = n465 ^ n445 ;
  assign n443 = n277 ^ x70 ;
  assign n444 = n235 & ~n443 ;
  assign n467 = n466 ^ n444 ;
  assign n469 = n468 ^ n467 ;
  assign n440 = n409 ^ n400 ;
  assign n441 = n406 & ~n440 ;
  assign n442 = n441 ^ n409 ;
  assign n470 = n469 ^ n442 ;
  assign n422 = x71 & ~x72 ;
  assign n425 = ~n317 & n422 ;
  assign n420 = x72 ^ x71 ;
  assign n423 = n422 ^ n420 ;
  assign n424 = ~n316 & n423 ;
  assign n426 = n425 ^ n424 ;
  assign n430 = ~n426 & n10145 ;
  assign n428 = x73 ^ x1 ;
  assign n431 = n430 ^ n428 ;
  assign n471 = n470 ^ n431 ;
  assign n435 = x2 & x71 ;
  assign n436 = n435 ^ x72 ;
  assign n437 = ~x1 & n436 ;
  assign n363 = x72 ^ x2 ;
  assign n432 = n431 ^ n363 ;
  assign n438 = n437 ^ n432 ;
  assign n439 = ~x0 & n438 ;
  assign n472 = n471 ^ n439 ;
  assign n417 = n415 ^ n410 ;
  assign n418 = n412 & ~n417 ;
  assign n419 = n418 ^ n415 ;
  assign n473 = n472 ^ n419 ;
  assign n536 = n470 ^ n419 ;
  assign n537 = n472 & n536 ;
  assign n538 = n537 ^ n470 ;
  assign n530 = n463 ^ n442 ;
  assign n531 = n469 & n530 ;
  assign n532 = n531 ^ n463 ;
  assign n528 = x70 & n231 ;
  assign n507 = ~n448 & ~n450 ;
  assign n521 = n461 & n507 ;
  assign n514 = ~x8 & ~x9 ;
  assign n515 = n514 ^ n449 ;
  assign n516 = n515 ^ x10 ;
  assign n517 = ~x64 & ~n516 ;
  assign n508 = x65 ^ x9 ;
  assign n511 = x65 ^ x8 ;
  assign n512 = ~n508 & n511 ;
  assign n509 = x10 ^ x8 ;
  assign n513 = n512 ^ n509 ;
  assign n518 = n517 ^ n513 ;
  assign n519 = n518 ^ n461 ;
  assign n522 = n521 ^ n519 ;
  assign n502 = x66 & n456 ;
  assign n501 = x68 & n384 ;
  assign n503 = n502 ^ n501 ;
  assign n504 = n503 ^ x8 ;
  assign n500 = ~n351 & n385 ;
  assign n505 = n504 ^ n500 ;
  assign n499 = x67 & n391 ;
  assign n506 = n505 ^ n499 ;
  assign n523 = n522 ^ n506 ;
  assign n524 = n523 ^ x5 ;
  assign n498 = x69 & n238 ;
  assign n525 = n524 ^ n498 ;
  assign n497 = x71 & n234 ;
  assign n526 = n525 ^ n497 ;
  assign n495 = n318 ^ x71 ;
  assign n496 = n235 & ~n495 ;
  assign n527 = n526 ^ n496 ;
  assign n529 = n528 ^ n527 ;
  assign n533 = n532 ^ n529 ;
  assign n478 = n425 ^ x72 ;
  assign n479 = x73 & n478 ;
  assign n480 = n479 ^ x73 ;
  assign n476 = x72 & ~x73 ;
  assign n477 = ~n424 & n476 ;
  assign n481 = n480 ^ n477 ;
  assign n485 = ~n481 & n10145 ;
  assign n483 = x74 ^ x1 ;
  assign n486 = n485 ^ n483 ;
  assign n534 = n533 ^ n486 ;
  assign n490 = x2 & x72 ;
  assign n491 = n490 ^ x73 ;
  assign n492 = ~x1 & n491 ;
  assign n427 = x73 ^ x2 ;
  assign n487 = n486 ^ n427 ;
  assign n493 = n492 ^ n487 ;
  assign n494 = ~x0 & n493 ;
  assign n535 = n534 ^ n494 ;
  assign n539 = n538 ^ n535 ;
  assign n612 = x71 & n231 ;
  assign n604 = n518 ^ n506 ;
  assign n605 = n522 & n604 ;
  assign n606 = n605 ^ n518 ;
  assign n602 = x68 & n391 ;
  assign n575 = ~x10 & ~n449 ;
  assign n584 = n575 ^ n514 ;
  assign n594 = n584 ^ n449 ;
  assign n595 = x64 & ~n594 ;
  assign n596 = ~x11 & n595 ;
  assign n588 = ~n450 & ~n518 ;
  assign n589 = x11 & n588 ;
  assign n591 = n589 ^ x11 ;
  assign n585 = x65 & n584 ;
  assign n576 = x11 ^ x10 ;
  assign n577 = n576 ^ n575 ;
  assign n574 = x11 & ~n449 ;
  assign n578 = n577 ^ n574 ;
  assign n579 = n578 ^ n449 ;
  assign n582 = ~n152 & ~n579 ;
  assign n581 = x66 & n449 ;
  assign n583 = n582 ^ n581 ;
  assign n586 = n585 ^ n583 ;
  assign n572 = ~x10 & x64 ;
  assign n573 = n514 & n572 ;
  assign n587 = n586 ^ n573 ;
  assign n592 = n591 ^ n587 ;
  assign n597 = n596 ^ n592 ;
  assign n598 = n597 ^ x8 ;
  assign n571 = x67 & n456 ;
  assign n599 = n598 ^ n571 ;
  assign n570 = x69 & n384 ;
  assign n600 = n599 ^ n570 ;
  assign n569 = ~n376 & n385 ;
  assign n601 = n600 ^ n569 ;
  assign n603 = n602 ^ n601 ;
  assign n607 = n606 ^ n603 ;
  assign n608 = n607 ^ x5 ;
  assign n568 = x70 & n238 ;
  assign n609 = n608 ^ n568 ;
  assign n567 = x72 & n234 ;
  assign n610 = n609 ^ n567 ;
  assign n565 = n362 ^ x72 ;
  assign n566 = n235 & n565 ;
  assign n611 = n610 ^ n566 ;
  assign n613 = n612 ^ n611 ;
  assign n562 = n532 ^ n523 ;
  assign n563 = ~n529 & n562 ;
  assign n564 = n563 ^ n532 ;
  assign n614 = n613 ^ n564 ;
  assign n547 = ~x74 & ~n479 ;
  assign n545 = n477 ^ x73 ;
  assign n546 = x74 & n545 ;
  assign n548 = n547 ^ n546 ;
  assign n552 = n548 & n10145 ;
  assign n550 = x75 ^ x1 ;
  assign n553 = n552 ^ n550 ;
  assign n615 = n614 ^ n553 ;
  assign n557 = x2 & x73 ;
  assign n558 = n557 ^ x74 ;
  assign n559 = ~x1 & n558 ;
  assign n482 = x74 ^ x2 ;
  assign n554 = n553 ^ n482 ;
  assign n560 = n559 ^ n554 ;
  assign n561 = ~x0 & n560 ;
  assign n616 = n615 ^ n561 ;
  assign n540 = n538 ^ n533 ;
  assign n541 = ~n535 & n540 ;
  assign n542 = n541 ^ n538 ;
  assign n617 = n616 ^ n542 ;
  assign n680 = n614 ^ n542 ;
  assign n681 = n616 & n680 ;
  assign n682 = n681 ^ n614 ;
  assign n674 = n607 ^ n564 ;
  assign n675 = n613 & n674 ;
  assign n676 = n675 ^ n607 ;
  assign n672 = x72 & n231 ;
  assign n661 = x68 & n456 ;
  assign n660 = x70 & n384 ;
  assign n662 = n661 ^ n660 ;
  assign n663 = n662 ^ x8 ;
  assign n659 = n385 & ~n443 ;
  assign n664 = n663 ^ n659 ;
  assign n658 = x69 & n391 ;
  assign n665 = n664 ^ n658 ;
  assign n649 = n574 ^ n515 ;
  assign n650 = n576 & ~n649 ;
  assign n651 = x65 & n650 ;
  assign n648 = x67 & ~n578 ;
  assign n652 = n651 ^ n648 ;
  assign n653 = n652 ^ x11 ;
  assign n647 = ~n295 & ~n579 ;
  assign n654 = n653 ^ n647 ;
  assign n646 = x66 & n584 ;
  assign n655 = n654 ^ n646 ;
  assign n644 = x12 ^ x11 ;
  assign n645 = x64 & n644 ;
  assign n656 = n655 ^ n645 ;
  assign n643 = ~n587 & n589 ;
  assign n657 = n656 ^ n643 ;
  assign n666 = n665 ^ n657 ;
  assign n640 = n606 ^ n597 ;
  assign n641 = ~n603 & n640 ;
  assign n642 = n641 ^ n606 ;
  assign n667 = n666 ^ n642 ;
  assign n668 = n667 ^ x5 ;
  assign n639 = x71 & n238 ;
  assign n669 = n668 ^ n639 ;
  assign n638 = x73 & n234 ;
  assign n670 = n669 ^ n638 ;
  assign n636 = n426 ^ x73 ;
  assign n637 = n235 & n636 ;
  assign n671 = n670 ^ n637 ;
  assign n673 = n672 ^ n671 ;
  assign n677 = n676 ^ n673 ;
  assign n621 = x75 & ~n547 ;
  assign n620 = ~x75 & ~n546 ;
  assign n622 = n621 ^ n620 ;
  assign n626 = n622 & n10145 ;
  assign n624 = x76 ^ x1 ;
  assign n627 = n626 ^ n624 ;
  assign n678 = n677 ^ n627 ;
  assign n631 = x2 & x74 ;
  assign n632 = n631 ^ x75 ;
  assign n633 = ~x1 & n632 ;
  assign n549 = x75 ^ x2 ;
  assign n628 = n627 ^ n549 ;
  assign n634 = n633 ^ n628 ;
  assign n635 = ~x0 & n634 ;
  assign n679 = n678 ^ n635 ;
  assign n683 = n682 ^ n679 ;
  assign n754 = x73 & n231 ;
  assign n746 = n665 ^ n642 ;
  assign n747 = n666 & n746 ;
  assign n748 = n747 ^ n665 ;
  assign n744 = x70 & n391 ;
  assign n723 = ~n643 & ~n645 ;
  assign n737 = n655 & n723 ;
  assign n733 = ~n152 & n644 ;
  assign n724 = x13 ^ x12 ;
  assign n725 = n724 ^ x65 ;
  assign n726 = n725 ^ x12 ;
  assign n727 = n726 ^ n724 ;
  assign n730 = n644 & n727 ;
  assign n731 = n730 ^ n724 ;
  assign n732 = x64 & n731 ;
  assign n734 = n733 ^ n732 ;
  assign n735 = n734 ^ n655 ;
  assign n738 = n737 ^ n735 ;
  assign n718 = x66 & n650 ;
  assign n717 = x68 & ~n578 ;
  assign n719 = n718 ^ n717 ;
  assign n720 = n719 ^ x11 ;
  assign n716 = ~n351 & ~n579 ;
  assign n721 = n720 ^ n716 ;
  assign n715 = x67 & n584 ;
  assign n722 = n721 ^ n715 ;
  assign n739 = n738 ^ n722 ;
  assign n740 = n739 ^ x8 ;
  assign n714 = x69 & n456 ;
  assign n741 = n740 ^ n714 ;
  assign n713 = x71 & n384 ;
  assign n742 = n741 ^ n713 ;
  assign n712 = n385 & ~n495 ;
  assign n743 = n742 ^ n712 ;
  assign n745 = n744 ^ n743 ;
  assign n749 = n748 ^ n745 ;
  assign n750 = n749 ^ x5 ;
  assign n711 = x72 & n238 ;
  assign n751 = n750 ^ n711 ;
  assign n710 = x74 & n234 ;
  assign n752 = n751 ^ n710 ;
  assign n708 = n481 ^ x74 ;
  assign n709 = n235 & n708 ;
  assign n753 = n752 ^ n709 ;
  assign n755 = n754 ^ n753 ;
  assign n705 = n676 ^ n667 ;
  assign n706 = ~n673 & n705 ;
  assign n707 = n706 ^ n676 ;
  assign n756 = n755 ^ n707 ;
  assign n690 = ~x76 & ~n621 ;
  assign n689 = x76 & ~n620 ;
  assign n691 = n690 ^ n689 ;
  assign n695 = n691 & n10145 ;
  assign n693 = x77 ^ x1 ;
  assign n696 = n695 ^ n693 ;
  assign n757 = n756 ^ n696 ;
  assign n700 = x2 & x75 ;
  assign n701 = n700 ^ x76 ;
  assign n702 = ~x1 & n701 ;
  assign n623 = x76 ^ x2 ;
  assign n697 = n696 ^ n623 ;
  assign n703 = n702 ^ n697 ;
  assign n704 = ~x0 & n703 ;
  assign n758 = n757 ^ n704 ;
  assign n684 = n682 ^ n677 ;
  assign n685 = ~n679 & n684 ;
  assign n686 = n685 ^ n682 ;
  assign n759 = n758 ^ n686 ;
  assign n837 = n756 ^ n686 ;
  assign n838 = n758 & n837 ;
  assign n839 = n838 ^ n756 ;
  assign n831 = n749 ^ n707 ;
  assign n832 = n755 & n831 ;
  assign n833 = n832 ^ n749 ;
  assign n829 = x74 & n231 ;
  assign n822 = x71 & n391 ;
  assign n814 = n734 ^ n722 ;
  assign n815 = n738 & n814 ;
  assign n816 = n815 ^ n734 ;
  assign n811 = n733 ^ x64 ;
  assign n812 = x14 & n811 ;
  assign n807 = x11 & x12 ;
  assign n808 = x13 & x64 ;
  assign n809 = n807 & n808 ;
  assign n801 = x67 & n650 ;
  assign n800 = x69 & ~n578 ;
  assign n802 = n801 ^ n800 ;
  assign n803 = n802 ^ x11 ;
  assign n799 = ~n376 & ~n579 ;
  assign n804 = n803 ^ n799 ;
  assign n798 = x68 & n584 ;
  assign n805 = n804 ^ n798 ;
  assign n795 = ~n644 & n724 ;
  assign n796 = x65 & n795 ;
  assign n788 = x14 ^ x13 ;
  assign n789 = n644 & ~n788 ;
  assign n790 = n789 ^ n644 ;
  assign n793 = ~n152 & n790 ;
  assign n792 = x66 & n644 ;
  assign n794 = n793 ^ n792 ;
  assign n797 = n796 ^ n794 ;
  assign n806 = n805 ^ n797 ;
  assign n810 = n809 ^ n806 ;
  assign n813 = n812 ^ n810 ;
  assign n817 = n816 ^ n813 ;
  assign n818 = n817 ^ x8 ;
  assign n787 = x70 & n456 ;
  assign n819 = n818 ^ n787 ;
  assign n786 = x72 & n384 ;
  assign n820 = n819 ^ n786 ;
  assign n785 = n385 & n565 ;
  assign n821 = n820 ^ n785 ;
  assign n823 = n822 ^ n821 ;
  assign n782 = n748 ^ n739 ;
  assign n783 = ~n745 & n782 ;
  assign n784 = n783 ^ n748 ;
  assign n824 = n823 ^ n784 ;
  assign n825 = n824 ^ x5 ;
  assign n781 = x73 & n238 ;
  assign n826 = n825 ^ n781 ;
  assign n780 = x75 & n234 ;
  assign n827 = n826 ^ n780 ;
  assign n778 = n548 ^ x75 ;
  assign n779 = n235 & ~n778 ;
  assign n828 = n827 ^ n779 ;
  assign n830 = n829 ^ n828 ;
  assign n834 = n833 ^ n830 ;
  assign n763 = x77 & ~n690 ;
  assign n762 = ~x77 & ~n689 ;
  assign n764 = n763 ^ n762 ;
  assign n768 = n764 & n10145 ;
  assign n766 = x78 ^ x1 ;
  assign n769 = n768 ^ n766 ;
  assign n835 = n834 ^ n769 ;
  assign n773 = x2 & x76 ;
  assign n774 = n773 ^ x77 ;
  assign n775 = ~x1 & n774 ;
  assign n692 = x77 ^ x2 ;
  assign n770 = n769 ^ n692 ;
  assign n776 = n775 ^ n770 ;
  assign n777 = ~x0 & n776 ;
  assign n836 = n835 ^ n777 ;
  assign n840 = n839 ^ n836 ;
  assign n915 = x75 & n231 ;
  assign n907 = n817 ^ n784 ;
  assign n908 = n823 & n907 ;
  assign n909 = n908 ^ n817 ;
  assign n905 = x72 & n391 ;
  assign n894 = x68 & n650 ;
  assign n893 = x70 & ~n578 ;
  assign n895 = n894 ^ n893 ;
  assign n896 = n895 ^ x11 ;
  assign n892 = ~n443 & ~n579 ;
  assign n897 = n896 ^ n892 ;
  assign n891 = x69 & n584 ;
  assign n898 = n897 ^ n891 ;
  assign n882 = x14 ^ x12 ;
  assign n883 = ~n644 & n882 ;
  assign n884 = n788 & n883 ;
  assign n885 = x65 & n884 ;
  assign n881 = x67 & n789 ;
  assign n886 = n885 ^ n881 ;
  assign n887 = n886 ^ x14 ;
  assign n880 = ~n295 & n790 ;
  assign n888 = n887 ^ n880 ;
  assign n879 = x66 & n795 ;
  assign n889 = n888 ^ n879 ;
  assign n875 = n811 ^ n809 ;
  assign n876 = x14 & ~n875 ;
  assign n877 = ~n797 & n876 ;
  assign n873 = x15 ^ x14 ;
  assign n874 = x64 & n873 ;
  assign n878 = n877 ^ n874 ;
  assign n890 = n889 ^ n878 ;
  assign n899 = n898 ^ n890 ;
  assign n870 = n816 ^ n805 ;
  assign n871 = ~n813 & n870 ;
  assign n872 = n871 ^ n816 ;
  assign n900 = n899 ^ n872 ;
  assign n901 = n900 ^ x8 ;
  assign n869 = x71 & n456 ;
  assign n902 = n901 ^ n869 ;
  assign n868 = x73 & n384 ;
  assign n903 = n902 ^ n868 ;
  assign n867 = n385 & n636 ;
  assign n904 = n903 ^ n867 ;
  assign n906 = n905 ^ n904 ;
  assign n910 = n909 ^ n906 ;
  assign n911 = n910 ^ x5 ;
  assign n866 = x74 & n238 ;
  assign n912 = n911 ^ n866 ;
  assign n865 = x76 & n234 ;
  assign n913 = n912 ^ n865 ;
  assign n863 = n622 ^ x76 ;
  assign n864 = n235 & ~n863 ;
  assign n914 = n913 ^ n864 ;
  assign n916 = n915 ^ n914 ;
  assign n860 = n833 ^ n824 ;
  assign n861 = ~n830 & n860 ;
  assign n862 = n861 ^ n833 ;
  assign n917 = n916 ^ n862 ;
  assign n844 = x78 ^ x77 ;
  assign n846 = n764 & n844 ;
  assign n850 = ~n846 & n10145 ;
  assign n848 = x79 ^ x1 ;
  assign n851 = n850 ^ n848 ;
  assign n918 = n917 ^ n851 ;
  assign n855 = x2 & x77 ;
  assign n856 = n855 ^ x78 ;
  assign n857 = ~x1 & n856 ;
  assign n765 = x78 ^ x2 ;
  assign n852 = n851 ^ n765 ;
  assign n858 = n857 ^ n852 ;
  assign n859 = ~x0 & n858 ;
  assign n919 = n918 ^ n859 ;
  assign n841 = n839 ^ n834 ;
  assign n842 = ~n836 & n841 ;
  assign n843 = n842 ^ n839 ;
  assign n920 = n919 ^ n843 ;
  assign n1010 = n917 ^ n843 ;
  assign n1011 = n919 & n1010 ;
  assign n1012 = n1011 ^ n917 ;
  assign n1004 = n910 ^ n862 ;
  assign n1005 = n916 & n1004 ;
  assign n1006 = n1005 ^ n910 ;
  assign n1002 = x76 & n231 ;
  assign n995 = x73 & n391 ;
  assign n987 = n898 ^ n872 ;
  assign n988 = n899 & n987 ;
  assign n989 = n988 ^ n898 ;
  assign n985 = x70 & n584 ;
  assign n964 = ~n874 & ~n877 ;
  assign n978 = n889 & n964 ;
  assign n971 = x14 & x15 ;
  assign n972 = n971 ^ x16 ;
  assign n973 = ~x64 & n972 ;
  assign n967 = x16 ^ x14 ;
  assign n974 = n973 ^ n967 ;
  assign n965 = x65 ^ x15 ;
  assign n966 = n873 & ~n965 ;
  assign n975 = n974 ^ n966 ;
  assign n976 = n975 ^ n889 ;
  assign n979 = n978 ^ n976 ;
  assign n959 = x66 & n884 ;
  assign n958 = x68 & n789 ;
  assign n960 = n959 ^ n958 ;
  assign n961 = n960 ^ x14 ;
  assign n957 = ~n351 & n790 ;
  assign n962 = n961 ^ n957 ;
  assign n956 = x67 & n795 ;
  assign n963 = n962 ^ n956 ;
  assign n980 = n979 ^ n963 ;
  assign n981 = n980 ^ x11 ;
  assign n955 = x69 & n650 ;
  assign n982 = n981 ^ n955 ;
  assign n954 = x71 & ~n578 ;
  assign n983 = n982 ^ n954 ;
  assign n953 = ~n495 & ~n579 ;
  assign n984 = n983 ^ n953 ;
  assign n986 = n985 ^ n984 ;
  assign n990 = n989 ^ n986 ;
  assign n991 = n990 ^ x8 ;
  assign n952 = x72 & n456 ;
  assign n992 = n991 ^ n952 ;
  assign n951 = x74 & n384 ;
  assign n993 = n992 ^ n951 ;
  assign n950 = n385 & n708 ;
  assign n994 = n993 ^ n950 ;
  assign n996 = n995 ^ n994 ;
  assign n947 = n909 ^ n900 ;
  assign n948 = ~n906 & n947 ;
  assign n949 = n948 ^ n909 ;
  assign n997 = n996 ^ n949 ;
  assign n998 = n997 ^ x5 ;
  assign n946 = x75 & n238 ;
  assign n999 = n998 ^ n946 ;
  assign n945 = x77 & n234 ;
  assign n1000 = n999 ^ n945 ;
  assign n943 = n691 ^ x77 ;
  assign n944 = n235 & ~n943 ;
  assign n1001 = n1000 ^ n944 ;
  assign n1003 = n1002 ^ n1001 ;
  assign n1007 = n1006 ^ n1003 ;
  assign n921 = x79 ^ x78 ;
  assign n927 = ~x79 & n764 ;
  assign n928 = n927 ^ n763 ;
  assign n929 = n921 & ~n928 ;
  assign n933 = ~n929 & n10145 ;
  assign n931 = x80 ^ x1 ;
  assign n934 = n933 ^ n931 ;
  assign n1008 = n1007 ^ n934 ;
  assign n938 = x2 & x78 ;
  assign n939 = n938 ^ x79 ;
  assign n940 = ~x1 & n939 ;
  assign n847 = x79 ^ x2 ;
  assign n935 = n934 ^ n847 ;
  assign n941 = n940 ^ n935 ;
  assign n942 = ~x0 & n941 ;
  assign n1009 = n1008 ^ n942 ;
  assign n1013 = n1012 ^ n1009 ;
  assign n1101 = x77 & n231 ;
  assign n1093 = n990 ^ n949 ;
  assign n1094 = n996 & n1093 ;
  assign n1095 = n1094 ^ n990 ;
  assign n1091 = x74 & n391 ;
  assign n1084 = x71 & n584 ;
  assign n1077 = x68 & n795 ;
  assign n969 = x16 ^ x15 ;
  assign n1068 = ~n873 & n969 ;
  assign n1069 = x65 & n1068 ;
  assign n1057 = x17 ^ x16 ;
  assign n1063 = n873 & ~n1057 ;
  assign n1064 = n1063 ^ n873 ;
  assign n1065 = ~n152 & n1064 ;
  assign n1062 = x66 & n873 ;
  assign n1066 = n1065 ^ n1062 ;
  assign n1067 = n1066 ^ x17 ;
  assign n1070 = n1069 ^ n1067 ;
  assign n1058 = x17 ^ x15 ;
  assign n1059 = ~n873 & n1058 ;
  assign n1060 = n1057 & n1059 ;
  assign n1061 = x64 & n1060 ;
  assign n1071 = n1070 ^ n1061 ;
  assign n1055 = ~n874 & ~n975 ;
  assign n1056 = x17 & n1055 ;
  assign n1072 = n1071 ^ n1056 ;
  assign n1073 = n1072 ^ x14 ;
  assign n1054 = x67 & n884 ;
  assign n1074 = n1073 ^ n1054 ;
  assign n1053 = x69 & n789 ;
  assign n1075 = n1074 ^ n1053 ;
  assign n1052 = ~n376 & n790 ;
  assign n1076 = n1075 ^ n1052 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1049 = n975 ^ n963 ;
  assign n1050 = n979 & n1049 ;
  assign n1051 = n1050 ^ n975 ;
  assign n1079 = n1078 ^ n1051 ;
  assign n1080 = n1079 ^ x11 ;
  assign n1048 = x70 & n650 ;
  assign n1081 = n1080 ^ n1048 ;
  assign n1047 = x72 & ~n578 ;
  assign n1082 = n1081 ^ n1047 ;
  assign n1046 = n565 & ~n579 ;
  assign n1083 = n1082 ^ n1046 ;
  assign n1085 = n1084 ^ n1083 ;
  assign n1043 = n989 ^ n980 ;
  assign n1044 = ~n986 & n1043 ;
  assign n1045 = n1044 ^ n989 ;
  assign n1086 = n1085 ^ n1045 ;
  assign n1087 = n1086 ^ x8 ;
  assign n1042 = x73 & n456 ;
  assign n1088 = n1087 ^ n1042 ;
  assign n1041 = x75 & n384 ;
  assign n1089 = n1088 ^ n1041 ;
  assign n1040 = n385 & ~n778 ;
  assign n1090 = n1089 ^ n1040 ;
  assign n1092 = n1091 ^ n1090 ;
  assign n1096 = n1095 ^ n1092 ;
  assign n1097 = n1096 ^ x5 ;
  assign n1039 = x76 & n238 ;
  assign n1098 = n1097 ^ n1039 ;
  assign n1038 = x78 & n234 ;
  assign n1099 = n1098 ^ n1038 ;
  assign n1036 = n764 ^ x78 ;
  assign n1037 = n235 & ~n1036 ;
  assign n1100 = n1099 ^ n1037 ;
  assign n1102 = n1101 ^ n1100 ;
  assign n1033 = n1006 ^ n997 ;
  assign n1034 = ~n1003 & n1033 ;
  assign n1035 = n1034 ^ n1006 ;
  assign n1103 = n1102 ^ n1035 ;
  assign n1017 = x80 ^ x79 ;
  assign n1019 = ~n929 & n1017 ;
  assign n1023 = ~n1019 & n10145 ;
  assign n1021 = x81 ^ x1 ;
  assign n1024 = n1023 ^ n1021 ;
  assign n1104 = n1103 ^ n1024 ;
  assign n1028 = x2 & x79 ;
  assign n1029 = n1028 ^ x80 ;
  assign n1030 = ~n259 & n1029 ;
  assign n930 = x80 ^ x2 ;
  assign n1025 = n1024 ^ n930 ;
  assign n1031 = n1030 ^ n1025 ;
  assign n1032 = ~x0 & n1031 ;
  assign n1105 = n1104 ^ n1032 ;
  assign n1014 = n1012 ^ n1007 ;
  assign n1015 = ~n1009 & n1014 ;
  assign n1016 = n1015 ^ n1012 ;
  assign n1106 = n1105 ^ n1016 ;
  assign n1191 = n1103 ^ n1016 ;
  assign n1192 = n1105 & n1191 ;
  assign n1193 = n1192 ^ n1103 ;
  assign n1185 = n1096 ^ n1035 ;
  assign n1186 = n1102 & n1185 ;
  assign n1187 = n1186 ^ n1096 ;
  assign n1183 = x78 & n231 ;
  assign n1176 = x75 & n391 ;
  assign n1168 = n1079 ^ n1045 ;
  assign n1169 = n1085 & n1168 ;
  assign n1170 = n1169 ^ n1079 ;
  assign n1166 = x72 & n584 ;
  assign n1159 = x69 & n795 ;
  assign n1148 = x65 & n1060 ;
  assign n1147 = x67 & n1063 ;
  assign n1149 = n1148 ^ n1147 ;
  assign n1150 = n1149 ^ x17 ;
  assign n1146 = ~n295 & n1064 ;
  assign n1151 = n1150 ^ n1146 ;
  assign n1145 = x66 & n1068 ;
  assign n1152 = n1151 ^ n1145 ;
  assign n1143 = x18 ^ x17 ;
  assign n1144 = x64 & n1143 ;
  assign n1153 = n1152 ^ n1144 ;
  assign n1142 = n1056 & n1071 ;
  assign n1154 = n1153 ^ n1142 ;
  assign n1155 = n1154 ^ x14 ;
  assign n1141 = x68 & n884 ;
  assign n1156 = n1155 ^ n1141 ;
  assign n1140 = x70 & n789 ;
  assign n1157 = n1156 ^ n1140 ;
  assign n1139 = ~n443 & n790 ;
  assign n1158 = n1157 ^ n1139 ;
  assign n1160 = n1159 ^ n1158 ;
  assign n1136 = n1072 ^ n1051 ;
  assign n1137 = n1078 & n1136 ;
  assign n1138 = n1137 ^ n1072 ;
  assign n1161 = n1160 ^ n1138 ;
  assign n1162 = n1161 ^ x11 ;
  assign n1135 = x71 & n650 ;
  assign n1163 = n1162 ^ n1135 ;
  assign n1134 = x73 & ~n578 ;
  assign n1164 = n1163 ^ n1134 ;
  assign n1133 = ~n579 & n636 ;
  assign n1165 = n1164 ^ n1133 ;
  assign n1167 = n1166 ^ n1165 ;
  assign n1171 = n1170 ^ n1167 ;
  assign n1172 = n1171 ^ x8 ;
  assign n1132 = x74 & n456 ;
  assign n1173 = n1172 ^ n1132 ;
  assign n1131 = x76 & n384 ;
  assign n1174 = n1173 ^ n1131 ;
  assign n1130 = n385 & ~n863 ;
  assign n1175 = n1174 ^ n1130 ;
  assign n1177 = n1176 ^ n1175 ;
  assign n1127 = n1095 ^ n1086 ;
  assign n1128 = ~n1092 & n1127 ;
  assign n1129 = n1128 ^ n1095 ;
  assign n1178 = n1177 ^ n1129 ;
  assign n1179 = n1178 ^ x5 ;
  assign n1126 = x77 & n238 ;
  assign n1180 = n1179 ^ n1126 ;
  assign n1125 = x79 & n234 ;
  assign n1181 = n1180 ^ n1125 ;
  assign n1123 = n846 ^ x79 ;
  assign n1124 = n235 & n1123 ;
  assign n1182 = n1181 ^ n1124 ;
  assign n1184 = n1183 ^ n1182 ;
  assign n1188 = n1187 ^ n1184 ;
  assign n1107 = x81 ^ x80 ;
  assign n1109 = ~n1019 & n1107 ;
  assign n1113 = ~n1109 & n10145 ;
  assign n1111 = x82 ^ x1 ;
  assign n1114 = n1113 ^ n1111 ;
  assign n1189 = n1188 ^ n1114 ;
  assign n1118 = x2 & x80 ;
  assign n1119 = n1118 ^ x81 ;
  assign n1120 = ~x1 & n1119 ;
  assign n1020 = x81 ^ x2 ;
  assign n1115 = n1114 ^ n1020 ;
  assign n1121 = n1120 ^ n1115 ;
  assign n1122 = ~x0 & n1121 ;
  assign n1190 = n1189 ^ n1122 ;
  assign n1194 = n1193 ^ n1190 ;
  assign n1288 = x79 & n231 ;
  assign n1280 = n1171 ^ n1129 ;
  assign n1281 = n1177 & n1280 ;
  assign n1282 = n1281 ^ n1171 ;
  assign n1278 = x76 & n391 ;
  assign n1271 = x73 & n584 ;
  assign n1263 = n1154 ^ n1138 ;
  assign n1264 = n1160 & n1263 ;
  assign n1265 = n1264 ^ n1154 ;
  assign n1261 = x70 & n795 ;
  assign n1254 = x67 & n1068 ;
  assign n1252 = ~n351 & n1064 ;
  assign n1246 = x17 & x18 ;
  assign n1247 = n1246 ^ x19 ;
  assign n1248 = ~x64 & n1247 ;
  assign n1242 = x19 ^ x17 ;
  assign n1249 = n1248 ^ n1242 ;
  assign n1240 = x65 ^ x18 ;
  assign n1241 = n1143 & ~n1240 ;
  assign n1250 = n1249 ^ n1241 ;
  assign n1237 = x66 & n1060 ;
  assign n1236 = x68 & n1063 ;
  assign n1238 = n1237 ^ n1236 ;
  assign n1239 = n1238 ^ x17 ;
  assign n1251 = n1250 ^ n1239 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1255 = n1254 ^ n1253 ;
  assign n1233 = ~n1144 & n1152 ;
  assign n1234 = ~n1142 & n1233 ;
  assign n1235 = n1234 ^ n1152 ;
  assign n1256 = n1255 ^ n1235 ;
  assign n1257 = n1256 ^ x14 ;
  assign n1232 = x69 & n884 ;
  assign n1258 = n1257 ^ n1232 ;
  assign n1231 = x71 & n789 ;
  assign n1259 = n1258 ^ n1231 ;
  assign n1230 = ~n495 & n790 ;
  assign n1260 = n1259 ^ n1230 ;
  assign n1262 = n1261 ^ n1260 ;
  assign n1266 = n1265 ^ n1262 ;
  assign n1267 = n1266 ^ x11 ;
  assign n1229 = x72 & n650 ;
  assign n1268 = n1267 ^ n1229 ;
  assign n1228 = x74 & ~n578 ;
  assign n1269 = n1268 ^ n1228 ;
  assign n1227 = ~n579 & n708 ;
  assign n1270 = n1269 ^ n1227 ;
  assign n1272 = n1271 ^ n1270 ;
  assign n1224 = n1170 ^ n1161 ;
  assign n1225 = ~n1167 & n1224 ;
  assign n1226 = n1225 ^ n1170 ;
  assign n1273 = n1272 ^ n1226 ;
  assign n1274 = n1273 ^ x8 ;
  assign n1223 = x75 & n456 ;
  assign n1275 = n1274 ^ n1223 ;
  assign n1222 = x77 & n384 ;
  assign n1276 = n1275 ^ n1222 ;
  assign n1221 = n385 & ~n943 ;
  assign n1277 = n1276 ^ n1221 ;
  assign n1279 = n1278 ^ n1277 ;
  assign n1283 = n1282 ^ n1279 ;
  assign n1284 = n1283 ^ x5 ;
  assign n1220 = x78 & n238 ;
  assign n1285 = n1284 ^ n1220 ;
  assign n1219 = x80 & n234 ;
  assign n1286 = n1285 ^ n1219 ;
  assign n1217 = n929 ^ x80 ;
  assign n1218 = n235 & n1217 ;
  assign n1287 = n1286 ^ n1218 ;
  assign n1289 = n1288 ^ n1287 ;
  assign n1214 = n1187 ^ n1178 ;
  assign n1215 = ~n1184 & n1214 ;
  assign n1216 = n1215 ^ n1187 ;
  assign n1290 = n1289 ^ n1216 ;
  assign n1198 = x82 ^ x81 ;
  assign n1200 = ~n1109 & n1198 ;
  assign n1204 = ~n1200 & n10145 ;
  assign n1202 = x83 ^ x1 ;
  assign n1205 = n1204 ^ n1202 ;
  assign n1291 = n1290 ^ n1205 ;
  assign n1209 = x2 & x81 ;
  assign n1210 = n1209 ^ x82 ;
  assign n1211 = ~x1 & n1210 ;
  assign n1110 = x82 ^ x2 ;
  assign n1206 = n1205 ^ n1110 ;
  assign n1212 = n1211 ^ n1206 ;
  assign n1213 = ~x0 & n1212 ;
  assign n1292 = n1291 ^ n1213 ;
  assign n1195 = n1193 ^ n1188 ;
  assign n1196 = ~n1190 & n1195 ;
  assign n1197 = n1196 ^ n1193 ;
  assign n1293 = n1292 ^ n1197 ;
  assign n1396 = n1290 ^ n1197 ;
  assign n1397 = n1292 & n1396 ;
  assign n1398 = n1397 ^ n1290 ;
  assign n1390 = n1283 ^ n1216 ;
  assign n1391 = n1289 & n1390 ;
  assign n1392 = n1391 ^ n1283 ;
  assign n1388 = x80 & n231 ;
  assign n1381 = x77 & n391 ;
  assign n1373 = n1266 ^ n1226 ;
  assign n1374 = n1272 & n1373 ;
  assign n1375 = n1374 ^ n1266 ;
  assign n1371 = x74 & n584 ;
  assign n1364 = x71 & n795 ;
  assign n1357 = x68 & n1068 ;
  assign n1244 = x19 ^ x18 ;
  assign n1348 = ~n1143 & n1244 ;
  assign n1349 = x65 & n1348 ;
  assign n1337 = x20 ^ x19 ;
  assign n1343 = n1143 & ~n1337 ;
  assign n1344 = n1343 ^ n1143 ;
  assign n1345 = ~n152 & n1344 ;
  assign n1342 = x66 & n1143 ;
  assign n1346 = n1345 ^ n1342 ;
  assign n1347 = n1346 ^ x20 ;
  assign n1350 = n1349 ^ n1347 ;
  assign n1338 = x20 ^ x18 ;
  assign n1339 = ~n1143 & n1338 ;
  assign n1340 = n1337 & n1339 ;
  assign n1341 = x64 & n1340 ;
  assign n1351 = n1350 ^ n1341 ;
  assign n1335 = ~n1144 & ~n1250 ;
  assign n1336 = x20 & n1335 ;
  assign n1352 = n1351 ^ n1336 ;
  assign n1353 = n1352 ^ x17 ;
  assign n1334 = x67 & n1060 ;
  assign n1354 = n1353 ^ n1334 ;
  assign n1333 = x69 & n1063 ;
  assign n1355 = n1354 ^ n1333 ;
  assign n1332 = ~n376 & n1064 ;
  assign n1356 = n1355 ^ n1332 ;
  assign n1358 = n1357 ^ n1356 ;
  assign n1329 = n1250 ^ n1235 ;
  assign n1330 = n1255 & n1329 ;
  assign n1331 = n1330 ^ n1250 ;
  assign n1359 = n1358 ^ n1331 ;
  assign n1360 = n1359 ^ x14 ;
  assign n1328 = x70 & n884 ;
  assign n1361 = n1360 ^ n1328 ;
  assign n1327 = x72 & n789 ;
  assign n1362 = n1361 ^ n1327 ;
  assign n1326 = n565 & n790 ;
  assign n1363 = n1362 ^ n1326 ;
  assign n1365 = n1364 ^ n1363 ;
  assign n1323 = n1265 ^ n1256 ;
  assign n1324 = ~n1262 & n1323 ;
  assign n1325 = n1324 ^ n1265 ;
  assign n1366 = n1365 ^ n1325 ;
  assign n1367 = n1366 ^ x11 ;
  assign n1322 = x73 & n650 ;
  assign n1368 = n1367 ^ n1322 ;
  assign n1321 = x75 & ~n578 ;
  assign n1369 = n1368 ^ n1321 ;
  assign n1320 = ~n579 & ~n778 ;
  assign n1370 = n1369 ^ n1320 ;
  assign n1372 = n1371 ^ n1370 ;
  assign n1376 = n1375 ^ n1372 ;
  assign n1377 = n1376 ^ x8 ;
  assign n1319 = x76 & n456 ;
  assign n1378 = n1377 ^ n1319 ;
  assign n1318 = x78 & n384 ;
  assign n1379 = n1378 ^ n1318 ;
  assign n1317 = n385 & ~n1036 ;
  assign n1380 = n1379 ^ n1317 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1314 = n1282 ^ n1273 ;
  assign n1315 = ~n1279 & n1314 ;
  assign n1316 = n1315 ^ n1282 ;
  assign n1383 = n1382 ^ n1316 ;
  assign n1384 = n1383 ^ x5 ;
  assign n1313 = x79 & n238 ;
  assign n1385 = n1384 ^ n1313 ;
  assign n1312 = x81 & n234 ;
  assign n1386 = n1385 ^ n1312 ;
  assign n1310 = n1019 ^ x81 ;
  assign n1311 = n235 & n1310 ;
  assign n1387 = n1386 ^ n1311 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1393 = n1392 ^ n1389 ;
  assign n1294 = x83 ^ x82 ;
  assign n1296 = ~n1200 & n1294 ;
  assign n1300 = ~n1296 & n10145 ;
  assign n1298 = x84 ^ x1 ;
  assign n1301 = n1300 ^ n1298 ;
  assign n1394 = n1393 ^ n1301 ;
  assign n1305 = x2 & x82 ;
  assign n1306 = n1305 ^ x83 ;
  assign n1307 = ~n259 & n1306 ;
  assign n1201 = x83 ^ x2 ;
  assign n1302 = n1301 ^ n1201 ;
  assign n1308 = n1307 ^ n1302 ;
  assign n1309 = ~x0 & n1308 ;
  assign n1395 = n1394 ^ n1309 ;
  assign n1399 = n1398 ^ n1395 ;
  assign n1495 = x81 & n231 ;
  assign n1487 = n1376 ^ n1316 ;
  assign n1488 = n1382 & n1487 ;
  assign n1489 = n1488 ^ n1376 ;
  assign n1485 = x78 & n391 ;
  assign n1478 = x75 & n584 ;
  assign n1470 = n1359 ^ n1325 ;
  assign n1471 = n1365 & n1470 ;
  assign n1472 = n1471 ^ n1359 ;
  assign n1468 = x72 & n795 ;
  assign n1460 = n1352 ^ n1331 ;
  assign n1461 = n1358 & n1460 ;
  assign n1462 = n1461 ^ n1352 ;
  assign n1458 = x69 & n1068 ;
  assign n1447 = x65 & n1340 ;
  assign n1446 = x67 & n1343 ;
  assign n1448 = n1447 ^ n1446 ;
  assign n1449 = n1448 ^ x20 ;
  assign n1445 = ~n295 & n1344 ;
  assign n1450 = n1449 ^ n1445 ;
  assign n1444 = x66 & n1348 ;
  assign n1451 = n1450 ^ n1444 ;
  assign n1442 = x21 ^ x20 ;
  assign n1443 = x64 & n1442 ;
  assign n1452 = n1451 ^ n1443 ;
  assign n1441 = n1336 & n1351 ;
  assign n1453 = n1452 ^ n1441 ;
  assign n1454 = n1453 ^ x17 ;
  assign n1440 = x68 & n1060 ;
  assign n1455 = n1454 ^ n1440 ;
  assign n1439 = x70 & n1063 ;
  assign n1456 = n1455 ^ n1439 ;
  assign n1438 = ~n443 & n1064 ;
  assign n1457 = n1456 ^ n1438 ;
  assign n1459 = n1458 ^ n1457 ;
  assign n1463 = n1462 ^ n1459 ;
  assign n1464 = n1463 ^ x14 ;
  assign n1437 = x71 & n884 ;
  assign n1465 = n1464 ^ n1437 ;
  assign n1436 = x73 & n789 ;
  assign n1466 = n1465 ^ n1436 ;
  assign n1435 = n636 & n790 ;
  assign n1467 = n1466 ^ n1435 ;
  assign n1469 = n1468 ^ n1467 ;
  assign n1473 = n1472 ^ n1469 ;
  assign n1474 = n1473 ^ x11 ;
  assign n1434 = x74 & n650 ;
  assign n1475 = n1474 ^ n1434 ;
  assign n1433 = x76 & ~n578 ;
  assign n1476 = n1475 ^ n1433 ;
  assign n1432 = ~n579 & ~n863 ;
  assign n1477 = n1476 ^ n1432 ;
  assign n1479 = n1478 ^ n1477 ;
  assign n1429 = n1375 ^ n1366 ;
  assign n1430 = ~n1372 & n1429 ;
  assign n1431 = n1430 ^ n1375 ;
  assign n1480 = n1479 ^ n1431 ;
  assign n1481 = n1480 ^ x8 ;
  assign n1428 = x77 & n456 ;
  assign n1482 = n1481 ^ n1428 ;
  assign n1427 = x79 & n384 ;
  assign n1483 = n1482 ^ n1427 ;
  assign n1426 = n385 & n1123 ;
  assign n1484 = n1483 ^ n1426 ;
  assign n1486 = n1485 ^ n1484 ;
  assign n1490 = n1489 ^ n1486 ;
  assign n1491 = n1490 ^ x5 ;
  assign n1425 = x80 & n238 ;
  assign n1492 = n1491 ^ n1425 ;
  assign n1424 = x82 & n234 ;
  assign n1493 = n1492 ^ n1424 ;
  assign n1422 = n1109 ^ x82 ;
  assign n1423 = n235 & n1422 ;
  assign n1494 = n1493 ^ n1423 ;
  assign n1496 = n1495 ^ n1494 ;
  assign n1419 = n1392 ^ n1383 ;
  assign n1420 = ~n1389 & n1419 ;
  assign n1421 = n1420 ^ n1392 ;
  assign n1497 = n1496 ^ n1421 ;
  assign n1403 = x84 ^ x83 ;
  assign n1405 = ~n1296 & n1403 ;
  assign n1407 = x85 ^ x1 ;
  assign n1406 = x85 ^ x2 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1409 = ~n1405 & n1408 ;
  assign n1410 = n1409 ^ n1407 ;
  assign n1498 = n1497 ^ n1410 ;
  assign n1414 = x2 & x83 ;
  assign n1415 = n1414 ^ x84 ;
  assign n1416 = ~x1 & n1415 ;
  assign n1297 = x84 ^ x2 ;
  assign n1411 = n1410 ^ n1297 ;
  assign n1417 = n1416 ^ n1411 ;
  assign n1418 = ~x0 & n1417 ;
  assign n1499 = n1498 ^ n1418 ;
  assign n1400 = n1398 ^ n1393 ;
  assign n1401 = ~n1395 & n1400 ;
  assign n1402 = n1401 ^ n1398 ;
  assign n1500 = n1499 ^ n1402 ;
  assign n1609 = n1497 ^ n1402 ;
  assign n1610 = n1499 & n1609 ;
  assign n1611 = n1610 ^ n1497 ;
  assign n1603 = n1490 ^ n1421 ;
  assign n1604 = n1496 & n1603 ;
  assign n1605 = n1604 ^ n1490 ;
  assign n1601 = x82 & n231 ;
  assign n1594 = x79 & n391 ;
  assign n1586 = n1473 ^ n1431 ;
  assign n1587 = n1479 & n1586 ;
  assign n1588 = n1587 ^ n1473 ;
  assign n1584 = x76 & n584 ;
  assign n1577 = x73 & n795 ;
  assign n1570 = x70 & n1068 ;
  assign n1563 = x67 & n1348 ;
  assign n1561 = ~n351 & n1344 ;
  assign n1555 = x20 & x21 ;
  assign n1556 = n1555 ^ x22 ;
  assign n1557 = ~x64 & n1556 ;
  assign n1551 = x22 ^ x20 ;
  assign n1558 = n1557 ^ n1551 ;
  assign n1549 = x65 ^ x21 ;
  assign n1550 = n1442 & ~n1549 ;
  assign n1559 = n1558 ^ n1550 ;
  assign n1546 = x66 & n1340 ;
  assign n1545 = x68 & n1343 ;
  assign n1547 = n1546 ^ n1545 ;
  assign n1548 = n1547 ^ x20 ;
  assign n1560 = n1559 ^ n1548 ;
  assign n1562 = n1561 ^ n1560 ;
  assign n1564 = n1563 ^ n1562 ;
  assign n1542 = ~n1443 & n1451 ;
  assign n1543 = ~n1441 & n1542 ;
  assign n1544 = n1543 ^ n1451 ;
  assign n1565 = n1564 ^ n1544 ;
  assign n1566 = n1565 ^ x17 ;
  assign n1541 = x69 & n1060 ;
  assign n1567 = n1566 ^ n1541 ;
  assign n1540 = x71 & n1063 ;
  assign n1568 = n1567 ^ n1540 ;
  assign n1539 = ~n495 & n1064 ;
  assign n1569 = n1568 ^ n1539 ;
  assign n1571 = n1570 ^ n1569 ;
  assign n1536 = n1462 ^ n1453 ;
  assign n1537 = ~n1459 & n1536 ;
  assign n1538 = n1537 ^ n1462 ;
  assign n1572 = n1571 ^ n1538 ;
  assign n1573 = n1572 ^ x14 ;
  assign n1535 = x72 & n884 ;
  assign n1574 = n1573 ^ n1535 ;
  assign n1534 = x74 & n789 ;
  assign n1575 = n1574 ^ n1534 ;
  assign n1533 = n708 & n790 ;
  assign n1576 = n1575 ^ n1533 ;
  assign n1578 = n1577 ^ n1576 ;
  assign n1530 = n1472 ^ n1463 ;
  assign n1531 = ~n1469 & n1530 ;
  assign n1532 = n1531 ^ n1472 ;
  assign n1579 = n1578 ^ n1532 ;
  assign n1580 = n1579 ^ x11 ;
  assign n1529 = x75 & n650 ;
  assign n1581 = n1580 ^ n1529 ;
  assign n1528 = x77 & ~n578 ;
  assign n1582 = n1581 ^ n1528 ;
  assign n1527 = ~n579 & ~n943 ;
  assign n1583 = n1582 ^ n1527 ;
  assign n1585 = n1584 ^ n1583 ;
  assign n1589 = n1588 ^ n1585 ;
  assign n1590 = n1589 ^ x8 ;
  assign n1526 = x78 & n456 ;
  assign n1591 = n1590 ^ n1526 ;
  assign n1525 = x80 & n384 ;
  assign n1592 = n1591 ^ n1525 ;
  assign n1524 = n385 & n1217 ;
  assign n1593 = n1592 ^ n1524 ;
  assign n1595 = n1594 ^ n1593 ;
  assign n1521 = n1489 ^ n1480 ;
  assign n1522 = ~n1486 & n1521 ;
  assign n1523 = n1522 ^ n1489 ;
  assign n1596 = n1595 ^ n1523 ;
  assign n1597 = n1596 ^ x5 ;
  assign n1520 = x81 & n238 ;
  assign n1598 = n1597 ^ n1520 ;
  assign n1519 = x83 & n234 ;
  assign n1599 = n1598 ^ n1519 ;
  assign n1517 = n1200 ^ x83 ;
  assign n1518 = n235 & n1517 ;
  assign n1600 = n1599 ^ n1518 ;
  assign n1602 = n1601 ^ n1600 ;
  assign n1606 = n1605 ^ n1602 ;
  assign n1501 = x85 ^ x84 ;
  assign n1503 = ~n1405 & n1501 ;
  assign n1505 = x86 ^ x1 ;
  assign n1504 = x86 ^ x2 ;
  assign n1506 = n1505 ^ n1504 ;
  assign n1507 = ~n1503 & n1506 ;
  assign n1508 = n1507 ^ n1505 ;
  assign n1607 = n1606 ^ n1508 ;
  assign n1512 = x2 & x84 ;
  assign n1513 = n1512 ^ x85 ;
  assign n1514 = ~x1 & n1513 ;
  assign n1509 = n1508 ^ n1406 ;
  assign n1515 = n1514 ^ n1509 ;
  assign n1516 = ~x0 & n1515 ;
  assign n1608 = n1607 ^ n1516 ;
  assign n1612 = n1611 ^ n1608 ;
  assign n1726 = x83 & n231 ;
  assign n1718 = n1589 ^ n1523 ;
  assign n1719 = n1595 & n1718 ;
  assign n1720 = n1719 ^ n1589 ;
  assign n1716 = x80 & n391 ;
  assign n1709 = x77 & n584 ;
  assign n1701 = n1572 ^ n1532 ;
  assign n1702 = n1578 & n1701 ;
  assign n1703 = n1702 ^ n1572 ;
  assign n1699 = x74 & n795 ;
  assign n1691 = n1565 ^ n1538 ;
  assign n1692 = n1571 & n1691 ;
  assign n1693 = n1692 ^ n1565 ;
  assign n1689 = x71 & n1068 ;
  assign n1682 = x68 & n1348 ;
  assign n1553 = x22 ^ x21 ;
  assign n1673 = ~n1442 & n1553 ;
  assign n1674 = x65 & n1673 ;
  assign n1662 = x23 ^ x22 ;
  assign n1668 = n1442 & ~n1662 ;
  assign n1669 = n1668 ^ n1442 ;
  assign n1670 = ~n152 & n1669 ;
  assign n1667 = x66 & n1442 ;
  assign n1671 = n1670 ^ n1667 ;
  assign n1672 = n1671 ^ x23 ;
  assign n1675 = n1674 ^ n1672 ;
  assign n1663 = x23 ^ x21 ;
  assign n1664 = ~n1442 & n1663 ;
  assign n1665 = n1662 & n1664 ;
  assign n1666 = x64 & n1665 ;
  assign n1676 = n1675 ^ n1666 ;
  assign n1660 = ~n1443 & ~n1559 ;
  assign n1661 = x23 & n1660 ;
  assign n1677 = n1676 ^ n1661 ;
  assign n1678 = n1677 ^ x20 ;
  assign n1659 = x67 & n1340 ;
  assign n1679 = n1678 ^ n1659 ;
  assign n1658 = x69 & n1343 ;
  assign n1680 = n1679 ^ n1658 ;
  assign n1657 = ~n376 & n1344 ;
  assign n1681 = n1680 ^ n1657 ;
  assign n1683 = n1682 ^ n1681 ;
  assign n1654 = n1559 ^ n1544 ;
  assign n1655 = n1564 & n1654 ;
  assign n1656 = n1655 ^ n1559 ;
  assign n1684 = n1683 ^ n1656 ;
  assign n1685 = n1684 ^ x17 ;
  assign n1653 = x70 & n1060 ;
  assign n1686 = n1685 ^ n1653 ;
  assign n1652 = x72 & n1063 ;
  assign n1687 = n1686 ^ n1652 ;
  assign n1651 = n565 & n1064 ;
  assign n1688 = n1687 ^ n1651 ;
  assign n1690 = n1689 ^ n1688 ;
  assign n1694 = n1693 ^ n1690 ;
  assign n1695 = n1694 ^ x14 ;
  assign n1650 = x73 & n884 ;
  assign n1696 = n1695 ^ n1650 ;
  assign n1649 = x75 & n789 ;
  assign n1697 = n1696 ^ n1649 ;
  assign n1648 = ~n778 & n790 ;
  assign n1698 = n1697 ^ n1648 ;
  assign n1700 = n1699 ^ n1698 ;
  assign n1704 = n1703 ^ n1700 ;
  assign n1705 = n1704 ^ x11 ;
  assign n1647 = x76 & n650 ;
  assign n1706 = n1705 ^ n1647 ;
  assign n1646 = x78 & ~n578 ;
  assign n1707 = n1706 ^ n1646 ;
  assign n1645 = ~n579 & ~n1036 ;
  assign n1708 = n1707 ^ n1645 ;
  assign n1710 = n1709 ^ n1708 ;
  assign n1642 = n1588 ^ n1579 ;
  assign n1643 = ~n1585 & n1642 ;
  assign n1644 = n1643 ^ n1588 ;
  assign n1711 = n1710 ^ n1644 ;
  assign n1712 = n1711 ^ x8 ;
  assign n1641 = x79 & n456 ;
  assign n1713 = n1712 ^ n1641 ;
  assign n1640 = x81 & n384 ;
  assign n1714 = n1713 ^ n1640 ;
  assign n1639 = n385 & n1310 ;
  assign n1715 = n1714 ^ n1639 ;
  assign n1717 = n1716 ^ n1715 ;
  assign n1721 = n1720 ^ n1717 ;
  assign n1722 = n1721 ^ x5 ;
  assign n1638 = x82 & n238 ;
  assign n1723 = n1722 ^ n1638 ;
  assign n1637 = x84 & n234 ;
  assign n1724 = n1723 ^ n1637 ;
  assign n1635 = n1296 ^ x84 ;
  assign n1636 = n235 & n1635 ;
  assign n1725 = n1724 ^ n1636 ;
  assign n1727 = n1726 ^ n1725 ;
  assign n1632 = n1605 ^ n1596 ;
  assign n1633 = ~n1602 & n1632 ;
  assign n1634 = n1633 ^ n1605 ;
  assign n1728 = n1727 ^ n1634 ;
  assign n1616 = x86 ^ x85 ;
  assign n1618 = ~n1503 & n1616 ;
  assign n1620 = x87 ^ x1 ;
  assign n1619 = x87 ^ x2 ;
  assign n1621 = n1620 ^ n1619 ;
  assign n1622 = ~n1618 & n1621 ;
  assign n1623 = n1622 ^ n1620 ;
  assign n1729 = n1728 ^ n1623 ;
  assign n1627 = x2 & x85 ;
  assign n1628 = n1627 ^ x86 ;
  assign n1629 = ~x1 & n1628 ;
  assign n1624 = n1623 ^ n1504 ;
  assign n1630 = n1629 ^ n1624 ;
  assign n1631 = ~x0 & n1630 ;
  assign n1730 = n1729 ^ n1631 ;
  assign n1613 = n1611 ^ n1606 ;
  assign n1614 = ~n1608 & n1613 ;
  assign n1615 = n1614 ^ n1611 ;
  assign n1731 = n1730 ^ n1615 ;
  assign n1842 = n1728 ^ n1615 ;
  assign n1843 = n1730 & n1842 ;
  assign n1844 = n1843 ^ n1728 ;
  assign n1836 = n1721 ^ n1634 ;
  assign n1837 = n1727 & n1836 ;
  assign n1838 = n1837 ^ n1721 ;
  assign n1834 = x84 & n231 ;
  assign n1827 = x81 & n391 ;
  assign n1819 = n1704 ^ n1644 ;
  assign n1820 = n1710 & n1819 ;
  assign n1821 = n1820 ^ n1704 ;
  assign n1817 = x78 & n584 ;
  assign n1810 = x75 & n795 ;
  assign n1803 = x72 & n1068 ;
  assign n1795 = n1677 ^ n1656 ;
  assign n1796 = n1683 & n1795 ;
  assign n1797 = n1796 ^ n1677 ;
  assign n1793 = x69 & n1348 ;
  assign n1782 = x65 & n1665 ;
  assign n1781 = x67 & n1668 ;
  assign n1783 = n1782 ^ n1781 ;
  assign n1784 = n1783 ^ x23 ;
  assign n1780 = ~n295 & n1669 ;
  assign n1785 = n1784 ^ n1780 ;
  assign n1779 = x66 & n1673 ;
  assign n1786 = n1785 ^ n1779 ;
  assign n1777 = x24 ^ x23 ;
  assign n1778 = x64 & n1777 ;
  assign n1787 = n1786 ^ n1778 ;
  assign n1776 = n1661 & n1676 ;
  assign n1788 = n1787 ^ n1776 ;
  assign n1789 = n1788 ^ x20 ;
  assign n1775 = x68 & n1340 ;
  assign n1790 = n1789 ^ n1775 ;
  assign n1774 = x70 & n1343 ;
  assign n1791 = n1790 ^ n1774 ;
  assign n1773 = ~n443 & n1344 ;
  assign n1792 = n1791 ^ n1773 ;
  assign n1794 = n1793 ^ n1792 ;
  assign n1798 = n1797 ^ n1794 ;
  assign n1799 = n1798 ^ x17 ;
  assign n1772 = x71 & n1060 ;
  assign n1800 = n1799 ^ n1772 ;
  assign n1771 = x73 & n1063 ;
  assign n1801 = n1800 ^ n1771 ;
  assign n1770 = n636 & n1064 ;
  assign n1802 = n1801 ^ n1770 ;
  assign n1804 = n1803 ^ n1802 ;
  assign n1767 = n1693 ^ n1684 ;
  assign n1768 = ~n1690 & n1767 ;
  assign n1769 = n1768 ^ n1693 ;
  assign n1805 = n1804 ^ n1769 ;
  assign n1806 = n1805 ^ x14 ;
  assign n1766 = x74 & n884 ;
  assign n1807 = n1806 ^ n1766 ;
  assign n1765 = x76 & n789 ;
  assign n1808 = n1807 ^ n1765 ;
  assign n1764 = n790 & ~n863 ;
  assign n1809 = n1808 ^ n1764 ;
  assign n1811 = n1810 ^ n1809 ;
  assign n1761 = n1703 ^ n1694 ;
  assign n1762 = ~n1700 & n1761 ;
  assign n1763 = n1762 ^ n1703 ;
  assign n1812 = n1811 ^ n1763 ;
  assign n1813 = n1812 ^ x11 ;
  assign n1760 = x77 & n650 ;
  assign n1814 = n1813 ^ n1760 ;
  assign n1759 = x79 & ~n578 ;
  assign n1815 = n1814 ^ n1759 ;
  assign n1758 = ~n579 & n1123 ;
  assign n1816 = n1815 ^ n1758 ;
  assign n1818 = n1817 ^ n1816 ;
  assign n1822 = n1821 ^ n1818 ;
  assign n1823 = n1822 ^ x8 ;
  assign n1757 = x80 & n456 ;
  assign n1824 = n1823 ^ n1757 ;
  assign n1756 = x82 & n384 ;
  assign n1825 = n1824 ^ n1756 ;
  assign n1755 = n385 & n1422 ;
  assign n1826 = n1825 ^ n1755 ;
  assign n1828 = n1827 ^ n1826 ;
  assign n1752 = n1720 ^ n1711 ;
  assign n1753 = ~n1717 & n1752 ;
  assign n1754 = n1753 ^ n1720 ;
  assign n1829 = n1828 ^ n1754 ;
  assign n1830 = n1829 ^ x5 ;
  assign n1751 = x83 & n238 ;
  assign n1831 = n1830 ^ n1751 ;
  assign n1750 = x85 & n234 ;
  assign n1832 = n1831 ^ n1750 ;
  assign n1748 = n1405 ^ x85 ;
  assign n1749 = n235 & n1748 ;
  assign n1833 = n1832 ^ n1749 ;
  assign n1835 = n1834 ^ n1833 ;
  assign n1839 = n1838 ^ n1835 ;
  assign n1732 = x87 ^ x86 ;
  assign n1734 = ~n1618 & n1732 ;
  assign n1736 = x88 ^ x1 ;
  assign n1735 = x88 ^ x2 ;
  assign n1737 = n1736 ^ n1735 ;
  assign n1738 = ~n1734 & n1737 ;
  assign n1739 = n1738 ^ n1736 ;
  assign n1840 = n1839 ^ n1739 ;
  assign n1743 = x2 & x86 ;
  assign n1744 = n1743 ^ x87 ;
  assign n1745 = ~x1 & n1744 ;
  assign n1740 = n1739 ^ n1619 ;
  assign n1746 = n1745 ^ n1740 ;
  assign n1747 = ~x0 & n1746 ;
  assign n1841 = n1840 ^ n1747 ;
  assign n1845 = n1844 ^ n1841 ;
  assign n1965 = x85 & n231 ;
  assign n1957 = n1822 ^ n1754 ;
  assign n1958 = n1828 & n1957 ;
  assign n1959 = n1958 ^ n1822 ;
  assign n1955 = x82 & n391 ;
  assign n1948 = x79 & n584 ;
  assign n1940 = n1805 ^ n1763 ;
  assign n1941 = n1811 & n1940 ;
  assign n1942 = n1941 ^ n1805 ;
  assign n1938 = x76 & n795 ;
  assign n1930 = n1798 ^ n1769 ;
  assign n1931 = n1804 & n1930 ;
  assign n1932 = n1931 ^ n1798 ;
  assign n1928 = x73 & n1068 ;
  assign n1921 = x70 & n1348 ;
  assign n1910 = x66 & n1665 ;
  assign n1909 = x68 & n1668 ;
  assign n1911 = n1910 ^ n1909 ;
  assign n1912 = n1911 ^ x23 ;
  assign n1908 = ~n351 & n1669 ;
  assign n1913 = n1912 ^ n1908 ;
  assign n1907 = x67 & n1673 ;
  assign n1914 = n1913 ^ n1907 ;
  assign n1904 = x65 ^ x24 ;
  assign n1905 = n1777 & ~n1904 ;
  assign n1900 = x23 & x24 ;
  assign n1901 = n1900 ^ x25 ;
  assign n1902 = ~x64 & n1901 ;
  assign n1896 = x25 ^ x23 ;
  assign n1903 = n1902 ^ n1896 ;
  assign n1906 = n1905 ^ n1903 ;
  assign n1915 = n1914 ^ n1906 ;
  assign n1893 = ~n1778 & n1786 ;
  assign n1894 = ~n1776 & n1893 ;
  assign n1895 = n1894 ^ n1786 ;
  assign n1916 = n1915 ^ n1895 ;
  assign n1917 = n1916 ^ x20 ;
  assign n1892 = x69 & n1340 ;
  assign n1918 = n1917 ^ n1892 ;
  assign n1891 = x71 & n1343 ;
  assign n1919 = n1918 ^ n1891 ;
  assign n1890 = ~n495 & n1344 ;
  assign n1920 = n1919 ^ n1890 ;
  assign n1922 = n1921 ^ n1920 ;
  assign n1887 = n1797 ^ n1788 ;
  assign n1888 = ~n1794 & n1887 ;
  assign n1889 = n1888 ^ n1797 ;
  assign n1923 = n1922 ^ n1889 ;
  assign n1924 = n1923 ^ x17 ;
  assign n1886 = x72 & n1060 ;
  assign n1925 = n1924 ^ n1886 ;
  assign n1885 = x74 & n1063 ;
  assign n1926 = n1925 ^ n1885 ;
  assign n1884 = n708 & n1064 ;
  assign n1927 = n1926 ^ n1884 ;
  assign n1929 = n1928 ^ n1927 ;
  assign n1933 = n1932 ^ n1929 ;
  assign n1934 = n1933 ^ x14 ;
  assign n1883 = x75 & n884 ;
  assign n1935 = n1934 ^ n1883 ;
  assign n1882 = x77 & n789 ;
  assign n1936 = n1935 ^ n1882 ;
  assign n1881 = n790 & ~n943 ;
  assign n1937 = n1936 ^ n1881 ;
  assign n1939 = n1938 ^ n1937 ;
  assign n1943 = n1942 ^ n1939 ;
  assign n1944 = n1943 ^ x11 ;
  assign n1880 = x78 & n650 ;
  assign n1945 = n1944 ^ n1880 ;
  assign n1879 = x80 & ~n578 ;
  assign n1946 = n1945 ^ n1879 ;
  assign n1878 = ~n579 & n1217 ;
  assign n1947 = n1946 ^ n1878 ;
  assign n1949 = n1948 ^ n1947 ;
  assign n1875 = n1821 ^ n1812 ;
  assign n1876 = ~n1818 & n1875 ;
  assign n1877 = n1876 ^ n1821 ;
  assign n1950 = n1949 ^ n1877 ;
  assign n1951 = n1950 ^ x8 ;
  assign n1874 = x81 & n456 ;
  assign n1952 = n1951 ^ n1874 ;
  assign n1873 = x83 & n384 ;
  assign n1953 = n1952 ^ n1873 ;
  assign n1872 = n385 & n1517 ;
  assign n1954 = n1953 ^ n1872 ;
  assign n1956 = n1955 ^ n1954 ;
  assign n1960 = n1959 ^ n1956 ;
  assign n1961 = n1960 ^ x5 ;
  assign n1871 = x84 & n238 ;
  assign n1962 = n1961 ^ n1871 ;
  assign n1870 = x86 & n234 ;
  assign n1963 = n1962 ^ n1870 ;
  assign n1868 = n1503 ^ x86 ;
  assign n1869 = n235 & n1868 ;
  assign n1964 = n1963 ^ n1869 ;
  assign n1966 = n1965 ^ n1964 ;
  assign n1865 = n1838 ^ n1829 ;
  assign n1866 = ~n1835 & n1865 ;
  assign n1867 = n1866 ^ n1838 ;
  assign n1967 = n1966 ^ n1867 ;
  assign n1849 = x88 ^ x87 ;
  assign n1851 = ~n1734 & n1849 ;
  assign n1853 = x89 ^ x1 ;
  assign n1852 = x89 ^ x2 ;
  assign n1854 = n1853 ^ n1852 ;
  assign n1855 = ~n1851 & n1854 ;
  assign n1856 = n1855 ^ n1853 ;
  assign n1968 = n1967 ^ n1856 ;
  assign n1860 = x2 & x87 ;
  assign n1861 = n1860 ^ x88 ;
  assign n1862 = ~x1 & n1861 ;
  assign n1857 = n1856 ^ n1735 ;
  assign n1863 = n1862 ^ n1857 ;
  assign n1864 = ~x0 & n1863 ;
  assign n1969 = n1968 ^ n1864 ;
  assign n1846 = n1844 ^ n1839 ;
  assign n1847 = ~n1841 & n1846 ;
  assign n1848 = n1847 ^ n1844 ;
  assign n1970 = n1969 ^ n1848 ;
  assign n2105 = n1967 ^ n1848 ;
  assign n2106 = n1969 & n2105 ;
  assign n2107 = n2106 ^ n1967 ;
  assign n2099 = n1960 ^ n1867 ;
  assign n2100 = n1966 & n2099 ;
  assign n2101 = n2100 ^ n1960 ;
  assign n2097 = x86 & n231 ;
  assign n2090 = x83 & n391 ;
  assign n2082 = n1943 ^ n1877 ;
  assign n2083 = n1949 & n2082 ;
  assign n2084 = n2083 ^ n1943 ;
  assign n2080 = x80 & n584 ;
  assign n2073 = x77 & n795 ;
  assign n2064 = n1916 ^ n1889 ;
  assign n2065 = n1922 & n2064 ;
  assign n2066 = n2065 ^ n1916 ;
  assign n2062 = x71 & n1348 ;
  assign n2051 = x67 & n1665 ;
  assign n2050 = x69 & n1668 ;
  assign n2052 = n2051 ^ n2050 ;
  assign n2053 = n2052 ^ x23 ;
  assign n2049 = ~n376 & n1669 ;
  assign n2054 = n2053 ^ n2049 ;
  assign n2048 = x68 & n1673 ;
  assign n2055 = n2054 ^ n2048 ;
  assign n2044 = ~n1778 & ~n1906 ;
  assign n2045 = x26 & n2044 ;
  assign n2046 = n2045 ^ x26 ;
  assign n2041 = x66 & n1777 ;
  assign n2027 = x26 ^ x25 ;
  assign n2028 = n1777 & ~n2027 ;
  assign n2029 = n2028 ^ n1777 ;
  assign n2037 = x65 & n2029 ;
  assign n2030 = x26 ^ x24 ;
  assign n2031 = ~n1777 & n2030 ;
  assign n2032 = n2027 & n2031 ;
  assign n2038 = n2037 ^ n2032 ;
  assign n2039 = ~x64 & n2038 ;
  assign n2040 = n2039 ^ n2032 ;
  assign n2042 = n2041 ^ n2040 ;
  assign n1898 = x25 ^ x24 ;
  assign n2025 = ~n1777 & n1898 ;
  assign n2026 = x65 & n2025 ;
  assign n2043 = n2042 ^ n2026 ;
  assign n2047 = n2046 ^ n2043 ;
  assign n2056 = n2055 ^ n2047 ;
  assign n2022 = n1906 ^ n1895 ;
  assign n2023 = n1915 & ~n2022 ;
  assign n2024 = n2023 ^ n1914 ;
  assign n2057 = n2056 ^ n2024 ;
  assign n2058 = n2057 ^ x20 ;
  assign n2021 = x70 & n1340 ;
  assign n2059 = n2058 ^ n2021 ;
  assign n2020 = x72 & n1343 ;
  assign n2060 = n2059 ^ n2020 ;
  assign n2019 = n565 & n1344 ;
  assign n2061 = n2060 ^ n2019 ;
  assign n2063 = n2062 ^ n2061 ;
  assign n2067 = n2066 ^ n2063 ;
  assign n2009 = x73 & n1060 ;
  assign n2008 = x75 & n1063 ;
  assign n2010 = n2009 ^ n2008 ;
  assign n2011 = n2010 ^ x17 ;
  assign n2007 = ~n778 & n1064 ;
  assign n2012 = n2011 ^ n2007 ;
  assign n2006 = x74 & n1068 ;
  assign n2013 = n2012 ^ n2006 ;
  assign n2014 = n2013 ^ n1932 ;
  assign n2015 = n2014 ^ n1923 ;
  assign n2016 = n2015 ^ n2013 ;
  assign n2017 = ~n1929 & n2016 ;
  assign n2018 = n2017 ^ n2014 ;
  assign n2068 = n2067 ^ n2018 ;
  assign n2069 = n2068 ^ x14 ;
  assign n2005 = x76 & n884 ;
  assign n2070 = n2069 ^ n2005 ;
  assign n2004 = x78 & n789 ;
  assign n2071 = n2070 ^ n2004 ;
  assign n2003 = n790 & ~n1036 ;
  assign n2072 = n2071 ^ n2003 ;
  assign n2074 = n2073 ^ n2072 ;
  assign n2000 = n1942 ^ n1933 ;
  assign n2001 = ~n1939 & n2000 ;
  assign n2002 = n2001 ^ n1942 ;
  assign n2075 = n2074 ^ n2002 ;
  assign n2076 = n2075 ^ x11 ;
  assign n1999 = x79 & n650 ;
  assign n2077 = n2076 ^ n1999 ;
  assign n1998 = x81 & ~n578 ;
  assign n2078 = n2077 ^ n1998 ;
  assign n1997 = ~n579 & n1310 ;
  assign n2079 = n2078 ^ n1997 ;
  assign n2081 = n2080 ^ n2079 ;
  assign n2085 = n2084 ^ n2081 ;
  assign n2086 = n2085 ^ x8 ;
  assign n1996 = x82 & n456 ;
  assign n2087 = n2086 ^ n1996 ;
  assign n1995 = x84 & n384 ;
  assign n2088 = n2087 ^ n1995 ;
  assign n1994 = n385 & n1635 ;
  assign n2089 = n2088 ^ n1994 ;
  assign n2091 = n2090 ^ n2089 ;
  assign n1991 = n1959 ^ n1950 ;
  assign n1992 = ~n1956 & n1991 ;
  assign n1993 = n1992 ^ n1959 ;
  assign n2092 = n2091 ^ n1993 ;
  assign n2093 = n2092 ^ x5 ;
  assign n1990 = x85 & n238 ;
  assign n2094 = n2093 ^ n1990 ;
  assign n1989 = x87 & n234 ;
  assign n2095 = n2094 ^ n1989 ;
  assign n1987 = n1618 ^ x87 ;
  assign n1988 = n235 & n1987 ;
  assign n2096 = n2095 ^ n1988 ;
  assign n2098 = n2097 ^ n2096 ;
  assign n2102 = n2101 ^ n2098 ;
  assign n1971 = x89 ^ x88 ;
  assign n1973 = ~n1851 & n1971 ;
  assign n1975 = x90 ^ x1 ;
  assign n1974 = x90 ^ x2 ;
  assign n1976 = n1975 ^ n1974 ;
  assign n1977 = ~n1973 & n1976 ;
  assign n1978 = n1977 ^ n1975 ;
  assign n2103 = n2102 ^ n1978 ;
  assign n1982 = x2 & x88 ;
  assign n1983 = n1982 ^ x89 ;
  assign n1984 = ~x1 & n1983 ;
  assign n1979 = n1978 ^ n1852 ;
  assign n1985 = n1984 ^ n1979 ;
  assign n1986 = ~x0 & n1985 ;
  assign n2104 = n2103 ^ n1986 ;
  assign n2108 = n2107 ^ n2104 ;
  assign n2233 = x87 & n231 ;
  assign n2225 = n2085 ^ n1993 ;
  assign n2226 = n2091 & n2225 ;
  assign n2227 = n2226 ^ n2085 ;
  assign n2223 = x84 & n391 ;
  assign n2216 = x81 & n584 ;
  assign n2208 = n2068 ^ n2002 ;
  assign n2209 = n2074 & n2208 ;
  assign n2210 = n2209 ^ n2068 ;
  assign n2206 = x78 & n795 ;
  assign n2199 = x75 & n1068 ;
  assign n2192 = x72 & n1348 ;
  assign n2184 = n2055 ^ n2024 ;
  assign n2185 = n2056 & n2184 ;
  assign n2186 = n2185 ^ n2055 ;
  assign n2178 = x68 & n1665 ;
  assign n2177 = x70 & n1668 ;
  assign n2179 = n2178 ^ n2177 ;
  assign n2180 = n2179 ^ x23 ;
  assign n2176 = ~n443 & n1669 ;
  assign n2181 = n2180 ^ n2176 ;
  assign n2175 = x69 & n1673 ;
  assign n2182 = n2181 ^ n2175 ;
  assign n2172 = ~n2043 & n2045 ;
  assign n2170 = x27 ^ x26 ;
  assign n2171 = x64 & n2170 ;
  assign n2173 = n2172 ^ n2171 ;
  assign n2166 = x65 & n2032 ;
  assign n2165 = x66 & n2025 ;
  assign n2167 = n2166 ^ n2165 ;
  assign n2168 = n2167 ^ x26 ;
  assign n2162 = ~n155 & ~n2027 ;
  assign n2163 = n2162 ^ n295 ;
  assign n2164 = n1777 & ~n2163 ;
  assign n2169 = n2168 ^ n2164 ;
  assign n2174 = n2173 ^ n2169 ;
  assign n2183 = n2182 ^ n2174 ;
  assign n2187 = n2186 ^ n2183 ;
  assign n2188 = n2187 ^ x20 ;
  assign n2158 = x71 & n1340 ;
  assign n2189 = n2188 ^ n2158 ;
  assign n2157 = x73 & n1343 ;
  assign n2190 = n2189 ^ n2157 ;
  assign n2156 = n636 & n1344 ;
  assign n2191 = n2190 ^ n2156 ;
  assign n2193 = n2192 ^ n2191 ;
  assign n2153 = n2066 ^ n2057 ;
  assign n2154 = ~n2063 & n2153 ;
  assign n2155 = n2154 ^ n2066 ;
  assign n2194 = n2193 ^ n2155 ;
  assign n2195 = n2194 ^ x17 ;
  assign n2152 = x74 & n1060 ;
  assign n2196 = n2195 ^ n2152 ;
  assign n2151 = x76 & n1063 ;
  assign n2197 = n2196 ^ n2151 ;
  assign n2150 = ~n863 & n1064 ;
  assign n2198 = n2197 ^ n2150 ;
  assign n2200 = n2199 ^ n2198 ;
  assign n2147 = n2067 ^ n2013 ;
  assign n2148 = n2018 & n2147 ;
  assign n2149 = n2148 ^ n2013 ;
  assign n2201 = n2200 ^ n2149 ;
  assign n2202 = n2201 ^ x14 ;
  assign n2146 = x77 & n884 ;
  assign n2203 = n2202 ^ n2146 ;
  assign n2145 = x79 & n789 ;
  assign n2204 = n2203 ^ n2145 ;
  assign n2144 = n790 & n1123 ;
  assign n2205 = n2204 ^ n2144 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2211 = n2210 ^ n2207 ;
  assign n2212 = n2211 ^ x11 ;
  assign n2143 = x80 & n650 ;
  assign n2213 = n2212 ^ n2143 ;
  assign n2142 = x82 & ~n578 ;
  assign n2214 = n2213 ^ n2142 ;
  assign n2141 = ~n579 & n1422 ;
  assign n2215 = n2214 ^ n2141 ;
  assign n2217 = n2216 ^ n2215 ;
  assign n2138 = n2084 ^ n2075 ;
  assign n2139 = ~n2081 & n2138 ;
  assign n2140 = n2139 ^ n2084 ;
  assign n2218 = n2217 ^ n2140 ;
  assign n2219 = n2218 ^ x8 ;
  assign n2137 = x83 & n456 ;
  assign n2220 = n2219 ^ n2137 ;
  assign n2136 = x85 & n384 ;
  assign n2221 = n2220 ^ n2136 ;
  assign n2135 = n385 & n1748 ;
  assign n2222 = n2221 ^ n2135 ;
  assign n2224 = n2223 ^ n2222 ;
  assign n2228 = n2227 ^ n2224 ;
  assign n2229 = n2228 ^ x5 ;
  assign n2134 = x86 & n238 ;
  assign n2230 = n2229 ^ n2134 ;
  assign n2133 = x88 & n234 ;
  assign n2231 = n2230 ^ n2133 ;
  assign n2131 = n1734 ^ x88 ;
  assign n2132 = n235 & n2131 ;
  assign n2232 = n2231 ^ n2132 ;
  assign n2234 = n2233 ^ n2232 ;
  assign n2128 = n2101 ^ n2092 ;
  assign n2129 = ~n2098 & n2128 ;
  assign n2130 = n2129 ^ n2101 ;
  assign n2235 = n2234 ^ n2130 ;
  assign n2112 = x90 ^ x89 ;
  assign n2114 = ~n1973 & n2112 ;
  assign n2116 = x91 ^ x1 ;
  assign n2115 = x91 ^ x2 ;
  assign n2117 = n2116 ^ n2115 ;
  assign n2118 = ~n2114 & n2117 ;
  assign n2119 = n2118 ^ n2116 ;
  assign n2236 = n2235 ^ n2119 ;
  assign n2123 = x2 & x89 ;
  assign n2124 = n2123 ^ x90 ;
  assign n2125 = ~x1 & n2124 ;
  assign n2120 = n2119 ^ n1974 ;
  assign n2126 = n2125 ^ n2120 ;
  assign n2127 = ~x0 & n2126 ;
  assign n2237 = n2236 ^ n2127 ;
  assign n2109 = n2107 ^ n2102 ;
  assign n2110 = ~n2104 & n2109 ;
  assign n2111 = n2110 ^ n2107 ;
  assign n2238 = n2237 ^ n2111 ;
  assign n2372 = n2235 ^ n2111 ;
  assign n2373 = n2237 & n2372 ;
  assign n2374 = n2373 ^ n2235 ;
  assign n2366 = n2228 ^ n2130 ;
  assign n2367 = n2234 & n2366 ;
  assign n2368 = n2367 ^ n2228 ;
  assign n2364 = x88 & n231 ;
  assign n2357 = x85 & n391 ;
  assign n2349 = n2211 ^ n2140 ;
  assign n2350 = n2217 & n2349 ;
  assign n2351 = n2350 ^ n2211 ;
  assign n2347 = x82 & n584 ;
  assign n2340 = x79 & n795 ;
  assign n2333 = x76 & n1068 ;
  assign n2325 = n2187 ^ n2155 ;
  assign n2326 = n2193 & n2325 ;
  assign n2327 = n2326 ^ n2187 ;
  assign n2323 = x73 & n1348 ;
  assign n2312 = x69 & n1665 ;
  assign n2311 = x71 & n1668 ;
  assign n2313 = n2312 ^ n2311 ;
  assign n2314 = n2313 ^ x23 ;
  assign n2310 = ~n495 & n1669 ;
  assign n2315 = n2314 ^ n2310 ;
  assign n2309 = x70 & n1673 ;
  assign n2316 = n2315 ^ n2309 ;
  assign n2305 = ~n2171 & ~n2172 ;
  assign n2306 = n2169 & n2305 ;
  assign n2307 = n2306 ^ n2169 ;
  assign n2299 = x66 & n2032 ;
  assign n2298 = x68 & n2028 ;
  assign n2300 = n2299 ^ n2298 ;
  assign n2301 = n2300 ^ x26 ;
  assign n2297 = ~n351 & n2029 ;
  assign n2302 = n2301 ^ n2297 ;
  assign n2296 = x67 & n2025 ;
  assign n2303 = n2302 ^ n2296 ;
  assign n2292 = x26 & x27 ;
  assign n2293 = n2292 ^ x28 ;
  assign n2294 = ~x64 & n2293 ;
  assign n2286 = x65 ^ x27 ;
  assign n2289 = x65 ^ x26 ;
  assign n2290 = ~n2286 & n2289 ;
  assign n2287 = x28 ^ x26 ;
  assign n2291 = n2290 ^ n2287 ;
  assign n2295 = n2294 ^ n2291 ;
  assign n2304 = n2303 ^ n2295 ;
  assign n2308 = n2307 ^ n2304 ;
  assign n2317 = n2316 ^ n2308 ;
  assign n2283 = n2186 ^ n2182 ;
  assign n2284 = ~n2183 & n2283 ;
  assign n2285 = n2284 ^ n2186 ;
  assign n2318 = n2317 ^ n2285 ;
  assign n2319 = n2318 ^ x20 ;
  assign n2282 = x72 & n1340 ;
  assign n2320 = n2319 ^ n2282 ;
  assign n2281 = x74 & n1343 ;
  assign n2321 = n2320 ^ n2281 ;
  assign n2280 = n708 & n1344 ;
  assign n2322 = n2321 ^ n2280 ;
  assign n2324 = n2323 ^ n2322 ;
  assign n2328 = n2327 ^ n2324 ;
  assign n2329 = n2328 ^ x17 ;
  assign n2279 = x75 & n1060 ;
  assign n2330 = n2329 ^ n2279 ;
  assign n2278 = x77 & n1063 ;
  assign n2331 = n2330 ^ n2278 ;
  assign n2277 = ~n943 & n1064 ;
  assign n2332 = n2331 ^ n2277 ;
  assign n2334 = n2333 ^ n2332 ;
  assign n2274 = n2194 ^ n2149 ;
  assign n2275 = n2200 & n2274 ;
  assign n2276 = n2275 ^ n2194 ;
  assign n2335 = n2334 ^ n2276 ;
  assign n2336 = n2335 ^ x14 ;
  assign n2273 = x78 & n884 ;
  assign n2337 = n2336 ^ n2273 ;
  assign n2272 = x80 & n789 ;
  assign n2338 = n2337 ^ n2272 ;
  assign n2271 = n790 & n1217 ;
  assign n2339 = n2338 ^ n2271 ;
  assign n2341 = n2340 ^ n2339 ;
  assign n2268 = n2210 ^ n2201 ;
  assign n2269 = ~n2207 & n2268 ;
  assign n2270 = n2269 ^ n2210 ;
  assign n2342 = n2341 ^ n2270 ;
  assign n2343 = n2342 ^ x11 ;
  assign n2267 = x81 & n650 ;
  assign n2344 = n2343 ^ n2267 ;
  assign n2266 = x83 & ~n578 ;
  assign n2345 = n2344 ^ n2266 ;
  assign n2265 = ~n579 & n1517 ;
  assign n2346 = n2345 ^ n2265 ;
  assign n2348 = n2347 ^ n2346 ;
  assign n2352 = n2351 ^ n2348 ;
  assign n2353 = n2352 ^ x8 ;
  assign n2264 = x84 & n456 ;
  assign n2354 = n2353 ^ n2264 ;
  assign n2263 = x86 & n384 ;
  assign n2355 = n2354 ^ n2263 ;
  assign n2262 = n385 & n1868 ;
  assign n2356 = n2355 ^ n2262 ;
  assign n2358 = n2357 ^ n2356 ;
  assign n2259 = n2227 ^ n2218 ;
  assign n2260 = ~n2224 & n2259 ;
  assign n2261 = n2260 ^ n2227 ;
  assign n2359 = n2358 ^ n2261 ;
  assign n2360 = n2359 ^ x5 ;
  assign n2258 = x87 & n238 ;
  assign n2361 = n2360 ^ n2258 ;
  assign n2257 = x89 & n234 ;
  assign n2362 = n2361 ^ n2257 ;
  assign n2255 = n1851 ^ x89 ;
  assign n2256 = n235 & n2255 ;
  assign n2363 = n2362 ^ n2256 ;
  assign n2365 = n2364 ^ n2363 ;
  assign n2369 = n2368 ^ n2365 ;
  assign n2239 = x91 ^ x90 ;
  assign n2241 = ~n2114 & n2239 ;
  assign n2243 = x92 ^ x1 ;
  assign n2242 = x92 ^ x2 ;
  assign n2244 = n2243 ^ n2242 ;
  assign n2245 = ~n2241 & n2244 ;
  assign n2246 = n2245 ^ n2243 ;
  assign n2370 = n2369 ^ n2246 ;
  assign n2250 = x2 & x90 ;
  assign n2251 = n2250 ^ x91 ;
  assign n2252 = ~n259 & n2251 ;
  assign n2247 = n2246 ^ n2115 ;
  assign n2253 = n2252 ^ n2247 ;
  assign n2254 = ~x0 & n2253 ;
  assign n2371 = n2370 ^ n2254 ;
  assign n2375 = n2374 ^ n2371 ;
  assign n2523 = x89 & n231 ;
  assign n2515 = n2352 ^ n2261 ;
  assign n2516 = n2358 & n2515 ;
  assign n2517 = n2516 ^ n2352 ;
  assign n2513 = x86 & n391 ;
  assign n2506 = x83 & n584 ;
  assign n2498 = n2335 ^ n2270 ;
  assign n2499 = n2341 & n2498 ;
  assign n2500 = n2499 ^ n2335 ;
  assign n2496 = x80 & n795 ;
  assign n2488 = n2328 ^ n2276 ;
  assign n2489 = n2334 & n2488 ;
  assign n2490 = n2489 ^ n2328 ;
  assign n2486 = x77 & n1068 ;
  assign n2479 = x74 & n1348 ;
  assign n2471 = n2316 ^ n2285 ;
  assign n2472 = n2317 & n2471 ;
  assign n2473 = n2472 ^ n2316 ;
  assign n2465 = x70 & n1665 ;
  assign n2464 = x72 & n1668 ;
  assign n2466 = n2465 ^ n2464 ;
  assign n2467 = n2466 ^ x23 ;
  assign n2463 = n565 & n1669 ;
  assign n2468 = n2467 ^ n2463 ;
  assign n2462 = x71 & n1673 ;
  assign n2469 = n2468 ^ n2462 ;
  assign n2459 = x68 & n2025 ;
  assign n2456 = x69 & n2028 ;
  assign n2454 = x67 & n2032 ;
  assign n2434 = x28 ^ x27 ;
  assign n2435 = ~n2170 & n2434 ;
  assign n2436 = x65 & n2435 ;
  assign n2427 = x29 ^ x28 ;
  assign n2428 = n2170 & ~n2427 ;
  assign n2429 = n2428 ^ n2170 ;
  assign n2432 = ~n152 & n2429 ;
  assign n2431 = x66 & n2170 ;
  assign n2433 = n2432 ^ n2431 ;
  assign n2437 = n2436 ^ n2433 ;
  assign n2439 = ~n2171 & ~n2295 ;
  assign n2442 = x28 & x64 ;
  assign n2448 = n2442 ^ x64 ;
  assign n2449 = x29 & ~n2448 ;
  assign n2450 = n2439 & n2449 ;
  assign n2451 = ~n2437 & n2450 ;
  assign n2438 = n2437 ^ x29 ;
  assign n2443 = n2292 & n2442 ;
  assign n2444 = n2443 ^ n2439 ;
  assign n2445 = ~n2437 & n2444 ;
  assign n2446 = n2445 ^ n2439 ;
  assign n2447 = ~n2438 & ~n2446 ;
  assign n2452 = n2451 ^ n2447 ;
  assign n2453 = n2452 ^ x26 ;
  assign n2455 = n2454 ^ n2453 ;
  assign n2457 = n2456 ^ n2455 ;
  assign n2426 = ~n376 & n2029 ;
  assign n2458 = n2457 ^ n2426 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2423 = n2307 ^ n2303 ;
  assign n2424 = ~n2304 & n2423 ;
  assign n2425 = n2424 ^ n2307 ;
  assign n2461 = n2460 ^ n2425 ;
  assign n2470 = n2469 ^ n2461 ;
  assign n2474 = n2473 ^ n2470 ;
  assign n2475 = n2474 ^ x20 ;
  assign n2422 = x73 & n1340 ;
  assign n2476 = n2475 ^ n2422 ;
  assign n2421 = x75 & n1343 ;
  assign n2477 = n2476 ^ n2421 ;
  assign n2420 = ~n778 & n1344 ;
  assign n2478 = n2477 ^ n2420 ;
  assign n2480 = n2479 ^ n2478 ;
  assign n2417 = n2327 ^ n2318 ;
  assign n2418 = ~n2324 & n2417 ;
  assign n2419 = n2418 ^ n2327 ;
  assign n2481 = n2480 ^ n2419 ;
  assign n2482 = n2481 ^ x17 ;
  assign n2416 = x76 & n1060 ;
  assign n2483 = n2482 ^ n2416 ;
  assign n2415 = x78 & n1063 ;
  assign n2484 = n2483 ^ n2415 ;
  assign n2414 = ~n1036 & n1064 ;
  assign n2485 = n2484 ^ n2414 ;
  assign n2487 = n2486 ^ n2485 ;
  assign n2491 = n2490 ^ n2487 ;
  assign n2492 = n2491 ^ x14 ;
  assign n2413 = x79 & n884 ;
  assign n2493 = n2492 ^ n2413 ;
  assign n2412 = x81 & n789 ;
  assign n2494 = n2493 ^ n2412 ;
  assign n2411 = n790 & n1310 ;
  assign n2495 = n2494 ^ n2411 ;
  assign n2497 = n2496 ^ n2495 ;
  assign n2501 = n2500 ^ n2497 ;
  assign n2502 = n2501 ^ x11 ;
  assign n2410 = x82 & n650 ;
  assign n2503 = n2502 ^ n2410 ;
  assign n2409 = x84 & ~n578 ;
  assign n2504 = n2503 ^ n2409 ;
  assign n2408 = ~n579 & n1635 ;
  assign n2505 = n2504 ^ n2408 ;
  assign n2507 = n2506 ^ n2505 ;
  assign n2405 = n2351 ^ n2342 ;
  assign n2406 = ~n2348 & n2405 ;
  assign n2407 = n2406 ^ n2351 ;
  assign n2508 = n2507 ^ n2407 ;
  assign n2509 = n2508 ^ x8 ;
  assign n2404 = x85 & n456 ;
  assign n2510 = n2509 ^ n2404 ;
  assign n2403 = x87 & n384 ;
  assign n2511 = n2510 ^ n2403 ;
  assign n2402 = n385 & n1987 ;
  assign n2512 = n2511 ^ n2402 ;
  assign n2514 = n2513 ^ n2512 ;
  assign n2518 = n2517 ^ n2514 ;
  assign n2519 = n2518 ^ x5 ;
  assign n2401 = x88 & n238 ;
  assign n2520 = n2519 ^ n2401 ;
  assign n2400 = x90 & n234 ;
  assign n2521 = n2520 ^ n2400 ;
  assign n2398 = n1973 ^ x90 ;
  assign n2399 = n235 & n2398 ;
  assign n2522 = n2521 ^ n2399 ;
  assign n2524 = n2523 ^ n2522 ;
  assign n2395 = n2368 ^ n2359 ;
  assign n2396 = ~n2365 & n2395 ;
  assign n2397 = n2396 ^ n2368 ;
  assign n2525 = n2524 ^ n2397 ;
  assign n2379 = x92 ^ x91 ;
  assign n2381 = ~n2241 & n2379 ;
  assign n2383 = x93 ^ x1 ;
  assign n2382 = x93 ^ x2 ;
  assign n2384 = n2383 ^ n2382 ;
  assign n2385 = ~n2381 & n2384 ;
  assign n2386 = n2385 ^ n2383 ;
  assign n2526 = n2525 ^ n2386 ;
  assign n2390 = x2 & x91 ;
  assign n2391 = n2390 ^ x92 ;
  assign n2392 = ~n259 & n2391 ;
  assign n2387 = n2386 ^ n2242 ;
  assign n2393 = n2392 ^ n2387 ;
  assign n2394 = ~x0 & n2393 ;
  assign n2527 = n2526 ^ n2394 ;
  assign n2376 = n2374 ^ n2369 ;
  assign n2377 = ~n2371 & n2376 ;
  assign n2378 = n2377 ^ n2374 ;
  assign n2528 = n2527 ^ n2378 ;
  assign n2670 = n2525 ^ n2378 ;
  assign n2671 = ~n2527 & ~n2670 ;
  assign n2672 = n2671 ^ n2525 ;
  assign n2664 = n2518 ^ n2397 ;
  assign n2665 = ~n2524 & ~n2664 ;
  assign n2666 = n2665 ^ n2518 ;
  assign n2662 = x90 & n231 ;
  assign n2655 = x87 & n391 ;
  assign n2647 = n2501 ^ n2407 ;
  assign n2648 = ~n2507 & ~n2647 ;
  assign n2649 = n2648 ^ n2501 ;
  assign n2645 = x84 & n584 ;
  assign n2638 = x81 & n795 ;
  assign n2631 = x78 & n1068 ;
  assign n2623 = n2474 ^ n2419 ;
  assign n2624 = ~n2480 & ~n2623 ;
  assign n2625 = n2624 ^ n2474 ;
  assign n2621 = x75 & n1348 ;
  assign n2614 = x72 & n1673 ;
  assign n2603 = x68 & n2032 ;
  assign n2602 = x70 & n2028 ;
  assign n2604 = n2603 ^ n2602 ;
  assign n2605 = n2604 ^ x26 ;
  assign n2601 = ~n443 & n2029 ;
  assign n2606 = n2605 ^ n2601 ;
  assign n2600 = x69 & n2025 ;
  assign n2607 = n2606 ^ n2600 ;
  assign n2591 = x29 ^ x27 ;
  assign n2592 = ~n2170 & n2591 ;
  assign n2593 = n2427 & n2592 ;
  assign n2594 = x65 & n2593 ;
  assign n2590 = x67 & n2428 ;
  assign n2595 = n2594 ^ n2590 ;
  assign n2596 = n2595 ^ x29 ;
  assign n2589 = ~n295 & n2429 ;
  assign n2597 = n2596 ^ n2589 ;
  assign n2588 = x66 & n2435 ;
  assign n2598 = n2597 ^ n2588 ;
  assign n2585 = x30 ^ x29 ;
  assign n2586 = x64 & n2585 ;
  assign n2587 = n2586 ^ n2451 ;
  assign n2599 = n2598 ^ n2587 ;
  assign n2608 = n2607 ^ n2599 ;
  assign n2582 = n2452 ^ n2425 ;
  assign n2583 = n2460 & ~n2582 ;
  assign n2584 = n2583 ^ n2425 ;
  assign n2609 = n2608 ^ n2584 ;
  assign n2610 = n2609 ^ x23 ;
  assign n2581 = x71 & n1665 ;
  assign n2611 = n2610 ^ n2581 ;
  assign n2580 = x73 & n1668 ;
  assign n2612 = n2611 ^ n2580 ;
  assign n2579 = n636 & n1669 ;
  assign n2613 = n2612 ^ n2579 ;
  assign n2615 = n2614 ^ n2613 ;
  assign n2576 = n2473 ^ n2469 ;
  assign n2577 = n2470 & n2576 ;
  assign n2578 = n2577 ^ n2473 ;
  assign n2616 = n2615 ^ n2578 ;
  assign n2617 = n2616 ^ x20 ;
  assign n2575 = x74 & n1340 ;
  assign n2618 = n2617 ^ n2575 ;
  assign n2574 = x76 & n1343 ;
  assign n2619 = n2618 ^ n2574 ;
  assign n2573 = ~n863 & n1344 ;
  assign n2620 = n2619 ^ n2573 ;
  assign n2622 = n2621 ^ n2620 ;
  assign n2626 = n2625 ^ n2622 ;
  assign n2627 = n2626 ^ x17 ;
  assign n2572 = x77 & n1060 ;
  assign n2628 = n2627 ^ n2572 ;
  assign n2571 = x79 & n1063 ;
  assign n2629 = n2628 ^ n2571 ;
  assign n2570 = n1064 & n1123 ;
  assign n2630 = n2629 ^ n2570 ;
  assign n2632 = n2631 ^ n2630 ;
  assign n2567 = n2490 ^ n2481 ;
  assign n2568 = n2487 & ~n2567 ;
  assign n2569 = n2568 ^ n2490 ;
  assign n2633 = n2632 ^ n2569 ;
  assign n2634 = n2633 ^ x14 ;
  assign n2566 = x80 & n884 ;
  assign n2635 = n2634 ^ n2566 ;
  assign n2565 = x82 & n789 ;
  assign n2636 = n2635 ^ n2565 ;
  assign n2564 = n790 & n1422 ;
  assign n2637 = n2636 ^ n2564 ;
  assign n2639 = n2638 ^ n2637 ;
  assign n2561 = n2500 ^ n2491 ;
  assign n2562 = n2497 & ~n2561 ;
  assign n2563 = n2562 ^ n2500 ;
  assign n2640 = n2639 ^ n2563 ;
  assign n2641 = n2640 ^ x11 ;
  assign n2560 = x83 & n650 ;
  assign n2642 = n2641 ^ n2560 ;
  assign n2559 = x85 & ~n578 ;
  assign n2643 = n2642 ^ n2559 ;
  assign n2558 = ~n579 & n1748 ;
  assign n2644 = n2643 ^ n2558 ;
  assign n2646 = n2645 ^ n2644 ;
  assign n2650 = n2649 ^ n2646 ;
  assign n2651 = n2650 ^ x8 ;
  assign n2557 = x86 & n456 ;
  assign n2652 = n2651 ^ n2557 ;
  assign n2556 = x88 & n384 ;
  assign n2653 = n2652 ^ n2556 ;
  assign n2555 = n385 & n2131 ;
  assign n2654 = n2653 ^ n2555 ;
  assign n2656 = n2655 ^ n2654 ;
  assign n2552 = n2517 ^ n2508 ;
  assign n2553 = n2514 & ~n2552 ;
  assign n2554 = n2553 ^ n2517 ;
  assign n2657 = n2656 ^ n2554 ;
  assign n2658 = n2657 ^ x5 ;
  assign n2551 = x89 & n238 ;
  assign n2659 = n2658 ^ n2551 ;
  assign n2550 = x91 & n234 ;
  assign n2660 = n2659 ^ n2550 ;
  assign n2548 = n2114 ^ x91 ;
  assign n2549 = n235 & n2548 ;
  assign n2661 = n2660 ^ n2549 ;
  assign n2663 = n2662 ^ n2661 ;
  assign n2667 = n2666 ^ n2663 ;
  assign n2531 = x93 ^ x91 ;
  assign n2529 = x93 ^ x92 ;
  assign n2532 = ~n2241 & n2529 ;
  assign n2533 = ~n2531 & n2532 ;
  assign n2534 = n2533 ^ n2529 ;
  assign n2536 = x94 ^ x1 ;
  assign n2535 = x94 ^ x2 ;
  assign n2537 = n2536 ^ n2535 ;
  assign n2538 = ~n2534 & n2537 ;
  assign n2539 = n2538 ^ n2536 ;
  assign n2668 = n2667 ^ n2539 ;
  assign n2543 = x2 & x92 ;
  assign n2544 = n2543 ^ x93 ;
  assign n2545 = ~x1 & n2544 ;
  assign n2540 = n2539 ^ n2382 ;
  assign n2546 = n2545 ^ n2540 ;
  assign n2547 = ~x0 & n2546 ;
  assign n2669 = n2668 ^ n2547 ;
  assign n2673 = n2672 ^ n2669 ;
  assign n2820 = x91 & n231 ;
  assign n2812 = n2650 ^ n2554 ;
  assign n2813 = n2656 & n2812 ;
  assign n2814 = n2813 ^ n2650 ;
  assign n2810 = x88 & n391 ;
  assign n2803 = x85 & n584 ;
  assign n2795 = n2633 ^ n2563 ;
  assign n2796 = ~n2639 & ~n2795 ;
  assign n2797 = n2796 ^ n2633 ;
  assign n2793 = x82 & n795 ;
  assign n2785 = n2626 ^ n2569 ;
  assign n2786 = ~n2632 & ~n2785 ;
  assign n2787 = n2786 ^ n2626 ;
  assign n2783 = x79 & n1068 ;
  assign n2776 = x76 & n1348 ;
  assign n2768 = n2609 ^ n2578 ;
  assign n2769 = n2615 & n2768 ;
  assign n2770 = n2769 ^ n2609 ;
  assign n2766 = x73 & n1673 ;
  assign n2758 = x67 & n2435 ;
  assign n2756 = ~n351 & n2429 ;
  assign n2752 = x66 & n2593 ;
  assign n2751 = x68 & n2428 ;
  assign n2753 = n2752 ^ n2751 ;
  assign n2754 = n2753 ^ x29 ;
  assign n2746 = ~x29 & ~x30 ;
  assign n2747 = n2746 ^ n2585 ;
  assign n2748 = n2747 ^ x31 ;
  assign n2749 = ~x64 & ~n2748 ;
  assign n2740 = x65 ^ x30 ;
  assign n2743 = x65 ^ x29 ;
  assign n2744 = ~n2740 & n2743 ;
  assign n2741 = x31 ^ x29 ;
  assign n2745 = n2744 ^ n2741 ;
  assign n2750 = n2749 ^ n2745 ;
  assign n2755 = n2754 ^ n2750 ;
  assign n2757 = n2756 ^ n2755 ;
  assign n2759 = n2758 ^ n2757 ;
  assign n2737 = ~n2451 & n2598 ;
  assign n2738 = ~n2586 & n2737 ;
  assign n2739 = n2738 ^ n2598 ;
  assign n2760 = n2759 ^ n2739 ;
  assign n2727 = x69 & n2032 ;
  assign n2726 = x71 & n2028 ;
  assign n2728 = n2727 ^ n2726 ;
  assign n2729 = n2728 ^ x26 ;
  assign n2725 = ~n495 & n2029 ;
  assign n2730 = n2729 ^ n2725 ;
  assign n2724 = x70 & n2025 ;
  assign n2731 = n2730 ^ n2724 ;
  assign n2732 = n2731 ^ n2607 ;
  assign n2733 = n2732 ^ n2584 ;
  assign n2734 = n2733 ^ n2731 ;
  assign n2735 = n2608 & n2734 ;
  assign n2736 = n2735 ^ n2732 ;
  assign n2761 = n2760 ^ n2736 ;
  assign n2762 = n2761 ^ x23 ;
  assign n2723 = x72 & n1665 ;
  assign n2763 = n2762 ^ n2723 ;
  assign n2722 = x74 & n1668 ;
  assign n2764 = n2763 ^ n2722 ;
  assign n2721 = n708 & n1669 ;
  assign n2765 = n2764 ^ n2721 ;
  assign n2767 = n2766 ^ n2765 ;
  assign n2771 = n2770 ^ n2767 ;
  assign n2772 = n2771 ^ x20 ;
  assign n2720 = x75 & n1340 ;
  assign n2773 = n2772 ^ n2720 ;
  assign n2719 = x77 & n1343 ;
  assign n2774 = n2773 ^ n2719 ;
  assign n2718 = ~n943 & n1344 ;
  assign n2775 = n2774 ^ n2718 ;
  assign n2777 = n2776 ^ n2775 ;
  assign n2715 = n2625 ^ n2616 ;
  assign n2716 = ~n2622 & ~n2715 ;
  assign n2717 = n2716 ^ n2625 ;
  assign n2778 = n2777 ^ n2717 ;
  assign n2779 = n2778 ^ x17 ;
  assign n2714 = x78 & n1060 ;
  assign n2780 = n2779 ^ n2714 ;
  assign n2713 = x80 & n1063 ;
  assign n2781 = n2780 ^ n2713 ;
  assign n2712 = n1064 & n1217 ;
  assign n2782 = n2781 ^ n2712 ;
  assign n2784 = n2783 ^ n2782 ;
  assign n2788 = n2787 ^ n2784 ;
  assign n2789 = n2788 ^ x14 ;
  assign n2711 = x81 & n884 ;
  assign n2790 = n2789 ^ n2711 ;
  assign n2710 = x83 & n789 ;
  assign n2791 = n2790 ^ n2710 ;
  assign n2709 = n790 & n1517 ;
  assign n2792 = n2791 ^ n2709 ;
  assign n2794 = n2793 ^ n2792 ;
  assign n2798 = n2797 ^ n2794 ;
  assign n2799 = n2798 ^ x11 ;
  assign n2708 = x84 & n650 ;
  assign n2800 = n2799 ^ n2708 ;
  assign n2707 = x86 & ~n578 ;
  assign n2801 = n2800 ^ n2707 ;
  assign n2706 = ~n579 & n1868 ;
  assign n2802 = n2801 ^ n2706 ;
  assign n2804 = n2803 ^ n2802 ;
  assign n2703 = n2649 ^ n2640 ;
  assign n2704 = n2646 & n2703 ;
  assign n2705 = n2704 ^ n2649 ;
  assign n2805 = n2804 ^ n2705 ;
  assign n2806 = n2805 ^ x8 ;
  assign n2702 = x87 & n456 ;
  assign n2807 = n2806 ^ n2702 ;
  assign n2701 = x89 & n384 ;
  assign n2808 = n2807 ^ n2701 ;
  assign n2700 = n385 & n2255 ;
  assign n2809 = n2808 ^ n2700 ;
  assign n2811 = n2810 ^ n2809 ;
  assign n2815 = n2814 ^ n2811 ;
  assign n2816 = n2815 ^ x5 ;
  assign n2699 = x90 & n238 ;
  assign n2817 = n2816 ^ n2699 ;
  assign n2698 = x92 & n234 ;
  assign n2818 = n2817 ^ n2698 ;
  assign n2696 = n2241 ^ x92 ;
  assign n2697 = n235 & n2696 ;
  assign n2819 = n2818 ^ n2697 ;
  assign n2821 = n2820 ^ n2819 ;
  assign n2693 = n2666 ^ n2657 ;
  assign n2694 = ~n2663 & ~n2693 ;
  assign n2695 = n2694 ^ n2666 ;
  assign n2822 = n2821 ^ n2695 ;
  assign n2677 = x94 ^ x93 ;
  assign n2679 = ~n2534 & n2677 ;
  assign n2681 = x95 ^ x1 ;
  assign n2680 = x95 ^ x2 ;
  assign n2682 = n2681 ^ n2680 ;
  assign n2683 = ~n2679 & n2682 ;
  assign n2684 = n2683 ^ n2681 ;
  assign n2823 = n2822 ^ n2684 ;
  assign n2688 = x2 & x93 ;
  assign n2689 = n2688 ^ x94 ;
  assign n2690 = ~n259 & n2689 ;
  assign n2685 = n2684 ^ n2535 ;
  assign n2691 = n2690 ^ n2685 ;
  assign n2692 = ~x0 & n2691 ;
  assign n2824 = n2823 ^ n2692 ;
  assign n2674 = n2672 ^ n2667 ;
  assign n2675 = n2669 & n2674 ;
  assign n2676 = n2675 ^ n2672 ;
  assign n2825 = n2824 ^ n2676 ;
  assign n2981 = n2822 ^ n2676 ;
  assign n2982 = ~n2824 & n2981 ;
  assign n2983 = n2982 ^ n2822 ;
  assign n2975 = n2815 ^ n2695 ;
  assign n2976 = n2821 & ~n2975 ;
  assign n2977 = n2976 ^ n2815 ;
  assign n2973 = x92 & n231 ;
  assign n2966 = x89 & n391 ;
  assign n2958 = n2798 ^ n2705 ;
  assign n2959 = ~n2804 & n2958 ;
  assign n2960 = n2959 ^ n2798 ;
  assign n2956 = x86 & n584 ;
  assign n2949 = x83 & n795 ;
  assign n2942 = x80 & n1068 ;
  assign n2934 = n2771 ^ n2717 ;
  assign n2935 = n2777 & ~n2934 ;
  assign n2936 = n2935 ^ n2771 ;
  assign n2932 = x77 & n1348 ;
  assign n2925 = x74 & n1673 ;
  assign n2918 = x71 & n2025 ;
  assign n2910 = n2750 ^ n2739 ;
  assign n2911 = n2759 & n2910 ;
  assign n2912 = n2911 ^ n2750 ;
  assign n2908 = x68 & n2435 ;
  assign n2898 = x31 ^ x30 ;
  assign n2899 = ~n2585 & n2898 ;
  assign n2900 = x65 & n2899 ;
  assign n2887 = x32 ^ x31 ;
  assign n2893 = n2585 & ~n2887 ;
  assign n2894 = n2893 ^ n2585 ;
  assign n2895 = ~n152 & n2894 ;
  assign n2892 = x66 & n2585 ;
  assign n2896 = n2895 ^ n2892 ;
  assign n2897 = n2896 ^ x32 ;
  assign n2901 = n2900 ^ n2897 ;
  assign n2888 = x32 ^ x30 ;
  assign n2889 = ~n2585 & n2888 ;
  assign n2890 = n2887 & n2889 ;
  assign n2891 = x64 & n2890 ;
  assign n2902 = n2901 ^ n2891 ;
  assign n2885 = ~n2586 & ~n2750 ;
  assign n2886 = x32 & n2885 ;
  assign n2903 = n2902 ^ n2886 ;
  assign n2904 = n2903 ^ x29 ;
  assign n2884 = x67 & n2593 ;
  assign n2905 = n2904 ^ n2884 ;
  assign n2883 = x69 & n2428 ;
  assign n2906 = n2905 ^ n2883 ;
  assign n2882 = ~n376 & n2429 ;
  assign n2907 = n2906 ^ n2882 ;
  assign n2909 = n2908 ^ n2907 ;
  assign n2913 = n2912 ^ n2909 ;
  assign n2914 = n2913 ^ x26 ;
  assign n2881 = x70 & n2032 ;
  assign n2915 = n2914 ^ n2881 ;
  assign n2880 = x72 & n2028 ;
  assign n2916 = n2915 ^ n2880 ;
  assign n2879 = n565 & n2029 ;
  assign n2917 = n2916 ^ n2879 ;
  assign n2919 = n2918 ^ n2917 ;
  assign n2876 = n2760 ^ n2731 ;
  assign n2877 = n2736 & n2876 ;
  assign n2878 = n2877 ^ n2731 ;
  assign n2920 = n2919 ^ n2878 ;
  assign n2921 = n2920 ^ x23 ;
  assign n2875 = x73 & n1665 ;
  assign n2922 = n2921 ^ n2875 ;
  assign n2874 = x75 & n1668 ;
  assign n2923 = n2922 ^ n2874 ;
  assign n2873 = ~n778 & n1669 ;
  assign n2924 = n2923 ^ n2873 ;
  assign n2926 = n2925 ^ n2924 ;
  assign n2870 = n2770 ^ n2761 ;
  assign n2871 = ~n2767 & n2870 ;
  assign n2872 = n2871 ^ n2770 ;
  assign n2927 = n2926 ^ n2872 ;
  assign n2928 = n2927 ^ x20 ;
  assign n2869 = x76 & n1340 ;
  assign n2929 = n2928 ^ n2869 ;
  assign n2868 = x78 & n1343 ;
  assign n2930 = n2929 ^ n2868 ;
  assign n2867 = ~n1036 & n1344 ;
  assign n2931 = n2930 ^ n2867 ;
  assign n2933 = n2932 ^ n2931 ;
  assign n2937 = n2936 ^ n2933 ;
  assign n2938 = n2937 ^ x17 ;
  assign n2866 = x79 & n1060 ;
  assign n2939 = n2938 ^ n2866 ;
  assign n2865 = x81 & n1063 ;
  assign n2940 = n2939 ^ n2865 ;
  assign n2864 = n1064 & n1310 ;
  assign n2941 = n2940 ^ n2864 ;
  assign n2943 = n2942 ^ n2941 ;
  assign n2861 = n2787 ^ n2778 ;
  assign n2862 = n2784 & n2861 ;
  assign n2863 = n2862 ^ n2787 ;
  assign n2944 = n2943 ^ n2863 ;
  assign n2945 = n2944 ^ x14 ;
  assign n2860 = x82 & n884 ;
  assign n2946 = n2945 ^ n2860 ;
  assign n2859 = x84 & n789 ;
  assign n2947 = n2946 ^ n2859 ;
  assign n2858 = n790 & n1635 ;
  assign n2948 = n2947 ^ n2858 ;
  assign n2950 = n2949 ^ n2948 ;
  assign n2855 = n2797 ^ n2788 ;
  assign n2856 = ~n2794 & ~n2855 ;
  assign n2857 = n2856 ^ n2797 ;
  assign n2951 = n2950 ^ n2857 ;
  assign n2952 = n2951 ^ x11 ;
  assign n2854 = x85 & n650 ;
  assign n2953 = n2952 ^ n2854 ;
  assign n2853 = x87 & ~n578 ;
  assign n2954 = n2953 ^ n2853 ;
  assign n2852 = ~n579 & n1987 ;
  assign n2955 = n2954 ^ n2852 ;
  assign n2957 = n2956 ^ n2955 ;
  assign n2961 = n2960 ^ n2957 ;
  assign n2962 = n2961 ^ x8 ;
  assign n2851 = x88 & n456 ;
  assign n2963 = n2962 ^ n2851 ;
  assign n2850 = x90 & n384 ;
  assign n2964 = n2963 ^ n2850 ;
  assign n2849 = n385 & n2398 ;
  assign n2965 = n2964 ^ n2849 ;
  assign n2967 = n2966 ^ n2965 ;
  assign n2846 = n2814 ^ n2805 ;
  assign n2847 = ~n2811 & n2846 ;
  assign n2848 = n2847 ^ n2814 ;
  assign n2968 = n2967 ^ n2848 ;
  assign n2969 = n2968 ^ x5 ;
  assign n2845 = x91 & n238 ;
  assign n2970 = n2969 ^ n2845 ;
  assign n2844 = x93 & n234 ;
  assign n2971 = n2970 ^ n2844 ;
  assign n2842 = n2381 ^ x93 ;
  assign n2843 = n235 & n2842 ;
  assign n2972 = n2971 ^ n2843 ;
  assign n2974 = n2973 ^ n2972 ;
  assign n2978 = n2977 ^ n2974 ;
  assign n2826 = x95 ^ x94 ;
  assign n2828 = ~n2679 & n2826 ;
  assign n2830 = x96 ^ x1 ;
  assign n2829 = x96 ^ x2 ;
  assign n2831 = n2830 ^ n2829 ;
  assign n2832 = ~n2828 & n2831 ;
  assign n2833 = n2832 ^ n2830 ;
  assign n2979 = n2978 ^ n2833 ;
  assign n2837 = x2 & x94 ;
  assign n2838 = n2837 ^ x95 ;
  assign n2839 = ~x1 & n2838 ;
  assign n2834 = n2833 ^ n2680 ;
  assign n2840 = n2839 ^ n2834 ;
  assign n2841 = ~x0 & n2840 ;
  assign n2980 = n2979 ^ n2841 ;
  assign n2984 = n2983 ^ n2980 ;
  assign n3135 = x93 & n231 ;
  assign n3127 = n2961 ^ n2848 ;
  assign n3128 = ~n2967 & ~n3127 ;
  assign n3129 = n3128 ^ n2961 ;
  assign n3125 = x90 & n391 ;
  assign n3118 = x87 & n584 ;
  assign n3110 = n2944 ^ n2857 ;
  assign n3111 = ~n2950 & n3110 ;
  assign n3112 = n3111 ^ n2944 ;
  assign n3108 = x84 & n795 ;
  assign n3100 = n2937 ^ n2863 ;
  assign n3101 = n2943 & ~n3100 ;
  assign n3102 = n3101 ^ n2937 ;
  assign n3098 = x81 & n1068 ;
  assign n3091 = x78 & n1348 ;
  assign n3083 = n2920 ^ n2872 ;
  assign n3084 = n2926 & n3083 ;
  assign n3085 = n3084 ^ n2920 ;
  assign n3081 = x75 & n1673 ;
  assign n3074 = x72 & n2025 ;
  assign n3067 = x69 & n2435 ;
  assign n3056 = x65 & n2890 ;
  assign n3055 = x67 & n2893 ;
  assign n3057 = n3056 ^ n3055 ;
  assign n3058 = n3057 ^ x32 ;
  assign n3054 = ~n295 & n2894 ;
  assign n3059 = n3058 ^ n3054 ;
  assign n3053 = x66 & n2899 ;
  assign n3060 = n3059 ^ n3053 ;
  assign n3051 = x33 ^ x32 ;
  assign n3052 = x64 & n3051 ;
  assign n3061 = n3060 ^ n3052 ;
  assign n3050 = n2886 & n2902 ;
  assign n3062 = n3061 ^ n3050 ;
  assign n3063 = n3062 ^ x29 ;
  assign n3049 = x68 & n2593 ;
  assign n3064 = n3063 ^ n3049 ;
  assign n3048 = x70 & n2428 ;
  assign n3065 = n3064 ^ n3048 ;
  assign n3047 = ~n443 & n2429 ;
  assign n3066 = n3065 ^ n3047 ;
  assign n3068 = n3067 ^ n3066 ;
  assign n3044 = n2912 ^ n2903 ;
  assign n3045 = ~n2909 & n3044 ;
  assign n3046 = n3045 ^ n2912 ;
  assign n3069 = n3068 ^ n3046 ;
  assign n3070 = n3069 ^ x26 ;
  assign n3043 = x71 & n2032 ;
  assign n3071 = n3070 ^ n3043 ;
  assign n3042 = x73 & n2028 ;
  assign n3072 = n3071 ^ n3042 ;
  assign n3041 = n636 & n2029 ;
  assign n3073 = n3072 ^ n3041 ;
  assign n3075 = n3074 ^ n3073 ;
  assign n3038 = n2913 ^ n2878 ;
  assign n3039 = n2919 & n3038 ;
  assign n3040 = n3039 ^ n2913 ;
  assign n3076 = n3075 ^ n3040 ;
  assign n3077 = n3076 ^ x23 ;
  assign n3037 = x74 & n1665 ;
  assign n3078 = n3077 ^ n3037 ;
  assign n3036 = x76 & n1668 ;
  assign n3079 = n3078 ^ n3036 ;
  assign n3035 = ~n863 & n1669 ;
  assign n3080 = n3079 ^ n3035 ;
  assign n3082 = n3081 ^ n3080 ;
  assign n3086 = n3085 ^ n3082 ;
  assign n3087 = n3086 ^ x20 ;
  assign n3034 = x77 & n1340 ;
  assign n3088 = n3087 ^ n3034 ;
  assign n3033 = x79 & n1343 ;
  assign n3089 = n3088 ^ n3033 ;
  assign n3032 = n1123 & n1344 ;
  assign n3090 = n3089 ^ n3032 ;
  assign n3092 = n3091 ^ n3090 ;
  assign n3029 = n2936 ^ n2927 ;
  assign n3030 = ~n2933 & n3029 ;
  assign n3031 = n3030 ^ n2936 ;
  assign n3093 = n3092 ^ n3031 ;
  assign n3094 = n3093 ^ x17 ;
  assign n3028 = x80 & n1060 ;
  assign n3095 = n3094 ^ n3028 ;
  assign n3027 = x82 & n1063 ;
  assign n3096 = n3095 ^ n3027 ;
  assign n3026 = n1064 & n1422 ;
  assign n3097 = n3096 ^ n3026 ;
  assign n3099 = n3098 ^ n3097 ;
  assign n3103 = n3102 ^ n3099 ;
  assign n3104 = n3103 ^ x14 ;
  assign n3025 = x83 & n884 ;
  assign n3105 = n3104 ^ n3025 ;
  assign n3024 = x85 & n789 ;
  assign n3106 = n3105 ^ n3024 ;
  assign n3023 = n790 & n1748 ;
  assign n3107 = n3106 ^ n3023 ;
  assign n3109 = n3108 ^ n3107 ;
  assign n3113 = n3112 ^ n3109 ;
  assign n3114 = n3113 ^ x11 ;
  assign n3022 = x86 & n650 ;
  assign n3115 = n3114 ^ n3022 ;
  assign n3021 = x88 & ~n578 ;
  assign n3116 = n3115 ^ n3021 ;
  assign n3020 = ~n579 & n2131 ;
  assign n3117 = n3116 ^ n3020 ;
  assign n3119 = n3118 ^ n3117 ;
  assign n3017 = n2960 ^ n2951 ;
  assign n3018 = ~n2957 & ~n3017 ;
  assign n3019 = n3018 ^ n2960 ;
  assign n3120 = n3119 ^ n3019 ;
  assign n3121 = n3120 ^ x8 ;
  assign n3016 = x89 & n456 ;
  assign n3122 = n3121 ^ n3016 ;
  assign n3015 = x91 & n384 ;
  assign n3123 = n3122 ^ n3015 ;
  assign n3014 = n385 & n2548 ;
  assign n3124 = n3123 ^ n3014 ;
  assign n3126 = n3125 ^ n3124 ;
  assign n3130 = n3129 ^ n3126 ;
  assign n3131 = n3130 ^ x5 ;
  assign n3013 = x92 & n238 ;
  assign n3132 = n3131 ^ n3013 ;
  assign n3012 = x94 & n234 ;
  assign n3133 = n3132 ^ n3012 ;
  assign n3010 = n2534 ^ x94 ;
  assign n3011 = n235 & n3010 ;
  assign n3134 = n3133 ^ n3011 ;
  assign n3136 = n3135 ^ n3134 ;
  assign n3007 = n2977 ^ n2968 ;
  assign n3008 = n2974 & ~n3007 ;
  assign n3009 = n3008 ^ n2977 ;
  assign n3137 = n3136 ^ n3009 ;
  assign n2990 = x96 ^ x94 ;
  assign n2988 = x96 ^ x95 ;
  assign n2991 = ~n2679 & n2988 ;
  assign n2992 = ~n2990 & n2991 ;
  assign n2993 = n2992 ^ n2988 ;
  assign n2995 = x97 ^ x1 ;
  assign n2994 = x97 ^ x2 ;
  assign n2996 = n2995 ^ n2994 ;
  assign n2997 = ~n2993 & n2996 ;
  assign n2998 = n2997 ^ n2995 ;
  assign n3138 = n3137 ^ n2998 ;
  assign n3002 = x2 & x95 ;
  assign n3003 = n3002 ^ x96 ;
  assign n3004 = ~x1 & n3003 ;
  assign n2999 = n2998 ^ n2829 ;
  assign n3005 = n3004 ^ n2999 ;
  assign n3006 = ~x0 & n3005 ;
  assign n3139 = n3138 ^ n3006 ;
  assign n2985 = n2983 ^ n2978 ;
  assign n2986 = n2980 & n2985 ;
  assign n2987 = n2986 ^ n2983 ;
  assign n3140 = n3139 ^ n2987 ;
  assign n3310 = n3137 ^ n2987 ;
  assign n3311 = ~n3139 & n3310 ;
  assign n3312 = n3311 ^ n3137 ;
  assign n3304 = n3130 ^ n3009 ;
  assign n3305 = ~n3136 & ~n3304 ;
  assign n3306 = n3305 ^ n3130 ;
  assign n3302 = x94 & n231 ;
  assign n3295 = x91 & n391 ;
  assign n3287 = n3113 ^ n3019 ;
  assign n3288 = ~n3119 & n3287 ;
  assign n3289 = n3288 ^ n3113 ;
  assign n3285 = x88 & n584 ;
  assign n3278 = x85 & n795 ;
  assign n3271 = x82 & n1068 ;
  assign n3263 = n3086 ^ n3031 ;
  assign n3264 = n3092 & n3263 ;
  assign n3265 = n3264 ^ n3086 ;
  assign n3261 = x79 & n1348 ;
  assign n3254 = x76 & n1673 ;
  assign n3246 = n3069 ^ n3040 ;
  assign n3247 = n3075 & n3246 ;
  assign n3248 = n3247 ^ n3069 ;
  assign n3244 = x73 & n2025 ;
  assign n3236 = n3062 ^ n3046 ;
  assign n3237 = n3068 & n3236 ;
  assign n3238 = n3237 ^ n3062 ;
  assign n3234 = x70 & n2435 ;
  assign n3227 = x67 & n2899 ;
  assign n3225 = ~n351 & n2894 ;
  assign n3219 = x32 & x33 ;
  assign n3220 = n3219 ^ x34 ;
  assign n3221 = ~x64 & n3220 ;
  assign n3215 = x34 ^ x32 ;
  assign n3222 = n3221 ^ n3215 ;
  assign n3213 = x65 ^ x33 ;
  assign n3214 = n3051 & ~n3213 ;
  assign n3223 = n3222 ^ n3214 ;
  assign n3210 = x66 & n2890 ;
  assign n3209 = x68 & n2893 ;
  assign n3211 = n3210 ^ n3209 ;
  assign n3212 = n3211 ^ x32 ;
  assign n3224 = n3223 ^ n3212 ;
  assign n3226 = n3225 ^ n3224 ;
  assign n3228 = n3227 ^ n3226 ;
  assign n3206 = ~n3052 & n3060 ;
  assign n3207 = ~n3050 & n3206 ;
  assign n3208 = n3207 ^ n3060 ;
  assign n3229 = n3228 ^ n3208 ;
  assign n3230 = n3229 ^ x29 ;
  assign n3205 = x69 & n2593 ;
  assign n3231 = n3230 ^ n3205 ;
  assign n3204 = x71 & n2428 ;
  assign n3232 = n3231 ^ n3204 ;
  assign n3203 = ~n495 & n2429 ;
  assign n3233 = n3232 ^ n3203 ;
  assign n3235 = n3234 ^ n3233 ;
  assign n3239 = n3238 ^ n3235 ;
  assign n3240 = n3239 ^ x26 ;
  assign n3202 = x72 & n2032 ;
  assign n3241 = n3240 ^ n3202 ;
  assign n3201 = x74 & n2028 ;
  assign n3242 = n3241 ^ n3201 ;
  assign n3200 = n708 & n2029 ;
  assign n3243 = n3242 ^ n3200 ;
  assign n3245 = n3244 ^ n3243 ;
  assign n3249 = n3248 ^ n3245 ;
  assign n3250 = n3249 ^ x23 ;
  assign n3199 = x75 & n1665 ;
  assign n3251 = n3250 ^ n3199 ;
  assign n3198 = x77 & n1668 ;
  assign n3252 = n3251 ^ n3198 ;
  assign n3197 = ~n943 & n1669 ;
  assign n3253 = n3252 ^ n3197 ;
  assign n3255 = n3254 ^ n3253 ;
  assign n3194 = n3085 ^ n3076 ;
  assign n3195 = ~n3082 & n3194 ;
  assign n3196 = n3195 ^ n3085 ;
  assign n3256 = n3255 ^ n3196 ;
  assign n3257 = n3256 ^ x20 ;
  assign n3193 = x78 & n1340 ;
  assign n3258 = n3257 ^ n3193 ;
  assign n3192 = x80 & n1343 ;
  assign n3259 = n3258 ^ n3192 ;
  assign n3191 = n1217 & n1344 ;
  assign n3260 = n3259 ^ n3191 ;
  assign n3262 = n3261 ^ n3260 ;
  assign n3266 = n3265 ^ n3262 ;
  assign n3267 = n3266 ^ x17 ;
  assign n3190 = x81 & n1060 ;
  assign n3268 = n3267 ^ n3190 ;
  assign n3189 = x83 & n1063 ;
  assign n3269 = n3268 ^ n3189 ;
  assign n3188 = n1064 & n1517 ;
  assign n3270 = n3269 ^ n3188 ;
  assign n3272 = n3271 ^ n3270 ;
  assign n3185 = n3102 ^ n3093 ;
  assign n3186 = ~n3099 & n3185 ;
  assign n3187 = n3186 ^ n3102 ;
  assign n3273 = n3272 ^ n3187 ;
  assign n3274 = n3273 ^ x14 ;
  assign n3184 = x84 & n884 ;
  assign n3275 = n3274 ^ n3184 ;
  assign n3183 = x86 & n789 ;
  assign n3276 = n3275 ^ n3183 ;
  assign n3182 = n790 & n1868 ;
  assign n3277 = n3276 ^ n3182 ;
  assign n3279 = n3278 ^ n3277 ;
  assign n3179 = n3112 ^ n3103 ;
  assign n3180 = ~n3109 & ~n3179 ;
  assign n3181 = n3180 ^ n3112 ;
  assign n3280 = n3279 ^ n3181 ;
  assign n3281 = n3280 ^ x11 ;
  assign n3178 = x87 & n650 ;
  assign n3282 = n3281 ^ n3178 ;
  assign n3177 = x89 & ~n578 ;
  assign n3283 = n3282 ^ n3177 ;
  assign n3176 = ~n579 & n2255 ;
  assign n3284 = n3283 ^ n3176 ;
  assign n3286 = n3285 ^ n3284 ;
  assign n3290 = n3289 ^ n3286 ;
  assign n3291 = n3290 ^ x8 ;
  assign n3175 = x90 & n456 ;
  assign n3292 = n3291 ^ n3175 ;
  assign n3174 = x92 & n384 ;
  assign n3293 = n3292 ^ n3174 ;
  assign n3173 = n385 & n2696 ;
  assign n3294 = n3293 ^ n3173 ;
  assign n3296 = n3295 ^ n3294 ;
  assign n3170 = n3129 ^ n3120 ;
  assign n3171 = ~n3126 & ~n3170 ;
  assign n3172 = n3171 ^ n3129 ;
  assign n3297 = n3296 ^ n3172 ;
  assign n3298 = n3297 ^ x5 ;
  assign n3169 = x93 & n238 ;
  assign n3299 = n3298 ^ n3169 ;
  assign n3168 = x95 & n234 ;
  assign n3300 = n3299 ^ n3168 ;
  assign n3166 = n2679 ^ x95 ;
  assign n3167 = n235 & n3166 ;
  assign n3301 = n3300 ^ n3167 ;
  assign n3303 = n3302 ^ n3301 ;
  assign n3307 = n3306 ^ n3303 ;
  assign n3141 = x97 ^ x96 ;
  assign n3145 = n2988 ^ x94 ;
  assign n3146 = n3145 ^ x97 ;
  assign n3147 = n3146 ^ n2988 ;
  assign n3148 = n2991 & n3147 ;
  assign n3149 = n3148 ^ n2988 ;
  assign n3150 = n3141 & n3149 ;
  assign n3151 = n3150 ^ x96 ;
  assign n3152 = n3151 ^ x97 ;
  assign n3154 = x98 ^ x1 ;
  assign n3153 = x98 ^ x2 ;
  assign n3155 = n3154 ^ n3153 ;
  assign n3156 = ~n3152 & n3155 ;
  assign n3157 = n3156 ^ n3154 ;
  assign n3308 = n3307 ^ n3157 ;
  assign n3161 = x2 & x96 ;
  assign n3162 = n3161 ^ x97 ;
  assign n3163 = ~x1 & n3162 ;
  assign n3158 = n3157 ^ n2994 ;
  assign n3164 = n3163 ^ n3158 ;
  assign n3165 = ~x0 & n3164 ;
  assign n3309 = n3308 ^ n3165 ;
  assign n3313 = n3312 ^ n3309 ;
  assign n3479 = x95 & n231 ;
  assign n3471 = n3290 ^ n3172 ;
  assign n3472 = n3296 & ~n3471 ;
  assign n3473 = n3472 ^ n3290 ;
  assign n3469 = x92 & n391 ;
  assign n3462 = x89 & n584 ;
  assign n3454 = n3273 ^ n3181 ;
  assign n3455 = n3279 & ~n3454 ;
  assign n3456 = n3455 ^ n3273 ;
  assign n3452 = x86 & n795 ;
  assign n3444 = n3266 ^ n3187 ;
  assign n3445 = n3272 & n3444 ;
  assign n3446 = n3445 ^ n3266 ;
  assign n3442 = x83 & n1068 ;
  assign n3435 = x80 & n1348 ;
  assign n3427 = n3249 ^ n3196 ;
  assign n3428 = n3255 & n3427 ;
  assign n3429 = n3428 ^ n3249 ;
  assign n3425 = x77 & n1673 ;
  assign n3418 = x74 & n2025 ;
  assign n3411 = x71 & n2435 ;
  assign n3404 = x68 & n2899 ;
  assign n3217 = x34 ^ x33 ;
  assign n3395 = ~n3051 & n3217 ;
  assign n3396 = x65 & n3395 ;
  assign n3384 = x35 ^ x34 ;
  assign n3390 = n3051 & ~n3384 ;
  assign n3391 = n3390 ^ n3051 ;
  assign n3392 = ~n152 & n3391 ;
  assign n3389 = x66 & n3051 ;
  assign n3393 = n3392 ^ n3389 ;
  assign n3394 = n3393 ^ x35 ;
  assign n3397 = n3396 ^ n3394 ;
  assign n3385 = x35 ^ x33 ;
  assign n3386 = ~n3051 & n3385 ;
  assign n3387 = n3384 & n3386 ;
  assign n3388 = x64 & n3387 ;
  assign n3398 = n3397 ^ n3388 ;
  assign n3382 = ~n3052 & ~n3223 ;
  assign n3383 = x35 & n3382 ;
  assign n3399 = n3398 ^ n3383 ;
  assign n3400 = n3399 ^ x32 ;
  assign n3381 = x67 & n2890 ;
  assign n3401 = n3400 ^ n3381 ;
  assign n3380 = x69 & n2893 ;
  assign n3402 = n3401 ^ n3380 ;
  assign n3379 = ~n376 & n2894 ;
  assign n3403 = n3402 ^ n3379 ;
  assign n3405 = n3404 ^ n3403 ;
  assign n3376 = n3223 ^ n3208 ;
  assign n3377 = n3228 & n3376 ;
  assign n3378 = n3377 ^ n3223 ;
  assign n3406 = n3405 ^ n3378 ;
  assign n3407 = n3406 ^ x29 ;
  assign n3375 = x70 & n2593 ;
  assign n3408 = n3407 ^ n3375 ;
  assign n3374 = x72 & n2428 ;
  assign n3409 = n3408 ^ n3374 ;
  assign n3373 = n565 & n2429 ;
  assign n3410 = n3409 ^ n3373 ;
  assign n3412 = n3411 ^ n3410 ;
  assign n3370 = n3238 ^ n3229 ;
  assign n3371 = ~n3235 & n3370 ;
  assign n3372 = n3371 ^ n3238 ;
  assign n3413 = n3412 ^ n3372 ;
  assign n3414 = n3413 ^ x26 ;
  assign n3369 = x73 & n2032 ;
  assign n3415 = n3414 ^ n3369 ;
  assign n3368 = x75 & n2028 ;
  assign n3416 = n3415 ^ n3368 ;
  assign n3367 = ~n778 & n2029 ;
  assign n3417 = n3416 ^ n3367 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n3364 = n3248 ^ n3239 ;
  assign n3365 = ~n3245 & n3364 ;
  assign n3366 = n3365 ^ n3248 ;
  assign n3420 = n3419 ^ n3366 ;
  assign n3421 = n3420 ^ x23 ;
  assign n3363 = x76 & n1665 ;
  assign n3422 = n3421 ^ n3363 ;
  assign n3362 = x78 & n1668 ;
  assign n3423 = n3422 ^ n3362 ;
  assign n3361 = ~n1036 & n1669 ;
  assign n3424 = n3423 ^ n3361 ;
  assign n3426 = n3425 ^ n3424 ;
  assign n3430 = n3429 ^ n3426 ;
  assign n3431 = n3430 ^ x20 ;
  assign n3360 = x79 & n1340 ;
  assign n3432 = n3431 ^ n3360 ;
  assign n3359 = x81 & n1343 ;
  assign n3433 = n3432 ^ n3359 ;
  assign n3358 = n1310 & n1344 ;
  assign n3434 = n3433 ^ n3358 ;
  assign n3436 = n3435 ^ n3434 ;
  assign n3355 = n3265 ^ n3256 ;
  assign n3356 = ~n3262 & n3355 ;
  assign n3357 = n3356 ^ n3265 ;
  assign n3437 = n3436 ^ n3357 ;
  assign n3438 = n3437 ^ x17 ;
  assign n3354 = x82 & n1060 ;
  assign n3439 = n3438 ^ n3354 ;
  assign n3353 = x84 & n1063 ;
  assign n3440 = n3439 ^ n3353 ;
  assign n3352 = n1064 & n1635 ;
  assign n3441 = n3440 ^ n3352 ;
  assign n3443 = n3442 ^ n3441 ;
  assign n3447 = n3446 ^ n3443 ;
  assign n3448 = n3447 ^ x14 ;
  assign n3351 = x85 & n884 ;
  assign n3449 = n3448 ^ n3351 ;
  assign n3350 = x87 & n789 ;
  assign n3450 = n3449 ^ n3350 ;
  assign n3349 = n790 & n1987 ;
  assign n3451 = n3450 ^ n3349 ;
  assign n3453 = n3452 ^ n3451 ;
  assign n3457 = n3456 ^ n3453 ;
  assign n3458 = n3457 ^ x11 ;
  assign n3348 = x88 & n650 ;
  assign n3459 = n3458 ^ n3348 ;
  assign n3347 = x90 & ~n578 ;
  assign n3460 = n3459 ^ n3347 ;
  assign n3346 = ~n579 & n2398 ;
  assign n3461 = n3460 ^ n3346 ;
  assign n3463 = n3462 ^ n3461 ;
  assign n3343 = n3289 ^ n3280 ;
  assign n3344 = n3286 & n3343 ;
  assign n3345 = n3344 ^ n3289 ;
  assign n3464 = n3463 ^ n3345 ;
  assign n3465 = n3464 ^ x8 ;
  assign n3342 = x91 & n456 ;
  assign n3466 = n3465 ^ n3342 ;
  assign n3341 = x93 & n384 ;
  assign n3467 = n3466 ^ n3341 ;
  assign n3340 = n385 & n2842 ;
  assign n3468 = n3467 ^ n3340 ;
  assign n3470 = n3469 ^ n3468 ;
  assign n3474 = n3473 ^ n3470 ;
  assign n3475 = n3474 ^ x5 ;
  assign n3339 = x94 & n238 ;
  assign n3476 = n3475 ^ n3339 ;
  assign n3338 = x96 & n234 ;
  assign n3477 = n3476 ^ n3338 ;
  assign n3336 = n2828 ^ x96 ;
  assign n3337 = n235 & n3336 ;
  assign n3478 = n3477 ^ n3337 ;
  assign n3480 = n3479 ^ n3478 ;
  assign n3333 = n3306 ^ n3297 ;
  assign n3334 = n3303 & n3333 ;
  assign n3335 = n3334 ^ n3306 ;
  assign n3481 = n3480 ^ n3335 ;
  assign n3317 = x98 ^ x97 ;
  assign n3319 = ~n3152 & n3317 ;
  assign n3321 = x99 ^ x1 ;
  assign n3320 = x99 ^ x2 ;
  assign n3322 = n3321 ^ n3320 ;
  assign n3323 = ~n3319 & n3322 ;
  assign n3324 = n3323 ^ n3321 ;
  assign n3482 = n3481 ^ n3324 ;
  assign n3328 = x2 & x97 ;
  assign n3329 = n3328 ^ x98 ;
  assign n3330 = ~x1 & n3329 ;
  assign n3325 = n3324 ^ n3153 ;
  assign n3331 = n3330 ^ n3325 ;
  assign n3332 = ~x0 & n3331 ;
  assign n3483 = n3482 ^ n3332 ;
  assign n3314 = n3312 ^ n3307 ;
  assign n3315 = ~n3309 & ~n3314 ;
  assign n3316 = n3315 ^ n3312 ;
  assign n3484 = n3483 ^ n3316 ;
  assign n3647 = n3481 ^ n3316 ;
  assign n3648 = n3483 & ~n3647 ;
  assign n3649 = n3648 ^ n3481 ;
  assign n3641 = n3474 ^ n3335 ;
  assign n3642 = ~n3480 & n3641 ;
  assign n3643 = n3642 ^ n3474 ;
  assign n3639 = x96 & n231 ;
  assign n3632 = x93 & n391 ;
  assign n3624 = n3457 ^ n3345 ;
  assign n3625 = n3463 & ~n3624 ;
  assign n3626 = n3625 ^ n3457 ;
  assign n3622 = x90 & n584 ;
  assign n3615 = x87 & n795 ;
  assign n3608 = x84 & n1068 ;
  assign n3600 = n3430 ^ n3357 ;
  assign n3601 = n3436 & n3600 ;
  assign n3602 = n3601 ^ n3430 ;
  assign n3598 = x81 & n1348 ;
  assign n3591 = x78 & n1673 ;
  assign n3583 = n3413 ^ n3366 ;
  assign n3584 = n3419 & n3583 ;
  assign n3585 = n3584 ^ n3413 ;
  assign n3581 = x75 & n2025 ;
  assign n3573 = n3406 ^ n3372 ;
  assign n3574 = n3412 & n3573 ;
  assign n3575 = n3574 ^ n3406 ;
  assign n3567 = x71 & n2593 ;
  assign n3566 = x73 & n2428 ;
  assign n3568 = n3567 ^ n3566 ;
  assign n3569 = n3568 ^ x29 ;
  assign n3565 = n636 & n2429 ;
  assign n3570 = n3569 ^ n3565 ;
  assign n3564 = x72 & n2435 ;
  assign n3571 = n3570 ^ n3564 ;
  assign n3560 = n3399 ^ n3378 ;
  assign n3561 = n3405 & n3560 ;
  assign n3562 = n3561 ^ n3399 ;
  assign n3558 = x69 & n2899 ;
  assign n3547 = x65 & n3387 ;
  assign n3546 = x67 & n3390 ;
  assign n3548 = n3547 ^ n3546 ;
  assign n3549 = n3548 ^ x35 ;
  assign n3545 = ~n295 & n3391 ;
  assign n3550 = n3549 ^ n3545 ;
  assign n3544 = x66 & n3395 ;
  assign n3551 = n3550 ^ n3544 ;
  assign n3542 = x36 ^ x35 ;
  assign n3543 = x64 & n3542 ;
  assign n3552 = n3551 ^ n3543 ;
  assign n3541 = n3383 & n3398 ;
  assign n3553 = n3552 ^ n3541 ;
  assign n3554 = n3553 ^ x32 ;
  assign n3540 = x68 & n2890 ;
  assign n3555 = n3554 ^ n3540 ;
  assign n3539 = x70 & n2893 ;
  assign n3556 = n3555 ^ n3539 ;
  assign n3538 = ~n443 & n2894 ;
  assign n3557 = n3556 ^ n3538 ;
  assign n3559 = n3558 ^ n3557 ;
  assign n3563 = n3562 ^ n3559 ;
  assign n3572 = n3571 ^ n3563 ;
  assign n3576 = n3575 ^ n3572 ;
  assign n3577 = n3576 ^ x26 ;
  assign n3537 = x74 & n2032 ;
  assign n3578 = n3577 ^ n3537 ;
  assign n3536 = x76 & n2028 ;
  assign n3579 = n3578 ^ n3536 ;
  assign n3535 = ~n863 & n2029 ;
  assign n3580 = n3579 ^ n3535 ;
  assign n3582 = n3581 ^ n3580 ;
  assign n3586 = n3585 ^ n3582 ;
  assign n3587 = n3586 ^ x23 ;
  assign n3534 = x77 & n1665 ;
  assign n3588 = n3587 ^ n3534 ;
  assign n3533 = x79 & n1668 ;
  assign n3589 = n3588 ^ n3533 ;
  assign n3532 = n1123 & n1669 ;
  assign n3590 = n3589 ^ n3532 ;
  assign n3592 = n3591 ^ n3590 ;
  assign n3529 = n3429 ^ n3420 ;
  assign n3530 = ~n3426 & n3529 ;
  assign n3531 = n3530 ^ n3429 ;
  assign n3593 = n3592 ^ n3531 ;
  assign n3594 = n3593 ^ x20 ;
  assign n3528 = x80 & n1340 ;
  assign n3595 = n3594 ^ n3528 ;
  assign n3527 = x82 & n1343 ;
  assign n3596 = n3595 ^ n3527 ;
  assign n3526 = n1344 & n1422 ;
  assign n3597 = n3596 ^ n3526 ;
  assign n3599 = n3598 ^ n3597 ;
  assign n3603 = n3602 ^ n3599 ;
  assign n3604 = n3603 ^ x17 ;
  assign n3525 = x83 & n1060 ;
  assign n3605 = n3604 ^ n3525 ;
  assign n3524 = x85 & n1063 ;
  assign n3606 = n3605 ^ n3524 ;
  assign n3523 = n1064 & n1748 ;
  assign n3607 = n3606 ^ n3523 ;
  assign n3609 = n3608 ^ n3607 ;
  assign n3520 = n3446 ^ n3437 ;
  assign n3521 = ~n3443 & n3520 ;
  assign n3522 = n3521 ^ n3446 ;
  assign n3610 = n3609 ^ n3522 ;
  assign n3611 = n3610 ^ x14 ;
  assign n3519 = x86 & n884 ;
  assign n3612 = n3611 ^ n3519 ;
  assign n3518 = x88 & n789 ;
  assign n3613 = n3612 ^ n3518 ;
  assign n3517 = n790 & n2131 ;
  assign n3614 = n3613 ^ n3517 ;
  assign n3616 = n3615 ^ n3614 ;
  assign n3514 = n3456 ^ n3447 ;
  assign n3515 = ~n3453 & n3514 ;
  assign n3516 = n3515 ^ n3456 ;
  assign n3617 = n3616 ^ n3516 ;
  assign n3618 = n3617 ^ x11 ;
  assign n3513 = x89 & n650 ;
  assign n3619 = n3618 ^ n3513 ;
  assign n3512 = x91 & ~n578 ;
  assign n3620 = n3619 ^ n3512 ;
  assign n3511 = ~n579 & n2548 ;
  assign n3621 = n3620 ^ n3511 ;
  assign n3623 = n3622 ^ n3621 ;
  assign n3627 = n3626 ^ n3623 ;
  assign n3628 = n3627 ^ x8 ;
  assign n3510 = x92 & n456 ;
  assign n3629 = n3628 ^ n3510 ;
  assign n3509 = x94 & n384 ;
  assign n3630 = n3629 ^ n3509 ;
  assign n3508 = n385 & n3010 ;
  assign n3631 = n3630 ^ n3508 ;
  assign n3633 = n3632 ^ n3631 ;
  assign n3505 = n3473 ^ n3464 ;
  assign n3506 = n3470 & ~n3505 ;
  assign n3507 = n3506 ^ n3473 ;
  assign n3634 = n3633 ^ n3507 ;
  assign n3635 = n3634 ^ x5 ;
  assign n3504 = x95 & n238 ;
  assign n3636 = n3635 ^ n3504 ;
  assign n3503 = x97 & n234 ;
  assign n3637 = n3636 ^ n3503 ;
  assign n3501 = n2993 ^ x97 ;
  assign n3502 = n235 & n3501 ;
  assign n3638 = n3637 ^ n3502 ;
  assign n3640 = n3639 ^ n3638 ;
  assign n3644 = n3643 ^ n3640 ;
  assign n3485 = x99 ^ x98 ;
  assign n3487 = ~n3319 & n3485 ;
  assign n3489 = x100 ^ x1 ;
  assign n3488 = x100 ^ x2 ;
  assign n3490 = n3489 ^ n3488 ;
  assign n3491 = ~n3487 & n3490 ;
  assign n3492 = n3491 ^ n3489 ;
  assign n3645 = n3644 ^ n3492 ;
  assign n3496 = x2 & x98 ;
  assign n3497 = n3496 ^ x99 ;
  assign n3498 = ~x1 & n3497 ;
  assign n3493 = n3492 ^ n3320 ;
  assign n3499 = n3498 ^ n3493 ;
  assign n3500 = ~x0 & n3499 ;
  assign n3646 = n3645 ^ n3500 ;
  assign n3650 = n3649 ^ n3646 ;
  assign n3823 = x97 & n231 ;
  assign n3815 = n3627 ^ n3507 ;
  assign n3816 = n3633 & n3815 ;
  assign n3817 = n3816 ^ n3627 ;
  assign n3813 = x94 & n391 ;
  assign n3806 = x91 & n584 ;
  assign n3798 = n3610 ^ n3516 ;
  assign n3799 = n3616 & n3798 ;
  assign n3800 = n3799 ^ n3610 ;
  assign n3796 = x88 & n795 ;
  assign n3788 = n3603 ^ n3522 ;
  assign n3789 = n3609 & n3788 ;
  assign n3790 = n3789 ^ n3603 ;
  assign n3786 = x85 & n1068 ;
  assign n3779 = x82 & n1348 ;
  assign n3771 = n3586 ^ n3531 ;
  assign n3772 = n3592 & n3771 ;
  assign n3773 = n3772 ^ n3586 ;
  assign n3769 = x79 & n1673 ;
  assign n3762 = x76 & n2025 ;
  assign n3755 = x73 & n2435 ;
  assign n3748 = x70 & n2899 ;
  assign n3727 = ~n3541 & ~n3543 ;
  assign n3741 = n3551 & n3727 ;
  assign n3734 = x35 & x36 ;
  assign n3735 = n3734 ^ x37 ;
  assign n3736 = ~x64 & n3735 ;
  assign n3730 = x37 ^ x35 ;
  assign n3737 = n3736 ^ n3730 ;
  assign n3728 = x65 ^ x36 ;
  assign n3729 = n3542 & ~n3728 ;
  assign n3738 = n3737 ^ n3729 ;
  assign n3739 = n3738 ^ n3551 ;
  assign n3742 = n3741 ^ n3739 ;
  assign n3722 = x66 & n3387 ;
  assign n3721 = x68 & n3390 ;
  assign n3723 = n3722 ^ n3721 ;
  assign n3724 = n3723 ^ x35 ;
  assign n3720 = ~n351 & n3391 ;
  assign n3725 = n3724 ^ n3720 ;
  assign n3719 = x67 & n3395 ;
  assign n3726 = n3725 ^ n3719 ;
  assign n3743 = n3742 ^ n3726 ;
  assign n3744 = n3743 ^ x32 ;
  assign n3718 = x69 & n2890 ;
  assign n3745 = n3744 ^ n3718 ;
  assign n3717 = x71 & n2893 ;
  assign n3746 = n3745 ^ n3717 ;
  assign n3716 = ~n495 & n2894 ;
  assign n3747 = n3746 ^ n3716 ;
  assign n3749 = n3748 ^ n3747 ;
  assign n3713 = n3562 ^ n3553 ;
  assign n3714 = ~n3559 & n3713 ;
  assign n3715 = n3714 ^ n3562 ;
  assign n3750 = n3749 ^ n3715 ;
  assign n3751 = n3750 ^ x29 ;
  assign n3712 = x72 & n2593 ;
  assign n3752 = n3751 ^ n3712 ;
  assign n3711 = x74 & n2428 ;
  assign n3753 = n3752 ^ n3711 ;
  assign n3710 = n708 & n2429 ;
  assign n3754 = n3753 ^ n3710 ;
  assign n3756 = n3755 ^ n3754 ;
  assign n3707 = n3575 ^ n3571 ;
  assign n3708 = ~n3572 & n3707 ;
  assign n3709 = n3708 ^ n3575 ;
  assign n3757 = n3756 ^ n3709 ;
  assign n3758 = n3757 ^ x26 ;
  assign n3706 = x75 & n2032 ;
  assign n3759 = n3758 ^ n3706 ;
  assign n3705 = x77 & n2028 ;
  assign n3760 = n3759 ^ n3705 ;
  assign n3704 = ~n943 & n2029 ;
  assign n3761 = n3760 ^ n3704 ;
  assign n3763 = n3762 ^ n3761 ;
  assign n3701 = n3585 ^ n3576 ;
  assign n3702 = ~n3582 & n3701 ;
  assign n3703 = n3702 ^ n3585 ;
  assign n3764 = n3763 ^ n3703 ;
  assign n3765 = n3764 ^ x23 ;
  assign n3700 = x78 & n1665 ;
  assign n3766 = n3765 ^ n3700 ;
  assign n3699 = x80 & n1668 ;
  assign n3767 = n3766 ^ n3699 ;
  assign n3698 = n1217 & n1669 ;
  assign n3768 = n3767 ^ n3698 ;
  assign n3770 = n3769 ^ n3768 ;
  assign n3774 = n3773 ^ n3770 ;
  assign n3775 = n3774 ^ x20 ;
  assign n3697 = x81 & n1340 ;
  assign n3776 = n3775 ^ n3697 ;
  assign n3696 = x83 & n1343 ;
  assign n3777 = n3776 ^ n3696 ;
  assign n3695 = n1344 & n1517 ;
  assign n3778 = n3777 ^ n3695 ;
  assign n3780 = n3779 ^ n3778 ;
  assign n3692 = n3602 ^ n3593 ;
  assign n3693 = ~n3599 & n3692 ;
  assign n3694 = n3693 ^ n3602 ;
  assign n3781 = n3780 ^ n3694 ;
  assign n3782 = n3781 ^ x17 ;
  assign n3691 = x84 & n1060 ;
  assign n3783 = n3782 ^ n3691 ;
  assign n3690 = x86 & n1063 ;
  assign n3784 = n3783 ^ n3690 ;
  assign n3689 = n1064 & n1868 ;
  assign n3785 = n3784 ^ n3689 ;
  assign n3787 = n3786 ^ n3785 ;
  assign n3791 = n3790 ^ n3787 ;
  assign n3792 = n3791 ^ x14 ;
  assign n3688 = x87 & n884 ;
  assign n3793 = n3792 ^ n3688 ;
  assign n3687 = x89 & n789 ;
  assign n3794 = n3793 ^ n3687 ;
  assign n3686 = n790 & n2255 ;
  assign n3795 = n3794 ^ n3686 ;
  assign n3797 = n3796 ^ n3795 ;
  assign n3801 = n3800 ^ n3797 ;
  assign n3802 = n3801 ^ x11 ;
  assign n3685 = x90 & n650 ;
  assign n3803 = n3802 ^ n3685 ;
  assign n3684 = x92 & ~n578 ;
  assign n3804 = n3803 ^ n3684 ;
  assign n3683 = ~n579 & n2696 ;
  assign n3805 = n3804 ^ n3683 ;
  assign n3807 = n3806 ^ n3805 ;
  assign n3680 = n3626 ^ n3617 ;
  assign n3681 = ~n3623 & n3680 ;
  assign n3682 = n3681 ^ n3626 ;
  assign n3808 = n3807 ^ n3682 ;
  assign n3809 = n3808 ^ x8 ;
  assign n3679 = x93 & n456 ;
  assign n3810 = n3809 ^ n3679 ;
  assign n3678 = x95 & n384 ;
  assign n3811 = n3810 ^ n3678 ;
  assign n3677 = n385 & n3166 ;
  assign n3812 = n3811 ^ n3677 ;
  assign n3814 = n3813 ^ n3812 ;
  assign n3818 = n3817 ^ n3814 ;
  assign n3819 = n3818 ^ x5 ;
  assign n3676 = x96 & n238 ;
  assign n3820 = n3819 ^ n3676 ;
  assign n3675 = x98 & n234 ;
  assign n3821 = n3820 ^ n3675 ;
  assign n3673 = n3317 ^ n3151 ;
  assign n3674 = n235 & n3673 ;
  assign n3822 = n3821 ^ n3674 ;
  assign n3824 = n3823 ^ n3822 ;
  assign n3670 = n3643 ^ n3634 ;
  assign n3671 = ~n3640 & ~n3670 ;
  assign n3672 = n3671 ^ n3643 ;
  assign n3825 = n3824 ^ n3672 ;
  assign n3654 = x100 ^ x99 ;
  assign n3656 = ~n3487 & n3654 ;
  assign n3658 = x101 ^ x1 ;
  assign n3657 = x101 ^ x2 ;
  assign n3659 = n3658 ^ n3657 ;
  assign n3660 = ~n3656 & n3659 ;
  assign n3661 = n3660 ^ n3658 ;
  assign n3826 = n3825 ^ n3661 ;
  assign n3665 = x2 & x99 ;
  assign n3666 = n3665 ^ x100 ;
  assign n3667 = ~n259 & n3666 ;
  assign n3662 = n3661 ^ n3488 ;
  assign n3668 = n3667 ^ n3662 ;
  assign n3669 = ~x0 & n3668 ;
  assign n3827 = n3826 ^ n3669 ;
  assign n3651 = n3649 ^ n3644 ;
  assign n3652 = n3646 & ~n3651 ;
  assign n3653 = n3652 ^ n3649 ;
  assign n3828 = n3827 ^ n3653 ;
  assign n4018 = n3825 ^ n3653 ;
  assign n4019 = ~n3827 & ~n4018 ;
  assign n4020 = n4019 ^ n3825 ;
  assign n4012 = n3818 ^ n3672 ;
  assign n4013 = n3824 & ~n4012 ;
  assign n4014 = n4013 ^ n3818 ;
  assign n4010 = x98 & n231 ;
  assign n4003 = x95 & n391 ;
  assign n3995 = n3801 ^ n3682 ;
  assign n3996 = n3807 & n3995 ;
  assign n3997 = n3996 ^ n3801 ;
  assign n3993 = x92 & n584 ;
  assign n3986 = x89 & n795 ;
  assign n3979 = x86 & n1068 ;
  assign n3971 = n3774 ^ n3694 ;
  assign n3972 = n3780 & n3971 ;
  assign n3973 = n3972 ^ n3774 ;
  assign n3969 = x83 & n1348 ;
  assign n3958 = n3743 ^ n3715 ;
  assign n3959 = n3749 & n3958 ;
  assign n3960 = n3959 ^ n3743 ;
  assign n3956 = x71 & n2899 ;
  assign n3949 = x68 & n3395 ;
  assign n3732 = x37 ^ x36 ;
  assign n3940 = ~n3542 & n3732 ;
  assign n3941 = x65 & n3940 ;
  assign n3929 = x38 ^ x37 ;
  assign n3935 = n3542 & ~n3929 ;
  assign n3936 = n3935 ^ n3542 ;
  assign n3937 = ~n152 & n3936 ;
  assign n3934 = x66 & n3542 ;
  assign n3938 = n3937 ^ n3934 ;
  assign n3939 = n3938 ^ x38 ;
  assign n3942 = n3941 ^ n3939 ;
  assign n3930 = x38 ^ x36 ;
  assign n3931 = ~n3542 & n3930 ;
  assign n3932 = n3929 & n3931 ;
  assign n3933 = x64 & n3932 ;
  assign n3943 = n3942 ^ n3933 ;
  assign n3927 = ~n3543 & ~n3738 ;
  assign n3928 = x38 & n3927 ;
  assign n3944 = n3943 ^ n3928 ;
  assign n3945 = n3944 ^ x35 ;
  assign n3926 = x67 & n3387 ;
  assign n3946 = n3945 ^ n3926 ;
  assign n3925 = x69 & n3390 ;
  assign n3947 = n3946 ^ n3925 ;
  assign n3924 = ~n376 & n3391 ;
  assign n3948 = n3947 ^ n3924 ;
  assign n3950 = n3949 ^ n3948 ;
  assign n3921 = n3738 ^ n3726 ;
  assign n3922 = n3742 & n3921 ;
  assign n3923 = n3922 ^ n3738 ;
  assign n3951 = n3950 ^ n3923 ;
  assign n3952 = n3951 ^ x32 ;
  assign n3920 = x70 & n2890 ;
  assign n3953 = n3952 ^ n3920 ;
  assign n3919 = x72 & n2893 ;
  assign n3954 = n3953 ^ n3919 ;
  assign n3918 = n565 & n2894 ;
  assign n3955 = n3954 ^ n3918 ;
  assign n3957 = n3956 ^ n3955 ;
  assign n3961 = n3960 ^ n3957 ;
  assign n3915 = n3750 ^ n3709 ;
  assign n3916 = n3756 & n3915 ;
  assign n3908 = x73 & n2593 ;
  assign n3907 = x75 & n2428 ;
  assign n3909 = n3908 ^ n3907 ;
  assign n3910 = n3909 ^ x29 ;
  assign n3906 = ~n778 & n2429 ;
  assign n3911 = n3910 ^ n3906 ;
  assign n3905 = x74 & n2435 ;
  assign n3912 = n3911 ^ n3905 ;
  assign n3913 = n3912 ^ n3750 ;
  assign n3917 = n3916 ^ n3913 ;
  assign n3962 = n3961 ^ n3917 ;
  assign n3902 = n3757 ^ n3703 ;
  assign n3903 = n3763 & n3902 ;
  assign n3895 = x76 & n2032 ;
  assign n3894 = x78 & n2028 ;
  assign n3896 = n3895 ^ n3894 ;
  assign n3897 = n3896 ^ x26 ;
  assign n3893 = ~n1036 & n2029 ;
  assign n3898 = n3897 ^ n3893 ;
  assign n3892 = x77 & n2025 ;
  assign n3899 = n3898 ^ n3892 ;
  assign n3900 = n3899 ^ n3757 ;
  assign n3904 = n3903 ^ n3900 ;
  assign n3963 = n3962 ^ n3904 ;
  assign n3882 = x79 & n1665 ;
  assign n3881 = x81 & n1668 ;
  assign n3883 = n3882 ^ n3881 ;
  assign n3884 = n3883 ^ x23 ;
  assign n3880 = n1310 & n1669 ;
  assign n3885 = n3884 ^ n3880 ;
  assign n3879 = x80 & n1673 ;
  assign n3886 = n3885 ^ n3879 ;
  assign n3887 = n3886 ^ n3773 ;
  assign n3888 = n3887 ^ n3764 ;
  assign n3889 = n3888 ^ n3886 ;
  assign n3890 = ~n3770 & n3889 ;
  assign n3891 = n3890 ^ n3887 ;
  assign n3964 = n3963 ^ n3891 ;
  assign n3965 = n3964 ^ x20 ;
  assign n3878 = x82 & n1340 ;
  assign n3966 = n3965 ^ n3878 ;
  assign n3877 = x84 & n1343 ;
  assign n3967 = n3966 ^ n3877 ;
  assign n3876 = n1344 & n1635 ;
  assign n3968 = n3967 ^ n3876 ;
  assign n3970 = n3969 ^ n3968 ;
  assign n3974 = n3973 ^ n3970 ;
  assign n3975 = n3974 ^ x17 ;
  assign n3875 = x85 & n1060 ;
  assign n3976 = n3975 ^ n3875 ;
  assign n3874 = x87 & n1063 ;
  assign n3977 = n3976 ^ n3874 ;
  assign n3873 = n1064 & n1987 ;
  assign n3978 = n3977 ^ n3873 ;
  assign n3980 = n3979 ^ n3978 ;
  assign n3870 = n3790 ^ n3781 ;
  assign n3871 = ~n3787 & n3870 ;
  assign n3872 = n3871 ^ n3790 ;
  assign n3981 = n3980 ^ n3872 ;
  assign n3982 = n3981 ^ x14 ;
  assign n3869 = x88 & n884 ;
  assign n3983 = n3982 ^ n3869 ;
  assign n3868 = x90 & n789 ;
  assign n3984 = n3983 ^ n3868 ;
  assign n3867 = n790 & n2398 ;
  assign n3985 = n3984 ^ n3867 ;
  assign n3987 = n3986 ^ n3985 ;
  assign n3864 = n3800 ^ n3791 ;
  assign n3865 = ~n3797 & n3864 ;
  assign n3866 = n3865 ^ n3800 ;
  assign n3988 = n3987 ^ n3866 ;
  assign n3989 = n3988 ^ x11 ;
  assign n3863 = x91 & n650 ;
  assign n3990 = n3989 ^ n3863 ;
  assign n3862 = x93 & ~n578 ;
  assign n3991 = n3990 ^ n3862 ;
  assign n3861 = ~n579 & n2842 ;
  assign n3992 = n3991 ^ n3861 ;
  assign n3994 = n3993 ^ n3992 ;
  assign n3998 = n3997 ^ n3994 ;
  assign n3999 = n3998 ^ x8 ;
  assign n3860 = x94 & n456 ;
  assign n4000 = n3999 ^ n3860 ;
  assign n3859 = x96 & n384 ;
  assign n4001 = n4000 ^ n3859 ;
  assign n3858 = n385 & n3336 ;
  assign n4002 = n4001 ^ n3858 ;
  assign n4004 = n4003 ^ n4002 ;
  assign n3855 = n3817 ^ n3808 ;
  assign n3856 = ~n3814 & n3855 ;
  assign n3857 = n3856 ^ n3817 ;
  assign n4005 = n4004 ^ n3857 ;
  assign n4006 = n4005 ^ x5 ;
  assign n3854 = x97 & n238 ;
  assign n4007 = n4006 ^ n3854 ;
  assign n3853 = x99 & n234 ;
  assign n4008 = n4007 ^ n3853 ;
  assign n3851 = n3319 ^ x99 ;
  assign n3852 = n235 & n3851 ;
  assign n4009 = n4008 ^ n3852 ;
  assign n4011 = n4010 ^ n4009 ;
  assign n4015 = n4014 ^ n4011 ;
  assign n3831 = x101 ^ x98 ;
  assign n3829 = x101 ^ x100 ;
  assign n3832 = n3654 & n3829 ;
  assign n3833 = ~n3319 & n3832 ;
  assign n3834 = n3831 & n3833 ;
  assign n3835 = n3834 ^ n3832 ;
  assign n3836 = n3835 ^ x100 ;
  assign n3837 = n3836 ^ x101 ;
  assign n3839 = x102 ^ x1 ;
  assign n3838 = x102 ^ x2 ;
  assign n3840 = n3839 ^ n3838 ;
  assign n3841 = ~n3837 & n3840 ;
  assign n3842 = n3841 ^ n3839 ;
  assign n4016 = n4015 ^ n3842 ;
  assign n3846 = x2 & x100 ;
  assign n3847 = n3846 ^ x101 ;
  assign n3848 = ~x1 & n3847 ;
  assign n3843 = n3842 ^ n3657 ;
  assign n3849 = n3848 ^ n3843 ;
  assign n3850 = ~x0 & n3849 ;
  assign n4017 = n4016 ^ n3850 ;
  assign n4021 = n4020 ^ n4017 ;
  assign n4199 = x99 & n231 ;
  assign n4191 = n3998 ^ n3857 ;
  assign n4192 = n4004 & n4191 ;
  assign n4193 = n4192 ^ n3998 ;
  assign n4189 = x96 & n391 ;
  assign n4182 = x93 & n584 ;
  assign n4174 = n3981 ^ n3866 ;
  assign n4175 = n3987 & n4174 ;
  assign n4176 = n4175 ^ n3981 ;
  assign n4172 = x90 & n795 ;
  assign n4164 = n3974 ^ n3872 ;
  assign n4165 = n3980 & n4164 ;
  assign n4166 = n4165 ^ n3974 ;
  assign n4162 = x87 & n1068 ;
  assign n4155 = x84 & n1348 ;
  assign n4148 = x81 & n1673 ;
  assign n4141 = x78 & n2025 ;
  assign n4134 = x75 & n2435 ;
  assign n4127 = x72 & n2899 ;
  assign n4120 = x69 & n3395 ;
  assign n4109 = x65 & n3932 ;
  assign n4108 = x67 & n3935 ;
  assign n4110 = n4109 ^ n4108 ;
  assign n4111 = n4110 ^ x38 ;
  assign n4107 = ~n295 & n3936 ;
  assign n4112 = n4111 ^ n4107 ;
  assign n4106 = x66 & n3940 ;
  assign n4113 = n4112 ^ n4106 ;
  assign n4104 = x39 ^ x38 ;
  assign n4105 = x64 & n4104 ;
  assign n4114 = n4113 ^ n4105 ;
  assign n4103 = n3928 & n3943 ;
  assign n4115 = n4114 ^ n4103 ;
  assign n4116 = n4115 ^ x35 ;
  assign n4102 = x68 & n3387 ;
  assign n4117 = n4116 ^ n4102 ;
  assign n4101 = x70 & n3390 ;
  assign n4118 = n4117 ^ n4101 ;
  assign n4100 = ~n443 & n3391 ;
  assign n4119 = n4118 ^ n4100 ;
  assign n4121 = n4120 ^ n4119 ;
  assign n4097 = n3944 ^ n3923 ;
  assign n4098 = n3950 & n4097 ;
  assign n4099 = n4098 ^ n3944 ;
  assign n4122 = n4121 ^ n4099 ;
  assign n4123 = n4122 ^ x32 ;
  assign n4096 = x71 & n2890 ;
  assign n4124 = n4123 ^ n4096 ;
  assign n4095 = x73 & n2893 ;
  assign n4125 = n4124 ^ n4095 ;
  assign n4094 = n636 & n2894 ;
  assign n4126 = n4125 ^ n4094 ;
  assign n4128 = n4127 ^ n4126 ;
  assign n4091 = n3960 ^ n3951 ;
  assign n4092 = ~n3957 & n4091 ;
  assign n4093 = n4092 ^ n3960 ;
  assign n4129 = n4128 ^ n4093 ;
  assign n4130 = n4129 ^ x29 ;
  assign n4090 = x74 & n2593 ;
  assign n4131 = n4130 ^ n4090 ;
  assign n4089 = x76 & n2428 ;
  assign n4132 = n4131 ^ n4089 ;
  assign n4088 = ~n863 & n2429 ;
  assign n4133 = n4132 ^ n4088 ;
  assign n4135 = n4134 ^ n4133 ;
  assign n4085 = n3961 ^ n3912 ;
  assign n4086 = n3917 & n4085 ;
  assign n4087 = n4086 ^ n3912 ;
  assign n4136 = n4135 ^ n4087 ;
  assign n4137 = n4136 ^ x26 ;
  assign n4084 = x77 & n2032 ;
  assign n4138 = n4137 ^ n4084 ;
  assign n4083 = x79 & n2028 ;
  assign n4139 = n4138 ^ n4083 ;
  assign n4082 = n1123 & n2029 ;
  assign n4140 = n4139 ^ n4082 ;
  assign n4142 = n4141 ^ n4140 ;
  assign n4079 = n3962 ^ n3899 ;
  assign n4080 = n3904 & n4079 ;
  assign n4081 = n4080 ^ n3899 ;
  assign n4143 = n4142 ^ n4081 ;
  assign n4144 = n4143 ^ x23 ;
  assign n4078 = x80 & n1665 ;
  assign n4145 = n4144 ^ n4078 ;
  assign n4077 = x82 & n1668 ;
  assign n4146 = n4145 ^ n4077 ;
  assign n4076 = n1422 & n1669 ;
  assign n4147 = n4146 ^ n4076 ;
  assign n4149 = n4148 ^ n4147 ;
  assign n4073 = n3963 ^ n3886 ;
  assign n4074 = n3891 & n4073 ;
  assign n4075 = n4074 ^ n3886 ;
  assign n4150 = n4149 ^ n4075 ;
  assign n4151 = n4150 ^ x20 ;
  assign n4072 = x83 & n1340 ;
  assign n4152 = n4151 ^ n4072 ;
  assign n4071 = x85 & n1343 ;
  assign n4153 = n4152 ^ n4071 ;
  assign n4070 = n1344 & n1748 ;
  assign n4154 = n4153 ^ n4070 ;
  assign n4156 = n4155 ^ n4154 ;
  assign n4067 = n3973 ^ n3964 ;
  assign n4068 = ~n3970 & n4067 ;
  assign n4069 = n4068 ^ n3973 ;
  assign n4157 = n4156 ^ n4069 ;
  assign n4158 = n4157 ^ x17 ;
  assign n4066 = x86 & n1060 ;
  assign n4159 = n4158 ^ n4066 ;
  assign n4065 = x88 & n1063 ;
  assign n4160 = n4159 ^ n4065 ;
  assign n4064 = n1064 & n2131 ;
  assign n4161 = n4160 ^ n4064 ;
  assign n4163 = n4162 ^ n4161 ;
  assign n4167 = n4166 ^ n4163 ;
  assign n4168 = n4167 ^ x14 ;
  assign n4063 = x89 & n884 ;
  assign n4169 = n4168 ^ n4063 ;
  assign n4062 = x91 & n789 ;
  assign n4170 = n4169 ^ n4062 ;
  assign n4061 = n790 & n2548 ;
  assign n4171 = n4170 ^ n4061 ;
  assign n4173 = n4172 ^ n4171 ;
  assign n4177 = n4176 ^ n4173 ;
  assign n4178 = n4177 ^ x11 ;
  assign n4060 = x92 & n650 ;
  assign n4179 = n4178 ^ n4060 ;
  assign n4059 = x94 & ~n578 ;
  assign n4180 = n4179 ^ n4059 ;
  assign n4058 = ~n579 & n3010 ;
  assign n4181 = n4180 ^ n4058 ;
  assign n4183 = n4182 ^ n4181 ;
  assign n4055 = n3997 ^ n3988 ;
  assign n4056 = ~n3994 & n4055 ;
  assign n4057 = n4056 ^ n3997 ;
  assign n4184 = n4183 ^ n4057 ;
  assign n4185 = n4184 ^ x8 ;
  assign n4054 = x95 & n456 ;
  assign n4186 = n4185 ^ n4054 ;
  assign n4053 = x97 & n384 ;
  assign n4187 = n4186 ^ n4053 ;
  assign n4052 = n385 & n3501 ;
  assign n4188 = n4187 ^ n4052 ;
  assign n4190 = n4189 ^ n4188 ;
  assign n4194 = n4193 ^ n4190 ;
  assign n4195 = n4194 ^ x5 ;
  assign n4051 = x98 & n238 ;
  assign n4196 = n4195 ^ n4051 ;
  assign n4050 = x100 & n234 ;
  assign n4197 = n4196 ^ n4050 ;
  assign n4048 = n3487 ^ x100 ;
  assign n4049 = n235 & n4048 ;
  assign n4198 = n4197 ^ n4049 ;
  assign n4200 = n4199 ^ n4198 ;
  assign n4045 = n4014 ^ n4005 ;
  assign n4046 = ~n4011 & n4045 ;
  assign n4047 = n4046 ^ n4014 ;
  assign n4201 = n4200 ^ n4047 ;
  assign n4027 = x101 & n3836 ;
  assign n4029 = n4027 ^ n3837 ;
  assign n4030 = x102 & n4029 ;
  assign n4028 = ~x102 & ~n4027 ;
  assign n4031 = n4030 ^ n4028 ;
  assign n4033 = x103 ^ x1 ;
  assign n4032 = x103 ^ x2 ;
  assign n4034 = n4033 ^ n4032 ;
  assign n4035 = n4031 & n4034 ;
  assign n4036 = n4035 ^ n4033 ;
  assign n4202 = n4201 ^ n4036 ;
  assign n4040 = x2 & x101 ;
  assign n4041 = n4040 ^ x102 ;
  assign n4042 = ~x1 & n4041 ;
  assign n4037 = n4036 ^ n3838 ;
  assign n4043 = n4042 ^ n4037 ;
  assign n4044 = ~x0 & n4043 ;
  assign n4203 = n4202 ^ n4044 ;
  assign n4022 = n4020 ^ n4015 ;
  assign n4023 = ~n4017 & ~n4022 ;
  assign n4024 = n4023 ^ n4020 ;
  assign n4204 = n4203 ^ n4024 ;
  assign n4397 = n4201 ^ n4024 ;
  assign n4398 = n4203 & ~n4397 ;
  assign n4399 = n4398 ^ n4201 ;
  assign n4391 = n4194 ^ n4047 ;
  assign n4392 = n4200 & n4391 ;
  assign n4393 = n4392 ^ n4194 ;
  assign n4389 = x100 & n231 ;
  assign n4382 = x97 & n391 ;
  assign n4374 = n4177 ^ n4057 ;
  assign n4375 = n4183 & n4374 ;
  assign n4376 = n4375 ^ n4177 ;
  assign n4372 = x94 & n584 ;
  assign n4365 = x91 & n795 ;
  assign n4358 = x88 & n1068 ;
  assign n4350 = n4150 ^ n4069 ;
  assign n4351 = n4156 & n4350 ;
  assign n4352 = n4351 ^ n4150 ;
  assign n4348 = x85 & n1348 ;
  assign n4341 = x82 & n1673 ;
  assign n4334 = x79 & n2025 ;
  assign n4327 = x76 & n2435 ;
  assign n4319 = n4122 ^ n4093 ;
  assign n4320 = n4128 & n4319 ;
  assign n4321 = n4320 ^ n4122 ;
  assign n4317 = x73 & n2899 ;
  assign n4293 = ~n4103 & ~n4105 ;
  assign n4309 = n4113 & n4293 ;
  assign n4300 = ~x38 & ~x39 ;
  assign n4301 = n4300 ^ x40 ;
  assign n4302 = ~x64 & ~n4301 ;
  assign n4303 = n4302 ^ n4104 ;
  assign n4304 = n4303 ^ n4105 ;
  assign n4296 = x40 ^ x38 ;
  assign n4305 = n4304 ^ n4296 ;
  assign n4294 = x65 ^ x39 ;
  assign n4295 = n4104 & ~n4294 ;
  assign n4306 = n4305 ^ n4295 ;
  assign n4307 = n4306 ^ n4113 ;
  assign n4310 = n4309 ^ n4307 ;
  assign n4288 = x66 & n3932 ;
  assign n4287 = x68 & n3935 ;
  assign n4289 = n4288 ^ n4287 ;
  assign n4290 = n4289 ^ x38 ;
  assign n4286 = ~n351 & n3936 ;
  assign n4291 = n4290 ^ n4286 ;
  assign n4285 = x67 & n3940 ;
  assign n4292 = n4291 ^ n4285 ;
  assign n4311 = n4310 ^ n4292 ;
  assign n4282 = n4115 ^ n4099 ;
  assign n4283 = n4121 & n4282 ;
  assign n4275 = x69 & n3387 ;
  assign n4274 = x71 & n3390 ;
  assign n4276 = n4275 ^ n4274 ;
  assign n4277 = n4276 ^ x35 ;
  assign n4273 = ~n495 & n3391 ;
  assign n4278 = n4277 ^ n4273 ;
  assign n4272 = x70 & n3395 ;
  assign n4279 = n4278 ^ n4272 ;
  assign n4280 = n4279 ^ n4115 ;
  assign n4284 = n4283 ^ n4280 ;
  assign n4312 = n4311 ^ n4284 ;
  assign n4313 = n4312 ^ x32 ;
  assign n4271 = x72 & n2890 ;
  assign n4314 = n4313 ^ n4271 ;
  assign n4270 = x74 & n2893 ;
  assign n4315 = n4314 ^ n4270 ;
  assign n4269 = n708 & n2894 ;
  assign n4316 = n4315 ^ n4269 ;
  assign n4318 = n4317 ^ n4316 ;
  assign n4322 = n4321 ^ n4318 ;
  assign n4323 = n4322 ^ x29 ;
  assign n4268 = x75 & n2593 ;
  assign n4324 = n4323 ^ n4268 ;
  assign n4267 = x77 & n2428 ;
  assign n4325 = n4324 ^ n4267 ;
  assign n4266 = ~n943 & n2429 ;
  assign n4326 = n4325 ^ n4266 ;
  assign n4328 = n4327 ^ n4326 ;
  assign n4263 = n4129 ^ n4087 ;
  assign n4264 = n4135 & n4263 ;
  assign n4265 = n4264 ^ n4129 ;
  assign n4329 = n4328 ^ n4265 ;
  assign n4330 = n4329 ^ x26 ;
  assign n4262 = x78 & n2032 ;
  assign n4331 = n4330 ^ n4262 ;
  assign n4261 = x80 & n2028 ;
  assign n4332 = n4331 ^ n4261 ;
  assign n4260 = n1217 & n2029 ;
  assign n4333 = n4332 ^ n4260 ;
  assign n4335 = n4334 ^ n4333 ;
  assign n4257 = n4136 ^ n4081 ;
  assign n4258 = n4142 & n4257 ;
  assign n4259 = n4258 ^ n4136 ;
  assign n4336 = n4335 ^ n4259 ;
  assign n4337 = n4336 ^ x23 ;
  assign n4256 = x81 & n1665 ;
  assign n4338 = n4337 ^ n4256 ;
  assign n4255 = x83 & n1668 ;
  assign n4339 = n4338 ^ n4255 ;
  assign n4254 = n1517 & n1669 ;
  assign n4340 = n4339 ^ n4254 ;
  assign n4342 = n4341 ^ n4340 ;
  assign n4251 = n4143 ^ n4075 ;
  assign n4252 = n4149 & n4251 ;
  assign n4253 = n4252 ^ n4143 ;
  assign n4343 = n4342 ^ n4253 ;
  assign n4344 = n4343 ^ x20 ;
  assign n4250 = x84 & n1340 ;
  assign n4345 = n4344 ^ n4250 ;
  assign n4249 = x86 & n1343 ;
  assign n4346 = n4345 ^ n4249 ;
  assign n4248 = n1344 & n1868 ;
  assign n4347 = n4346 ^ n4248 ;
  assign n4349 = n4348 ^ n4347 ;
  assign n4353 = n4352 ^ n4349 ;
  assign n4354 = n4353 ^ x17 ;
  assign n4247 = x87 & n1060 ;
  assign n4355 = n4354 ^ n4247 ;
  assign n4246 = x89 & n1063 ;
  assign n4356 = n4355 ^ n4246 ;
  assign n4245 = n1064 & n2255 ;
  assign n4357 = n4356 ^ n4245 ;
  assign n4359 = n4358 ^ n4357 ;
  assign n4242 = n4166 ^ n4157 ;
  assign n4243 = ~n4163 & n4242 ;
  assign n4244 = n4243 ^ n4166 ;
  assign n4360 = n4359 ^ n4244 ;
  assign n4361 = n4360 ^ x14 ;
  assign n4241 = x90 & n884 ;
  assign n4362 = n4361 ^ n4241 ;
  assign n4240 = x92 & n789 ;
  assign n4363 = n4362 ^ n4240 ;
  assign n4239 = n790 & n2696 ;
  assign n4364 = n4363 ^ n4239 ;
  assign n4366 = n4365 ^ n4364 ;
  assign n4236 = n4176 ^ n4167 ;
  assign n4237 = ~n4173 & n4236 ;
  assign n4238 = n4237 ^ n4176 ;
  assign n4367 = n4366 ^ n4238 ;
  assign n4368 = n4367 ^ x11 ;
  assign n4235 = x93 & n650 ;
  assign n4369 = n4368 ^ n4235 ;
  assign n4234 = x95 & ~n578 ;
  assign n4370 = n4369 ^ n4234 ;
  assign n4233 = ~n579 & n3166 ;
  assign n4371 = n4370 ^ n4233 ;
  assign n4373 = n4372 ^ n4371 ;
  assign n4377 = n4376 ^ n4373 ;
  assign n4378 = n4377 ^ x8 ;
  assign n4232 = x96 & n456 ;
  assign n4379 = n4378 ^ n4232 ;
  assign n4231 = x98 & n384 ;
  assign n4380 = n4379 ^ n4231 ;
  assign n4230 = n385 & n3673 ;
  assign n4381 = n4380 ^ n4230 ;
  assign n4383 = n4382 ^ n4381 ;
  assign n4227 = n4193 ^ n4184 ;
  assign n4228 = ~n4190 & n4227 ;
  assign n4229 = n4228 ^ n4193 ;
  assign n4384 = n4383 ^ n4229 ;
  assign n4385 = n4384 ^ x5 ;
  assign n4226 = x99 & n238 ;
  assign n4386 = n4385 ^ n4226 ;
  assign n4225 = x101 & n234 ;
  assign n4387 = n4386 ^ n4225 ;
  assign n4223 = n3656 ^ x101 ;
  assign n4224 = n235 & n4223 ;
  assign n4388 = n4387 ^ n4224 ;
  assign n4390 = n4389 ^ n4388 ;
  assign n4394 = n4393 ^ n4390 ;
  assign n4208 = ~x103 & ~n4030 ;
  assign n4207 = x103 & ~n4028 ;
  assign n4209 = n4208 ^ n4207 ;
  assign n4211 = x104 ^ x1 ;
  assign n4210 = x104 ^ x2 ;
  assign n4212 = n4211 ^ n4210 ;
  assign n4213 = n4209 & n4212 ;
  assign n4214 = n4213 ^ n4211 ;
  assign n4395 = n4394 ^ n4214 ;
  assign n4218 = x2 & x102 ;
  assign n4219 = n4218 ^ x103 ;
  assign n4220 = ~x1 & n4219 ;
  assign n4215 = n4214 ^ n4032 ;
  assign n4221 = n4220 ^ n4215 ;
  assign n4222 = ~x0 & n4221 ;
  assign n4396 = n4395 ^ n4222 ;
  assign n4400 = n4399 ^ n4396 ;
  assign n4600 = x101 & n231 ;
  assign n4592 = n4377 ^ n4229 ;
  assign n4593 = n4383 & n4592 ;
  assign n4594 = n4593 ^ n4377 ;
  assign n4590 = x98 & n391 ;
  assign n4583 = x95 & n584 ;
  assign n4575 = n4360 ^ n4238 ;
  assign n4576 = n4366 & n4575 ;
  assign n4577 = n4576 ^ n4360 ;
  assign n4573 = x92 & n795 ;
  assign n4565 = n4353 ^ n4244 ;
  assign n4566 = n4359 & n4565 ;
  assign n4567 = n4566 ^ n4353 ;
  assign n4563 = x89 & n1068 ;
  assign n4556 = x86 & n1348 ;
  assign n4548 = n4336 ^ n4253 ;
  assign n4549 = n4342 & n4548 ;
  assign n4550 = n4549 ^ n4336 ;
  assign n4546 = x83 & n1673 ;
  assign n4538 = n4329 ^ n4259 ;
  assign n4539 = n4335 & n4538 ;
  assign n4540 = n4539 ^ n4329 ;
  assign n4536 = x80 & n2025 ;
  assign n4528 = n4322 ^ n4265 ;
  assign n4529 = n4328 & n4528 ;
  assign n4530 = n4529 ^ n4322 ;
  assign n4526 = x77 & n2435 ;
  assign n4519 = x74 & n2899 ;
  assign n4512 = x71 & n3395 ;
  assign n4504 = n4306 ^ n4292 ;
  assign n4505 = n4310 & n4504 ;
  assign n4506 = n4505 ^ n4306 ;
  assign n4498 = x67 & n3932 ;
  assign n4497 = x69 & n3935 ;
  assign n4499 = n4498 ^ n4497 ;
  assign n4500 = n4499 ^ x38 ;
  assign n4496 = ~n376 & n3936 ;
  assign n4501 = n4500 ^ n4496 ;
  assign n4495 = x68 & n3940 ;
  assign n4502 = n4501 ^ n4495 ;
  assign n4491 = x66 & n4104 ;
  assign n4477 = x41 ^ x40 ;
  assign n4478 = n4104 & ~n4477 ;
  assign n4479 = n4478 ^ n4104 ;
  assign n4487 = x65 & n4479 ;
  assign n4480 = x41 ^ x39 ;
  assign n4481 = ~n4104 & n4480 ;
  assign n4482 = n4477 & n4481 ;
  assign n4488 = n4487 ^ n4482 ;
  assign n4489 = ~x64 & n4488 ;
  assign n4490 = n4489 ^ n4482 ;
  assign n4492 = n4491 ^ n4490 ;
  assign n4298 = x40 ^ x39 ;
  assign n4475 = ~n4104 & n4298 ;
  assign n4476 = x65 & n4475 ;
  assign n4493 = n4492 ^ n4476 ;
  assign n4471 = x41 & ~n151 ;
  assign n4472 = n4302 ^ n4298 ;
  assign n4473 = ~n4104 & ~n4472 ;
  assign n4474 = n4471 & ~n4473 ;
  assign n4494 = n4493 ^ n4474 ;
  assign n4503 = n4502 ^ n4494 ;
  assign n4507 = n4506 ^ n4503 ;
  assign n4508 = n4507 ^ x35 ;
  assign n4470 = x70 & n3387 ;
  assign n4509 = n4508 ^ n4470 ;
  assign n4469 = x72 & n3390 ;
  assign n4510 = n4509 ^ n4469 ;
  assign n4468 = n565 & n3391 ;
  assign n4511 = n4510 ^ n4468 ;
  assign n4513 = n4512 ^ n4511 ;
  assign n4465 = n4311 ^ n4279 ;
  assign n4466 = n4284 & n4465 ;
  assign n4467 = n4466 ^ n4279 ;
  assign n4514 = n4513 ^ n4467 ;
  assign n4515 = n4514 ^ x32 ;
  assign n4464 = x73 & n2890 ;
  assign n4516 = n4515 ^ n4464 ;
  assign n4463 = x75 & n2893 ;
  assign n4517 = n4516 ^ n4463 ;
  assign n4462 = ~n778 & n2894 ;
  assign n4518 = n4517 ^ n4462 ;
  assign n4520 = n4519 ^ n4518 ;
  assign n4459 = n4321 ^ n4312 ;
  assign n4460 = ~n4318 & n4459 ;
  assign n4461 = n4460 ^ n4321 ;
  assign n4521 = n4520 ^ n4461 ;
  assign n4522 = n4521 ^ x29 ;
  assign n4458 = x76 & n2593 ;
  assign n4523 = n4522 ^ n4458 ;
  assign n4457 = x78 & n2428 ;
  assign n4524 = n4523 ^ n4457 ;
  assign n4456 = ~n1036 & n2429 ;
  assign n4525 = n4524 ^ n4456 ;
  assign n4527 = n4526 ^ n4525 ;
  assign n4531 = n4530 ^ n4527 ;
  assign n4532 = n4531 ^ x26 ;
  assign n4455 = x79 & n2032 ;
  assign n4533 = n4532 ^ n4455 ;
  assign n4454 = x81 & n2028 ;
  assign n4534 = n4533 ^ n4454 ;
  assign n4453 = n1310 & n2029 ;
  assign n4535 = n4534 ^ n4453 ;
  assign n4537 = n4536 ^ n4535 ;
  assign n4541 = n4540 ^ n4537 ;
  assign n4542 = n4541 ^ x23 ;
  assign n4452 = x82 & n1665 ;
  assign n4543 = n4542 ^ n4452 ;
  assign n4451 = x84 & n1668 ;
  assign n4544 = n4543 ^ n4451 ;
  assign n4450 = n1635 & n1669 ;
  assign n4545 = n4544 ^ n4450 ;
  assign n4547 = n4546 ^ n4545 ;
  assign n4551 = n4550 ^ n4547 ;
  assign n4552 = n4551 ^ x20 ;
  assign n4449 = x85 & n1340 ;
  assign n4553 = n4552 ^ n4449 ;
  assign n4448 = x87 & n1343 ;
  assign n4554 = n4553 ^ n4448 ;
  assign n4447 = n1344 & n1987 ;
  assign n4555 = n4554 ^ n4447 ;
  assign n4557 = n4556 ^ n4555 ;
  assign n4444 = n4352 ^ n4343 ;
  assign n4445 = ~n4349 & n4444 ;
  assign n4446 = n4445 ^ n4352 ;
  assign n4558 = n4557 ^ n4446 ;
  assign n4559 = n4558 ^ x17 ;
  assign n4443 = x88 & n1060 ;
  assign n4560 = n4559 ^ n4443 ;
  assign n4442 = x90 & n1063 ;
  assign n4561 = n4560 ^ n4442 ;
  assign n4441 = n1064 & n2398 ;
  assign n4562 = n4561 ^ n4441 ;
  assign n4564 = n4563 ^ n4562 ;
  assign n4568 = n4567 ^ n4564 ;
  assign n4569 = n4568 ^ x14 ;
  assign n4440 = x91 & n884 ;
  assign n4570 = n4569 ^ n4440 ;
  assign n4439 = x93 & n789 ;
  assign n4571 = n4570 ^ n4439 ;
  assign n4438 = n790 & n2842 ;
  assign n4572 = n4571 ^ n4438 ;
  assign n4574 = n4573 ^ n4572 ;
  assign n4578 = n4577 ^ n4574 ;
  assign n4579 = n4578 ^ x11 ;
  assign n4437 = x94 & n650 ;
  assign n4580 = n4579 ^ n4437 ;
  assign n4436 = x96 & ~n578 ;
  assign n4581 = n4580 ^ n4436 ;
  assign n4435 = ~n579 & n3336 ;
  assign n4582 = n4581 ^ n4435 ;
  assign n4584 = n4583 ^ n4582 ;
  assign n4432 = n4376 ^ n4367 ;
  assign n4433 = ~n4373 & n4432 ;
  assign n4434 = n4433 ^ n4376 ;
  assign n4585 = n4584 ^ n4434 ;
  assign n4586 = n4585 ^ x8 ;
  assign n4431 = x97 & n456 ;
  assign n4587 = n4586 ^ n4431 ;
  assign n4430 = x99 & n384 ;
  assign n4588 = n4587 ^ n4430 ;
  assign n4429 = n385 & n3851 ;
  assign n4589 = n4588 ^ n4429 ;
  assign n4591 = n4590 ^ n4589 ;
  assign n4595 = n4594 ^ n4591 ;
  assign n4596 = n4595 ^ x5 ;
  assign n4428 = x100 & n238 ;
  assign n4597 = n4596 ^ n4428 ;
  assign n4427 = x102 & n234 ;
  assign n4598 = n4597 ^ n4427 ;
  assign n4425 = n3837 ^ x102 ;
  assign n4426 = n235 & n4425 ;
  assign n4599 = n4598 ^ n4426 ;
  assign n4601 = n4600 ^ n4599 ;
  assign n4422 = n4393 ^ n4384 ;
  assign n4423 = ~n4390 & n4422 ;
  assign n4424 = n4423 ^ n4393 ;
  assign n4602 = n4601 ^ n4424 ;
  assign n4407 = x104 & ~n4208 ;
  assign n4406 = ~x104 & ~n4207 ;
  assign n4408 = n4407 ^ n4406 ;
  assign n4410 = x105 ^ x1 ;
  assign n4409 = x105 ^ x2 ;
  assign n4411 = n4410 ^ n4409 ;
  assign n4412 = n4408 & n4411 ;
  assign n4413 = n4412 ^ n4410 ;
  assign n4603 = n4602 ^ n4413 ;
  assign n4417 = x2 & x103 ;
  assign n4418 = n4417 ^ x104 ;
  assign n4419 = ~x1 & n4418 ;
  assign n4414 = n4413 ^ n4210 ;
  assign n4420 = n4419 ^ n4414 ;
  assign n4421 = ~x0 & n4420 ;
  assign n4604 = n4603 ^ n4421 ;
  assign n4401 = n4399 ^ n4394 ;
  assign n4402 = ~n4396 & n4401 ;
  assign n4403 = n4402 ^ n4399 ;
  assign n4605 = n4604 ^ n4403 ;
  assign n4802 = n4602 ^ n4403 ;
  assign n4803 = n4604 & n4802 ;
  assign n4804 = n4803 ^ n4602 ;
  assign n4796 = n4595 ^ n4424 ;
  assign n4797 = n4601 & n4796 ;
  assign n4798 = n4797 ^ n4595 ;
  assign n4794 = x102 & n231 ;
  assign n4787 = x99 & n391 ;
  assign n4779 = n4578 ^ n4434 ;
  assign n4780 = n4584 & n4779 ;
  assign n4781 = n4780 ^ n4578 ;
  assign n4777 = x96 & n584 ;
  assign n4770 = x93 & n795 ;
  assign n4763 = x90 & n1068 ;
  assign n4755 = n4551 ^ n4446 ;
  assign n4756 = n4557 & n4755 ;
  assign n4757 = n4756 ^ n4551 ;
  assign n4753 = x87 & n1348 ;
  assign n4746 = x84 & n1673 ;
  assign n4739 = x81 & n2025 ;
  assign n4732 = x78 & n2435 ;
  assign n4724 = n4514 ^ n4461 ;
  assign n4725 = n4520 & n4724 ;
  assign n4726 = n4725 ^ n4514 ;
  assign n4722 = x75 & n2899 ;
  assign n4715 = x72 & n3395 ;
  assign n4708 = x69 & n3940 ;
  assign n4700 = ~n4474 & ~n4493 ;
  assign n4701 = x41 & n4700 ;
  assign n4695 = x65 & n4482 ;
  assign n4694 = x66 & n4475 ;
  assign n4696 = n4695 ^ n4694 ;
  assign n4691 = ~n155 & n4477 ;
  assign n4692 = n4691 ^ x67 ;
  assign n4693 = n4104 & n4692 ;
  assign n4697 = n4696 ^ n4693 ;
  assign n4698 = n4697 ^ x41 ;
  assign n4702 = n4701 ^ n4698 ;
  assign n4685 = x42 ^ x41 ;
  assign n4686 = x64 & n4685 ;
  assign n4703 = n4702 ^ n4686 ;
  assign n4704 = n4703 ^ x38 ;
  assign n4684 = x68 & n3932 ;
  assign n4705 = n4704 ^ n4684 ;
  assign n4683 = x70 & n3935 ;
  assign n4706 = n4705 ^ n4683 ;
  assign n4682 = ~n443 & n3936 ;
  assign n4707 = n4706 ^ n4682 ;
  assign n4709 = n4708 ^ n4707 ;
  assign n4679 = n4506 ^ n4502 ;
  assign n4680 = ~n4503 & n4679 ;
  assign n4681 = n4680 ^ n4506 ;
  assign n4710 = n4709 ^ n4681 ;
  assign n4711 = n4710 ^ x35 ;
  assign n4678 = x71 & n3387 ;
  assign n4712 = n4711 ^ n4678 ;
  assign n4677 = x73 & n3390 ;
  assign n4713 = n4712 ^ n4677 ;
  assign n4676 = n636 & n3391 ;
  assign n4714 = n4713 ^ n4676 ;
  assign n4716 = n4715 ^ n4714 ;
  assign n4673 = n4507 ^ n4467 ;
  assign n4674 = n4513 & n4673 ;
  assign n4675 = n4674 ^ n4507 ;
  assign n4717 = n4716 ^ n4675 ;
  assign n4718 = n4717 ^ x32 ;
  assign n4672 = x74 & n2890 ;
  assign n4719 = n4718 ^ n4672 ;
  assign n4671 = x76 & n2893 ;
  assign n4720 = n4719 ^ n4671 ;
  assign n4670 = ~n863 & n2894 ;
  assign n4721 = n4720 ^ n4670 ;
  assign n4723 = n4722 ^ n4721 ;
  assign n4727 = n4726 ^ n4723 ;
  assign n4728 = n4727 ^ x29 ;
  assign n4669 = x77 & n2593 ;
  assign n4729 = n4728 ^ n4669 ;
  assign n4668 = x79 & n2428 ;
  assign n4730 = n4729 ^ n4668 ;
  assign n4667 = n1123 & n2429 ;
  assign n4731 = n4730 ^ n4667 ;
  assign n4733 = n4732 ^ n4731 ;
  assign n4664 = n4530 ^ n4521 ;
  assign n4665 = ~n4527 & n4664 ;
  assign n4666 = n4665 ^ n4530 ;
  assign n4734 = n4733 ^ n4666 ;
  assign n4735 = n4734 ^ x26 ;
  assign n4663 = x80 & n2032 ;
  assign n4736 = n4735 ^ n4663 ;
  assign n4662 = x82 & n2028 ;
  assign n4737 = n4736 ^ n4662 ;
  assign n4661 = n1422 & n2029 ;
  assign n4738 = n4737 ^ n4661 ;
  assign n4740 = n4739 ^ n4738 ;
  assign n4658 = n4540 ^ n4531 ;
  assign n4659 = ~n4537 & n4658 ;
  assign n4660 = n4659 ^ n4540 ;
  assign n4741 = n4740 ^ n4660 ;
  assign n4742 = n4741 ^ x23 ;
  assign n4657 = x83 & n1665 ;
  assign n4743 = n4742 ^ n4657 ;
  assign n4656 = x85 & n1668 ;
  assign n4744 = n4743 ^ n4656 ;
  assign n4655 = n1669 & n1748 ;
  assign n4745 = n4744 ^ n4655 ;
  assign n4747 = n4746 ^ n4745 ;
  assign n4652 = n4550 ^ n4541 ;
  assign n4653 = ~n4547 & n4652 ;
  assign n4654 = n4653 ^ n4550 ;
  assign n4748 = n4747 ^ n4654 ;
  assign n4749 = n4748 ^ x20 ;
  assign n4651 = x86 & n1340 ;
  assign n4750 = n4749 ^ n4651 ;
  assign n4650 = x88 & n1343 ;
  assign n4751 = n4750 ^ n4650 ;
  assign n4649 = n1344 & n2131 ;
  assign n4752 = n4751 ^ n4649 ;
  assign n4754 = n4753 ^ n4752 ;
  assign n4758 = n4757 ^ n4754 ;
  assign n4759 = n4758 ^ x17 ;
  assign n4648 = x89 & n1060 ;
  assign n4760 = n4759 ^ n4648 ;
  assign n4647 = x91 & n1063 ;
  assign n4761 = n4760 ^ n4647 ;
  assign n4646 = n1064 & n2548 ;
  assign n4762 = n4761 ^ n4646 ;
  assign n4764 = n4763 ^ n4762 ;
  assign n4643 = n4567 ^ n4558 ;
  assign n4644 = ~n4564 & n4643 ;
  assign n4645 = n4644 ^ n4567 ;
  assign n4765 = n4764 ^ n4645 ;
  assign n4766 = n4765 ^ x14 ;
  assign n4642 = x92 & n884 ;
  assign n4767 = n4766 ^ n4642 ;
  assign n4641 = x94 & n789 ;
  assign n4768 = n4767 ^ n4641 ;
  assign n4640 = n790 & n3010 ;
  assign n4769 = n4768 ^ n4640 ;
  assign n4771 = n4770 ^ n4769 ;
  assign n4637 = n4577 ^ n4568 ;
  assign n4638 = ~n4574 & n4637 ;
  assign n4639 = n4638 ^ n4577 ;
  assign n4772 = n4771 ^ n4639 ;
  assign n4773 = n4772 ^ x11 ;
  assign n4636 = x95 & n650 ;
  assign n4774 = n4773 ^ n4636 ;
  assign n4635 = x97 & ~n578 ;
  assign n4775 = n4774 ^ n4635 ;
  assign n4634 = ~n579 & n3501 ;
  assign n4776 = n4775 ^ n4634 ;
  assign n4778 = n4777 ^ n4776 ;
  assign n4782 = n4781 ^ n4778 ;
  assign n4783 = n4782 ^ x8 ;
  assign n4633 = x98 & n456 ;
  assign n4784 = n4783 ^ n4633 ;
  assign n4632 = x100 & n384 ;
  assign n4785 = n4784 ^ n4632 ;
  assign n4631 = n385 & n4048 ;
  assign n4786 = n4785 ^ n4631 ;
  assign n4788 = n4787 ^ n4786 ;
  assign n4628 = n4594 ^ n4585 ;
  assign n4629 = ~n4591 & n4628 ;
  assign n4630 = n4629 ^ n4594 ;
  assign n4789 = n4788 ^ n4630 ;
  assign n4790 = n4789 ^ x5 ;
  assign n4627 = x101 & n238 ;
  assign n4791 = n4790 ^ n4627 ;
  assign n4626 = x103 & n234 ;
  assign n4792 = n4791 ^ n4626 ;
  assign n4624 = n4031 ^ x103 ;
  assign n4625 = n235 & ~n4624 ;
  assign n4793 = n4792 ^ n4625 ;
  assign n4795 = n4794 ^ n4793 ;
  assign n4799 = n4798 ^ n4795 ;
  assign n4609 = ~x105 & ~n4407 ;
  assign n4608 = x105 & ~n4406 ;
  assign n4610 = n4609 ^ n4608 ;
  assign n4612 = x106 ^ x1 ;
  assign n4611 = x106 ^ x2 ;
  assign n4613 = n4612 ^ n4611 ;
  assign n4614 = n4610 & n4613 ;
  assign n4615 = n4614 ^ n4612 ;
  assign n4800 = n4799 ^ n4615 ;
  assign n4619 = x2 & x104 ;
  assign n4620 = n4619 ^ x105 ;
  assign n4621 = ~x1 & n4620 ;
  assign n4616 = n4615 ^ n4409 ;
  assign n4622 = n4621 ^ n4616 ;
  assign n4623 = ~x0 & n4622 ;
  assign n4801 = n4800 ^ n4623 ;
  assign n4805 = n4804 ^ n4801 ;
  assign n5006 = x103 & n231 ;
  assign n4998 = n4782 ^ n4630 ;
  assign n4999 = n4788 & n4998 ;
  assign n5000 = n4999 ^ n4782 ;
  assign n4996 = x100 & n391 ;
  assign n4989 = x97 & n584 ;
  assign n4981 = n4765 ^ n4639 ;
  assign n4982 = n4771 & n4981 ;
  assign n4983 = n4982 ^ n4765 ;
  assign n4979 = x94 & n795 ;
  assign n4971 = n4758 ^ n4645 ;
  assign n4972 = n4764 & n4971 ;
  assign n4973 = n4972 ^ n4758 ;
  assign n4969 = x91 & n1068 ;
  assign n4962 = x88 & n1348 ;
  assign n4954 = n4741 ^ n4654 ;
  assign n4955 = n4747 & n4954 ;
  assign n4956 = n4955 ^ n4741 ;
  assign n4952 = x85 & n1673 ;
  assign n4944 = n4734 ^ n4660 ;
  assign n4945 = n4740 & n4944 ;
  assign n4946 = n4945 ^ n4734 ;
  assign n4942 = x82 & n2025 ;
  assign n4934 = n4727 ^ n4666 ;
  assign n4935 = n4733 & n4934 ;
  assign n4936 = n4935 ^ n4727 ;
  assign n4932 = x79 & n2435 ;
  assign n4925 = x76 & n2899 ;
  assign n4917 = n4710 ^ n4675 ;
  assign n4918 = n4716 & n4917 ;
  assign n4919 = n4918 ^ n4710 ;
  assign n4915 = x73 & n3395 ;
  assign n4907 = n4703 ^ n4681 ;
  assign n4908 = n4709 & n4907 ;
  assign n4909 = n4908 ^ n4703 ;
  assign n4905 = x70 & n3940 ;
  assign n4897 = ~n4686 & n4702 ;
  assign n4898 = n4698 & n4897 ;
  assign n4890 = x41 & x42 ;
  assign n4891 = n4890 ^ x43 ;
  assign n4892 = ~x64 & n4891 ;
  assign n4886 = x43 ^ x41 ;
  assign n4893 = n4892 ^ n4886 ;
  assign n4884 = x65 ^ x42 ;
  assign n4885 = n4685 & ~n4884 ;
  assign n4894 = n4893 ^ n4885 ;
  assign n4895 = n4894 ^ n4698 ;
  assign n4899 = n4898 ^ n4895 ;
  assign n4879 = x66 & n4482 ;
  assign n4878 = x68 & n4478 ;
  assign n4880 = n4879 ^ n4878 ;
  assign n4881 = n4880 ^ x41 ;
  assign n4877 = ~n351 & n4479 ;
  assign n4882 = n4881 ^ n4877 ;
  assign n4876 = x67 & n4475 ;
  assign n4883 = n4882 ^ n4876 ;
  assign n4900 = n4899 ^ n4883 ;
  assign n4901 = n4900 ^ x38 ;
  assign n4875 = x69 & n3932 ;
  assign n4902 = n4901 ^ n4875 ;
  assign n4874 = x71 & n3935 ;
  assign n4903 = n4902 ^ n4874 ;
  assign n4873 = ~n495 & n3936 ;
  assign n4904 = n4903 ^ n4873 ;
  assign n4906 = n4905 ^ n4904 ;
  assign n4910 = n4909 ^ n4906 ;
  assign n4911 = n4910 ^ x35 ;
  assign n4872 = x72 & n3387 ;
  assign n4912 = n4911 ^ n4872 ;
  assign n4871 = x74 & n3390 ;
  assign n4913 = n4912 ^ n4871 ;
  assign n4870 = n708 & n3391 ;
  assign n4914 = n4913 ^ n4870 ;
  assign n4916 = n4915 ^ n4914 ;
  assign n4920 = n4919 ^ n4916 ;
  assign n4921 = n4920 ^ x32 ;
  assign n4869 = x75 & n2890 ;
  assign n4922 = n4921 ^ n4869 ;
  assign n4868 = x77 & n2893 ;
  assign n4923 = n4922 ^ n4868 ;
  assign n4867 = ~n943 & n2894 ;
  assign n4924 = n4923 ^ n4867 ;
  assign n4926 = n4925 ^ n4924 ;
  assign n4864 = n4726 ^ n4717 ;
  assign n4865 = ~n4723 & n4864 ;
  assign n4866 = n4865 ^ n4726 ;
  assign n4927 = n4926 ^ n4866 ;
  assign n4928 = n4927 ^ x29 ;
  assign n4863 = x78 & n2593 ;
  assign n4929 = n4928 ^ n4863 ;
  assign n4862 = x80 & n2428 ;
  assign n4930 = n4929 ^ n4862 ;
  assign n4861 = n1217 & n2429 ;
  assign n4931 = n4930 ^ n4861 ;
  assign n4933 = n4932 ^ n4931 ;
  assign n4937 = n4936 ^ n4933 ;
  assign n4938 = n4937 ^ x26 ;
  assign n4860 = x81 & n2032 ;
  assign n4939 = n4938 ^ n4860 ;
  assign n4859 = x83 & n2028 ;
  assign n4940 = n4939 ^ n4859 ;
  assign n4858 = n1517 & n2029 ;
  assign n4941 = n4940 ^ n4858 ;
  assign n4943 = n4942 ^ n4941 ;
  assign n4947 = n4946 ^ n4943 ;
  assign n4948 = n4947 ^ x23 ;
  assign n4857 = x84 & n1665 ;
  assign n4949 = n4948 ^ n4857 ;
  assign n4856 = x86 & n1668 ;
  assign n4950 = n4949 ^ n4856 ;
  assign n4855 = n1669 & n1868 ;
  assign n4951 = n4950 ^ n4855 ;
  assign n4953 = n4952 ^ n4951 ;
  assign n4957 = n4956 ^ n4953 ;
  assign n4958 = n4957 ^ x20 ;
  assign n4854 = x87 & n1340 ;
  assign n4959 = n4958 ^ n4854 ;
  assign n4853 = x89 & n1343 ;
  assign n4960 = n4959 ^ n4853 ;
  assign n4852 = n1344 & n2255 ;
  assign n4961 = n4960 ^ n4852 ;
  assign n4963 = n4962 ^ n4961 ;
  assign n4849 = n4757 ^ n4748 ;
  assign n4850 = ~n4754 & n4849 ;
  assign n4851 = n4850 ^ n4757 ;
  assign n4964 = n4963 ^ n4851 ;
  assign n4965 = n4964 ^ x17 ;
  assign n4848 = x90 & n1060 ;
  assign n4966 = n4965 ^ n4848 ;
  assign n4847 = x92 & n1063 ;
  assign n4967 = n4966 ^ n4847 ;
  assign n4846 = n1064 & n2696 ;
  assign n4968 = n4967 ^ n4846 ;
  assign n4970 = n4969 ^ n4968 ;
  assign n4974 = n4973 ^ n4970 ;
  assign n4975 = n4974 ^ x14 ;
  assign n4845 = x93 & n884 ;
  assign n4976 = n4975 ^ n4845 ;
  assign n4844 = x95 & n789 ;
  assign n4977 = n4976 ^ n4844 ;
  assign n4843 = n790 & n3166 ;
  assign n4978 = n4977 ^ n4843 ;
  assign n4980 = n4979 ^ n4978 ;
  assign n4984 = n4983 ^ n4980 ;
  assign n4985 = n4984 ^ x11 ;
  assign n4842 = x96 & n650 ;
  assign n4986 = n4985 ^ n4842 ;
  assign n4841 = x98 & ~n578 ;
  assign n4987 = n4986 ^ n4841 ;
  assign n4840 = ~n579 & n3673 ;
  assign n4988 = n4987 ^ n4840 ;
  assign n4990 = n4989 ^ n4988 ;
  assign n4837 = n4781 ^ n4772 ;
  assign n4838 = ~n4778 & n4837 ;
  assign n4839 = n4838 ^ n4781 ;
  assign n4991 = n4990 ^ n4839 ;
  assign n4992 = n4991 ^ x8 ;
  assign n4836 = x99 & n456 ;
  assign n4993 = n4992 ^ n4836 ;
  assign n4835 = x101 & n384 ;
  assign n4994 = n4993 ^ n4835 ;
  assign n4834 = n385 & n4223 ;
  assign n4995 = n4994 ^ n4834 ;
  assign n4997 = n4996 ^ n4995 ;
  assign n5001 = n5000 ^ n4997 ;
  assign n5002 = n5001 ^ x5 ;
  assign n4833 = x102 & n238 ;
  assign n5003 = n5002 ^ n4833 ;
  assign n4832 = x104 & n234 ;
  assign n5004 = n5003 ^ n4832 ;
  assign n4830 = n4209 ^ x104 ;
  assign n4831 = n235 & ~n4830 ;
  assign n5005 = n5004 ^ n4831 ;
  assign n5007 = n5006 ^ n5005 ;
  assign n4827 = n4798 ^ n4789 ;
  assign n4828 = ~n4795 & n4827 ;
  assign n4829 = n4828 ^ n4798 ;
  assign n5008 = n5007 ^ n4829 ;
  assign n4812 = x106 & ~n4609 ;
  assign n4811 = ~x106 & ~n4608 ;
  assign n4813 = n4812 ^ n4811 ;
  assign n4815 = x107 ^ x1 ;
  assign n4814 = x107 ^ x2 ;
  assign n4816 = n4815 ^ n4814 ;
  assign n4817 = n4813 & n4816 ;
  assign n4818 = n4817 ^ n4815 ;
  assign n5009 = n5008 ^ n4818 ;
  assign n4822 = x2 & x105 ;
  assign n4823 = n4822 ^ x106 ;
  assign n4824 = ~x1 & n4823 ;
  assign n4819 = n4818 ^ n4611 ;
  assign n4825 = n4824 ^ n4819 ;
  assign n4826 = ~x0 & n4825 ;
  assign n5010 = n5009 ^ n4826 ;
  assign n4806 = n4804 ^ n4799 ;
  assign n4807 = ~n4801 & n4806 ;
  assign n4808 = n4807 ^ n4804 ;
  assign n5011 = n5010 ^ n4808 ;
  assign n5225 = n5008 ^ n4808 ;
  assign n5226 = n5010 & n5225 ;
  assign n5227 = n5226 ^ n5008 ;
  assign n5219 = n5001 ^ n4829 ;
  assign n5220 = n5007 & n5219 ;
  assign n5221 = n5220 ^ n5001 ;
  assign n5217 = x104 & n231 ;
  assign n5210 = x101 & n391 ;
  assign n5202 = n4984 ^ n4839 ;
  assign n5203 = n4990 & n5202 ;
  assign n5204 = n5203 ^ n4984 ;
  assign n5200 = x98 & n584 ;
  assign n5193 = x95 & n795 ;
  assign n5186 = x92 & n1068 ;
  assign n5178 = n4957 ^ n4851 ;
  assign n5179 = n4963 & n5178 ;
  assign n5180 = n5179 ^ n4957 ;
  assign n5176 = x89 & n1348 ;
  assign n5169 = x86 & n1673 ;
  assign n5162 = x83 & n2025 ;
  assign n5155 = x80 & n2435 ;
  assign n5147 = n4920 ^ n4866 ;
  assign n5148 = n4926 & n5147 ;
  assign n5149 = n5148 ^ n4920 ;
  assign n5145 = x77 & n2899 ;
  assign n5137 = x71 & n3940 ;
  assign n5130 = x68 & n4475 ;
  assign n4888 = x43 ^ x42 ;
  assign n5121 = ~n4685 & n4888 ;
  assign n5122 = x65 & n5121 ;
  assign n5110 = x44 ^ x43 ;
  assign n5116 = n4685 & ~n5110 ;
  assign n5117 = n5116 ^ n4685 ;
  assign n5118 = ~n152 & n5117 ;
  assign n5115 = x66 & n4685 ;
  assign n5119 = n5118 ^ n5115 ;
  assign n5120 = n5119 ^ x44 ;
  assign n5123 = n5122 ^ n5120 ;
  assign n5111 = x44 ^ x42 ;
  assign n5112 = ~n4685 & n5111 ;
  assign n5113 = n5110 & n5112 ;
  assign n5114 = x64 & n5113 ;
  assign n5124 = n5123 ^ n5114 ;
  assign n5108 = ~n4686 & ~n4894 ;
  assign n5109 = x44 & n5108 ;
  assign n5125 = n5124 ^ n5109 ;
  assign n5126 = n5125 ^ x41 ;
  assign n5107 = x67 & n4482 ;
  assign n5127 = n5126 ^ n5107 ;
  assign n5106 = x69 & n4478 ;
  assign n5128 = n5127 ^ n5106 ;
  assign n5105 = ~n376 & n4479 ;
  assign n5129 = n5128 ^ n5105 ;
  assign n5131 = n5130 ^ n5129 ;
  assign n5102 = n4894 ^ n4883 ;
  assign n5103 = n4899 & n5102 ;
  assign n5104 = n5103 ^ n4894 ;
  assign n5132 = n5131 ^ n5104 ;
  assign n5133 = n5132 ^ x38 ;
  assign n5101 = x70 & n3932 ;
  assign n5134 = n5133 ^ n5101 ;
  assign n5100 = x72 & n3935 ;
  assign n5135 = n5134 ^ n5100 ;
  assign n5099 = n565 & n3936 ;
  assign n5136 = n5135 ^ n5099 ;
  assign n5138 = n5137 ^ n5136 ;
  assign n5096 = n4909 ^ n4900 ;
  assign n5097 = ~n4906 & n5096 ;
  assign n5098 = n5097 ^ n4909 ;
  assign n5139 = n5138 ^ n5098 ;
  assign n5086 = x73 & n3387 ;
  assign n5085 = x75 & n3390 ;
  assign n5087 = n5086 ^ n5085 ;
  assign n5088 = n5087 ^ x35 ;
  assign n5084 = ~n778 & n3391 ;
  assign n5089 = n5088 ^ n5084 ;
  assign n5083 = x74 & n3395 ;
  assign n5090 = n5089 ^ n5083 ;
  assign n5091 = n5090 ^ n4919 ;
  assign n5092 = n5091 ^ n4910 ;
  assign n5093 = n5092 ^ n5090 ;
  assign n5094 = ~n4916 & n5093 ;
  assign n5095 = n5094 ^ n5091 ;
  assign n5140 = n5139 ^ n5095 ;
  assign n5141 = n5140 ^ x32 ;
  assign n5082 = x76 & n2890 ;
  assign n5142 = n5141 ^ n5082 ;
  assign n5081 = x78 & n2893 ;
  assign n5143 = n5142 ^ n5081 ;
  assign n5080 = ~n1036 & n2894 ;
  assign n5144 = n5143 ^ n5080 ;
  assign n5146 = n5145 ^ n5144 ;
  assign n5150 = n5149 ^ n5146 ;
  assign n5151 = n5150 ^ x29 ;
  assign n5079 = x79 & n2593 ;
  assign n5152 = n5151 ^ n5079 ;
  assign n5078 = x81 & n2428 ;
  assign n5153 = n5152 ^ n5078 ;
  assign n5077 = n1310 & n2429 ;
  assign n5154 = n5153 ^ n5077 ;
  assign n5156 = n5155 ^ n5154 ;
  assign n5074 = n4936 ^ n4927 ;
  assign n5075 = ~n4933 & n5074 ;
  assign n5076 = n5075 ^ n4936 ;
  assign n5157 = n5156 ^ n5076 ;
  assign n5158 = n5157 ^ x26 ;
  assign n5073 = x82 & n2032 ;
  assign n5159 = n5158 ^ n5073 ;
  assign n5072 = x84 & n2028 ;
  assign n5160 = n5159 ^ n5072 ;
  assign n5071 = n1635 & n2029 ;
  assign n5161 = n5160 ^ n5071 ;
  assign n5163 = n5162 ^ n5161 ;
  assign n5068 = n4946 ^ n4937 ;
  assign n5069 = ~n4943 & n5068 ;
  assign n5070 = n5069 ^ n4946 ;
  assign n5164 = n5163 ^ n5070 ;
  assign n5165 = n5164 ^ x23 ;
  assign n5067 = x85 & n1665 ;
  assign n5166 = n5165 ^ n5067 ;
  assign n5066 = x87 & n1668 ;
  assign n5167 = n5166 ^ n5066 ;
  assign n5065 = n1669 & n1987 ;
  assign n5168 = n5167 ^ n5065 ;
  assign n5170 = n5169 ^ n5168 ;
  assign n5062 = n4956 ^ n4947 ;
  assign n5063 = ~n4953 & n5062 ;
  assign n5064 = n5063 ^ n4956 ;
  assign n5171 = n5170 ^ n5064 ;
  assign n5172 = n5171 ^ x20 ;
  assign n5061 = x88 & n1340 ;
  assign n5173 = n5172 ^ n5061 ;
  assign n5060 = x90 & n1343 ;
  assign n5174 = n5173 ^ n5060 ;
  assign n5059 = n1344 & n2398 ;
  assign n5175 = n5174 ^ n5059 ;
  assign n5177 = n5176 ^ n5175 ;
  assign n5181 = n5180 ^ n5177 ;
  assign n5182 = n5181 ^ x17 ;
  assign n5058 = x91 & n1060 ;
  assign n5183 = n5182 ^ n5058 ;
  assign n5057 = x93 & n1063 ;
  assign n5184 = n5183 ^ n5057 ;
  assign n5056 = n1064 & n2842 ;
  assign n5185 = n5184 ^ n5056 ;
  assign n5187 = n5186 ^ n5185 ;
  assign n5053 = n4973 ^ n4964 ;
  assign n5054 = ~n4970 & n5053 ;
  assign n5055 = n5054 ^ n4973 ;
  assign n5188 = n5187 ^ n5055 ;
  assign n5189 = n5188 ^ x14 ;
  assign n5052 = x94 & n884 ;
  assign n5190 = n5189 ^ n5052 ;
  assign n5051 = x96 & n789 ;
  assign n5191 = n5190 ^ n5051 ;
  assign n5050 = n790 & n3336 ;
  assign n5192 = n5191 ^ n5050 ;
  assign n5194 = n5193 ^ n5192 ;
  assign n5047 = n4983 ^ n4974 ;
  assign n5048 = ~n4980 & n5047 ;
  assign n5049 = n5048 ^ n4983 ;
  assign n5195 = n5194 ^ n5049 ;
  assign n5196 = n5195 ^ x11 ;
  assign n5046 = x97 & n650 ;
  assign n5197 = n5196 ^ n5046 ;
  assign n5045 = x99 & ~n578 ;
  assign n5198 = n5197 ^ n5045 ;
  assign n5044 = ~n579 & n3851 ;
  assign n5199 = n5198 ^ n5044 ;
  assign n5201 = n5200 ^ n5199 ;
  assign n5205 = n5204 ^ n5201 ;
  assign n5206 = n5205 ^ x8 ;
  assign n5043 = x100 & n456 ;
  assign n5207 = n5206 ^ n5043 ;
  assign n5042 = x102 & n384 ;
  assign n5208 = n5207 ^ n5042 ;
  assign n5041 = n385 & n4425 ;
  assign n5209 = n5208 ^ n5041 ;
  assign n5211 = n5210 ^ n5209 ;
  assign n5038 = n5000 ^ n4991 ;
  assign n5039 = ~n4997 & n5038 ;
  assign n5040 = n5039 ^ n5000 ;
  assign n5212 = n5211 ^ n5040 ;
  assign n5213 = n5212 ^ x5 ;
  assign n5037 = x103 & n238 ;
  assign n5214 = n5213 ^ n5037 ;
  assign n5036 = x105 & n234 ;
  assign n5215 = n5214 ^ n5036 ;
  assign n5034 = n4408 ^ x105 ;
  assign n5035 = n235 & ~n5034 ;
  assign n5216 = n5215 ^ n5035 ;
  assign n5218 = n5217 ^ n5216 ;
  assign n5222 = n5221 ^ n5218 ;
  assign n5012 = x107 ^ x106 ;
  assign n5018 = x107 & n4610 ;
  assign n5019 = n5018 ^ n4609 ;
  assign n5020 = n5012 & ~n5019 ;
  assign n5022 = x108 ^ x1 ;
  assign n5021 = x108 ^ x2 ;
  assign n5023 = n5022 ^ n5021 ;
  assign n5024 = ~n5020 & n5023 ;
  assign n5025 = n5024 ^ n5022 ;
  assign n5223 = n5222 ^ n5025 ;
  assign n5029 = x2 & x106 ;
  assign n5030 = n5029 ^ x107 ;
  assign n5031 = ~x1 & n5030 ;
  assign n5026 = n5025 ^ n4814 ;
  assign n5032 = n5031 ^ n5026 ;
  assign n5033 = ~x0 & n5032 ;
  assign n5224 = n5223 ^ n5033 ;
  assign n5228 = n5227 ^ n5224 ;
  assign n5435 = x105 & n231 ;
  assign n5427 = n5205 ^ n5040 ;
  assign n5428 = n5211 & n5427 ;
  assign n5429 = n5428 ^ n5205 ;
  assign n5425 = x102 & n391 ;
  assign n5418 = x99 & n584 ;
  assign n5410 = n5188 ^ n5049 ;
  assign n5411 = n5194 & n5410 ;
  assign n5412 = n5411 ^ n5188 ;
  assign n5408 = x96 & n795 ;
  assign n5400 = n5181 ^ n5055 ;
  assign n5401 = n5187 & n5400 ;
  assign n5402 = n5401 ^ n5181 ;
  assign n5398 = x93 & n1068 ;
  assign n5391 = x90 & n1348 ;
  assign n5383 = n5164 ^ n5064 ;
  assign n5384 = n5170 & n5383 ;
  assign n5385 = n5384 ^ n5164 ;
  assign n5381 = x87 & n1673 ;
  assign n5373 = n5157 ^ n5070 ;
  assign n5374 = n5163 & n5373 ;
  assign n5375 = n5374 ^ n5157 ;
  assign n5371 = x84 & n2025 ;
  assign n5363 = n5150 ^ n5076 ;
  assign n5364 = n5156 & n5363 ;
  assign n5365 = n5364 ^ n5150 ;
  assign n5361 = x81 & n2435 ;
  assign n5354 = x78 & n2899 ;
  assign n5347 = x75 & n3395 ;
  assign n5339 = x69 & n4475 ;
  assign n5328 = x65 & n5113 ;
  assign n5327 = x67 & n5116 ;
  assign n5329 = n5328 ^ n5327 ;
  assign n5330 = n5329 ^ x44 ;
  assign n5326 = ~n295 & n5117 ;
  assign n5331 = n5330 ^ n5326 ;
  assign n5325 = x66 & n5121 ;
  assign n5332 = n5331 ^ n5325 ;
  assign n5323 = x45 ^ x44 ;
  assign n5324 = x64 & n5323 ;
  assign n5333 = n5332 ^ n5324 ;
  assign n5322 = n5109 & n5124 ;
  assign n5334 = n5333 ^ n5322 ;
  assign n5335 = n5334 ^ x41 ;
  assign n5321 = x68 & n4482 ;
  assign n5336 = n5335 ^ n5321 ;
  assign n5320 = x70 & n4478 ;
  assign n5337 = n5336 ^ n5320 ;
  assign n5319 = ~n443 & n4479 ;
  assign n5338 = n5337 ^ n5319 ;
  assign n5340 = n5339 ^ n5338 ;
  assign n5316 = n5125 ^ n5104 ;
  assign n5317 = n5131 & n5316 ;
  assign n5318 = n5317 ^ n5125 ;
  assign n5341 = n5340 ^ n5318 ;
  assign n5313 = n5132 ^ n5098 ;
  assign n5314 = n5138 & n5313 ;
  assign n5306 = x71 & n3932 ;
  assign n5305 = x73 & n3935 ;
  assign n5307 = n5306 ^ n5305 ;
  assign n5308 = n5307 ^ x38 ;
  assign n5304 = n636 & n3936 ;
  assign n5309 = n5308 ^ n5304 ;
  assign n5303 = x72 & n3940 ;
  assign n5310 = n5309 ^ n5303 ;
  assign n5311 = n5310 ^ n5132 ;
  assign n5315 = n5314 ^ n5311 ;
  assign n5342 = n5341 ^ n5315 ;
  assign n5343 = n5342 ^ x35 ;
  assign n5302 = x74 & n3387 ;
  assign n5344 = n5343 ^ n5302 ;
  assign n5301 = x76 & n3390 ;
  assign n5345 = n5344 ^ n5301 ;
  assign n5300 = ~n863 & n3391 ;
  assign n5346 = n5345 ^ n5300 ;
  assign n5348 = n5347 ^ n5346 ;
  assign n5297 = n5139 ^ n5090 ;
  assign n5298 = n5095 & n5297 ;
  assign n5299 = n5298 ^ n5090 ;
  assign n5349 = n5348 ^ n5299 ;
  assign n5350 = n5349 ^ x32 ;
  assign n5296 = x77 & n2890 ;
  assign n5351 = n5350 ^ n5296 ;
  assign n5295 = x79 & n2893 ;
  assign n5352 = n5351 ^ n5295 ;
  assign n5294 = n1123 & n2894 ;
  assign n5353 = n5352 ^ n5294 ;
  assign n5355 = n5354 ^ n5353 ;
  assign n5291 = n5149 ^ n5140 ;
  assign n5292 = ~n5146 & n5291 ;
  assign n5293 = n5292 ^ n5149 ;
  assign n5356 = n5355 ^ n5293 ;
  assign n5357 = n5356 ^ x29 ;
  assign n5290 = x80 & n2593 ;
  assign n5358 = n5357 ^ n5290 ;
  assign n5289 = x82 & n2428 ;
  assign n5359 = n5358 ^ n5289 ;
  assign n5288 = n1422 & n2429 ;
  assign n5360 = n5359 ^ n5288 ;
  assign n5362 = n5361 ^ n5360 ;
  assign n5366 = n5365 ^ n5362 ;
  assign n5367 = n5366 ^ x26 ;
  assign n5287 = x83 & n2032 ;
  assign n5368 = n5367 ^ n5287 ;
  assign n5286 = x85 & n2028 ;
  assign n5369 = n5368 ^ n5286 ;
  assign n5285 = n1748 & n2029 ;
  assign n5370 = n5369 ^ n5285 ;
  assign n5372 = n5371 ^ n5370 ;
  assign n5376 = n5375 ^ n5372 ;
  assign n5377 = n5376 ^ x23 ;
  assign n5284 = x86 & n1665 ;
  assign n5378 = n5377 ^ n5284 ;
  assign n5283 = x88 & n1668 ;
  assign n5379 = n5378 ^ n5283 ;
  assign n5282 = n1669 & n2131 ;
  assign n5380 = n5379 ^ n5282 ;
  assign n5382 = n5381 ^ n5380 ;
  assign n5386 = n5385 ^ n5382 ;
  assign n5387 = n5386 ^ x20 ;
  assign n5281 = x89 & n1340 ;
  assign n5388 = n5387 ^ n5281 ;
  assign n5280 = x91 & n1343 ;
  assign n5389 = n5388 ^ n5280 ;
  assign n5279 = n1344 & n2548 ;
  assign n5390 = n5389 ^ n5279 ;
  assign n5392 = n5391 ^ n5390 ;
  assign n5276 = n5180 ^ n5171 ;
  assign n5277 = ~n5177 & n5276 ;
  assign n5278 = n5277 ^ n5180 ;
  assign n5393 = n5392 ^ n5278 ;
  assign n5394 = n5393 ^ x17 ;
  assign n5275 = x92 & n1060 ;
  assign n5395 = n5394 ^ n5275 ;
  assign n5274 = x94 & n1063 ;
  assign n5396 = n5395 ^ n5274 ;
  assign n5273 = n1064 & n3010 ;
  assign n5397 = n5396 ^ n5273 ;
  assign n5399 = n5398 ^ n5397 ;
  assign n5403 = n5402 ^ n5399 ;
  assign n5404 = n5403 ^ x14 ;
  assign n5272 = x95 & n884 ;
  assign n5405 = n5404 ^ n5272 ;
  assign n5271 = x97 & n789 ;
  assign n5406 = n5405 ^ n5271 ;
  assign n5270 = n790 & n3501 ;
  assign n5407 = n5406 ^ n5270 ;
  assign n5409 = n5408 ^ n5407 ;
  assign n5413 = n5412 ^ n5409 ;
  assign n5414 = n5413 ^ x11 ;
  assign n5269 = x98 & n650 ;
  assign n5415 = n5414 ^ n5269 ;
  assign n5268 = x100 & ~n578 ;
  assign n5416 = n5415 ^ n5268 ;
  assign n5267 = ~n579 & n4048 ;
  assign n5417 = n5416 ^ n5267 ;
  assign n5419 = n5418 ^ n5417 ;
  assign n5264 = n5204 ^ n5195 ;
  assign n5265 = ~n5201 & n5264 ;
  assign n5266 = n5265 ^ n5204 ;
  assign n5420 = n5419 ^ n5266 ;
  assign n5421 = n5420 ^ x8 ;
  assign n5263 = x101 & n456 ;
  assign n5422 = n5421 ^ n5263 ;
  assign n5262 = x103 & n384 ;
  assign n5423 = n5422 ^ n5262 ;
  assign n5261 = n385 & ~n4624 ;
  assign n5424 = n5423 ^ n5261 ;
  assign n5426 = n5425 ^ n5424 ;
  assign n5430 = n5429 ^ n5426 ;
  assign n5431 = n5430 ^ x5 ;
  assign n5260 = x104 & n238 ;
  assign n5432 = n5431 ^ n5260 ;
  assign n5259 = x106 & n234 ;
  assign n5433 = n5432 ^ n5259 ;
  assign n5257 = n4610 ^ x106 ;
  assign n5258 = n235 & ~n5257 ;
  assign n5434 = n5433 ^ n5258 ;
  assign n5436 = n5435 ^ n5434 ;
  assign n5254 = n5221 ^ n5212 ;
  assign n5255 = ~n5218 & n5254 ;
  assign n5256 = n5255 ^ n5221 ;
  assign n5437 = n5436 ^ n5256 ;
  assign n5232 = x108 ^ x107 ;
  assign n5238 = x108 & n4813 ;
  assign n5239 = n5238 ^ n4811 ;
  assign n5240 = n5232 & ~n5239 ;
  assign n5242 = x109 ^ x1 ;
  assign n5241 = x109 ^ x2 ;
  assign n5243 = n5242 ^ n5241 ;
  assign n5244 = ~n5240 & n5243 ;
  assign n5245 = n5244 ^ n5242 ;
  assign n5438 = n5437 ^ n5245 ;
  assign n5249 = x2 & x107 ;
  assign n5250 = n5249 ^ x108 ;
  assign n5251 = ~n259 & n5250 ;
  assign n5246 = n5245 ^ n5021 ;
  assign n5252 = n5251 ^ n5246 ;
  assign n5253 = ~x0 & n5252 ;
  assign n5439 = n5438 ^ n5253 ;
  assign n5229 = n5227 ^ n5222 ;
  assign n5230 = ~n5224 & n5229 ;
  assign n5231 = n5230 ^ n5227 ;
  assign n5440 = n5439 ^ n5231 ;
  assign n5657 = n5437 ^ n5231 ;
  assign n5658 = n5439 & n5657 ;
  assign n5659 = n5658 ^ n5437 ;
  assign n5651 = n5430 ^ n5256 ;
  assign n5652 = n5436 & n5651 ;
  assign n5653 = n5652 ^ n5430 ;
  assign n5649 = x106 & n231 ;
  assign n5642 = x103 & n391 ;
  assign n5634 = n5413 ^ n5266 ;
  assign n5635 = n5419 & n5634 ;
  assign n5636 = n5635 ^ n5413 ;
  assign n5632 = x100 & n584 ;
  assign n5625 = x97 & n795 ;
  assign n5618 = x94 & n1068 ;
  assign n5610 = n5386 ^ n5278 ;
  assign n5611 = n5392 & n5610 ;
  assign n5612 = n5611 ^ n5386 ;
  assign n5608 = x91 & n1348 ;
  assign n5601 = x88 & n1673 ;
  assign n5594 = x85 & n2025 ;
  assign n5587 = x82 & n2435 ;
  assign n5579 = n5349 ^ n5293 ;
  assign n5580 = n5355 & n5579 ;
  assign n5581 = n5580 ^ n5349 ;
  assign n5577 = x79 & n2899 ;
  assign n5569 = x73 & n3940 ;
  assign n5561 = x67 & n5121 ;
  assign n5559 = ~n351 & n5117 ;
  assign n5555 = x66 & n5113 ;
  assign n5554 = x68 & n5116 ;
  assign n5556 = n5555 ^ n5554 ;
  assign n5557 = n5556 ^ x44 ;
  assign n5549 = ~x44 & ~x45 ;
  assign n5550 = n5549 ^ n5323 ;
  assign n5551 = n5550 ^ x46 ;
  assign n5552 = ~x64 & ~n5551 ;
  assign n5543 = x65 ^ x45 ;
  assign n5546 = x65 ^ x44 ;
  assign n5547 = ~n5543 & n5546 ;
  assign n5544 = x46 ^ x44 ;
  assign n5548 = n5547 ^ n5544 ;
  assign n5553 = n5552 ^ n5548 ;
  assign n5558 = n5557 ^ n5553 ;
  assign n5560 = n5559 ^ n5558 ;
  assign n5562 = n5561 ^ n5560 ;
  assign n5540 = ~n5324 & n5332 ;
  assign n5541 = ~n5322 & n5540 ;
  assign n5542 = n5541 ^ n5332 ;
  assign n5563 = n5562 ^ n5542 ;
  assign n5537 = n5334 ^ n5318 ;
  assign n5538 = n5340 & n5537 ;
  assign n5530 = x69 & n4482 ;
  assign n5529 = x71 & n4478 ;
  assign n5531 = n5530 ^ n5529 ;
  assign n5532 = n5531 ^ x41 ;
  assign n5528 = ~n495 & n4479 ;
  assign n5533 = n5532 ^ n5528 ;
  assign n5527 = x70 & n4475 ;
  assign n5534 = n5533 ^ n5527 ;
  assign n5535 = n5534 ^ n5334 ;
  assign n5539 = n5538 ^ n5535 ;
  assign n5564 = n5563 ^ n5539 ;
  assign n5565 = n5564 ^ x38 ;
  assign n5526 = x72 & n3932 ;
  assign n5566 = n5565 ^ n5526 ;
  assign n5525 = x74 & n3935 ;
  assign n5567 = n5566 ^ n5525 ;
  assign n5524 = n708 & n3936 ;
  assign n5568 = n5567 ^ n5524 ;
  assign n5570 = n5569 ^ n5568 ;
  assign n5521 = n5341 ^ n5310 ;
  assign n5522 = n5315 & n5521 ;
  assign n5523 = n5522 ^ n5310 ;
  assign n5571 = n5570 ^ n5523 ;
  assign n5511 = x75 & n3387 ;
  assign n5510 = x77 & n3390 ;
  assign n5512 = n5511 ^ n5510 ;
  assign n5513 = n5512 ^ x35 ;
  assign n5509 = ~n943 & n3391 ;
  assign n5514 = n5513 ^ n5509 ;
  assign n5508 = x76 & n3395 ;
  assign n5515 = n5514 ^ n5508 ;
  assign n5516 = n5515 ^ n5342 ;
  assign n5517 = n5516 ^ n5299 ;
  assign n5518 = n5517 ^ n5515 ;
  assign n5519 = n5348 & n5518 ;
  assign n5520 = n5519 ^ n5516 ;
  assign n5572 = n5571 ^ n5520 ;
  assign n5573 = n5572 ^ x32 ;
  assign n5507 = x78 & n2890 ;
  assign n5574 = n5573 ^ n5507 ;
  assign n5506 = x80 & n2893 ;
  assign n5575 = n5574 ^ n5506 ;
  assign n5505 = n1217 & n2894 ;
  assign n5576 = n5575 ^ n5505 ;
  assign n5578 = n5577 ^ n5576 ;
  assign n5582 = n5581 ^ n5578 ;
  assign n5583 = n5582 ^ x29 ;
  assign n5504 = x81 & n2593 ;
  assign n5584 = n5583 ^ n5504 ;
  assign n5503 = x83 & n2428 ;
  assign n5585 = n5584 ^ n5503 ;
  assign n5502 = n1517 & n2429 ;
  assign n5586 = n5585 ^ n5502 ;
  assign n5588 = n5587 ^ n5586 ;
  assign n5499 = n5365 ^ n5356 ;
  assign n5500 = ~n5362 & n5499 ;
  assign n5501 = n5500 ^ n5365 ;
  assign n5589 = n5588 ^ n5501 ;
  assign n5590 = n5589 ^ x26 ;
  assign n5498 = x84 & n2032 ;
  assign n5591 = n5590 ^ n5498 ;
  assign n5497 = x86 & n2028 ;
  assign n5592 = n5591 ^ n5497 ;
  assign n5496 = n1868 & n2029 ;
  assign n5593 = n5592 ^ n5496 ;
  assign n5595 = n5594 ^ n5593 ;
  assign n5493 = n5375 ^ n5366 ;
  assign n5494 = ~n5372 & n5493 ;
  assign n5495 = n5494 ^ n5375 ;
  assign n5596 = n5595 ^ n5495 ;
  assign n5597 = n5596 ^ x23 ;
  assign n5492 = x87 & n1665 ;
  assign n5598 = n5597 ^ n5492 ;
  assign n5491 = x89 & n1668 ;
  assign n5599 = n5598 ^ n5491 ;
  assign n5490 = n1669 & n2255 ;
  assign n5600 = n5599 ^ n5490 ;
  assign n5602 = n5601 ^ n5600 ;
  assign n5487 = n5385 ^ n5376 ;
  assign n5488 = ~n5382 & n5487 ;
  assign n5489 = n5488 ^ n5385 ;
  assign n5603 = n5602 ^ n5489 ;
  assign n5604 = n5603 ^ x20 ;
  assign n5486 = x90 & n1340 ;
  assign n5605 = n5604 ^ n5486 ;
  assign n5485 = x92 & n1343 ;
  assign n5606 = n5605 ^ n5485 ;
  assign n5484 = n1344 & n2696 ;
  assign n5607 = n5606 ^ n5484 ;
  assign n5609 = n5608 ^ n5607 ;
  assign n5613 = n5612 ^ n5609 ;
  assign n5614 = n5613 ^ x17 ;
  assign n5483 = x93 & n1060 ;
  assign n5615 = n5614 ^ n5483 ;
  assign n5482 = x95 & n1063 ;
  assign n5616 = n5615 ^ n5482 ;
  assign n5481 = n1064 & n3166 ;
  assign n5617 = n5616 ^ n5481 ;
  assign n5619 = n5618 ^ n5617 ;
  assign n5478 = n5402 ^ n5393 ;
  assign n5479 = ~n5399 & n5478 ;
  assign n5480 = n5479 ^ n5402 ;
  assign n5620 = n5619 ^ n5480 ;
  assign n5621 = n5620 ^ x14 ;
  assign n5477 = x96 & n884 ;
  assign n5622 = n5621 ^ n5477 ;
  assign n5476 = x98 & n789 ;
  assign n5623 = n5622 ^ n5476 ;
  assign n5475 = n790 & n3673 ;
  assign n5624 = n5623 ^ n5475 ;
  assign n5626 = n5625 ^ n5624 ;
  assign n5472 = n5412 ^ n5403 ;
  assign n5473 = ~n5409 & n5472 ;
  assign n5474 = n5473 ^ n5412 ;
  assign n5627 = n5626 ^ n5474 ;
  assign n5628 = n5627 ^ x11 ;
  assign n5471 = x99 & n650 ;
  assign n5629 = n5628 ^ n5471 ;
  assign n5470 = x101 & ~n578 ;
  assign n5630 = n5629 ^ n5470 ;
  assign n5469 = ~n579 & n4223 ;
  assign n5631 = n5630 ^ n5469 ;
  assign n5633 = n5632 ^ n5631 ;
  assign n5637 = n5636 ^ n5633 ;
  assign n5638 = n5637 ^ x8 ;
  assign n5468 = x102 & n456 ;
  assign n5639 = n5638 ^ n5468 ;
  assign n5467 = x104 & n384 ;
  assign n5640 = n5639 ^ n5467 ;
  assign n5466 = n385 & ~n4830 ;
  assign n5641 = n5640 ^ n5466 ;
  assign n5643 = n5642 ^ n5641 ;
  assign n5463 = n5429 ^ n5420 ;
  assign n5464 = ~n5426 & n5463 ;
  assign n5465 = n5464 ^ n5429 ;
  assign n5644 = n5643 ^ n5465 ;
  assign n5645 = n5644 ^ x5 ;
  assign n5462 = x105 & n238 ;
  assign n5646 = n5645 ^ n5462 ;
  assign n5461 = x107 & n234 ;
  assign n5647 = n5646 ^ n5461 ;
  assign n5459 = n4813 ^ x107 ;
  assign n5460 = n235 & ~n5459 ;
  assign n5648 = n5647 ^ n5460 ;
  assign n5650 = n5649 ^ n5648 ;
  assign n5654 = n5653 ^ n5650 ;
  assign n5441 = x109 ^ x108 ;
  assign n5443 = n5240 & n5441 ;
  assign n5444 = n5443 ^ x108 ;
  assign n5445 = n5444 ^ x109 ;
  assign n5447 = x110 ^ x1 ;
  assign n5446 = x110 ^ x2 ;
  assign n5448 = n5447 ^ n5446 ;
  assign n5449 = ~n5445 & n5448 ;
  assign n5450 = n5449 ^ n5447 ;
  assign n5655 = n5654 ^ n5450 ;
  assign n5454 = x2 & x108 ;
  assign n5455 = n5454 ^ x109 ;
  assign n5456 = ~n259 & n5455 ;
  assign n5451 = n5450 ^ n5241 ;
  assign n5457 = n5456 ^ n5451 ;
  assign n5458 = ~x0 & n5457 ;
  assign n5656 = n5655 ^ n5458 ;
  assign n5660 = n5659 ^ n5656 ;
  assign n5888 = x107 & n231 ;
  assign n5880 = n5637 ^ n5465 ;
  assign n5881 = n5643 & n5880 ;
  assign n5882 = n5881 ^ n5637 ;
  assign n5878 = x104 & n391 ;
  assign n5871 = x101 & n584 ;
  assign n5863 = n5620 ^ n5474 ;
  assign n5864 = n5626 & n5863 ;
  assign n5865 = n5864 ^ n5620 ;
  assign n5861 = x98 & n795 ;
  assign n5853 = n5613 ^ n5480 ;
  assign n5854 = n5619 & n5853 ;
  assign n5855 = n5854 ^ n5613 ;
  assign n5851 = x95 & n1068 ;
  assign n5844 = x92 & n1348 ;
  assign n5836 = n5596 ^ n5489 ;
  assign n5837 = n5602 & n5836 ;
  assign n5838 = n5837 ^ n5596 ;
  assign n5834 = x89 & n1673 ;
  assign n5826 = n5589 ^ n5495 ;
  assign n5827 = n5595 & n5826 ;
  assign n5828 = n5827 ^ n5589 ;
  assign n5824 = x86 & n2025 ;
  assign n5816 = n5582 ^ n5501 ;
  assign n5817 = n5588 & n5816 ;
  assign n5818 = n5817 ^ n5582 ;
  assign n5814 = x83 & n2435 ;
  assign n5807 = x80 & n2899 ;
  assign n5800 = x77 & n3395 ;
  assign n5790 = x73 & n3932 ;
  assign n5789 = x75 & n3935 ;
  assign n5791 = n5790 ^ n5789 ;
  assign n5792 = n5791 ^ x38 ;
  assign n5788 = ~n778 & n3936 ;
  assign n5793 = n5792 ^ n5788 ;
  assign n5787 = x74 & n3940 ;
  assign n5794 = n5793 ^ n5787 ;
  assign n5780 = x70 & n4482 ;
  assign n5779 = x72 & n4478 ;
  assign n5781 = n5780 ^ n5779 ;
  assign n5782 = n5781 ^ x41 ;
  assign n5778 = n565 & n4479 ;
  assign n5783 = n5782 ^ n5778 ;
  assign n5777 = x71 & n4475 ;
  assign n5784 = n5783 ^ n5777 ;
  assign n5766 = n5553 ^ n5542 ;
  assign n5767 = n5562 & n5766 ;
  assign n5768 = n5767 ^ n5553 ;
  assign n5758 = ~x46 & x47 ;
  assign n5759 = x64 & n5549 ;
  assign n5760 = n5758 & n5759 ;
  assign n5754 = x46 ^ x45 ;
  assign n5755 = ~n5323 & n5754 ;
  assign n5756 = x65 & n5755 ;
  assign n5747 = x47 ^ x46 ;
  assign n5748 = n5323 & ~n5747 ;
  assign n5749 = n5748 ^ n5323 ;
  assign n5752 = ~n152 & n5749 ;
  assign n5751 = x66 & n5323 ;
  assign n5753 = n5752 ^ n5751 ;
  assign n5757 = n5756 ^ n5753 ;
  assign n5761 = n5760 ^ n5757 ;
  assign n5746 = ~n5324 & ~n5553 ;
  assign n5762 = n5761 ^ n5746 ;
  assign n5769 = n5768 ^ n5762 ;
  assign n5763 = n5762 ^ n5757 ;
  assign n5744 = x46 & x64 ;
  assign n5745 = ~n5550 & n5744 ;
  assign n5764 = n5763 ^ n5745 ;
  assign n5765 = ~x47 & ~n5764 ;
  assign n5770 = n5769 ^ n5765 ;
  assign n5739 = x67 & n5113 ;
  assign n5738 = x69 & n5116 ;
  assign n5740 = n5739 ^ n5738 ;
  assign n5741 = n5740 ^ x44 ;
  assign n5737 = ~n376 & n5117 ;
  assign n5742 = n5741 ^ n5737 ;
  assign n5736 = x68 & n5121 ;
  assign n5743 = n5742 ^ n5736 ;
  assign n5771 = n5770 ^ n5743 ;
  assign n5773 = n5771 ^ n5534 ;
  assign n5772 = n5771 ^ n5563 ;
  assign n5774 = n5773 ^ n5772 ;
  assign n5775 = n5539 & n5774 ;
  assign n5776 = n5775 ^ n5773 ;
  assign n5785 = n5784 ^ n5776 ;
  assign n5733 = n5564 ^ n5523 ;
  assign n5734 = n5570 & n5733 ;
  assign n5735 = n5734 ^ n5564 ;
  assign n5786 = n5785 ^ n5735 ;
  assign n5795 = n5794 ^ n5786 ;
  assign n5796 = n5795 ^ x35 ;
  assign n5732 = x76 & n3387 ;
  assign n5797 = n5796 ^ n5732 ;
  assign n5731 = x78 & n3390 ;
  assign n5798 = n5797 ^ n5731 ;
  assign n5730 = ~n1036 & n3391 ;
  assign n5799 = n5798 ^ n5730 ;
  assign n5801 = n5800 ^ n5799 ;
  assign n5727 = n5571 ^ n5515 ;
  assign n5728 = n5520 & n5727 ;
  assign n5729 = n5728 ^ n5515 ;
  assign n5802 = n5801 ^ n5729 ;
  assign n5803 = n5802 ^ x32 ;
  assign n5726 = x79 & n2890 ;
  assign n5804 = n5803 ^ n5726 ;
  assign n5725 = x81 & n2893 ;
  assign n5805 = n5804 ^ n5725 ;
  assign n5724 = n1310 & n2894 ;
  assign n5806 = n5805 ^ n5724 ;
  assign n5808 = n5807 ^ n5806 ;
  assign n5721 = n5581 ^ n5572 ;
  assign n5722 = ~n5578 & n5721 ;
  assign n5723 = n5722 ^ n5581 ;
  assign n5809 = n5808 ^ n5723 ;
  assign n5810 = n5809 ^ x29 ;
  assign n5720 = x82 & n2593 ;
  assign n5811 = n5810 ^ n5720 ;
  assign n5719 = x84 & n2428 ;
  assign n5812 = n5811 ^ n5719 ;
  assign n5718 = n1635 & n2429 ;
  assign n5813 = n5812 ^ n5718 ;
  assign n5815 = n5814 ^ n5813 ;
  assign n5819 = n5818 ^ n5815 ;
  assign n5820 = n5819 ^ x26 ;
  assign n5717 = x85 & n2032 ;
  assign n5821 = n5820 ^ n5717 ;
  assign n5716 = x87 & n2028 ;
  assign n5822 = n5821 ^ n5716 ;
  assign n5715 = n1987 & n2029 ;
  assign n5823 = n5822 ^ n5715 ;
  assign n5825 = n5824 ^ n5823 ;
  assign n5829 = n5828 ^ n5825 ;
  assign n5830 = n5829 ^ x23 ;
  assign n5714 = x88 & n1665 ;
  assign n5831 = n5830 ^ n5714 ;
  assign n5713 = x90 & n1668 ;
  assign n5832 = n5831 ^ n5713 ;
  assign n5712 = n1669 & n2398 ;
  assign n5833 = n5832 ^ n5712 ;
  assign n5835 = n5834 ^ n5833 ;
  assign n5839 = n5838 ^ n5835 ;
  assign n5840 = n5839 ^ x20 ;
  assign n5711 = x91 & n1340 ;
  assign n5841 = n5840 ^ n5711 ;
  assign n5710 = x93 & n1343 ;
  assign n5842 = n5841 ^ n5710 ;
  assign n5709 = n1344 & n2842 ;
  assign n5843 = n5842 ^ n5709 ;
  assign n5845 = n5844 ^ n5843 ;
  assign n5706 = n5612 ^ n5603 ;
  assign n5707 = ~n5609 & n5706 ;
  assign n5708 = n5707 ^ n5612 ;
  assign n5846 = n5845 ^ n5708 ;
  assign n5847 = n5846 ^ x17 ;
  assign n5705 = x94 & n1060 ;
  assign n5848 = n5847 ^ n5705 ;
  assign n5704 = x96 & n1063 ;
  assign n5849 = n5848 ^ n5704 ;
  assign n5703 = n1064 & n3336 ;
  assign n5850 = n5849 ^ n5703 ;
  assign n5852 = n5851 ^ n5850 ;
  assign n5856 = n5855 ^ n5852 ;
  assign n5857 = n5856 ^ x14 ;
  assign n5702 = x97 & n884 ;
  assign n5858 = n5857 ^ n5702 ;
  assign n5701 = x99 & n789 ;
  assign n5859 = n5858 ^ n5701 ;
  assign n5700 = n790 & n3851 ;
  assign n5860 = n5859 ^ n5700 ;
  assign n5862 = n5861 ^ n5860 ;
  assign n5866 = n5865 ^ n5862 ;
  assign n5867 = n5866 ^ x11 ;
  assign n5699 = x100 & n650 ;
  assign n5868 = n5867 ^ n5699 ;
  assign n5698 = x102 & ~n578 ;
  assign n5869 = n5868 ^ n5698 ;
  assign n5697 = ~n579 & n4425 ;
  assign n5870 = n5869 ^ n5697 ;
  assign n5872 = n5871 ^ n5870 ;
  assign n5694 = n5636 ^ n5627 ;
  assign n5695 = ~n5633 & n5694 ;
  assign n5696 = n5695 ^ n5636 ;
  assign n5873 = n5872 ^ n5696 ;
  assign n5874 = n5873 ^ x8 ;
  assign n5693 = x103 & n456 ;
  assign n5875 = n5874 ^ n5693 ;
  assign n5692 = x105 & n384 ;
  assign n5876 = n5875 ^ n5692 ;
  assign n5691 = n385 & ~n5034 ;
  assign n5877 = n5876 ^ n5691 ;
  assign n5879 = n5878 ^ n5877 ;
  assign n5883 = n5882 ^ n5879 ;
  assign n5884 = n5883 ^ x5 ;
  assign n5690 = x106 & n238 ;
  assign n5885 = n5884 ^ n5690 ;
  assign n5689 = x108 & n234 ;
  assign n5886 = n5885 ^ n5689 ;
  assign n5687 = n5020 ^ x108 ;
  assign n5688 = n235 & n5687 ;
  assign n5887 = n5886 ^ n5688 ;
  assign n5889 = n5888 ^ n5887 ;
  assign n5684 = n5653 ^ n5644 ;
  assign n5685 = ~n5650 & n5684 ;
  assign n5686 = n5685 ^ n5653 ;
  assign n5890 = n5889 ^ n5686 ;
  assign n5666 = x109 & n5444 ;
  assign n5668 = n5666 ^ n5445 ;
  assign n5669 = x110 & n5668 ;
  assign n5667 = ~x110 & ~n5666 ;
  assign n5670 = n5669 ^ n5667 ;
  assign n5672 = x111 ^ x1 ;
  assign n5671 = x111 ^ x2 ;
  assign n5673 = n5672 ^ n5671 ;
  assign n5674 = n5670 & n5673 ;
  assign n5675 = n5674 ^ n5672 ;
  assign n5891 = n5890 ^ n5675 ;
  assign n5679 = x2 & x109 ;
  assign n5680 = n5679 ^ x110 ;
  assign n5681 = ~x1 & n5680 ;
  assign n5676 = n5675 ^ n5446 ;
  assign n5682 = n5681 ^ n5676 ;
  assign n5683 = ~x0 & n5682 ;
  assign n5892 = n5891 ^ n5683 ;
  assign n5661 = n5659 ^ n5654 ;
  assign n5662 = ~n5656 & n5661 ;
  assign n5663 = n5662 ^ n5659 ;
  assign n5893 = n5892 ^ n5663 ;
  assign n6117 = n5890 ^ n5663 ;
  assign n6118 = ~n5892 & ~n6117 ;
  assign n6119 = n6118 ^ n5890 ;
  assign n6111 = n5883 ^ n5686 ;
  assign n6112 = ~n5889 & ~n6111 ;
  assign n6113 = n6112 ^ n5883 ;
  assign n6109 = x108 & n231 ;
  assign n6102 = x105 & n391 ;
  assign n6094 = n5866 ^ n5696 ;
  assign n6095 = ~n5872 & ~n6094 ;
  assign n6096 = n6095 ^ n5866 ;
  assign n6092 = x102 & n584 ;
  assign n6085 = x99 & n795 ;
  assign n6078 = x96 & n1068 ;
  assign n6070 = n5839 ^ n5708 ;
  assign n6071 = ~n5845 & ~n6070 ;
  assign n6072 = n6071 ^ n5839 ;
  assign n6068 = x93 & n1348 ;
  assign n6061 = x90 & n1673 ;
  assign n6054 = x87 & n2025 ;
  assign n6047 = x84 & n2435 ;
  assign n6039 = n5802 ^ n5723 ;
  assign n6040 = ~n5808 & ~n6039 ;
  assign n6041 = n6040 ^ n5802 ;
  assign n6037 = x81 & n2899 ;
  assign n6027 = x77 & n3387 ;
  assign n6026 = x79 & n3390 ;
  assign n6028 = n6027 ^ n6026 ;
  assign n6029 = n6028 ^ x35 ;
  assign n6025 = n1123 & n3391 ;
  assign n6030 = n6029 ^ n6025 ;
  assign n6024 = x78 & n3395 ;
  assign n6031 = n6030 ^ n6024 ;
  assign n6020 = x75 & n3940 ;
  assign n6010 = x71 & n4482 ;
  assign n6009 = x73 & n4478 ;
  assign n6011 = n6010 ^ n6009 ;
  assign n6012 = n6011 ^ x41 ;
  assign n6008 = n636 & n4479 ;
  assign n6013 = n6012 ^ n6008 ;
  assign n6007 = x72 & n4475 ;
  assign n6014 = n6013 ^ n6007 ;
  assign n5998 = n5768 ^ n5743 ;
  assign n5999 = ~n5770 & n5998 ;
  assign n6000 = n5999 ^ n5768 ;
  assign n5996 = x69 & n5121 ;
  assign n5988 = n5746 & ~n5761 ;
  assign n5989 = x47 & n5988 ;
  assign n5986 = x48 ^ x47 ;
  assign n5987 = x64 & n5986 ;
  assign n5990 = n5989 ^ n5987 ;
  assign n5979 = x47 ^ x45 ;
  assign n5980 = ~n5323 & n5979 ;
  assign n5981 = n5747 & n5980 ;
  assign n5982 = x65 & n5981 ;
  assign n5978 = x66 & n5755 ;
  assign n5983 = n5982 ^ n5978 ;
  assign n5984 = n5983 ^ x47 ;
  assign n5975 = ~n155 & ~n5747 ;
  assign n5976 = n5975 ^ n295 ;
  assign n5977 = n5323 & ~n5976 ;
  assign n5985 = n5984 ^ n5977 ;
  assign n5991 = n5990 ^ n5985 ;
  assign n5992 = n5991 ^ x44 ;
  assign n5972 = x68 & n5113 ;
  assign n5993 = n5992 ^ n5972 ;
  assign n5971 = x70 & n5116 ;
  assign n5994 = n5993 ^ n5971 ;
  assign n5970 = ~n443 & n5117 ;
  assign n5995 = n5994 ^ n5970 ;
  assign n5997 = n5996 ^ n5995 ;
  assign n6001 = n6000 ^ n5997 ;
  assign n6003 = n6001 ^ n5771 ;
  assign n6002 = n6001 ^ n5784 ;
  assign n6004 = n6003 ^ n6002 ;
  assign n6005 = ~n5776 & ~n6004 ;
  assign n6006 = n6005 ^ n6003 ;
  assign n6015 = n6014 ^ n6006 ;
  assign n6016 = n6015 ^ x38 ;
  assign n5969 = x74 & n3932 ;
  assign n6017 = n6016 ^ n5969 ;
  assign n5968 = x76 & n3935 ;
  assign n6018 = n6017 ^ n5968 ;
  assign n5967 = ~n863 & n3936 ;
  assign n6019 = n6018 ^ n5967 ;
  assign n6021 = n6020 ^ n6019 ;
  assign n5964 = n5794 ^ n5735 ;
  assign n5965 = n5786 & n5964 ;
  assign n5966 = n5965 ^ n5794 ;
  assign n6022 = n6021 ^ n5966 ;
  assign n5961 = n5795 ^ n5729 ;
  assign n5962 = ~n5801 & ~n5961 ;
  assign n5963 = n5962 ^ n5795 ;
  assign n6023 = n6022 ^ n5963 ;
  assign n6032 = n6031 ^ n6023 ;
  assign n6033 = n6032 ^ x32 ;
  assign n5960 = x80 & n2890 ;
  assign n6034 = n6033 ^ n5960 ;
  assign n5959 = x82 & n2893 ;
  assign n6035 = n6034 ^ n5959 ;
  assign n5958 = n1422 & n2894 ;
  assign n6036 = n6035 ^ n5958 ;
  assign n6038 = n6037 ^ n6036 ;
  assign n6042 = n6041 ^ n6038 ;
  assign n6043 = n6042 ^ x29 ;
  assign n5957 = x83 & n2593 ;
  assign n6044 = n6043 ^ n5957 ;
  assign n5956 = x85 & n2428 ;
  assign n6045 = n6044 ^ n5956 ;
  assign n5955 = n1748 & n2429 ;
  assign n6046 = n6045 ^ n5955 ;
  assign n6048 = n6047 ^ n6046 ;
  assign n5952 = n5818 ^ n5809 ;
  assign n5953 = n5815 & ~n5952 ;
  assign n5954 = n5953 ^ n5818 ;
  assign n6049 = n6048 ^ n5954 ;
  assign n6050 = n6049 ^ x26 ;
  assign n5951 = x86 & n2032 ;
  assign n6051 = n6050 ^ n5951 ;
  assign n5950 = x88 & n2028 ;
  assign n6052 = n6051 ^ n5950 ;
  assign n5949 = n2029 & n2131 ;
  assign n6053 = n6052 ^ n5949 ;
  assign n6055 = n6054 ^ n6053 ;
  assign n5946 = n5828 ^ n5819 ;
  assign n5947 = n5825 & ~n5946 ;
  assign n5948 = n5947 ^ n5828 ;
  assign n6056 = n6055 ^ n5948 ;
  assign n6057 = n6056 ^ x23 ;
  assign n5945 = x89 & n1665 ;
  assign n6058 = n6057 ^ n5945 ;
  assign n5944 = x91 & n1668 ;
  assign n6059 = n6058 ^ n5944 ;
  assign n5943 = n1669 & n2548 ;
  assign n6060 = n6059 ^ n5943 ;
  assign n6062 = n6061 ^ n6060 ;
  assign n5940 = n5838 ^ n5829 ;
  assign n5941 = n5835 & ~n5940 ;
  assign n5942 = n5941 ^ n5838 ;
  assign n6063 = n6062 ^ n5942 ;
  assign n6064 = n6063 ^ x20 ;
  assign n5939 = x92 & n1340 ;
  assign n6065 = n6064 ^ n5939 ;
  assign n5938 = x94 & n1343 ;
  assign n6066 = n6065 ^ n5938 ;
  assign n5937 = n1344 & n3010 ;
  assign n6067 = n6066 ^ n5937 ;
  assign n6069 = n6068 ^ n6067 ;
  assign n6073 = n6072 ^ n6069 ;
  assign n6074 = n6073 ^ x17 ;
  assign n5936 = x95 & n1060 ;
  assign n6075 = n6074 ^ n5936 ;
  assign n5935 = x97 & n1063 ;
  assign n6076 = n6075 ^ n5935 ;
  assign n5934 = n1064 & n3501 ;
  assign n6077 = n6076 ^ n5934 ;
  assign n6079 = n6078 ^ n6077 ;
  assign n5931 = n5855 ^ n5846 ;
  assign n5932 = n5852 & ~n5931 ;
  assign n5933 = n5932 ^ n5855 ;
  assign n6080 = n6079 ^ n5933 ;
  assign n6081 = n6080 ^ x14 ;
  assign n5930 = x98 & n884 ;
  assign n6082 = n6081 ^ n5930 ;
  assign n5929 = x100 & n789 ;
  assign n6083 = n6082 ^ n5929 ;
  assign n5928 = n790 & n4048 ;
  assign n6084 = n6083 ^ n5928 ;
  assign n6086 = n6085 ^ n6084 ;
  assign n5925 = n5865 ^ n5856 ;
  assign n5926 = n5862 & ~n5925 ;
  assign n5927 = n5926 ^ n5865 ;
  assign n6087 = n6086 ^ n5927 ;
  assign n6088 = n6087 ^ x11 ;
  assign n5924 = x101 & n650 ;
  assign n6089 = n6088 ^ n5924 ;
  assign n5923 = x103 & ~n578 ;
  assign n6090 = n6089 ^ n5923 ;
  assign n5922 = ~n579 & ~n4624 ;
  assign n6091 = n6090 ^ n5922 ;
  assign n6093 = n6092 ^ n6091 ;
  assign n6097 = n6096 ^ n6093 ;
  assign n6098 = n6097 ^ x8 ;
  assign n5921 = x104 & n456 ;
  assign n6099 = n6098 ^ n5921 ;
  assign n5920 = x106 & n384 ;
  assign n6100 = n6099 ^ n5920 ;
  assign n5919 = n385 & ~n5257 ;
  assign n6101 = n6100 ^ n5919 ;
  assign n6103 = n6102 ^ n6101 ;
  assign n5916 = n5882 ^ n5873 ;
  assign n5917 = n5879 & ~n5916 ;
  assign n5918 = n5917 ^ n5882 ;
  assign n6104 = n6103 ^ n5918 ;
  assign n6105 = n6104 ^ x5 ;
  assign n5915 = x107 & n238 ;
  assign n6106 = n6105 ^ n5915 ;
  assign n5914 = x109 & n234 ;
  assign n6107 = n6106 ^ n5914 ;
  assign n5912 = n5240 ^ x109 ;
  assign n5913 = n235 & n5912 ;
  assign n6108 = n6107 ^ n5913 ;
  assign n6110 = n6109 ^ n6108 ;
  assign n6114 = n6113 ^ n6110 ;
  assign n5897 = ~x111 & ~n5669 ;
  assign n5896 = x111 & ~n5667 ;
  assign n5898 = n5897 ^ n5896 ;
  assign n5900 = x112 ^ x1 ;
  assign n5899 = x112 ^ x2 ;
  assign n5901 = n5900 ^ n5899 ;
  assign n5902 = n5898 & n5901 ;
  assign n5903 = n5902 ^ n5900 ;
  assign n6115 = n6114 ^ n5903 ;
  assign n5907 = x2 & x110 ;
  assign n5908 = n5907 ^ x111 ;
  assign n5909 = ~x1 & n5908 ;
  assign n5904 = n5903 ^ n5671 ;
  assign n5910 = n5909 ^ n5904 ;
  assign n5911 = ~x0 & n5910 ;
  assign n6116 = n6115 ^ n5911 ;
  assign n6120 = n6119 ^ n6116 ;
  assign n6346 = x109 & n231 ;
  assign n6338 = n6097 ^ n5918 ;
  assign n6339 = ~n6103 & ~n6338 ;
  assign n6340 = n6339 ^ n6097 ;
  assign n6336 = x106 & n391 ;
  assign n6329 = x103 & n584 ;
  assign n6321 = n6080 ^ n5927 ;
  assign n6322 = n6086 & n6321 ;
  assign n6323 = n6322 ^ n6080 ;
  assign n6319 = x100 & n795 ;
  assign n6311 = n6073 ^ n5933 ;
  assign n6312 = n6079 & n6311 ;
  assign n6313 = n6312 ^ n6073 ;
  assign n6309 = x97 & n1068 ;
  assign n6302 = x94 & n1348 ;
  assign n6294 = n6056 ^ n5942 ;
  assign n6295 = ~n6062 & ~n6294 ;
  assign n6296 = n6295 ^ n6056 ;
  assign n6292 = x91 & n1673 ;
  assign n6284 = n6049 ^ n5948 ;
  assign n6285 = ~n6055 & ~n6284 ;
  assign n6286 = n6285 ^ n6049 ;
  assign n6282 = x88 & n2025 ;
  assign n6274 = n6042 ^ n5954 ;
  assign n6275 = ~n6048 & ~n6274 ;
  assign n6276 = n6275 ^ n6042 ;
  assign n6272 = x85 & n2435 ;
  assign n6265 = x82 & n2899 ;
  assign n6258 = x79 & n3395 ;
  assign n6251 = x76 & n3940 ;
  assign n6243 = n6014 ^ n6001 ;
  assign n6244 = ~n6006 & n6243 ;
  assign n6245 = n6244 ^ n6001 ;
  assign n6241 = x73 & n4475 ;
  assign n6234 = x70 & n5121 ;
  assign n6224 = x66 & n5981 ;
  assign n6223 = x68 & n5748 ;
  assign n6225 = n6224 ^ n6223 ;
  assign n6226 = n6225 ^ x47 ;
  assign n6222 = ~n351 & n5749 ;
  assign n6227 = n6226 ^ n6222 ;
  assign n6221 = x67 & n5755 ;
  assign n6228 = n6227 ^ n6221 ;
  assign n6217 = ~n5987 & ~n5989 ;
  assign n6218 = n5985 & n6217 ;
  assign n6219 = n6218 ^ n5985 ;
  assign n6214 = x65 ^ x48 ;
  assign n6215 = n5986 & ~n6214 ;
  assign n6210 = x47 & x48 ;
  assign n6211 = n6210 ^ x49 ;
  assign n6212 = ~x64 & n6211 ;
  assign n6206 = x49 ^ x47 ;
  assign n6213 = n6212 ^ n6206 ;
  assign n6216 = n6215 ^ n6213 ;
  assign n6220 = n6219 ^ n6216 ;
  assign n6229 = n6228 ^ n6220 ;
  assign n6230 = n6229 ^ x44 ;
  assign n6205 = x69 & n5113 ;
  assign n6231 = n6230 ^ n6205 ;
  assign n6204 = x71 & n5116 ;
  assign n6232 = n6231 ^ n6204 ;
  assign n6203 = ~n495 & n5117 ;
  assign n6233 = n6232 ^ n6203 ;
  assign n6235 = n6234 ^ n6233 ;
  assign n6200 = n6000 ^ n5991 ;
  assign n6201 = ~n5997 & n6200 ;
  assign n6202 = n6201 ^ n6000 ;
  assign n6236 = n6235 ^ n6202 ;
  assign n6237 = n6236 ^ x41 ;
  assign n6199 = x72 & n4482 ;
  assign n6238 = n6237 ^ n6199 ;
  assign n6198 = x74 & n4478 ;
  assign n6239 = n6238 ^ n6198 ;
  assign n6197 = n708 & n4479 ;
  assign n6240 = n6239 ^ n6197 ;
  assign n6242 = n6241 ^ n6240 ;
  assign n6246 = n6245 ^ n6242 ;
  assign n6247 = n6246 ^ x38 ;
  assign n6196 = x75 & n3932 ;
  assign n6248 = n6247 ^ n6196 ;
  assign n6195 = x77 & n3935 ;
  assign n6249 = n6248 ^ n6195 ;
  assign n6194 = ~n943 & n3936 ;
  assign n6250 = n6249 ^ n6194 ;
  assign n6252 = n6251 ^ n6250 ;
  assign n6191 = n6015 ^ n5966 ;
  assign n6192 = ~n6021 & ~n6191 ;
  assign n6193 = n6192 ^ n6015 ;
  assign n6253 = n6252 ^ n6193 ;
  assign n6254 = n6253 ^ x35 ;
  assign n6190 = x78 & n3387 ;
  assign n6255 = n6254 ^ n6190 ;
  assign n6189 = x80 & n3390 ;
  assign n6256 = n6255 ^ n6189 ;
  assign n6188 = n1217 & n3391 ;
  assign n6257 = n6256 ^ n6188 ;
  assign n6259 = n6258 ^ n6257 ;
  assign n6185 = n6031 ^ n5963 ;
  assign n6186 = ~n6023 & ~n6185 ;
  assign n6187 = n6186 ^ n6031 ;
  assign n6260 = n6259 ^ n6187 ;
  assign n6261 = n6260 ^ x32 ;
  assign n6184 = x81 & n2890 ;
  assign n6262 = n6261 ^ n6184 ;
  assign n6183 = x83 & n2893 ;
  assign n6263 = n6262 ^ n6183 ;
  assign n6182 = n1517 & n2894 ;
  assign n6264 = n6263 ^ n6182 ;
  assign n6266 = n6265 ^ n6264 ;
  assign n6179 = n6041 ^ n6032 ;
  assign n6180 = ~n6038 & ~n6179 ;
  assign n6181 = n6180 ^ n6041 ;
  assign n6267 = n6266 ^ n6181 ;
  assign n6268 = n6267 ^ x29 ;
  assign n6178 = x84 & n2593 ;
  assign n6269 = n6268 ^ n6178 ;
  assign n6177 = x86 & n2428 ;
  assign n6270 = n6269 ^ n6177 ;
  assign n6176 = n1868 & n2429 ;
  assign n6271 = n6270 ^ n6176 ;
  assign n6273 = n6272 ^ n6271 ;
  assign n6277 = n6276 ^ n6273 ;
  assign n6278 = n6277 ^ x26 ;
  assign n6175 = x87 & n2032 ;
  assign n6279 = n6278 ^ n6175 ;
  assign n6174 = x89 & n2028 ;
  assign n6280 = n6279 ^ n6174 ;
  assign n6173 = n2029 & n2255 ;
  assign n6281 = n6280 ^ n6173 ;
  assign n6283 = n6282 ^ n6281 ;
  assign n6287 = n6286 ^ n6283 ;
  assign n6288 = n6287 ^ x23 ;
  assign n6172 = x90 & n1665 ;
  assign n6289 = n6288 ^ n6172 ;
  assign n6171 = x92 & n1668 ;
  assign n6290 = n6289 ^ n6171 ;
  assign n6170 = n1669 & n2696 ;
  assign n6291 = n6290 ^ n6170 ;
  assign n6293 = n6292 ^ n6291 ;
  assign n6297 = n6296 ^ n6293 ;
  assign n6298 = n6297 ^ x20 ;
  assign n6169 = x93 & n1340 ;
  assign n6299 = n6298 ^ n6169 ;
  assign n6168 = x95 & n1343 ;
  assign n6300 = n6299 ^ n6168 ;
  assign n6167 = n1344 & n3166 ;
  assign n6301 = n6300 ^ n6167 ;
  assign n6303 = n6302 ^ n6301 ;
  assign n6164 = n6072 ^ n6063 ;
  assign n6165 = n6069 & n6164 ;
  assign n6166 = n6165 ^ n6072 ;
  assign n6304 = n6303 ^ n6166 ;
  assign n6305 = n6304 ^ x17 ;
  assign n6163 = x96 & n1060 ;
  assign n6306 = n6305 ^ n6163 ;
  assign n6162 = x98 & n1063 ;
  assign n6307 = n6306 ^ n6162 ;
  assign n6161 = n1064 & n3673 ;
  assign n6308 = n6307 ^ n6161 ;
  assign n6310 = n6309 ^ n6308 ;
  assign n6314 = n6313 ^ n6310 ;
  assign n6315 = n6314 ^ x14 ;
  assign n6160 = x99 & n884 ;
  assign n6316 = n6315 ^ n6160 ;
  assign n6159 = x101 & n789 ;
  assign n6317 = n6316 ^ n6159 ;
  assign n6158 = n790 & n4223 ;
  assign n6318 = n6317 ^ n6158 ;
  assign n6320 = n6319 ^ n6318 ;
  assign n6324 = n6323 ^ n6320 ;
  assign n6325 = n6324 ^ x11 ;
  assign n6157 = x102 & n650 ;
  assign n6326 = n6325 ^ n6157 ;
  assign n6156 = x104 & ~n578 ;
  assign n6327 = n6326 ^ n6156 ;
  assign n6155 = ~n579 & ~n4830 ;
  assign n6328 = n6327 ^ n6155 ;
  assign n6330 = n6329 ^ n6328 ;
  assign n6152 = n6096 ^ n6087 ;
  assign n6153 = ~n6093 & ~n6152 ;
  assign n6154 = n6153 ^ n6096 ;
  assign n6331 = n6330 ^ n6154 ;
  assign n6332 = n6331 ^ x8 ;
  assign n6151 = x105 & n456 ;
  assign n6333 = n6332 ^ n6151 ;
  assign n6150 = x107 & n384 ;
  assign n6334 = n6333 ^ n6150 ;
  assign n6149 = n385 & ~n5459 ;
  assign n6335 = n6334 ^ n6149 ;
  assign n6337 = n6336 ^ n6335 ;
  assign n6341 = n6340 ^ n6337 ;
  assign n6342 = n6341 ^ x5 ;
  assign n6148 = x108 & n238 ;
  assign n6343 = n6342 ^ n6148 ;
  assign n6147 = x110 & n234 ;
  assign n6344 = n6343 ^ n6147 ;
  assign n5664 = x110 ^ x109 ;
  assign n6145 = n5664 ^ n5444 ;
  assign n6146 = n235 & n6145 ;
  assign n6345 = n6344 ^ n6146 ;
  assign n6347 = n6346 ^ n6345 ;
  assign n6142 = n6113 ^ n6104 ;
  assign n6143 = n6110 & n6142 ;
  assign n6144 = n6143 ^ n6113 ;
  assign n6348 = n6347 ^ n6144 ;
  assign n6127 = x112 & ~n5897 ;
  assign n6126 = ~x112 & ~n5896 ;
  assign n6128 = n6127 ^ n6126 ;
  assign n6130 = x113 ^ x1 ;
  assign n6129 = x113 ^ x2 ;
  assign n6131 = n6130 ^ n6129 ;
  assign n6132 = n6128 & n6131 ;
  assign n6133 = n6132 ^ n6130 ;
  assign n6349 = n6348 ^ n6133 ;
  assign n6137 = x2 & x111 ;
  assign n6138 = n6137 ^ x112 ;
  assign n6139 = ~x1 & n6138 ;
  assign n6134 = n6133 ^ n5899 ;
  assign n6140 = n6139 ^ n6134 ;
  assign n6141 = ~x0 & n6140 ;
  assign n6350 = n6349 ^ n6141 ;
  assign n6121 = n6119 ^ n6114 ;
  assign n6122 = ~n6116 & ~n6121 ;
  assign n6123 = n6122 ^ n6119 ;
  assign n6351 = n6350 ^ n6123 ;
  assign n6588 = n6348 ^ n6123 ;
  assign n6589 = ~n6350 & n6588 ;
  assign n6590 = n6589 ^ n6348 ;
  assign n6582 = n6341 ^ n6144 ;
  assign n6583 = n6347 & ~n6582 ;
  assign n6584 = n6583 ^ n6341 ;
  assign n6580 = x110 & n231 ;
  assign n6573 = x107 & n391 ;
  assign n6565 = n6324 ^ n6154 ;
  assign n6566 = n6330 & ~n6565 ;
  assign n6567 = n6566 ^ n6324 ;
  assign n6563 = x104 & n584 ;
  assign n6556 = x101 & n795 ;
  assign n6549 = x98 & n1068 ;
  assign n6541 = n6297 ^ n6166 ;
  assign n6542 = ~n6303 & n6541 ;
  assign n6543 = n6542 ^ n6297 ;
  assign n6539 = x95 & n1348 ;
  assign n6532 = x92 & n1673 ;
  assign n6525 = x89 & n2025 ;
  assign n6518 = x86 & n2435 ;
  assign n6510 = n6260 ^ n6181 ;
  assign n6511 = ~n6266 & n6510 ;
  assign n6512 = n6511 ^ n6260 ;
  assign n6504 = x82 & n2890 ;
  assign n6503 = x84 & n2893 ;
  assign n6505 = n6504 ^ n6503 ;
  assign n6506 = n6505 ^ x32 ;
  assign n6502 = n1635 & n2894 ;
  assign n6507 = n6506 ^ n6502 ;
  assign n6501 = x83 & n2899 ;
  assign n6508 = n6507 ^ n6501 ;
  assign n6498 = x80 & n3395 ;
  assign n6490 = n6246 ^ n6193 ;
  assign n6491 = n6252 & ~n6490 ;
  assign n6492 = n6491 ^ n6246 ;
  assign n6488 = x77 & n3940 ;
  assign n6477 = x70 & n5113 ;
  assign n6476 = x72 & n5116 ;
  assign n6478 = n6477 ^ n6476 ;
  assign n6479 = n6478 ^ x44 ;
  assign n6475 = n565 & n5117 ;
  assign n6480 = n6479 ^ n6475 ;
  assign n6474 = x71 & n5121 ;
  assign n6481 = n6480 ^ n6474 ;
  assign n6471 = n6229 ^ n6202 ;
  assign n6472 = n6235 & n6471 ;
  assign n6461 = x67 & n5981 ;
  assign n6460 = x69 & n5748 ;
  assign n6462 = n6461 ^ n6460 ;
  assign n6463 = n6462 ^ x47 ;
  assign n6459 = ~n376 & n5749 ;
  assign n6464 = n6463 ^ n6459 ;
  assign n6458 = x68 & n5755 ;
  assign n6465 = n6464 ^ n6458 ;
  assign n6456 = ~n5987 & ~n6216 ;
  assign n6457 = x50 & n6456 ;
  assign n6466 = n6465 ^ n6457 ;
  assign n6441 = x64 & ~n6206 ;
  assign n6208 = x49 ^ x48 ;
  assign n6449 = ~n5986 & n6208 ;
  assign n6450 = x65 & n6449 ;
  assign n6443 = x50 ^ x49 ;
  assign n6444 = n5986 & ~n6443 ;
  assign n6445 = n6444 ^ n5986 ;
  assign n6446 = ~n152 & n6445 ;
  assign n6442 = x66 & n5986 ;
  assign n6447 = n6446 ^ n6442 ;
  assign n6448 = n6447 ^ x50 ;
  assign n6451 = n6450 ^ n6448 ;
  assign n6452 = n6451 ^ x47 ;
  assign n6453 = ~n6208 & n6452 ;
  assign n6454 = n6441 & n6453 ;
  assign n6455 = n6454 ^ n6451 ;
  assign n6467 = n6466 ^ n6455 ;
  assign n6438 = n6228 ^ n6219 ;
  assign n6439 = ~n6220 & n6438 ;
  assign n6440 = n6439 ^ n6228 ;
  assign n6468 = n6467 ^ n6440 ;
  assign n6469 = n6468 ^ n6229 ;
  assign n6473 = n6472 ^ n6469 ;
  assign n6482 = n6481 ^ n6473 ;
  assign n6428 = x73 & n4482 ;
  assign n6427 = x75 & n4478 ;
  assign n6429 = n6428 ^ n6427 ;
  assign n6430 = n6429 ^ x41 ;
  assign n6426 = ~n778 & n4479 ;
  assign n6431 = n6430 ^ n6426 ;
  assign n6425 = x74 & n4475 ;
  assign n6432 = n6431 ^ n6425 ;
  assign n6433 = n6432 ^ n6245 ;
  assign n6434 = n6433 ^ n6236 ;
  assign n6435 = n6434 ^ n6432 ;
  assign n6436 = ~n6242 & n6435 ;
  assign n6437 = n6436 ^ n6433 ;
  assign n6483 = n6482 ^ n6437 ;
  assign n6484 = n6483 ^ x38 ;
  assign n6424 = x76 & n3932 ;
  assign n6485 = n6484 ^ n6424 ;
  assign n6423 = x78 & n3935 ;
  assign n6486 = n6485 ^ n6423 ;
  assign n6422 = ~n1036 & n3936 ;
  assign n6487 = n6486 ^ n6422 ;
  assign n6489 = n6488 ^ n6487 ;
  assign n6493 = n6492 ^ n6489 ;
  assign n6494 = n6493 ^ x35 ;
  assign n6421 = x79 & n3387 ;
  assign n6495 = n6494 ^ n6421 ;
  assign n6420 = x81 & n3390 ;
  assign n6496 = n6495 ^ n6420 ;
  assign n6419 = n1310 & n3391 ;
  assign n6497 = n6496 ^ n6419 ;
  assign n6499 = n6498 ^ n6497 ;
  assign n6416 = n6253 ^ n6187 ;
  assign n6417 = ~n6259 & ~n6416 ;
  assign n6418 = n6417 ^ n6253 ;
  assign n6500 = n6499 ^ n6418 ;
  assign n6509 = n6508 ^ n6500 ;
  assign n6513 = n6512 ^ n6509 ;
  assign n6514 = n6513 ^ x29 ;
  assign n6415 = x85 & n2593 ;
  assign n6515 = n6514 ^ n6415 ;
  assign n6414 = x87 & n2428 ;
  assign n6516 = n6515 ^ n6414 ;
  assign n6413 = n1987 & n2429 ;
  assign n6517 = n6516 ^ n6413 ;
  assign n6519 = n6518 ^ n6517 ;
  assign n6410 = n6276 ^ n6267 ;
  assign n6411 = ~n6273 & ~n6410 ;
  assign n6412 = n6411 ^ n6276 ;
  assign n6520 = n6519 ^ n6412 ;
  assign n6521 = n6520 ^ x26 ;
  assign n6409 = x88 & n2032 ;
  assign n6522 = n6521 ^ n6409 ;
  assign n6408 = x90 & n2028 ;
  assign n6523 = n6522 ^ n6408 ;
  assign n6407 = n2029 & n2398 ;
  assign n6524 = n6523 ^ n6407 ;
  assign n6526 = n6525 ^ n6524 ;
  assign n6404 = n6286 ^ n6277 ;
  assign n6405 = n6283 & n6404 ;
  assign n6406 = n6405 ^ n6286 ;
  assign n6527 = n6526 ^ n6406 ;
  assign n6528 = n6527 ^ x23 ;
  assign n6403 = x91 & n1665 ;
  assign n6529 = n6528 ^ n6403 ;
  assign n6402 = x93 & n1668 ;
  assign n6530 = n6529 ^ n6402 ;
  assign n6401 = n1669 & n2842 ;
  assign n6531 = n6530 ^ n6401 ;
  assign n6533 = n6532 ^ n6531 ;
  assign n6398 = n6296 ^ n6287 ;
  assign n6399 = ~n6293 & ~n6398 ;
  assign n6400 = n6399 ^ n6296 ;
  assign n6534 = n6533 ^ n6400 ;
  assign n6535 = n6534 ^ x20 ;
  assign n6397 = x94 & n1340 ;
  assign n6536 = n6535 ^ n6397 ;
  assign n6396 = x96 & n1343 ;
  assign n6537 = n6536 ^ n6396 ;
  assign n6395 = n1344 & n3336 ;
  assign n6538 = n6537 ^ n6395 ;
  assign n6540 = n6539 ^ n6538 ;
  assign n6544 = n6543 ^ n6540 ;
  assign n6545 = n6544 ^ x17 ;
  assign n6394 = x97 & n1060 ;
  assign n6546 = n6545 ^ n6394 ;
  assign n6393 = x99 & n1063 ;
  assign n6547 = n6546 ^ n6393 ;
  assign n6392 = n1064 & n3851 ;
  assign n6548 = n6547 ^ n6392 ;
  assign n6550 = n6549 ^ n6548 ;
  assign n6389 = n6313 ^ n6304 ;
  assign n6390 = ~n6310 & n6389 ;
  assign n6391 = n6390 ^ n6313 ;
  assign n6551 = n6550 ^ n6391 ;
  assign n6552 = n6551 ^ x14 ;
  assign n6388 = x100 & n884 ;
  assign n6553 = n6552 ^ n6388 ;
  assign n6387 = x102 & n789 ;
  assign n6554 = n6553 ^ n6387 ;
  assign n6386 = n790 & n4425 ;
  assign n6555 = n6554 ^ n6386 ;
  assign n6557 = n6556 ^ n6555 ;
  assign n6383 = n6323 ^ n6314 ;
  assign n6384 = ~n6320 & n6383 ;
  assign n6385 = n6384 ^ n6323 ;
  assign n6558 = n6557 ^ n6385 ;
  assign n6559 = n6558 ^ x11 ;
  assign n6382 = x103 & n650 ;
  assign n6560 = n6559 ^ n6382 ;
  assign n6381 = x105 & ~n578 ;
  assign n6561 = n6560 ^ n6381 ;
  assign n6380 = ~n579 & ~n5034 ;
  assign n6562 = n6561 ^ n6380 ;
  assign n6564 = n6563 ^ n6562 ;
  assign n6568 = n6567 ^ n6564 ;
  assign n6569 = n6568 ^ x8 ;
  assign n6379 = x106 & n456 ;
  assign n6570 = n6569 ^ n6379 ;
  assign n6378 = x108 & n384 ;
  assign n6571 = n6570 ^ n6378 ;
  assign n6377 = n385 & n5687 ;
  assign n6572 = n6571 ^ n6377 ;
  assign n6574 = n6573 ^ n6572 ;
  assign n6374 = n6340 ^ n6331 ;
  assign n6375 = n6337 & n6374 ;
  assign n6376 = n6375 ^ n6340 ;
  assign n6575 = n6574 ^ n6376 ;
  assign n6576 = n6575 ^ x5 ;
  assign n6373 = x109 & n238 ;
  assign n6577 = n6576 ^ n6373 ;
  assign n6372 = x111 & n234 ;
  assign n6578 = n6577 ^ n6372 ;
  assign n6370 = n5670 ^ x111 ;
  assign n6371 = n235 & ~n6370 ;
  assign n6579 = n6578 ^ n6371 ;
  assign n6581 = n6580 ^ n6579 ;
  assign n6585 = n6584 ^ n6581 ;
  assign n6355 = ~x113 & ~n6127 ;
  assign n6354 = x113 & ~n6126 ;
  assign n6356 = n6355 ^ n6354 ;
  assign n6358 = x114 ^ x1 ;
  assign n6357 = x114 ^ x2 ;
  assign n6359 = n6358 ^ n6357 ;
  assign n6360 = n6356 & n6359 ;
  assign n6361 = n6360 ^ n6358 ;
  assign n6586 = n6585 ^ n6361 ;
  assign n6365 = x2 & x112 ;
  assign n6366 = n6365 ^ x113 ;
  assign n6367 = ~x1 & n6366 ;
  assign n6362 = n6361 ^ n6129 ;
  assign n6368 = n6367 ^ n6362 ;
  assign n6369 = ~x0 & n6368 ;
  assign n6587 = n6586 ^ n6369 ;
  assign n6591 = n6590 ^ n6587 ;
  assign n6825 = x111 & n231 ;
  assign n6817 = n6568 ^ n6376 ;
  assign n6818 = n6574 & ~n6817 ;
  assign n6819 = n6818 ^ n6568 ;
  assign n6815 = x108 & n391 ;
  assign n6808 = x105 & n584 ;
  assign n6800 = n6551 ^ n6385 ;
  assign n6801 = n6557 & n6800 ;
  assign n6802 = n6801 ^ n6551 ;
  assign n6798 = x102 & n795 ;
  assign n6790 = n6544 ^ n6391 ;
  assign n6791 = n6550 & n6790 ;
  assign n6792 = n6791 ^ n6544 ;
  assign n6788 = x99 & n1068 ;
  assign n6781 = x96 & n1348 ;
  assign n6773 = n6527 ^ n6400 ;
  assign n6774 = n6533 & ~n6773 ;
  assign n6775 = n6774 ^ n6527 ;
  assign n6771 = x93 & n1673 ;
  assign n6763 = n6520 ^ n6406 ;
  assign n6764 = ~n6526 & n6763 ;
  assign n6765 = n6764 ^ n6520 ;
  assign n6761 = x90 & n2025 ;
  assign n6753 = n6513 ^ n6412 ;
  assign n6754 = n6519 & ~n6753 ;
  assign n6755 = n6754 ^ n6513 ;
  assign n6751 = x87 & n2435 ;
  assign n6744 = x84 & n2899 ;
  assign n6742 = n1748 & n2894 ;
  assign n6738 = x83 & n2890 ;
  assign n6737 = x85 & n2893 ;
  assign n6739 = n6738 ^ n6737 ;
  assign n6740 = n6739 ^ x32 ;
  assign n6733 = n6493 ^ n6418 ;
  assign n6734 = n6499 & ~n6733 ;
  assign n6735 = n6734 ^ n6493 ;
  assign n6731 = x81 & n3395 ;
  assign n6723 = x75 & n4475 ;
  assign n6715 = n6481 ^ n6468 ;
  assign n6716 = n6473 & n6715 ;
  assign n6717 = n6716 ^ n6468 ;
  assign n6713 = x72 & n5121 ;
  assign n6702 = x68 & n5981 ;
  assign n6701 = x70 & n5748 ;
  assign n6703 = n6702 ^ n6701 ;
  assign n6704 = n6703 ^ x47 ;
  assign n6700 = ~n443 & n5749 ;
  assign n6705 = n6704 ^ n6700 ;
  assign n6699 = x69 & n5755 ;
  assign n6706 = n6705 ^ n6699 ;
  assign n6679 = n6468 ^ n6455 ;
  assign n6696 = n6457 ^ n6455 ;
  assign n6697 = n6679 & n6696 ;
  assign n6685 = x50 ^ x48 ;
  assign n6686 = ~n5986 & n6685 ;
  assign n6687 = n6443 & n6686 ;
  assign n6688 = x65 & n6687 ;
  assign n6684 = x67 & n6444 ;
  assign n6689 = n6688 ^ n6684 ;
  assign n6690 = n6689 ^ x50 ;
  assign n6683 = ~n295 & n6445 ;
  assign n6691 = n6690 ^ n6683 ;
  assign n6682 = x66 & n6449 ;
  assign n6692 = n6691 ^ n6682 ;
  assign n6680 = x51 ^ x50 ;
  assign n6681 = x64 & n6680 ;
  assign n6693 = n6692 ^ n6681 ;
  assign n6694 = n6693 ^ n6457 ;
  assign n6698 = n6697 ^ n6694 ;
  assign n6707 = n6706 ^ n6698 ;
  assign n6678 = n6440 & n6465 ;
  assign n6708 = n6707 ^ n6678 ;
  assign n6709 = n6708 ^ x44 ;
  assign n6677 = x71 & n5113 ;
  assign n6710 = n6709 ^ n6677 ;
  assign n6676 = x73 & n5116 ;
  assign n6711 = n6710 ^ n6676 ;
  assign n6675 = n636 & n5117 ;
  assign n6712 = n6711 ^ n6675 ;
  assign n6714 = n6713 ^ n6712 ;
  assign n6718 = n6717 ^ n6714 ;
  assign n6719 = n6718 ^ x41 ;
  assign n6674 = x74 & n4482 ;
  assign n6720 = n6719 ^ n6674 ;
  assign n6673 = x76 & n4478 ;
  assign n6721 = n6720 ^ n6673 ;
  assign n6672 = ~n863 & n4479 ;
  assign n6722 = n6721 ^ n6672 ;
  assign n6724 = n6723 ^ n6722 ;
  assign n6669 = n6482 ^ n6432 ;
  assign n6670 = n6437 & n6669 ;
  assign n6671 = n6670 ^ n6432 ;
  assign n6725 = n6724 ^ n6671 ;
  assign n6659 = x77 & n3932 ;
  assign n6658 = x79 & n3935 ;
  assign n6660 = n6659 ^ n6658 ;
  assign n6661 = n6660 ^ x38 ;
  assign n6657 = n1123 & n3936 ;
  assign n6662 = n6661 ^ n6657 ;
  assign n6656 = x78 & n3940 ;
  assign n6663 = n6662 ^ n6656 ;
  assign n6664 = n6663 ^ n6492 ;
  assign n6665 = n6664 ^ n6483 ;
  assign n6666 = n6665 ^ n6663 ;
  assign n6667 = ~n6489 & n6666 ;
  assign n6668 = n6667 ^ n6664 ;
  assign n6726 = n6725 ^ n6668 ;
  assign n6727 = n6726 ^ x35 ;
  assign n6655 = x80 & n3387 ;
  assign n6728 = n6727 ^ n6655 ;
  assign n6654 = x82 & n3390 ;
  assign n6729 = n6728 ^ n6654 ;
  assign n6653 = n1422 & n3391 ;
  assign n6730 = n6729 ^ n6653 ;
  assign n6732 = n6731 ^ n6730 ;
  assign n6736 = n6735 ^ n6732 ;
  assign n6741 = n6740 ^ n6736 ;
  assign n6743 = n6742 ^ n6741 ;
  assign n6745 = n6744 ^ n6743 ;
  assign n6650 = n6512 ^ n6508 ;
  assign n6651 = n6509 & ~n6650 ;
  assign n6652 = n6651 ^ n6512 ;
  assign n6746 = n6745 ^ n6652 ;
  assign n6747 = n6746 ^ x29 ;
  assign n6649 = x86 & n2593 ;
  assign n6748 = n6747 ^ n6649 ;
  assign n6648 = x88 & n2428 ;
  assign n6749 = n6748 ^ n6648 ;
  assign n6647 = n2131 & n2429 ;
  assign n6750 = n6749 ^ n6647 ;
  assign n6752 = n6751 ^ n6750 ;
  assign n6756 = n6755 ^ n6752 ;
  assign n6757 = n6756 ^ x26 ;
  assign n6646 = x89 & n2032 ;
  assign n6758 = n6757 ^ n6646 ;
  assign n6645 = x91 & n2028 ;
  assign n6759 = n6758 ^ n6645 ;
  assign n6644 = n2029 & n2548 ;
  assign n6760 = n6759 ^ n6644 ;
  assign n6762 = n6761 ^ n6760 ;
  assign n6766 = n6765 ^ n6762 ;
  assign n6767 = n6766 ^ x23 ;
  assign n6643 = x92 & n1665 ;
  assign n6768 = n6767 ^ n6643 ;
  assign n6642 = x94 & n1668 ;
  assign n6769 = n6768 ^ n6642 ;
  assign n6641 = n1669 & n3010 ;
  assign n6770 = n6769 ^ n6641 ;
  assign n6772 = n6771 ^ n6770 ;
  assign n6776 = n6775 ^ n6772 ;
  assign n6777 = n6776 ^ x20 ;
  assign n6640 = x95 & n1340 ;
  assign n6778 = n6777 ^ n6640 ;
  assign n6639 = x97 & n1343 ;
  assign n6779 = n6778 ^ n6639 ;
  assign n6638 = n1344 & n3501 ;
  assign n6780 = n6779 ^ n6638 ;
  assign n6782 = n6781 ^ n6780 ;
  assign n6635 = n6543 ^ n6534 ;
  assign n6636 = n6540 & n6635 ;
  assign n6637 = n6636 ^ n6543 ;
  assign n6783 = n6782 ^ n6637 ;
  assign n6784 = n6783 ^ x17 ;
  assign n6634 = x98 & n1060 ;
  assign n6785 = n6784 ^ n6634 ;
  assign n6633 = x100 & n1063 ;
  assign n6786 = n6785 ^ n6633 ;
  assign n6632 = n1064 & n4048 ;
  assign n6787 = n6786 ^ n6632 ;
  assign n6789 = n6788 ^ n6787 ;
  assign n6793 = n6792 ^ n6789 ;
  assign n6794 = n6793 ^ x14 ;
  assign n6631 = x101 & n884 ;
  assign n6795 = n6794 ^ n6631 ;
  assign n6630 = x103 & n789 ;
  assign n6796 = n6795 ^ n6630 ;
  assign n6629 = n790 & ~n4624 ;
  assign n6797 = n6796 ^ n6629 ;
  assign n6799 = n6798 ^ n6797 ;
  assign n6803 = n6802 ^ n6799 ;
  assign n6804 = n6803 ^ x11 ;
  assign n6628 = x104 & n650 ;
  assign n6805 = n6804 ^ n6628 ;
  assign n6627 = x106 & ~n578 ;
  assign n6806 = n6805 ^ n6627 ;
  assign n6626 = ~n579 & ~n5257 ;
  assign n6807 = n6806 ^ n6626 ;
  assign n6809 = n6808 ^ n6807 ;
  assign n6623 = n6567 ^ n6558 ;
  assign n6624 = ~n6564 & n6623 ;
  assign n6625 = n6624 ^ n6567 ;
  assign n6810 = n6809 ^ n6625 ;
  assign n6811 = n6810 ^ x8 ;
  assign n6622 = x107 & n456 ;
  assign n6812 = n6811 ^ n6622 ;
  assign n6621 = x109 & n384 ;
  assign n6813 = n6812 ^ n6621 ;
  assign n6620 = n385 & n5912 ;
  assign n6814 = n6813 ^ n6620 ;
  assign n6816 = n6815 ^ n6814 ;
  assign n6820 = n6819 ^ n6816 ;
  assign n6821 = n6820 ^ x5 ;
  assign n6619 = x110 & n238 ;
  assign n6822 = n6821 ^ n6619 ;
  assign n6618 = x112 & n234 ;
  assign n6823 = n6822 ^ n6618 ;
  assign n6616 = n5898 ^ x112 ;
  assign n6617 = n235 & ~n6616 ;
  assign n6824 = n6823 ^ n6617 ;
  assign n6826 = n6825 ^ n6824 ;
  assign n6613 = n6584 ^ n6575 ;
  assign n6614 = n6581 & ~n6613 ;
  assign n6615 = n6614 ^ n6584 ;
  assign n6827 = n6826 ^ n6615 ;
  assign n6598 = x114 & ~n6355 ;
  assign n6597 = ~x114 & ~n6354 ;
  assign n6599 = n6598 ^ n6597 ;
  assign n6601 = x115 ^ x1 ;
  assign n6600 = x115 ^ x2 ;
  assign n6602 = n6601 ^ n6600 ;
  assign n6603 = n6599 & n6602 ;
  assign n6604 = n6603 ^ n6601 ;
  assign n6828 = n6827 ^ n6604 ;
  assign n6608 = x2 & x113 ;
  assign n6609 = n6608 ^ x114 ;
  assign n6610 = ~x1 & n6609 ;
  assign n6605 = n6604 ^ n6357 ;
  assign n6611 = n6610 ^ n6605 ;
  assign n6612 = ~x0 & n6611 ;
  assign n6829 = n6828 ^ n6612 ;
  assign n6592 = n6590 ^ n6585 ;
  assign n6593 = n6587 & n6592 ;
  assign n6594 = n6593 ^ n6590 ;
  assign n6830 = n6829 ^ n6594 ;
  assign n7080 = n6827 ^ n6594 ;
  assign n7081 = ~n6829 & n7080 ;
  assign n7082 = n7081 ^ n6827 ;
  assign n7074 = n6820 ^ n6615 ;
  assign n7075 = ~n6826 & ~n7074 ;
  assign n7076 = n7075 ^ n6820 ;
  assign n7072 = x112 & n231 ;
  assign n7065 = x109 & n391 ;
  assign n7057 = n6803 ^ n6625 ;
  assign n7058 = ~n6809 & ~n7057 ;
  assign n7059 = n7058 ^ n6803 ;
  assign n7055 = x106 & n584 ;
  assign n7048 = x103 & n795 ;
  assign n7041 = x100 & n1068 ;
  assign n7033 = n6776 ^ n6637 ;
  assign n7034 = n6782 & ~n7033 ;
  assign n7035 = n7034 ^ n6776 ;
  assign n7031 = x97 & n1348 ;
  assign n7024 = x94 & n1673 ;
  assign n7017 = x91 & n2025 ;
  assign n7010 = x88 & n2435 ;
  assign n7002 = n6736 ^ n6652 ;
  assign n7003 = n6745 & ~n7002 ;
  assign n7004 = n7003 ^ n6736 ;
  assign n6996 = x84 & n2890 ;
  assign n6995 = x86 & n2893 ;
  assign n6997 = n6996 ^ n6995 ;
  assign n6998 = n6997 ^ x32 ;
  assign n6994 = n1868 & n2894 ;
  assign n6999 = n6998 ^ n6994 ;
  assign n6993 = x85 & n2899 ;
  assign n7000 = n6999 ^ n6993 ;
  assign n6990 = x82 & n3395 ;
  assign n6983 = x79 & n3940 ;
  assign n6975 = x73 & n5121 ;
  assign n6964 = x66 & n6687 ;
  assign n6963 = x68 & n6444 ;
  assign n6965 = n6964 ^ n6963 ;
  assign n6966 = n6965 ^ x50 ;
  assign n6962 = ~n351 & n6445 ;
  assign n6967 = n6966 ^ n6962 ;
  assign n6961 = x67 & n6449 ;
  assign n6968 = n6967 ^ n6961 ;
  assign n6955 = x50 & x51 ;
  assign n6956 = n6955 ^ x52 ;
  assign n6957 = ~x64 & n6956 ;
  assign n6951 = x52 ^ x50 ;
  assign n6958 = n6957 ^ n6951 ;
  assign n6949 = x65 ^ x51 ;
  assign n6950 = n6680 & ~n6949 ;
  assign n6959 = n6958 ^ n6950 ;
  assign n6939 = n6457 & n6693 ;
  assign n6940 = n6455 & n6939 ;
  assign n6941 = n6940 ^ n6693 ;
  assign n6948 = n6692 & ~n6941 ;
  assign n6960 = n6959 ^ n6948 ;
  assign n6969 = n6968 ^ n6960 ;
  assign n6932 = x69 & n5981 ;
  assign n6931 = x71 & n5748 ;
  assign n6933 = n6932 ^ n6931 ;
  assign n6934 = n6933 ^ x47 ;
  assign n6930 = ~n495 & n5749 ;
  assign n6935 = n6934 ^ n6930 ;
  assign n6929 = x70 & n5755 ;
  assign n6936 = n6935 ^ n6929 ;
  assign n6937 = n6936 ^ n6678 ;
  assign n6926 = n6706 ^ n6678 ;
  assign n6927 = n6926 ^ n6693 ;
  assign n6928 = n6698 & n6927 ;
  assign n6938 = n6937 ^ n6928 ;
  assign n6942 = n6941 ^ n6938 ;
  assign n6943 = n6942 ^ n6936 ;
  assign n6944 = n6943 ^ n6941 ;
  assign n6945 = ~n6706 & ~n6928 ;
  assign n6946 = n6944 & n6945 ;
  assign n6947 = n6946 ^ n6942 ;
  assign n6970 = n6969 ^ n6947 ;
  assign n6971 = n6970 ^ x44 ;
  assign n6925 = x72 & n5113 ;
  assign n6972 = n6971 ^ n6925 ;
  assign n6924 = x74 & n5116 ;
  assign n6973 = n6972 ^ n6924 ;
  assign n6923 = n708 & n5117 ;
  assign n6974 = n6973 ^ n6923 ;
  assign n6976 = n6975 ^ n6974 ;
  assign n6920 = n6717 ^ n6708 ;
  assign n6921 = ~n6714 & n6920 ;
  assign n6922 = n6921 ^ n6717 ;
  assign n6977 = n6976 ^ n6922 ;
  assign n6910 = x75 & n4482 ;
  assign n6909 = x77 & n4478 ;
  assign n6911 = n6910 ^ n6909 ;
  assign n6912 = n6911 ^ x41 ;
  assign n6908 = ~n943 & n4479 ;
  assign n6913 = n6912 ^ n6908 ;
  assign n6907 = x76 & n4475 ;
  assign n6914 = n6913 ^ n6907 ;
  assign n6915 = n6914 ^ n6718 ;
  assign n6916 = n6915 ^ n6671 ;
  assign n6917 = n6916 ^ n6914 ;
  assign n6918 = n6724 & n6917 ;
  assign n6919 = n6918 ^ n6915 ;
  assign n6978 = n6977 ^ n6919 ;
  assign n6979 = n6978 ^ x38 ;
  assign n6906 = x78 & n3932 ;
  assign n6980 = n6979 ^ n6906 ;
  assign n6905 = x80 & n3935 ;
  assign n6981 = n6980 ^ n6905 ;
  assign n6904 = n1217 & n3936 ;
  assign n6982 = n6981 ^ n6904 ;
  assign n6984 = n6983 ^ n6982 ;
  assign n6901 = n6725 ^ n6663 ;
  assign n6902 = n6668 & n6901 ;
  assign n6903 = n6902 ^ n6663 ;
  assign n6985 = n6984 ^ n6903 ;
  assign n6986 = n6985 ^ x35 ;
  assign n6900 = x81 & n3387 ;
  assign n6987 = n6986 ^ n6900 ;
  assign n6899 = x83 & n3390 ;
  assign n6988 = n6987 ^ n6899 ;
  assign n6898 = n1517 & n3391 ;
  assign n6989 = n6988 ^ n6898 ;
  assign n6991 = n6990 ^ n6989 ;
  assign n6895 = n6735 ^ n6726 ;
  assign n6896 = ~n6732 & n6895 ;
  assign n6897 = n6896 ^ n6735 ;
  assign n6992 = n6991 ^ n6897 ;
  assign n7001 = n7000 ^ n6992 ;
  assign n7005 = n7004 ^ n7001 ;
  assign n7006 = n7005 ^ x29 ;
  assign n6894 = x87 & n2593 ;
  assign n7007 = n7006 ^ n6894 ;
  assign n6893 = x89 & n2428 ;
  assign n7008 = n7007 ^ n6893 ;
  assign n6892 = n2255 & n2429 ;
  assign n7009 = n7008 ^ n6892 ;
  assign n7011 = n7010 ^ n7009 ;
  assign n6889 = n6755 ^ n6746 ;
  assign n6890 = n6752 & ~n6889 ;
  assign n6891 = n6890 ^ n6755 ;
  assign n7012 = n7011 ^ n6891 ;
  assign n7013 = n7012 ^ x26 ;
  assign n6888 = x90 & n2032 ;
  assign n7014 = n7013 ^ n6888 ;
  assign n6887 = x92 & n2028 ;
  assign n7015 = n7014 ^ n6887 ;
  assign n6886 = n2029 & n2696 ;
  assign n7016 = n7015 ^ n6886 ;
  assign n7018 = n7017 ^ n7016 ;
  assign n6883 = n6765 ^ n6756 ;
  assign n6884 = n6762 & n6883 ;
  assign n6885 = n6884 ^ n6765 ;
  assign n7019 = n7018 ^ n6885 ;
  assign n7020 = n7019 ^ x23 ;
  assign n6882 = x93 & n1665 ;
  assign n7021 = n7020 ^ n6882 ;
  assign n6881 = x95 & n1668 ;
  assign n7022 = n7021 ^ n6881 ;
  assign n6880 = n1669 & n3166 ;
  assign n7023 = n7022 ^ n6880 ;
  assign n7025 = n7024 ^ n7023 ;
  assign n6877 = n6775 ^ n6766 ;
  assign n6878 = ~n6772 & n6877 ;
  assign n6879 = n6878 ^ n6775 ;
  assign n7026 = n7025 ^ n6879 ;
  assign n7027 = n7026 ^ x20 ;
  assign n6876 = x96 & n1340 ;
  assign n7028 = n7027 ^ n6876 ;
  assign n6875 = x98 & n1343 ;
  assign n7029 = n7028 ^ n6875 ;
  assign n6874 = n1344 & n3673 ;
  assign n7030 = n7029 ^ n6874 ;
  assign n7032 = n7031 ^ n7030 ;
  assign n7036 = n7035 ^ n7032 ;
  assign n7037 = n7036 ^ x17 ;
  assign n6873 = x99 & n1060 ;
  assign n7038 = n7037 ^ n6873 ;
  assign n6872 = x101 & n1063 ;
  assign n7039 = n7038 ^ n6872 ;
  assign n6871 = n1064 & n4223 ;
  assign n7040 = n7039 ^ n6871 ;
  assign n7042 = n7041 ^ n7040 ;
  assign n6868 = n6792 ^ n6783 ;
  assign n6869 = n6789 & ~n6868 ;
  assign n6870 = n6869 ^ n6792 ;
  assign n7043 = n7042 ^ n6870 ;
  assign n7044 = n7043 ^ x14 ;
  assign n6867 = x102 & n884 ;
  assign n7045 = n7044 ^ n6867 ;
  assign n6866 = x104 & n789 ;
  assign n7046 = n7045 ^ n6866 ;
  assign n6865 = n790 & ~n4830 ;
  assign n7047 = n7046 ^ n6865 ;
  assign n7049 = n7048 ^ n7047 ;
  assign n6862 = n6802 ^ n6793 ;
  assign n6863 = n6799 & ~n6862 ;
  assign n6864 = n6863 ^ n6802 ;
  assign n7050 = n7049 ^ n6864 ;
  assign n7051 = n7050 ^ x11 ;
  assign n6861 = x105 & n650 ;
  assign n7052 = n7051 ^ n6861 ;
  assign n6860 = x107 & ~n578 ;
  assign n7053 = n7052 ^ n6860 ;
  assign n6859 = ~n579 & ~n5459 ;
  assign n7054 = n7053 ^ n6859 ;
  assign n7056 = n7055 ^ n7054 ;
  assign n7060 = n7059 ^ n7056 ;
  assign n7061 = n7060 ^ x8 ;
  assign n6858 = x108 & n456 ;
  assign n7062 = n7061 ^ n6858 ;
  assign n6857 = x110 & n384 ;
  assign n7063 = n7062 ^ n6857 ;
  assign n6856 = n385 & n6145 ;
  assign n7064 = n7063 ^ n6856 ;
  assign n7066 = n7065 ^ n7064 ;
  assign n6853 = n6819 ^ n6810 ;
  assign n6854 = n6816 & ~n6853 ;
  assign n6855 = n6854 ^ n6819 ;
  assign n7067 = n7066 ^ n6855 ;
  assign n7068 = n7067 ^ x5 ;
  assign n6852 = x111 & n238 ;
  assign n7069 = n7068 ^ n6852 ;
  assign n6851 = x113 & n234 ;
  assign n7070 = n7069 ^ n6851 ;
  assign n6849 = n6128 ^ x113 ;
  assign n6850 = n235 & ~n6849 ;
  assign n7071 = n7070 ^ n6850 ;
  assign n7073 = n7072 ^ n7071 ;
  assign n7077 = n7076 ^ n7073 ;
  assign n6834 = ~x115 & ~n6598 ;
  assign n6833 = x115 & ~n6597 ;
  assign n6835 = n6834 ^ n6833 ;
  assign n6837 = x116 ^ x1 ;
  assign n6836 = x116 ^ x2 ;
  assign n6838 = n6837 ^ n6836 ;
  assign n6839 = n6835 & n6838 ;
  assign n6840 = n6839 ^ n6837 ;
  assign n7078 = n7077 ^ n6840 ;
  assign n6844 = x2 & x114 ;
  assign n6845 = n6844 ^ x115 ;
  assign n6846 = ~n259 & n6845 ;
  assign n6841 = n6840 ^ n6600 ;
  assign n6847 = n6846 ^ n6841 ;
  assign n6848 = ~x0 & n6847 ;
  assign n7079 = n7078 ^ n6848 ;
  assign n7083 = n7082 ^ n7079 ;
  assign n7329 = x113 & n231 ;
  assign n7321 = n7060 ^ n6855 ;
  assign n7322 = n7066 & n7321 ;
  assign n7323 = n7322 ^ n7060 ;
  assign n7319 = x110 & n391 ;
  assign n7312 = x107 & n584 ;
  assign n7304 = n7043 ^ n6864 ;
  assign n7305 = ~n7049 & ~n7304 ;
  assign n7306 = n7305 ^ n7043 ;
  assign n7302 = x104 & n795 ;
  assign n7294 = n7036 ^ n6870 ;
  assign n7295 = ~n7042 & ~n7294 ;
  assign n7296 = n7295 ^ n7036 ;
  assign n7292 = x101 & n1068 ;
  assign n7285 = x98 & n1348 ;
  assign n7277 = n7019 ^ n6879 ;
  assign n7278 = ~n7025 & ~n7277 ;
  assign n7279 = n7278 ^ n7019 ;
  assign n7275 = x95 & n1673 ;
  assign n7267 = n7012 ^ n6885 ;
  assign n7268 = n7018 & ~n7267 ;
  assign n7269 = n7268 ^ n7012 ;
  assign n7265 = x92 & n2025 ;
  assign n7257 = n7005 ^ n6891 ;
  assign n7258 = n7011 & n7257 ;
  assign n7259 = n7258 ^ n7005 ;
  assign n7255 = x89 & n2435 ;
  assign n7248 = x86 & n2899 ;
  assign n7240 = n6985 ^ n6897 ;
  assign n7241 = n6991 & n7240 ;
  assign n7242 = n7241 ^ n6985 ;
  assign n7238 = x83 & n3395 ;
  assign n7228 = x79 & n3932 ;
  assign n7227 = x81 & n3935 ;
  assign n7229 = n7228 ^ n7227 ;
  assign n7230 = n7229 ^ x38 ;
  assign n7226 = n1310 & n3936 ;
  assign n7231 = n7230 ^ n7226 ;
  assign n7225 = x80 & n3940 ;
  assign n7232 = n7231 ^ n7225 ;
  assign n7221 = x77 & n4475 ;
  assign n7214 = x74 & n5121 ;
  assign n7207 = x71 & n5755 ;
  assign n7200 = x68 & n6449 ;
  assign n6953 = x52 ^ x51 ;
  assign n7191 = ~n6680 & n6953 ;
  assign n7192 = x65 & n7191 ;
  assign n7180 = x53 ^ x52 ;
  assign n7186 = n6680 & ~n7180 ;
  assign n7187 = n7186 ^ n6680 ;
  assign n7188 = ~n152 & n7187 ;
  assign n7185 = x66 & n6680 ;
  assign n7189 = n7188 ^ n7185 ;
  assign n7190 = n7189 ^ x53 ;
  assign n7193 = n7192 ^ n7190 ;
  assign n7181 = x53 ^ x51 ;
  assign n7182 = ~n6680 & n7181 ;
  assign n7183 = n7180 & n7182 ;
  assign n7184 = x64 & n7183 ;
  assign n7194 = n7193 ^ n7184 ;
  assign n7178 = ~n6681 & ~n6959 ;
  assign n7179 = x53 & n7178 ;
  assign n7195 = n7194 ^ n7179 ;
  assign n7196 = n7195 ^ x50 ;
  assign n7177 = x67 & n6687 ;
  assign n7197 = n7196 ^ n7177 ;
  assign n7176 = x69 & n6444 ;
  assign n7198 = n7197 ^ n7176 ;
  assign n7175 = ~n376 & n6445 ;
  assign n7199 = n7198 ^ n7175 ;
  assign n7201 = n7200 ^ n7199 ;
  assign n7172 = n6968 ^ n6959 ;
  assign n7173 = ~n6960 & n7172 ;
  assign n7174 = n7173 ^ n6968 ;
  assign n7202 = n7201 ^ n7174 ;
  assign n7203 = n7202 ^ x47 ;
  assign n7171 = x70 & n5981 ;
  assign n7204 = n7203 ^ n7171 ;
  assign n7170 = x72 & n5748 ;
  assign n7205 = n7204 ^ n7170 ;
  assign n7169 = n565 & n5749 ;
  assign n7206 = n7205 ^ n7169 ;
  assign n7208 = n7207 ^ n7206 ;
  assign n7166 = n6969 ^ n6936 ;
  assign n7167 = n6947 & n7166 ;
  assign n7168 = n7167 ^ n6936 ;
  assign n7209 = n7208 ^ n7168 ;
  assign n7210 = n7209 ^ x44 ;
  assign n7165 = x73 & n5113 ;
  assign n7211 = n7210 ^ n7165 ;
  assign n7164 = x75 & n5116 ;
  assign n7212 = n7211 ^ n7164 ;
  assign n7163 = ~n778 & n5117 ;
  assign n7213 = n7212 ^ n7163 ;
  assign n7215 = n7214 ^ n7213 ;
  assign n7160 = n6970 ^ n6922 ;
  assign n7161 = n6976 & n7160 ;
  assign n7162 = n7161 ^ n6970 ;
  assign n7216 = n7215 ^ n7162 ;
  assign n7217 = n7216 ^ x41 ;
  assign n7159 = x76 & n4482 ;
  assign n7218 = n7217 ^ n7159 ;
  assign n7158 = x78 & n4478 ;
  assign n7219 = n7218 ^ n7158 ;
  assign n7157 = ~n1036 & n4479 ;
  assign n7220 = n7219 ^ n7157 ;
  assign n7222 = n7221 ^ n7220 ;
  assign n7154 = n6977 ^ n6914 ;
  assign n7155 = n6919 & n7154 ;
  assign n7156 = n7155 ^ n6914 ;
  assign n7223 = n7222 ^ n7156 ;
  assign n7151 = n6978 ^ n6903 ;
  assign n7152 = n6984 & n7151 ;
  assign n7153 = n7152 ^ n6978 ;
  assign n7224 = n7223 ^ n7153 ;
  assign n7233 = n7232 ^ n7224 ;
  assign n7234 = n7233 ^ x35 ;
  assign n7150 = x82 & n3387 ;
  assign n7235 = n7234 ^ n7150 ;
  assign n7149 = x84 & n3390 ;
  assign n7236 = n7235 ^ n7149 ;
  assign n7148 = n1635 & n3391 ;
  assign n7237 = n7236 ^ n7148 ;
  assign n7239 = n7238 ^ n7237 ;
  assign n7243 = n7242 ^ n7239 ;
  assign n7244 = n7243 ^ x32 ;
  assign n7147 = x85 & n2890 ;
  assign n7245 = n7244 ^ n7147 ;
  assign n7146 = x87 & n2893 ;
  assign n7246 = n7245 ^ n7146 ;
  assign n7145 = n1987 & n2894 ;
  assign n7247 = n7246 ^ n7145 ;
  assign n7249 = n7248 ^ n7247 ;
  assign n7142 = n7004 ^ n7000 ;
  assign n7143 = ~n7001 & n7142 ;
  assign n7144 = n7143 ^ n7004 ;
  assign n7250 = n7249 ^ n7144 ;
  assign n7251 = n7250 ^ x29 ;
  assign n7141 = x88 & n2593 ;
  assign n7252 = n7251 ^ n7141 ;
  assign n7140 = x90 & n2428 ;
  assign n7253 = n7252 ^ n7140 ;
  assign n7139 = n2398 & n2429 ;
  assign n7254 = n7253 ^ n7139 ;
  assign n7256 = n7255 ^ n7254 ;
  assign n7260 = n7259 ^ n7256 ;
  assign n7261 = n7260 ^ x26 ;
  assign n7138 = x91 & n2032 ;
  assign n7262 = n7261 ^ n7138 ;
  assign n7137 = x93 & n2028 ;
  assign n7263 = n7262 ^ n7137 ;
  assign n7136 = n2029 & n2842 ;
  assign n7264 = n7263 ^ n7136 ;
  assign n7266 = n7265 ^ n7264 ;
  assign n7270 = n7269 ^ n7266 ;
  assign n7271 = n7270 ^ x23 ;
  assign n7135 = x94 & n1665 ;
  assign n7272 = n7271 ^ n7135 ;
  assign n7134 = x96 & n1668 ;
  assign n7273 = n7272 ^ n7134 ;
  assign n7133 = n1669 & n3336 ;
  assign n7274 = n7273 ^ n7133 ;
  assign n7276 = n7275 ^ n7274 ;
  assign n7280 = n7279 ^ n7276 ;
  assign n7281 = n7280 ^ x20 ;
  assign n7132 = x97 & n1340 ;
  assign n7282 = n7281 ^ n7132 ;
  assign n7131 = x99 & n1343 ;
  assign n7283 = n7282 ^ n7131 ;
  assign n7130 = n1344 & n3851 ;
  assign n7284 = n7283 ^ n7130 ;
  assign n7286 = n7285 ^ n7284 ;
  assign n7127 = n7035 ^ n7026 ;
  assign n7128 = n7032 & ~n7127 ;
  assign n7129 = n7128 ^ n7035 ;
  assign n7287 = n7286 ^ n7129 ;
  assign n7288 = n7287 ^ x17 ;
  assign n7126 = x100 & n1060 ;
  assign n7289 = n7288 ^ n7126 ;
  assign n7125 = x102 & n1063 ;
  assign n7290 = n7289 ^ n7125 ;
  assign n7124 = n1064 & n4425 ;
  assign n7291 = n7290 ^ n7124 ;
  assign n7293 = n7292 ^ n7291 ;
  assign n7297 = n7296 ^ n7293 ;
  assign n7298 = n7297 ^ x14 ;
  assign n7123 = x103 & n884 ;
  assign n7299 = n7298 ^ n7123 ;
  assign n7122 = x105 & n789 ;
  assign n7300 = n7299 ^ n7122 ;
  assign n7121 = n790 & ~n5034 ;
  assign n7301 = n7300 ^ n7121 ;
  assign n7303 = n7302 ^ n7301 ;
  assign n7307 = n7306 ^ n7303 ;
  assign n7308 = n7307 ^ x11 ;
  assign n7120 = x106 & n650 ;
  assign n7309 = n7308 ^ n7120 ;
  assign n7119 = x108 & ~n578 ;
  assign n7310 = n7309 ^ n7119 ;
  assign n7118 = ~n579 & n5687 ;
  assign n7311 = n7310 ^ n7118 ;
  assign n7313 = n7312 ^ n7311 ;
  assign n7115 = n7059 ^ n7050 ;
  assign n7116 = n7056 & n7115 ;
  assign n7117 = n7116 ^ n7059 ;
  assign n7314 = n7313 ^ n7117 ;
  assign n7315 = n7314 ^ x8 ;
  assign n7114 = x109 & n456 ;
  assign n7316 = n7315 ^ n7114 ;
  assign n7113 = x111 & n384 ;
  assign n7317 = n7316 ^ n7113 ;
  assign n7112 = n385 & ~n6370 ;
  assign n7318 = n7317 ^ n7112 ;
  assign n7320 = n7319 ^ n7318 ;
  assign n7324 = n7323 ^ n7320 ;
  assign n7325 = n7324 ^ x5 ;
  assign n7111 = x112 & n238 ;
  assign n7326 = n7325 ^ n7111 ;
  assign n7110 = x114 & n234 ;
  assign n7327 = n7326 ^ n7110 ;
  assign n7108 = n6356 ^ x114 ;
  assign n7109 = n235 & ~n7108 ;
  assign n7328 = n7327 ^ n7109 ;
  assign n7330 = n7329 ^ n7328 ;
  assign n7105 = n7076 ^ n7067 ;
  assign n7106 = ~n7073 & ~n7105 ;
  assign n7107 = n7106 ^ n7076 ;
  assign n7331 = n7330 ^ n7107 ;
  assign n7090 = x116 & ~n6834 ;
  assign n7089 = ~x116 & ~n6833 ;
  assign n7091 = n7090 ^ n7089 ;
  assign n7093 = x117 ^ x1 ;
  assign n7092 = x117 ^ x2 ;
  assign n7094 = n7093 ^ n7092 ;
  assign n7095 = n7091 & n7094 ;
  assign n7096 = n7095 ^ n7093 ;
  assign n7332 = n7331 ^ n7096 ;
  assign n7100 = x2 & x115 ;
  assign n7101 = n7100 ^ x116 ;
  assign n7102 = ~n259 & n7101 ;
  assign n7097 = n7096 ^ n6836 ;
  assign n7103 = n7102 ^ n7097 ;
  assign n7104 = ~x0 & n7103 ;
  assign n7333 = n7332 ^ n7104 ;
  assign n7084 = n7082 ^ n7077 ;
  assign n7085 = n7079 & n7084 ;
  assign n7086 = n7085 ^ n7082 ;
  assign n7334 = n7333 ^ n7086 ;
  assign n7578 = n7331 ^ n7086 ;
  assign n7579 = ~n7333 & n7578 ;
  assign n7580 = n7579 ^ n7331 ;
  assign n7572 = n7324 ^ n7107 ;
  assign n7573 = n7330 & ~n7572 ;
  assign n7574 = n7573 ^ n7324 ;
  assign n7570 = x114 & n231 ;
  assign n7563 = x111 & n391 ;
  assign n7555 = n7307 ^ n7117 ;
  assign n7556 = ~n7313 & n7555 ;
  assign n7557 = n7556 ^ n7307 ;
  assign n7549 = x107 & n650 ;
  assign n7548 = x109 & ~n578 ;
  assign n7550 = n7549 ^ n7548 ;
  assign n7551 = n7550 ^ x11 ;
  assign n7547 = ~n579 & n5912 ;
  assign n7552 = n7551 ^ n7547 ;
  assign n7546 = x108 & n584 ;
  assign n7553 = n7552 ^ n7546 ;
  assign n7543 = x105 & n795 ;
  assign n7536 = x102 & n1068 ;
  assign n7528 = n7280 ^ n7129 ;
  assign n7529 = ~n7286 & ~n7528 ;
  assign n7530 = n7529 ^ n7280 ;
  assign n7526 = x99 & n1348 ;
  assign n7519 = x96 & n1673 ;
  assign n7512 = x93 & n2025 ;
  assign n7505 = x90 & n2435 ;
  assign n7497 = n7243 ^ n7144 ;
  assign n7498 = n7249 & n7497 ;
  assign n7499 = n7498 ^ n7243 ;
  assign n7495 = x87 & n2899 ;
  assign n7488 = x84 & n3395 ;
  assign n7481 = x81 & n3940 ;
  assign n7473 = x75 & n5121 ;
  assign n7466 = x72 & n5755 ;
  assign n7458 = n7195 ^ n7174 ;
  assign n7459 = n7201 & n7458 ;
  assign n7460 = n7459 ^ n7195 ;
  assign n7456 = x69 & n6449 ;
  assign n7445 = x65 & n7183 ;
  assign n7444 = x67 & n7186 ;
  assign n7446 = n7445 ^ n7444 ;
  assign n7447 = n7446 ^ x53 ;
  assign n7443 = ~n295 & n7187 ;
  assign n7448 = n7447 ^ n7443 ;
  assign n7442 = x66 & n7191 ;
  assign n7449 = n7448 ^ n7442 ;
  assign n7440 = x54 ^ x53 ;
  assign n7441 = x64 & n7440 ;
  assign n7450 = n7449 ^ n7441 ;
  assign n7439 = n7179 & n7194 ;
  assign n7451 = n7450 ^ n7439 ;
  assign n7452 = n7451 ^ x50 ;
  assign n7438 = x68 & n6687 ;
  assign n7453 = n7452 ^ n7438 ;
  assign n7437 = x70 & n6444 ;
  assign n7454 = n7453 ^ n7437 ;
  assign n7436 = ~n443 & n6445 ;
  assign n7455 = n7454 ^ n7436 ;
  assign n7457 = n7456 ^ n7455 ;
  assign n7461 = n7460 ^ n7457 ;
  assign n7462 = n7461 ^ x47 ;
  assign n7435 = x71 & n5981 ;
  assign n7463 = n7462 ^ n7435 ;
  assign n7434 = x73 & n5748 ;
  assign n7464 = n7463 ^ n7434 ;
  assign n7433 = n636 & n5749 ;
  assign n7465 = n7464 ^ n7433 ;
  assign n7467 = n7466 ^ n7465 ;
  assign n7430 = n7202 ^ n7168 ;
  assign n7431 = n7208 & n7430 ;
  assign n7432 = n7431 ^ n7202 ;
  assign n7468 = n7467 ^ n7432 ;
  assign n7469 = n7468 ^ x44 ;
  assign n7429 = x74 & n5113 ;
  assign n7470 = n7469 ^ n7429 ;
  assign n7428 = x76 & n5116 ;
  assign n7471 = n7470 ^ n7428 ;
  assign n7427 = ~n863 & n5117 ;
  assign n7472 = n7471 ^ n7427 ;
  assign n7474 = n7473 ^ n7472 ;
  assign n7424 = n7209 ^ n7162 ;
  assign n7425 = n7215 & n7424 ;
  assign n7426 = n7425 ^ n7209 ;
  assign n7475 = n7474 ^ n7426 ;
  assign n7414 = x77 & n4482 ;
  assign n7413 = x79 & n4478 ;
  assign n7415 = n7414 ^ n7413 ;
  assign n7416 = n7415 ^ x41 ;
  assign n7412 = n1123 & n4479 ;
  assign n7417 = n7416 ^ n7412 ;
  assign n7411 = x78 & n4475 ;
  assign n7418 = n7417 ^ n7411 ;
  assign n7419 = n7418 ^ n7216 ;
  assign n7420 = n7419 ^ n7156 ;
  assign n7421 = n7420 ^ n7418 ;
  assign n7422 = n7222 & n7421 ;
  assign n7423 = n7422 ^ n7419 ;
  assign n7476 = n7475 ^ n7423 ;
  assign n7477 = n7476 ^ x38 ;
  assign n7410 = x80 & n3932 ;
  assign n7478 = n7477 ^ n7410 ;
  assign n7409 = x82 & n3935 ;
  assign n7479 = n7478 ^ n7409 ;
  assign n7408 = n1422 & n3936 ;
  assign n7480 = n7479 ^ n7408 ;
  assign n7482 = n7481 ^ n7480 ;
  assign n7405 = n7232 ^ n7153 ;
  assign n7406 = ~n7224 & n7405 ;
  assign n7407 = n7406 ^ n7232 ;
  assign n7483 = n7482 ^ n7407 ;
  assign n7484 = n7483 ^ x35 ;
  assign n7404 = x83 & n3387 ;
  assign n7485 = n7484 ^ n7404 ;
  assign n7403 = x85 & n3390 ;
  assign n7486 = n7485 ^ n7403 ;
  assign n7402 = n1748 & n3391 ;
  assign n7487 = n7486 ^ n7402 ;
  assign n7489 = n7488 ^ n7487 ;
  assign n7399 = n7242 ^ n7233 ;
  assign n7400 = ~n7239 & n7399 ;
  assign n7401 = n7400 ^ n7242 ;
  assign n7490 = n7489 ^ n7401 ;
  assign n7491 = n7490 ^ x32 ;
  assign n7398 = x86 & n2890 ;
  assign n7492 = n7491 ^ n7398 ;
  assign n7397 = x88 & n2893 ;
  assign n7493 = n7492 ^ n7397 ;
  assign n7396 = n2131 & n2894 ;
  assign n7494 = n7493 ^ n7396 ;
  assign n7496 = n7495 ^ n7494 ;
  assign n7500 = n7499 ^ n7496 ;
  assign n7501 = n7500 ^ x29 ;
  assign n7395 = x89 & n2593 ;
  assign n7502 = n7501 ^ n7395 ;
  assign n7394 = x91 & n2428 ;
  assign n7503 = n7502 ^ n7394 ;
  assign n7393 = n2429 & n2548 ;
  assign n7504 = n7503 ^ n7393 ;
  assign n7506 = n7505 ^ n7504 ;
  assign n7390 = n7259 ^ n7250 ;
  assign n7391 = ~n7256 & n7390 ;
  assign n7392 = n7391 ^ n7259 ;
  assign n7507 = n7506 ^ n7392 ;
  assign n7508 = n7507 ^ x26 ;
  assign n7389 = x92 & n2032 ;
  assign n7509 = n7508 ^ n7389 ;
  assign n7388 = x94 & n2028 ;
  assign n7510 = n7509 ^ n7388 ;
  assign n7387 = n2029 & n3010 ;
  assign n7511 = n7510 ^ n7387 ;
  assign n7513 = n7512 ^ n7511 ;
  assign n7384 = n7269 ^ n7260 ;
  assign n7385 = ~n7266 & n7384 ;
  assign n7386 = n7385 ^ n7269 ;
  assign n7514 = n7513 ^ n7386 ;
  assign n7515 = n7514 ^ x23 ;
  assign n7383 = x95 & n1665 ;
  assign n7516 = n7515 ^ n7383 ;
  assign n7382 = x97 & n1668 ;
  assign n7517 = n7516 ^ n7382 ;
  assign n7381 = n1669 & n3501 ;
  assign n7518 = n7517 ^ n7381 ;
  assign n7520 = n7519 ^ n7518 ;
  assign n7378 = n7279 ^ n7270 ;
  assign n7379 = ~n7276 & ~n7378 ;
  assign n7380 = n7379 ^ n7279 ;
  assign n7521 = n7520 ^ n7380 ;
  assign n7522 = n7521 ^ x20 ;
  assign n7377 = x98 & n1340 ;
  assign n7523 = n7522 ^ n7377 ;
  assign n7376 = x100 & n1343 ;
  assign n7524 = n7523 ^ n7376 ;
  assign n7375 = n1344 & n4048 ;
  assign n7525 = n7524 ^ n7375 ;
  assign n7527 = n7526 ^ n7525 ;
  assign n7531 = n7530 ^ n7527 ;
  assign n7532 = n7531 ^ x17 ;
  assign n7374 = x101 & n1060 ;
  assign n7533 = n7532 ^ n7374 ;
  assign n7373 = x103 & n1063 ;
  assign n7534 = n7533 ^ n7373 ;
  assign n7372 = n1064 & ~n4624 ;
  assign n7535 = n7534 ^ n7372 ;
  assign n7537 = n7536 ^ n7535 ;
  assign n7369 = n7296 ^ n7287 ;
  assign n7370 = n7293 & n7369 ;
  assign n7371 = n7370 ^ n7296 ;
  assign n7538 = n7537 ^ n7371 ;
  assign n7539 = n7538 ^ x14 ;
  assign n7368 = x104 & n884 ;
  assign n7540 = n7539 ^ n7368 ;
  assign n7367 = x106 & n789 ;
  assign n7541 = n7540 ^ n7367 ;
  assign n7366 = n790 & ~n5257 ;
  assign n7542 = n7541 ^ n7366 ;
  assign n7544 = n7543 ^ n7542 ;
  assign n7363 = n7306 ^ n7297 ;
  assign n7364 = ~n7303 & ~n7363 ;
  assign n7365 = n7364 ^ n7306 ;
  assign n7545 = n7544 ^ n7365 ;
  assign n7554 = n7553 ^ n7545 ;
  assign n7558 = n7557 ^ n7554 ;
  assign n7559 = n7558 ^ x8 ;
  assign n7362 = x110 & n456 ;
  assign n7560 = n7559 ^ n7362 ;
  assign n7361 = x112 & n384 ;
  assign n7561 = n7560 ^ n7361 ;
  assign n7360 = n385 & ~n6616 ;
  assign n7562 = n7561 ^ n7360 ;
  assign n7564 = n7563 ^ n7562 ;
  assign n7357 = n7323 ^ n7314 ;
  assign n7358 = ~n7320 & n7357 ;
  assign n7359 = n7358 ^ n7323 ;
  assign n7565 = n7564 ^ n7359 ;
  assign n7566 = n7565 ^ x5 ;
  assign n7356 = x113 & n238 ;
  assign n7567 = n7566 ^ n7356 ;
  assign n7355 = x115 & n234 ;
  assign n7568 = n7567 ^ n7355 ;
  assign n7353 = n6599 ^ x115 ;
  assign n7354 = n235 & ~n7353 ;
  assign n7569 = n7568 ^ n7354 ;
  assign n7571 = n7570 ^ n7569 ;
  assign n7575 = n7574 ^ n7571 ;
  assign n7338 = ~x117 & ~n7090 ;
  assign n7337 = x117 & ~n7089 ;
  assign n7339 = n7338 ^ n7337 ;
  assign n7341 = x118 ^ x1 ;
  assign n7340 = x118 ^ x2 ;
  assign n7342 = n7341 ^ n7340 ;
  assign n7343 = n7339 & n7342 ;
  assign n7344 = n7343 ^ n7341 ;
  assign n7576 = n7575 ^ n7344 ;
  assign n7348 = x2 & x116 ;
  assign n7349 = n7348 ^ x117 ;
  assign n7350 = ~x1 & n7349 ;
  assign n7345 = n7344 ^ n7092 ;
  assign n7351 = n7350 ^ n7345 ;
  assign n7352 = ~x0 & n7351 ;
  assign n7577 = n7576 ^ n7352 ;
  assign n7581 = n7580 ^ n7577 ;
  assign n7832 = x115 & n231 ;
  assign n7824 = n7558 ^ n7359 ;
  assign n7825 = ~n7564 & ~n7824 ;
  assign n7826 = n7825 ^ n7558 ;
  assign n7822 = x112 & n391 ;
  assign n7815 = x109 & n584 ;
  assign n7807 = n7538 ^ n7365 ;
  assign n7808 = ~n7544 & n7807 ;
  assign n7809 = n7808 ^ n7538 ;
  assign n7805 = x106 & n795 ;
  assign n7797 = n7531 ^ n7371 ;
  assign n7798 = n7537 & ~n7797 ;
  assign n7799 = n7798 ^ n7531 ;
  assign n7795 = x103 & n1068 ;
  assign n7788 = x100 & n1348 ;
  assign n7780 = n7514 ^ n7380 ;
  assign n7781 = n7520 & ~n7780 ;
  assign n7782 = n7781 ^ n7514 ;
  assign n7778 = x97 & n1673 ;
  assign n7770 = n7507 ^ n7386 ;
  assign n7771 = n7513 & n7770 ;
  assign n7772 = n7771 ^ n7507 ;
  assign n7768 = x94 & n2025 ;
  assign n7760 = n7500 ^ n7392 ;
  assign n7761 = n7506 & n7760 ;
  assign n7762 = n7761 ^ n7500 ;
  assign n7758 = x91 & n2435 ;
  assign n7751 = x88 & n2899 ;
  assign n7743 = n7483 ^ n7401 ;
  assign n7744 = n7489 & n7743 ;
  assign n7745 = n7744 ^ n7483 ;
  assign n7741 = x85 & n3395 ;
  assign n7734 = x82 & n3940 ;
  assign n7727 = x79 & n4475 ;
  assign n7718 = n7461 ^ n7432 ;
  assign n7719 = n7467 & n7718 ;
  assign n7720 = n7719 ^ n7461 ;
  assign n7716 = x73 & n5755 ;
  assign n7709 = x70 & n6449 ;
  assign n7698 = x66 & n7183 ;
  assign n7697 = x68 & n7186 ;
  assign n7699 = n7698 ^ n7697 ;
  assign n7700 = n7699 ^ x53 ;
  assign n7696 = ~n351 & n7187 ;
  assign n7701 = n7700 ^ n7696 ;
  assign n7695 = x67 & n7191 ;
  assign n7702 = n7701 ^ n7695 ;
  assign n7692 = x65 ^ x54 ;
  assign n7693 = n7440 & ~n7692 ;
  assign n7688 = x53 & x54 ;
  assign n7689 = n7688 ^ x55 ;
  assign n7690 = ~x64 & n7689 ;
  assign n7684 = x55 ^ x53 ;
  assign n7691 = n7690 ^ n7684 ;
  assign n7694 = n7693 ^ n7691 ;
  assign n7703 = n7702 ^ n7694 ;
  assign n7681 = ~n7441 & n7449 ;
  assign n7682 = ~n7439 & n7681 ;
  assign n7683 = n7682 ^ n7449 ;
  assign n7704 = n7703 ^ n7683 ;
  assign n7705 = n7704 ^ x50 ;
  assign n7680 = x69 & n6687 ;
  assign n7706 = n7705 ^ n7680 ;
  assign n7679 = x71 & n6444 ;
  assign n7707 = n7706 ^ n7679 ;
  assign n7678 = ~n495 & n6445 ;
  assign n7708 = n7707 ^ n7678 ;
  assign n7710 = n7709 ^ n7708 ;
  assign n7675 = n7460 ^ n7451 ;
  assign n7676 = ~n7457 & n7675 ;
  assign n7677 = n7676 ^ n7460 ;
  assign n7711 = n7710 ^ n7677 ;
  assign n7712 = n7711 ^ x47 ;
  assign n7674 = x72 & n5981 ;
  assign n7713 = n7712 ^ n7674 ;
  assign n7673 = x74 & n5748 ;
  assign n7714 = n7713 ^ n7673 ;
  assign n7672 = n708 & n5749 ;
  assign n7715 = n7714 ^ n7672 ;
  assign n7717 = n7716 ^ n7715 ;
  assign n7721 = n7720 ^ n7717 ;
  assign n7662 = x75 & n5113 ;
  assign n7661 = x77 & n5116 ;
  assign n7663 = n7662 ^ n7661 ;
  assign n7664 = n7663 ^ x44 ;
  assign n7660 = ~n943 & n5117 ;
  assign n7665 = n7664 ^ n7660 ;
  assign n7659 = x76 & n5121 ;
  assign n7666 = n7665 ^ n7659 ;
  assign n7667 = n7666 ^ n7468 ;
  assign n7668 = n7667 ^ n7426 ;
  assign n7669 = n7668 ^ n7666 ;
  assign n7670 = n7474 & n7669 ;
  assign n7671 = n7670 ^ n7667 ;
  assign n7722 = n7721 ^ n7671 ;
  assign n7723 = n7722 ^ x41 ;
  assign n7658 = x78 & n4482 ;
  assign n7724 = n7723 ^ n7658 ;
  assign n7657 = x80 & n4478 ;
  assign n7725 = n7724 ^ n7657 ;
  assign n7656 = n1217 & n4479 ;
  assign n7726 = n7725 ^ n7656 ;
  assign n7728 = n7727 ^ n7726 ;
  assign n7653 = n7475 ^ n7418 ;
  assign n7654 = n7423 & n7653 ;
  assign n7655 = n7654 ^ n7418 ;
  assign n7729 = n7728 ^ n7655 ;
  assign n7730 = n7729 ^ x38 ;
  assign n7652 = x81 & n3932 ;
  assign n7731 = n7730 ^ n7652 ;
  assign n7651 = x83 & n3935 ;
  assign n7732 = n7731 ^ n7651 ;
  assign n7650 = n1517 & n3936 ;
  assign n7733 = n7732 ^ n7650 ;
  assign n7735 = n7734 ^ n7733 ;
  assign n7647 = n7476 ^ n7407 ;
  assign n7648 = n7482 & n7647 ;
  assign n7649 = n7648 ^ n7476 ;
  assign n7736 = n7735 ^ n7649 ;
  assign n7737 = n7736 ^ x35 ;
  assign n7646 = x84 & n3387 ;
  assign n7738 = n7737 ^ n7646 ;
  assign n7645 = x86 & n3390 ;
  assign n7739 = n7738 ^ n7645 ;
  assign n7644 = n1868 & n3391 ;
  assign n7740 = n7739 ^ n7644 ;
  assign n7742 = n7741 ^ n7740 ;
  assign n7746 = n7745 ^ n7742 ;
  assign n7747 = n7746 ^ x32 ;
  assign n7643 = x87 & n2890 ;
  assign n7748 = n7747 ^ n7643 ;
  assign n7642 = x89 & n2893 ;
  assign n7749 = n7748 ^ n7642 ;
  assign n7641 = n2255 & n2894 ;
  assign n7750 = n7749 ^ n7641 ;
  assign n7752 = n7751 ^ n7750 ;
  assign n7638 = n7499 ^ n7490 ;
  assign n7639 = ~n7496 & n7638 ;
  assign n7640 = n7639 ^ n7499 ;
  assign n7753 = n7752 ^ n7640 ;
  assign n7754 = n7753 ^ x29 ;
  assign n7637 = x90 & n2593 ;
  assign n7755 = n7754 ^ n7637 ;
  assign n7636 = x92 & n2428 ;
  assign n7756 = n7755 ^ n7636 ;
  assign n7635 = n2429 & n2696 ;
  assign n7757 = n7756 ^ n7635 ;
  assign n7759 = n7758 ^ n7757 ;
  assign n7763 = n7762 ^ n7759 ;
  assign n7764 = n7763 ^ x26 ;
  assign n7634 = x93 & n2032 ;
  assign n7765 = n7764 ^ n7634 ;
  assign n7633 = x95 & n2028 ;
  assign n7766 = n7765 ^ n7633 ;
  assign n7632 = n2029 & n3166 ;
  assign n7767 = n7766 ^ n7632 ;
  assign n7769 = n7768 ^ n7767 ;
  assign n7773 = n7772 ^ n7769 ;
  assign n7774 = n7773 ^ x23 ;
  assign n7631 = x96 & n1665 ;
  assign n7775 = n7774 ^ n7631 ;
  assign n7630 = x98 & n1668 ;
  assign n7776 = n7775 ^ n7630 ;
  assign n7629 = n1669 & n3673 ;
  assign n7777 = n7776 ^ n7629 ;
  assign n7779 = n7778 ^ n7777 ;
  assign n7783 = n7782 ^ n7779 ;
  assign n7784 = n7783 ^ x20 ;
  assign n7628 = x99 & n1340 ;
  assign n7785 = n7784 ^ n7628 ;
  assign n7627 = x101 & n1343 ;
  assign n7786 = n7785 ^ n7627 ;
  assign n7626 = n1344 & n4223 ;
  assign n7787 = n7786 ^ n7626 ;
  assign n7789 = n7788 ^ n7787 ;
  assign n7623 = n7530 ^ n7521 ;
  assign n7624 = n7527 & n7623 ;
  assign n7625 = n7624 ^ n7530 ;
  assign n7790 = n7789 ^ n7625 ;
  assign n7791 = n7790 ^ x17 ;
  assign n7622 = x102 & n1060 ;
  assign n7792 = n7791 ^ n7622 ;
  assign n7621 = x104 & n1063 ;
  assign n7793 = n7792 ^ n7621 ;
  assign n7620 = n1064 & ~n4830 ;
  assign n7794 = n7793 ^ n7620 ;
  assign n7796 = n7795 ^ n7794 ;
  assign n7800 = n7799 ^ n7796 ;
  assign n7801 = n7800 ^ x14 ;
  assign n7619 = x105 & n884 ;
  assign n7802 = n7801 ^ n7619 ;
  assign n7618 = x107 & n789 ;
  assign n7803 = n7802 ^ n7618 ;
  assign n7617 = n790 & ~n5459 ;
  assign n7804 = n7803 ^ n7617 ;
  assign n7806 = n7805 ^ n7804 ;
  assign n7810 = n7809 ^ n7806 ;
  assign n7811 = n7810 ^ x11 ;
  assign n7616 = x108 & n650 ;
  assign n7812 = n7811 ^ n7616 ;
  assign n7615 = x110 & ~n578 ;
  assign n7813 = n7812 ^ n7615 ;
  assign n7614 = ~n579 & n6145 ;
  assign n7814 = n7813 ^ n7614 ;
  assign n7816 = n7815 ^ n7814 ;
  assign n7611 = n7557 ^ n7553 ;
  assign n7612 = ~n7554 & ~n7611 ;
  assign n7613 = n7612 ^ n7557 ;
  assign n7817 = n7816 ^ n7613 ;
  assign n7818 = n7817 ^ x8 ;
  assign n7610 = x111 & n456 ;
  assign n7819 = n7818 ^ n7610 ;
  assign n7609 = x113 & n384 ;
  assign n7820 = n7819 ^ n7609 ;
  assign n7608 = n385 & ~n6849 ;
  assign n7821 = n7820 ^ n7608 ;
  assign n7823 = n7822 ^ n7821 ;
  assign n7827 = n7826 ^ n7823 ;
  assign n7828 = n7827 ^ x5 ;
  assign n7607 = x114 & n238 ;
  assign n7829 = n7828 ^ n7607 ;
  assign n7606 = x116 & n234 ;
  assign n7830 = n7829 ^ n7606 ;
  assign n7604 = n6835 ^ x116 ;
  assign n7605 = n235 & ~n7604 ;
  assign n7831 = n7830 ^ n7605 ;
  assign n7833 = n7832 ^ n7831 ;
  assign n7601 = n7574 ^ n7565 ;
  assign n7602 = n7571 & ~n7601 ;
  assign n7603 = n7602 ^ n7574 ;
  assign n7834 = n7833 ^ n7603 ;
  assign n7585 = x118 ^ x117 ;
  assign n7587 = n7339 & n7585 ;
  assign n7589 = x119 ^ x1 ;
  assign n7588 = x119 ^ x2 ;
  assign n7590 = n7589 ^ n7588 ;
  assign n7591 = ~n7587 & n7590 ;
  assign n7592 = n7591 ^ n7589 ;
  assign n7835 = n7834 ^ n7592 ;
  assign n7596 = x2 & x117 ;
  assign n7597 = n7596 ^ x118 ;
  assign n7598 = ~x1 & n7597 ;
  assign n7593 = n7592 ^ n7340 ;
  assign n7599 = n7598 ^ n7593 ;
  assign n7600 = ~x0 & n7599 ;
  assign n7836 = n7835 ^ n7600 ;
  assign n7582 = n7580 ^ n7575 ;
  assign n7583 = n7577 & n7582 ;
  assign n7584 = n7583 ^ n7580 ;
  assign n7837 = n7836 ^ n7584 ;
  assign n8107 = n7834 ^ n7584 ;
  assign n8108 = n7836 & ~n8107 ;
  assign n8109 = n8108 ^ n7834 ;
  assign n8101 = n7827 ^ n7603 ;
  assign n8102 = n7833 & n8101 ;
  assign n8103 = n8102 ^ n7827 ;
  assign n8099 = x116 & n231 ;
  assign n8092 = x113 & n391 ;
  assign n8084 = n7810 ^ n7613 ;
  assign n8085 = n7816 & ~n8084 ;
  assign n8086 = n8085 ^ n7810 ;
  assign n8082 = x110 & n584 ;
  assign n8075 = x107 & n795 ;
  assign n8068 = x104 & n1068 ;
  assign n8060 = n7783 ^ n7625 ;
  assign n8061 = n7789 & ~n8060 ;
  assign n8062 = n8061 ^ n7783 ;
  assign n8058 = x101 & n1348 ;
  assign n8051 = x98 & n1673 ;
  assign n8044 = x95 & n2025 ;
  assign n8037 = x92 & n2435 ;
  assign n8029 = n7746 ^ n7640 ;
  assign n8030 = n7752 & n8029 ;
  assign n8031 = n8030 ^ n7746 ;
  assign n8027 = x89 & n2899 ;
  assign n8020 = x86 & n3395 ;
  assign n8012 = n7729 ^ n7649 ;
  assign n8013 = n7735 & n8012 ;
  assign n8014 = n8013 ^ n7729 ;
  assign n8010 = x83 & n3940 ;
  assign n8001 = x77 & n5121 ;
  assign n7994 = x74 & n5755 ;
  assign n7986 = n7704 ^ n7677 ;
  assign n7987 = n7710 & n7986 ;
  assign n7988 = n7987 ^ n7704 ;
  assign n7984 = x71 & n6449 ;
  assign n7973 = x67 & n7183 ;
  assign n7972 = x69 & n7186 ;
  assign n7974 = n7973 ^ n7972 ;
  assign n7975 = n7974 ^ x53 ;
  assign n7971 = ~n376 & n7187 ;
  assign n7976 = n7975 ^ n7971 ;
  assign n7970 = x68 & n7191 ;
  assign n7977 = n7976 ^ n7970 ;
  assign n7966 = ~n7441 & ~n7694 ;
  assign n7967 = x56 & n7966 ;
  assign n7968 = n7967 ^ x56 ;
  assign n7963 = x66 & n7440 ;
  assign n7949 = x56 ^ x55 ;
  assign n7950 = n7440 & ~n7949 ;
  assign n7951 = n7950 ^ n7440 ;
  assign n7959 = x65 & n7951 ;
  assign n7952 = x56 ^ x54 ;
  assign n7953 = ~n7440 & n7952 ;
  assign n7954 = n7949 & n7953 ;
  assign n7960 = n7959 ^ n7954 ;
  assign n7961 = ~x64 & n7960 ;
  assign n7962 = n7961 ^ n7954 ;
  assign n7964 = n7963 ^ n7962 ;
  assign n7686 = x55 ^ x54 ;
  assign n7947 = ~n7440 & n7686 ;
  assign n7948 = x65 & n7947 ;
  assign n7965 = n7964 ^ n7948 ;
  assign n7969 = n7968 ^ n7965 ;
  assign n7978 = n7977 ^ n7969 ;
  assign n7944 = n7694 ^ n7683 ;
  assign n7945 = n7703 & ~n7944 ;
  assign n7946 = n7945 ^ n7702 ;
  assign n7979 = n7978 ^ n7946 ;
  assign n7980 = n7979 ^ x50 ;
  assign n7943 = x70 & n6687 ;
  assign n7981 = n7980 ^ n7943 ;
  assign n7942 = x72 & n6444 ;
  assign n7982 = n7981 ^ n7942 ;
  assign n7941 = n565 & n6445 ;
  assign n7983 = n7982 ^ n7941 ;
  assign n7985 = n7984 ^ n7983 ;
  assign n7989 = n7988 ^ n7985 ;
  assign n7990 = n7989 ^ x47 ;
  assign n7940 = x73 & n5981 ;
  assign n7991 = n7990 ^ n7940 ;
  assign n7939 = x75 & n5748 ;
  assign n7992 = n7991 ^ n7939 ;
  assign n7938 = ~n778 & n5749 ;
  assign n7993 = n7992 ^ n7938 ;
  assign n7995 = n7994 ^ n7993 ;
  assign n7935 = n7720 ^ n7711 ;
  assign n7936 = ~n7717 & n7935 ;
  assign n7937 = n7936 ^ n7720 ;
  assign n7996 = n7995 ^ n7937 ;
  assign n7997 = n7996 ^ x44 ;
  assign n7934 = x76 & n5113 ;
  assign n7998 = n7997 ^ n7934 ;
  assign n7933 = x78 & n5116 ;
  assign n7999 = n7998 ^ n7933 ;
  assign n7932 = ~n1036 & n5117 ;
  assign n8000 = n7999 ^ n7932 ;
  assign n8002 = n8001 ^ n8000 ;
  assign n7927 = x79 & n4482 ;
  assign n7926 = x81 & n4478 ;
  assign n7928 = n7927 ^ n7926 ;
  assign n7929 = n7928 ^ x41 ;
  assign n7925 = n1310 & n4479 ;
  assign n7930 = n7929 ^ n7925 ;
  assign n7924 = x80 & n4475 ;
  assign n7931 = n7930 ^ n7924 ;
  assign n8003 = n8002 ^ n7931 ;
  assign n7921 = n7721 ^ n7666 ;
  assign n7922 = n7671 & n7921 ;
  assign n7923 = n7922 ^ n7666 ;
  assign n8004 = n8003 ^ n7923 ;
  assign n7918 = n7722 ^ n7655 ;
  assign n7919 = n7728 & n7918 ;
  assign n7920 = n7919 ^ n7722 ;
  assign n8005 = n8004 ^ n7920 ;
  assign n8006 = n8005 ^ x38 ;
  assign n7917 = x82 & n3932 ;
  assign n8007 = n8006 ^ n7917 ;
  assign n7916 = x84 & n3935 ;
  assign n8008 = n8007 ^ n7916 ;
  assign n7915 = n1635 & n3936 ;
  assign n8009 = n8008 ^ n7915 ;
  assign n8011 = n8010 ^ n8009 ;
  assign n8015 = n8014 ^ n8011 ;
  assign n8016 = n8015 ^ x35 ;
  assign n7914 = x85 & n3387 ;
  assign n8017 = n8016 ^ n7914 ;
  assign n7913 = x87 & n3390 ;
  assign n8018 = n8017 ^ n7913 ;
  assign n7912 = n1987 & n3391 ;
  assign n8019 = n8018 ^ n7912 ;
  assign n8021 = n8020 ^ n8019 ;
  assign n7909 = n7745 ^ n7736 ;
  assign n7910 = ~n7742 & n7909 ;
  assign n7911 = n7910 ^ n7745 ;
  assign n8022 = n8021 ^ n7911 ;
  assign n8023 = n8022 ^ x32 ;
  assign n7908 = x88 & n2890 ;
  assign n8024 = n8023 ^ n7908 ;
  assign n7907 = x90 & n2893 ;
  assign n8025 = n8024 ^ n7907 ;
  assign n7906 = n2398 & n2894 ;
  assign n8026 = n8025 ^ n7906 ;
  assign n8028 = n8027 ^ n8026 ;
  assign n8032 = n8031 ^ n8028 ;
  assign n8033 = n8032 ^ x29 ;
  assign n7905 = x91 & n2593 ;
  assign n8034 = n8033 ^ n7905 ;
  assign n7904 = x93 & n2428 ;
  assign n8035 = n8034 ^ n7904 ;
  assign n7903 = n2429 & n2842 ;
  assign n8036 = n8035 ^ n7903 ;
  assign n8038 = n8037 ^ n8036 ;
  assign n7900 = n7762 ^ n7753 ;
  assign n7901 = ~n7759 & n7900 ;
  assign n7902 = n7901 ^ n7762 ;
  assign n8039 = n8038 ^ n7902 ;
  assign n8040 = n8039 ^ x26 ;
  assign n7899 = x94 & n2032 ;
  assign n8041 = n8040 ^ n7899 ;
  assign n7898 = x96 & n2028 ;
  assign n8042 = n8041 ^ n7898 ;
  assign n7897 = n2029 & n3336 ;
  assign n8043 = n8042 ^ n7897 ;
  assign n8045 = n8044 ^ n8043 ;
  assign n7894 = n7772 ^ n7763 ;
  assign n7895 = ~n7769 & n7894 ;
  assign n7896 = n7895 ^ n7772 ;
  assign n8046 = n8045 ^ n7896 ;
  assign n8047 = n8046 ^ x23 ;
  assign n7893 = x97 & n1665 ;
  assign n8048 = n8047 ^ n7893 ;
  assign n7892 = x99 & n1668 ;
  assign n8049 = n8048 ^ n7892 ;
  assign n7891 = n1669 & n3851 ;
  assign n8050 = n8049 ^ n7891 ;
  assign n8052 = n8051 ^ n8050 ;
  assign n7888 = n7782 ^ n7773 ;
  assign n7889 = ~n7779 & n7888 ;
  assign n7890 = n7889 ^ n7782 ;
  assign n8053 = n8052 ^ n7890 ;
  assign n8054 = n8053 ^ x20 ;
  assign n7887 = x100 & n1340 ;
  assign n8055 = n8054 ^ n7887 ;
  assign n7886 = x102 & n1343 ;
  assign n8056 = n8055 ^ n7886 ;
  assign n7885 = n1344 & n4425 ;
  assign n8057 = n8056 ^ n7885 ;
  assign n8059 = n8058 ^ n8057 ;
  assign n8063 = n8062 ^ n8059 ;
  assign n8064 = n8063 ^ x17 ;
  assign n7884 = x103 & n1060 ;
  assign n8065 = n8064 ^ n7884 ;
  assign n7883 = x105 & n1063 ;
  assign n8066 = n8065 ^ n7883 ;
  assign n7882 = n1064 & ~n5034 ;
  assign n8067 = n8066 ^ n7882 ;
  assign n8069 = n8068 ^ n8067 ;
  assign n7879 = n7799 ^ n7790 ;
  assign n7880 = n7796 & ~n7879 ;
  assign n7881 = n7880 ^ n7799 ;
  assign n8070 = n8069 ^ n7881 ;
  assign n8071 = n8070 ^ x14 ;
  assign n7878 = x106 & n884 ;
  assign n8072 = n8071 ^ n7878 ;
  assign n7877 = x108 & n789 ;
  assign n8073 = n8072 ^ n7877 ;
  assign n7876 = n790 & n5687 ;
  assign n8074 = n8073 ^ n7876 ;
  assign n8076 = n8075 ^ n8074 ;
  assign n7873 = n7809 ^ n7800 ;
  assign n7874 = n7806 & n7873 ;
  assign n7875 = n7874 ^ n7809 ;
  assign n8077 = n8076 ^ n7875 ;
  assign n8078 = n8077 ^ x11 ;
  assign n7872 = x109 & n650 ;
  assign n8079 = n8078 ^ n7872 ;
  assign n7871 = x111 & ~n578 ;
  assign n8080 = n8079 ^ n7871 ;
  assign n7870 = ~n579 & ~n6370 ;
  assign n8081 = n8080 ^ n7870 ;
  assign n8083 = n8082 ^ n8081 ;
  assign n8087 = n8086 ^ n8083 ;
  assign n8088 = n8087 ^ x8 ;
  assign n7869 = x112 & n456 ;
  assign n8089 = n8088 ^ n7869 ;
  assign n7868 = x114 & n384 ;
  assign n8090 = n8089 ^ n7868 ;
  assign n7867 = n385 & ~n7108 ;
  assign n8091 = n8090 ^ n7867 ;
  assign n8093 = n8092 ^ n8091 ;
  assign n7864 = n7826 ^ n7817 ;
  assign n7865 = n7823 & n7864 ;
  assign n7866 = n7865 ^ n7826 ;
  assign n8094 = n8093 ^ n7866 ;
  assign n8095 = n8094 ^ x5 ;
  assign n7863 = x115 & n238 ;
  assign n8096 = n8095 ^ n7863 ;
  assign n7862 = x117 & n234 ;
  assign n8097 = n8096 ^ n7862 ;
  assign n7860 = n7091 ^ x117 ;
  assign n7861 = n235 & ~n7860 ;
  assign n8098 = n8097 ^ n7861 ;
  assign n8100 = n8099 ^ n8098 ;
  assign n8104 = n8103 ^ n8100 ;
  assign n7838 = x119 ^ x118 ;
  assign n7844 = ~x119 & n7339 ;
  assign n7845 = n7844 ^ n7337 ;
  assign n7846 = n7838 & ~n7845 ;
  assign n7848 = x120 ^ x1 ;
  assign n7847 = x120 ^ x2 ;
  assign n7849 = n7848 ^ n7847 ;
  assign n7850 = ~n7846 & n7849 ;
  assign n7851 = n7850 ^ n7848 ;
  assign n8105 = n8104 ^ n7851 ;
  assign n7855 = x2 & x118 ;
  assign n7856 = n7855 ^ x119 ;
  assign n7857 = ~x1 & n7856 ;
  assign n7852 = n7851 ^ n7588 ;
  assign n7858 = n7857 ^ n7852 ;
  assign n7859 = ~x0 & n7858 ;
  assign n8106 = n8105 ^ n7859 ;
  assign n8110 = n8109 ^ n8106 ;
  assign n8377 = x117 & n231 ;
  assign n8369 = n8087 ^ n7866 ;
  assign n8370 = ~n8093 & n8369 ;
  assign n8371 = n8370 ^ n8087 ;
  assign n8367 = x114 & n391 ;
  assign n8360 = x111 & n584 ;
  assign n8352 = n8070 ^ n7875 ;
  assign n8353 = n8076 & ~n8352 ;
  assign n8354 = n8353 ^ n8070 ;
  assign n8350 = x108 & n795 ;
  assign n8342 = n8063 ^ n7881 ;
  assign n8343 = n8069 & n8342 ;
  assign n8344 = n8343 ^ n8063 ;
  assign n8340 = x105 & n1068 ;
  assign n8333 = x102 & n1348 ;
  assign n8325 = n8046 ^ n7890 ;
  assign n8326 = n8052 & n8325 ;
  assign n8327 = n8326 ^ n8046 ;
  assign n8323 = x99 & n1673 ;
  assign n8315 = n8039 ^ n7896 ;
  assign n8316 = n8045 & n8315 ;
  assign n8317 = n8316 ^ n8039 ;
  assign n8313 = x96 & n2025 ;
  assign n8305 = n8032 ^ n7902 ;
  assign n8306 = n8038 & n8305 ;
  assign n8307 = n8306 ^ n8032 ;
  assign n8303 = x93 & n2435 ;
  assign n8296 = x90 & n2899 ;
  assign n8288 = n8015 ^ n7911 ;
  assign n8289 = n8021 & n8288 ;
  assign n8290 = n8289 ^ n8015 ;
  assign n8286 = x87 & n3395 ;
  assign n8279 = x84 & n3940 ;
  assign n8271 = n7931 ^ n7920 ;
  assign n8272 = n8004 & n8271 ;
  assign n8273 = n8272 ^ n7931 ;
  assign n8269 = x81 & n4475 ;
  assign n8260 = n7989 ^ n7937 ;
  assign n8261 = n7995 & n8260 ;
  assign n8262 = n8261 ^ n7989 ;
  assign n8258 = x75 & n5755 ;
  assign n8245 = x65 & n7954 ;
  assign n8244 = x66 & n7947 ;
  assign n8246 = n8245 ^ n8244 ;
  assign n8247 = n8246 ^ x56 ;
  assign n8241 = ~n155 & ~n7949 ;
  assign n8242 = n8241 ^ n295 ;
  assign n8243 = n7440 & ~n8242 ;
  assign n8248 = n8247 ^ n8243 ;
  assign n8234 = x57 ^ x56 ;
  assign n8235 = x64 & n8234 ;
  assign n8249 = n8248 ^ n8235 ;
  assign n8236 = ~n7965 & n7967 ;
  assign n8237 = ~n8235 & ~n8236 ;
  assign n8238 = n8237 ^ n8236 ;
  assign n8250 = n8249 ^ n8238 ;
  assign n8251 = n8250 ^ n8237 ;
  assign n8231 = n7977 ^ n7946 ;
  assign n8232 = n7978 & n8231 ;
  assign n8224 = x68 & n7183 ;
  assign n8223 = x70 & n7186 ;
  assign n8225 = n8224 ^ n8223 ;
  assign n8226 = n8225 ^ x53 ;
  assign n8222 = ~n443 & n7187 ;
  assign n8227 = n8226 ^ n8222 ;
  assign n8221 = x69 & n7191 ;
  assign n8228 = n8227 ^ n8221 ;
  assign n8229 = n8228 ^ n7977 ;
  assign n8233 = n8232 ^ n8229 ;
  assign n8252 = n8251 ^ n8233 ;
  assign n8211 = x71 & n6687 ;
  assign n8210 = x73 & n6444 ;
  assign n8212 = n8211 ^ n8210 ;
  assign n8213 = n8212 ^ x50 ;
  assign n8209 = n636 & n6445 ;
  assign n8214 = n8213 ^ n8209 ;
  assign n8208 = x72 & n6449 ;
  assign n8215 = n8214 ^ n8208 ;
  assign n8216 = n8215 ^ n7988 ;
  assign n8217 = n8216 ^ n7979 ;
  assign n8218 = n8217 ^ n8215 ;
  assign n8219 = ~n7985 & n8218 ;
  assign n8220 = n8219 ^ n8216 ;
  assign n8253 = n8252 ^ n8220 ;
  assign n8254 = n8253 ^ x47 ;
  assign n8207 = x74 & n5981 ;
  assign n8255 = n8254 ^ n8207 ;
  assign n8206 = x76 & n5748 ;
  assign n8256 = n8255 ^ n8206 ;
  assign n8205 = ~n863 & n5749 ;
  assign n8257 = n8256 ^ n8205 ;
  assign n8259 = n8258 ^ n8257 ;
  assign n8263 = n8262 ^ n8259 ;
  assign n8195 = x77 & n5113 ;
  assign n8194 = x79 & n5116 ;
  assign n8196 = n8195 ^ n8194 ;
  assign n8197 = n8196 ^ x44 ;
  assign n8193 = n1123 & n5117 ;
  assign n8198 = n8197 ^ n8193 ;
  assign n8192 = x78 & n5121 ;
  assign n8199 = n8198 ^ n8192 ;
  assign n8200 = n8199 ^ n7996 ;
  assign n8201 = n8200 ^ n7923 ;
  assign n8202 = n8201 ^ n8199 ;
  assign n8203 = n8002 & n8202 ;
  assign n8204 = n8203 ^ n8200 ;
  assign n8264 = n8263 ^ n8204 ;
  assign n8265 = n8264 ^ x41 ;
  assign n8191 = x80 & n4482 ;
  assign n8266 = n8265 ^ n8191 ;
  assign n8190 = x82 & n4478 ;
  assign n8267 = n8266 ^ n8190 ;
  assign n8189 = n1422 & n4479 ;
  assign n8268 = n8267 ^ n8189 ;
  assign n8270 = n8269 ^ n8268 ;
  assign n8274 = n8273 ^ n8270 ;
  assign n8275 = n8274 ^ x38 ;
  assign n8188 = x83 & n3932 ;
  assign n8276 = n8275 ^ n8188 ;
  assign n8187 = x85 & n3935 ;
  assign n8277 = n8276 ^ n8187 ;
  assign n8186 = n1748 & n3936 ;
  assign n8278 = n8277 ^ n8186 ;
  assign n8280 = n8279 ^ n8278 ;
  assign n8183 = n8014 ^ n8005 ;
  assign n8184 = ~n8011 & n8183 ;
  assign n8185 = n8184 ^ n8014 ;
  assign n8281 = n8280 ^ n8185 ;
  assign n8282 = n8281 ^ x35 ;
  assign n8182 = x86 & n3387 ;
  assign n8283 = n8282 ^ n8182 ;
  assign n8181 = x88 & n3390 ;
  assign n8284 = n8283 ^ n8181 ;
  assign n8180 = n2131 & n3391 ;
  assign n8285 = n8284 ^ n8180 ;
  assign n8287 = n8286 ^ n8285 ;
  assign n8291 = n8290 ^ n8287 ;
  assign n8292 = n8291 ^ x32 ;
  assign n8179 = x89 & n2890 ;
  assign n8293 = n8292 ^ n8179 ;
  assign n8178 = x91 & n2893 ;
  assign n8294 = n8293 ^ n8178 ;
  assign n8177 = n2548 & n2894 ;
  assign n8295 = n8294 ^ n8177 ;
  assign n8297 = n8296 ^ n8295 ;
  assign n8174 = n8031 ^ n8022 ;
  assign n8175 = ~n8028 & n8174 ;
  assign n8176 = n8175 ^ n8031 ;
  assign n8298 = n8297 ^ n8176 ;
  assign n8299 = n8298 ^ x29 ;
  assign n8173 = x92 & n2593 ;
  assign n8300 = n8299 ^ n8173 ;
  assign n8172 = x94 & n2428 ;
  assign n8301 = n8300 ^ n8172 ;
  assign n8171 = n2429 & n3010 ;
  assign n8302 = n8301 ^ n8171 ;
  assign n8304 = n8303 ^ n8302 ;
  assign n8308 = n8307 ^ n8304 ;
  assign n8309 = n8308 ^ x26 ;
  assign n8170 = x95 & n2032 ;
  assign n8310 = n8309 ^ n8170 ;
  assign n8169 = x97 & n2028 ;
  assign n8311 = n8310 ^ n8169 ;
  assign n8168 = n2029 & n3501 ;
  assign n8312 = n8311 ^ n8168 ;
  assign n8314 = n8313 ^ n8312 ;
  assign n8318 = n8317 ^ n8314 ;
  assign n8319 = n8318 ^ x23 ;
  assign n8167 = x98 & n1665 ;
  assign n8320 = n8319 ^ n8167 ;
  assign n8166 = x100 & n1668 ;
  assign n8321 = n8320 ^ n8166 ;
  assign n8165 = n1669 & n4048 ;
  assign n8322 = n8321 ^ n8165 ;
  assign n8324 = n8323 ^ n8322 ;
  assign n8328 = n8327 ^ n8324 ;
  assign n8329 = n8328 ^ x20 ;
  assign n8164 = x101 & n1340 ;
  assign n8330 = n8329 ^ n8164 ;
  assign n8163 = x103 & n1343 ;
  assign n8331 = n8330 ^ n8163 ;
  assign n8162 = n1344 & ~n4624 ;
  assign n8332 = n8331 ^ n8162 ;
  assign n8334 = n8333 ^ n8332 ;
  assign n8159 = n8062 ^ n8053 ;
  assign n8160 = ~n8059 & n8159 ;
  assign n8161 = n8160 ^ n8062 ;
  assign n8335 = n8334 ^ n8161 ;
  assign n8336 = n8335 ^ x17 ;
  assign n8158 = x104 & n1060 ;
  assign n8337 = n8336 ^ n8158 ;
  assign n8157 = x106 & n1063 ;
  assign n8338 = n8337 ^ n8157 ;
  assign n8156 = n1064 & ~n5257 ;
  assign n8339 = n8338 ^ n8156 ;
  assign n8341 = n8340 ^ n8339 ;
  assign n8345 = n8344 ^ n8341 ;
  assign n8346 = n8345 ^ x14 ;
  assign n8155 = x107 & n884 ;
  assign n8347 = n8346 ^ n8155 ;
  assign n8154 = x109 & n789 ;
  assign n8348 = n8347 ^ n8154 ;
  assign n8153 = n790 & n5912 ;
  assign n8349 = n8348 ^ n8153 ;
  assign n8351 = n8350 ^ n8349 ;
  assign n8355 = n8354 ^ n8351 ;
  assign n8356 = n8355 ^ x11 ;
  assign n8152 = x110 & n650 ;
  assign n8357 = n8356 ^ n8152 ;
  assign n8151 = x112 & ~n578 ;
  assign n8358 = n8357 ^ n8151 ;
  assign n8150 = ~n579 & ~n6616 ;
  assign n8359 = n8358 ^ n8150 ;
  assign n8361 = n8360 ^ n8359 ;
  assign n8147 = n8086 ^ n8077 ;
  assign n8148 = n8083 & ~n8147 ;
  assign n8149 = n8148 ^ n8086 ;
  assign n8362 = n8361 ^ n8149 ;
  assign n8363 = n8362 ^ x8 ;
  assign n8146 = x113 & n456 ;
  assign n8364 = n8363 ^ n8146 ;
  assign n8145 = x115 & n384 ;
  assign n8365 = n8364 ^ n8145 ;
  assign n8144 = n385 & ~n7353 ;
  assign n8366 = n8365 ^ n8144 ;
  assign n8368 = n8367 ^ n8366 ;
  assign n8372 = n8371 ^ n8368 ;
  assign n8373 = n8372 ^ x5 ;
  assign n8143 = x116 & n238 ;
  assign n8374 = n8373 ^ n8143 ;
  assign n8142 = x118 & n234 ;
  assign n8375 = n8374 ^ n8142 ;
  assign n8139 = n7339 ^ x117 ;
  assign n8140 = n8139 ^ n7585 ;
  assign n8141 = n235 & ~n8140 ;
  assign n8376 = n8375 ^ n8141 ;
  assign n8378 = n8377 ^ n8376 ;
  assign n8136 = n8103 ^ n8094 ;
  assign n8137 = ~n8100 & n8136 ;
  assign n8138 = n8137 ^ n8103 ;
  assign n8379 = n8378 ^ n8138 ;
  assign n8116 = x120 ^ x117 ;
  assign n8114 = x120 ^ x119 ;
  assign n8117 = n7838 & n8114 ;
  assign n8118 = n7339 & n8117 ;
  assign n8119 = n8116 & n8118 ;
  assign n8120 = n8119 ^ n8117 ;
  assign n8121 = n8120 ^ x119 ;
  assign n8122 = n8121 ^ x120 ;
  assign n8124 = x121 ^ x1 ;
  assign n8123 = x121 ^ x2 ;
  assign n8125 = n8124 ^ n8123 ;
  assign n8126 = ~n8122 & n8125 ;
  assign n8127 = n8126 ^ n8124 ;
  assign n8380 = n8379 ^ n8127 ;
  assign n8131 = x2 & x119 ;
  assign n8132 = n8131 ^ x120 ;
  assign n8133 = ~x1 & n8132 ;
  assign n8128 = n8127 ^ n7847 ;
  assign n8134 = n8133 ^ n8128 ;
  assign n8135 = ~x0 & n8134 ;
  assign n8381 = n8380 ^ n8135 ;
  assign n8111 = n8109 ^ n8104 ;
  assign n8112 = ~n8106 & n8111 ;
  assign n8113 = n8112 ^ n8109 ;
  assign n8382 = n8381 ^ n8113 ;
  assign n8649 = n8379 ^ n8113 ;
  assign n8650 = ~n8381 & ~n8649 ;
  assign n8651 = n8650 ^ n8379 ;
  assign n8645 = n8372 ^ n8138 ;
  assign n8646 = ~n8378 & ~n8645 ;
  assign n8647 = n8646 ^ n8372 ;
  assign n8641 = x115 & n391 ;
  assign n8633 = n8355 ^ n8149 ;
  assign n8634 = n8361 & n8633 ;
  assign n8635 = n8634 ^ n8355 ;
  assign n8631 = x112 & n584 ;
  assign n8624 = x109 & n795 ;
  assign n8617 = x106 & n1068 ;
  assign n8609 = n8328 ^ n8161 ;
  assign n8610 = n8334 & n8609 ;
  assign n8611 = n8610 ^ n8328 ;
  assign n8607 = x103 & n1348 ;
  assign n8600 = x100 & n1673 ;
  assign n8593 = x97 & n2025 ;
  assign n8582 = x93 & n2593 ;
  assign n8581 = x95 & n2428 ;
  assign n8583 = n8582 ^ n8581 ;
  assign n8584 = n8583 ^ x29 ;
  assign n8580 = n2429 & n3166 ;
  assign n8585 = n8584 ^ n8580 ;
  assign n8579 = x94 & n2435 ;
  assign n8586 = n8585 ^ n8579 ;
  assign n8575 = n8291 ^ n8176 ;
  assign n8576 = n8297 & n8575 ;
  assign n8577 = n8576 ^ n8291 ;
  assign n8573 = x91 & n2899 ;
  assign n8566 = x88 & n3395 ;
  assign n8558 = n8274 ^ n8185 ;
  assign n8559 = n8280 & n8558 ;
  assign n8560 = n8559 ^ n8274 ;
  assign n8556 = x85 & n3940 ;
  assign n8549 = x82 & n4475 ;
  assign n8542 = x79 & n5121 ;
  assign n8535 = x76 & n5755 ;
  assign n8528 = x73 & n6449 ;
  assign n8521 = x70 & n7191 ;
  assign n8511 = x66 & n7954 ;
  assign n8510 = x68 & n7950 ;
  assign n8512 = n8511 ^ n8510 ;
  assign n8513 = n8512 ^ x56 ;
  assign n8509 = ~n351 & n7951 ;
  assign n8514 = n8513 ^ n8509 ;
  assign n8508 = x67 & n7947 ;
  assign n8515 = n8514 ^ n8508 ;
  assign n8506 = ~n8237 & n8248 ;
  assign n8503 = x65 ^ x57 ;
  assign n8504 = n8234 & ~n8503 ;
  assign n8499 = x56 & x57 ;
  assign n8500 = n8499 ^ x58 ;
  assign n8501 = ~x64 & n8500 ;
  assign n8495 = x58 ^ x56 ;
  assign n8502 = n8501 ^ n8495 ;
  assign n8505 = n8504 ^ n8502 ;
  assign n8507 = n8506 ^ n8505 ;
  assign n8516 = n8515 ^ n8507 ;
  assign n8517 = n8516 ^ x53 ;
  assign n8494 = x69 & n7183 ;
  assign n8518 = n8517 ^ n8494 ;
  assign n8493 = x71 & n7186 ;
  assign n8519 = n8518 ^ n8493 ;
  assign n8492 = ~n495 & n7187 ;
  assign n8520 = n8519 ^ n8492 ;
  assign n8522 = n8521 ^ n8520 ;
  assign n8489 = n8251 ^ n8228 ;
  assign n8490 = n8233 & n8489 ;
  assign n8491 = n8490 ^ n8228 ;
  assign n8523 = n8522 ^ n8491 ;
  assign n8524 = n8523 ^ x50 ;
  assign n8488 = x72 & n6687 ;
  assign n8525 = n8524 ^ n8488 ;
  assign n8487 = x74 & n6444 ;
  assign n8526 = n8525 ^ n8487 ;
  assign n8486 = n708 & n6445 ;
  assign n8527 = n8526 ^ n8486 ;
  assign n8529 = n8528 ^ n8527 ;
  assign n8483 = n8252 ^ n8215 ;
  assign n8484 = n8220 & n8483 ;
  assign n8485 = n8484 ^ n8215 ;
  assign n8530 = n8529 ^ n8485 ;
  assign n8531 = n8530 ^ x47 ;
  assign n8482 = x75 & n5981 ;
  assign n8532 = n8531 ^ n8482 ;
  assign n8481 = x77 & n5748 ;
  assign n8533 = n8532 ^ n8481 ;
  assign n8480 = ~n943 & n5749 ;
  assign n8534 = n8533 ^ n8480 ;
  assign n8536 = n8535 ^ n8534 ;
  assign n8477 = n8262 ^ n8253 ;
  assign n8478 = ~n8259 & n8477 ;
  assign n8479 = n8478 ^ n8262 ;
  assign n8537 = n8536 ^ n8479 ;
  assign n8538 = n8537 ^ x44 ;
  assign n8476 = x78 & n5113 ;
  assign n8539 = n8538 ^ n8476 ;
  assign n8475 = x80 & n5116 ;
  assign n8540 = n8539 ^ n8475 ;
  assign n8474 = n1217 & n5117 ;
  assign n8541 = n8540 ^ n8474 ;
  assign n8543 = n8542 ^ n8541 ;
  assign n8471 = n8263 ^ n8199 ;
  assign n8472 = n8204 & n8471 ;
  assign n8473 = n8472 ^ n8199 ;
  assign n8544 = n8543 ^ n8473 ;
  assign n8545 = n8544 ^ x41 ;
  assign n8470 = x81 & n4482 ;
  assign n8546 = n8545 ^ n8470 ;
  assign n8469 = x83 & n4478 ;
  assign n8547 = n8546 ^ n8469 ;
  assign n8468 = n1517 & n4479 ;
  assign n8548 = n8547 ^ n8468 ;
  assign n8550 = n8549 ^ n8548 ;
  assign n8465 = n8273 ^ n8264 ;
  assign n8466 = ~n8270 & n8465 ;
  assign n8467 = n8466 ^ n8273 ;
  assign n8551 = n8550 ^ n8467 ;
  assign n8552 = n8551 ^ x38 ;
  assign n8464 = x84 & n3932 ;
  assign n8553 = n8552 ^ n8464 ;
  assign n8463 = x86 & n3935 ;
  assign n8554 = n8553 ^ n8463 ;
  assign n8462 = n1868 & n3936 ;
  assign n8555 = n8554 ^ n8462 ;
  assign n8557 = n8556 ^ n8555 ;
  assign n8561 = n8560 ^ n8557 ;
  assign n8562 = n8561 ^ x35 ;
  assign n8461 = x87 & n3387 ;
  assign n8563 = n8562 ^ n8461 ;
  assign n8460 = x89 & n3390 ;
  assign n8564 = n8563 ^ n8460 ;
  assign n8459 = n2255 & n3391 ;
  assign n8565 = n8564 ^ n8459 ;
  assign n8567 = n8566 ^ n8565 ;
  assign n8456 = n8290 ^ n8281 ;
  assign n8457 = ~n8287 & n8456 ;
  assign n8458 = n8457 ^ n8290 ;
  assign n8568 = n8567 ^ n8458 ;
  assign n8569 = n8568 ^ x32 ;
  assign n8455 = x90 & n2890 ;
  assign n8570 = n8569 ^ n8455 ;
  assign n8454 = x92 & n2893 ;
  assign n8571 = n8570 ^ n8454 ;
  assign n8453 = n2696 & n2894 ;
  assign n8572 = n8571 ^ n8453 ;
  assign n8574 = n8573 ^ n8572 ;
  assign n8578 = n8577 ^ n8574 ;
  assign n8587 = n8586 ^ n8578 ;
  assign n8450 = n8307 ^ n8298 ;
  assign n8451 = ~n8304 & n8450 ;
  assign n8452 = n8451 ^ n8307 ;
  assign n8588 = n8587 ^ n8452 ;
  assign n8589 = n8588 ^ x26 ;
  assign n8449 = x96 & n2032 ;
  assign n8590 = n8589 ^ n8449 ;
  assign n8448 = x98 & n2028 ;
  assign n8591 = n8590 ^ n8448 ;
  assign n8447 = n2029 & n3673 ;
  assign n8592 = n8591 ^ n8447 ;
  assign n8594 = n8593 ^ n8592 ;
  assign n8444 = n8317 ^ n8308 ;
  assign n8445 = ~n8314 & n8444 ;
  assign n8446 = n8445 ^ n8317 ;
  assign n8595 = n8594 ^ n8446 ;
  assign n8596 = n8595 ^ x23 ;
  assign n8443 = x99 & n1665 ;
  assign n8597 = n8596 ^ n8443 ;
  assign n8442 = x101 & n1668 ;
  assign n8598 = n8597 ^ n8442 ;
  assign n8441 = n1669 & n4223 ;
  assign n8599 = n8598 ^ n8441 ;
  assign n8601 = n8600 ^ n8599 ;
  assign n8438 = n8327 ^ n8318 ;
  assign n8439 = ~n8324 & n8438 ;
  assign n8440 = n8439 ^ n8327 ;
  assign n8602 = n8601 ^ n8440 ;
  assign n8603 = n8602 ^ x20 ;
  assign n8437 = x102 & n1340 ;
  assign n8604 = n8603 ^ n8437 ;
  assign n8436 = x104 & n1343 ;
  assign n8605 = n8604 ^ n8436 ;
  assign n8435 = n1344 & ~n4830 ;
  assign n8606 = n8605 ^ n8435 ;
  assign n8608 = n8607 ^ n8606 ;
  assign n8612 = n8611 ^ n8608 ;
  assign n8613 = n8612 ^ x17 ;
  assign n8434 = x105 & n1060 ;
  assign n8614 = n8613 ^ n8434 ;
  assign n8433 = x107 & n1063 ;
  assign n8615 = n8614 ^ n8433 ;
  assign n8432 = n1064 & ~n5459 ;
  assign n8616 = n8615 ^ n8432 ;
  assign n8618 = n8617 ^ n8616 ;
  assign n8429 = n8344 ^ n8335 ;
  assign n8430 = ~n8341 & n8429 ;
  assign n8431 = n8430 ^ n8344 ;
  assign n8619 = n8618 ^ n8431 ;
  assign n8620 = n8619 ^ x14 ;
  assign n8428 = x108 & n884 ;
  assign n8621 = n8620 ^ n8428 ;
  assign n8427 = x110 & n789 ;
  assign n8622 = n8621 ^ n8427 ;
  assign n8426 = n790 & n6145 ;
  assign n8623 = n8622 ^ n8426 ;
  assign n8625 = n8624 ^ n8623 ;
  assign n8423 = n8354 ^ n8345 ;
  assign n8424 = ~n8351 & n8423 ;
  assign n8425 = n8424 ^ n8354 ;
  assign n8626 = n8625 ^ n8425 ;
  assign n8627 = n8626 ^ x11 ;
  assign n8422 = x111 & n650 ;
  assign n8628 = n8627 ^ n8422 ;
  assign n8421 = x113 & ~n578 ;
  assign n8629 = n8628 ^ n8421 ;
  assign n8420 = ~n579 & ~n6849 ;
  assign n8630 = n8629 ^ n8420 ;
  assign n8632 = n8631 ^ n8630 ;
  assign n8636 = n8635 ^ n8632 ;
  assign n8637 = n8636 ^ x8 ;
  assign n8419 = x114 & n456 ;
  assign n8638 = n8637 ^ n8419 ;
  assign n8418 = x116 & n384 ;
  assign n8639 = n8638 ^ n8418 ;
  assign n8417 = n385 & ~n7604 ;
  assign n8640 = n8639 ^ n8417 ;
  assign n8642 = n8641 ^ n8640 ;
  assign n8414 = n8371 ^ n8362 ;
  assign n8415 = ~n8368 & ~n8414 ;
  assign n8416 = n8415 ^ n8371 ;
  assign n8643 = n8642 ^ n8416 ;
  assign n8408 = x117 & n238 ;
  assign n8407 = x119 & n234 ;
  assign n8409 = n8408 ^ n8407 ;
  assign n8410 = n8409 ^ x5 ;
  assign n8405 = n7587 ^ x119 ;
  assign n8406 = n235 & n8405 ;
  assign n8411 = n8410 ^ n8406 ;
  assign n8404 = x118 & n231 ;
  assign n8412 = n8411 ^ n8404 ;
  assign n8398 = x2 & x120 ;
  assign n8399 = n8398 ^ x121 ;
  assign n8400 = ~x1 & n8399 ;
  assign n8383 = x120 & n8121 ;
  assign n8385 = n8383 ^ n8122 ;
  assign n8386 = x121 & n8385 ;
  assign n8384 = ~x121 & ~n8383 ;
  assign n8387 = n8386 ^ n8384 ;
  assign n8389 = x122 ^ x1 ;
  assign n8388 = x122 ^ x2 ;
  assign n8390 = n8389 ^ n8388 ;
  assign n8391 = n8387 & n8390 ;
  assign n8392 = n8391 ^ n8389 ;
  assign n8395 = n8392 ^ n8123 ;
  assign n8401 = n8400 ^ n8395 ;
  assign n8402 = ~x0 & n8401 ;
  assign n8403 = n8402 ^ n8392 ;
  assign n8413 = n8412 ^ n8403 ;
  assign n8644 = n8643 ^ n8413 ;
  assign n8648 = n8647 ^ n8644 ;
  assign n8652 = n8651 ^ n8648 ;
  assign n8654 = n8647 ^ n8643 ;
  assign n8935 = n8651 ^ n8647 ;
  assign n8936 = ~n8654 & ~n8935 ;
  assign n8931 = x119 & n231 ;
  assign n8921 = x2 & x121 ;
  assign n8922 = n8921 ^ x122 ;
  assign n8923 = ~x1 & n8922 ;
  assign n8909 = ~x122 & ~n8386 ;
  assign n8908 = x122 & ~n8384 ;
  assign n8910 = n8909 ^ n8908 ;
  assign n8912 = x123 ^ x1 ;
  assign n8911 = x123 ^ x2 ;
  assign n8913 = n8912 ^ n8911 ;
  assign n8914 = n8910 & n8913 ;
  assign n8915 = n8914 ^ n8912 ;
  assign n8918 = n8915 ^ n8388 ;
  assign n8924 = n8923 ^ n8918 ;
  assign n8925 = ~x0 & n8924 ;
  assign n8926 = n8925 ^ n8915 ;
  assign n8927 = n8926 ^ x5 ;
  assign n8907 = x118 & n238 ;
  assign n8928 = n8927 ^ n8907 ;
  assign n8906 = x120 & n234 ;
  assign n8929 = n8928 ^ n8906 ;
  assign n8904 = n7846 ^ x120 ;
  assign n8905 = n235 & n8904 ;
  assign n8930 = n8929 ^ n8905 ;
  assign n8932 = n8931 ^ n8930 ;
  assign n8900 = n8636 ^ n8416 ;
  assign n8901 = n8642 & ~n8900 ;
  assign n8902 = n8901 ^ n8636 ;
  assign n8898 = x116 & n391 ;
  assign n8891 = x113 & n584 ;
  assign n8883 = n8619 ^ n8425 ;
  assign n8884 = n8625 & n8883 ;
  assign n8885 = n8884 ^ n8619 ;
  assign n8881 = x110 & n795 ;
  assign n8873 = n8612 ^ n8431 ;
  assign n8874 = n8618 & n8873 ;
  assign n8875 = n8874 ^ n8612 ;
  assign n8871 = x107 & n1068 ;
  assign n8864 = x104 & n1348 ;
  assign n8856 = n8595 ^ n8440 ;
  assign n8857 = n8601 & n8856 ;
  assign n8858 = n8857 ^ n8595 ;
  assign n8854 = x101 & n1673 ;
  assign n8846 = n8588 ^ n8446 ;
  assign n8847 = n8594 & n8846 ;
  assign n8848 = n8847 ^ n8588 ;
  assign n8844 = x98 & n2025 ;
  assign n8837 = x95 & n2435 ;
  assign n8835 = n2429 & n3336 ;
  assign n8831 = x94 & n2593 ;
  assign n8830 = x96 & n2428 ;
  assign n8832 = n8831 ^ n8830 ;
  assign n8833 = n8832 ^ x29 ;
  assign n8827 = x92 & n2899 ;
  assign n8819 = n8561 ^ n8458 ;
  assign n8820 = n8567 & n8819 ;
  assign n8821 = n8820 ^ n8561 ;
  assign n8817 = x89 & n3395 ;
  assign n8810 = x86 & n3940 ;
  assign n8802 = n8544 ^ n8467 ;
  assign n8803 = n8550 & n8802 ;
  assign n8804 = n8803 ^ n8544 ;
  assign n8800 = x83 & n4475 ;
  assign n8793 = x80 & n5121 ;
  assign n8784 = x71 & n7191 ;
  assign n8774 = x67 & n7954 ;
  assign n8773 = x69 & n7950 ;
  assign n8775 = n8774 ^ n8773 ;
  assign n8776 = n8775 ^ x56 ;
  assign n8772 = ~n376 & n7951 ;
  assign n8777 = n8776 ^ n8772 ;
  assign n8771 = x68 & n7947 ;
  assign n8778 = n8777 ^ n8771 ;
  assign n8762 = ~n8235 & ~n8505 ;
  assign n8763 = x59 & n8762 ;
  assign n8764 = n8763 ^ x59 ;
  assign n8759 = x66 & n8234 ;
  assign n8745 = x59 ^ x58 ;
  assign n8746 = n8234 & ~n8745 ;
  assign n8747 = n8746 ^ n8234 ;
  assign n8755 = x65 & n8747 ;
  assign n8748 = x59 ^ x57 ;
  assign n8749 = ~n8234 & n8748 ;
  assign n8750 = n8745 & n8749 ;
  assign n8756 = n8755 ^ n8750 ;
  assign n8757 = ~x64 & n8756 ;
  assign n8758 = n8757 ^ n8750 ;
  assign n8760 = n8759 ^ n8758 ;
  assign n8497 = x58 ^ x57 ;
  assign n8743 = ~n8234 & n8497 ;
  assign n8744 = x65 & n8743 ;
  assign n8761 = n8760 ^ n8744 ;
  assign n8765 = n8764 ^ n8761 ;
  assign n8766 = n8765 ^ n8515 ;
  assign n8767 = n8766 ^ n8505 ;
  assign n8768 = n8767 ^ n8765 ;
  assign n8769 = ~n8507 & n8768 ;
  assign n8770 = n8769 ^ n8766 ;
  assign n8779 = n8778 ^ n8770 ;
  assign n8780 = n8779 ^ x53 ;
  assign n8742 = x70 & n7183 ;
  assign n8781 = n8780 ^ n8742 ;
  assign n8741 = x72 & n7186 ;
  assign n8782 = n8781 ^ n8741 ;
  assign n8740 = n565 & n7187 ;
  assign n8783 = n8782 ^ n8740 ;
  assign n8785 = n8784 ^ n8783 ;
  assign n8737 = n8516 ^ n8491 ;
  assign n8738 = n8522 & n8737 ;
  assign n8739 = n8738 ^ n8516 ;
  assign n8786 = n8785 ^ n8739 ;
  assign n8727 = x73 & n6687 ;
  assign n8726 = x75 & n6444 ;
  assign n8728 = n8727 ^ n8726 ;
  assign n8729 = n8728 ^ x50 ;
  assign n8725 = ~n778 & n6445 ;
  assign n8730 = n8729 ^ n8725 ;
  assign n8724 = x74 & n6449 ;
  assign n8731 = n8730 ^ n8724 ;
  assign n8732 = n8731 ^ n8523 ;
  assign n8733 = n8732 ^ n8485 ;
  assign n8734 = n8733 ^ n8731 ;
  assign n8735 = n8529 & n8734 ;
  assign n8736 = n8735 ^ n8732 ;
  assign n8787 = n8786 ^ n8736 ;
  assign n8721 = n8530 ^ n8479 ;
  assign n8722 = n8536 & n8721 ;
  assign n8714 = x76 & n5981 ;
  assign n8713 = x78 & n5748 ;
  assign n8715 = n8714 ^ n8713 ;
  assign n8716 = n8715 ^ x47 ;
  assign n8712 = ~n1036 & n5749 ;
  assign n8717 = n8716 ^ n8712 ;
  assign n8711 = x77 & n5755 ;
  assign n8718 = n8717 ^ n8711 ;
  assign n8719 = n8718 ^ n8530 ;
  assign n8723 = n8722 ^ n8719 ;
  assign n8788 = n8787 ^ n8723 ;
  assign n8789 = n8788 ^ x44 ;
  assign n8710 = x79 & n5113 ;
  assign n8790 = n8789 ^ n8710 ;
  assign n8709 = x81 & n5116 ;
  assign n8791 = n8790 ^ n8709 ;
  assign n8708 = n1310 & n5117 ;
  assign n8792 = n8791 ^ n8708 ;
  assign n8794 = n8793 ^ n8792 ;
  assign n8705 = n8537 ^ n8473 ;
  assign n8706 = n8543 & n8705 ;
  assign n8707 = n8706 ^ n8537 ;
  assign n8795 = n8794 ^ n8707 ;
  assign n8796 = n8795 ^ x41 ;
  assign n8704 = x82 & n4482 ;
  assign n8797 = n8796 ^ n8704 ;
  assign n8703 = x84 & n4478 ;
  assign n8798 = n8797 ^ n8703 ;
  assign n8702 = n1635 & n4479 ;
  assign n8799 = n8798 ^ n8702 ;
  assign n8801 = n8800 ^ n8799 ;
  assign n8805 = n8804 ^ n8801 ;
  assign n8806 = n8805 ^ x38 ;
  assign n8701 = x85 & n3932 ;
  assign n8807 = n8806 ^ n8701 ;
  assign n8700 = x87 & n3935 ;
  assign n8808 = n8807 ^ n8700 ;
  assign n8699 = n1987 & n3936 ;
  assign n8809 = n8808 ^ n8699 ;
  assign n8811 = n8810 ^ n8809 ;
  assign n8696 = n8560 ^ n8551 ;
  assign n8697 = ~n8557 & n8696 ;
  assign n8698 = n8697 ^ n8560 ;
  assign n8812 = n8811 ^ n8698 ;
  assign n8813 = n8812 ^ x35 ;
  assign n8695 = x88 & n3387 ;
  assign n8814 = n8813 ^ n8695 ;
  assign n8694 = x90 & n3390 ;
  assign n8815 = n8814 ^ n8694 ;
  assign n8693 = n2398 & n3391 ;
  assign n8816 = n8815 ^ n8693 ;
  assign n8818 = n8817 ^ n8816 ;
  assign n8822 = n8821 ^ n8818 ;
  assign n8823 = n8822 ^ x32 ;
  assign n8692 = x91 & n2890 ;
  assign n8824 = n8823 ^ n8692 ;
  assign n8691 = x93 & n2893 ;
  assign n8825 = n8824 ^ n8691 ;
  assign n8690 = n2842 & n2894 ;
  assign n8826 = n8825 ^ n8690 ;
  assign n8828 = n8827 ^ n8826 ;
  assign n8687 = n8577 ^ n8568 ;
  assign n8688 = ~n8574 & n8687 ;
  assign n8689 = n8688 ^ n8577 ;
  assign n8829 = n8828 ^ n8689 ;
  assign n8834 = n8833 ^ n8829 ;
  assign n8836 = n8835 ^ n8834 ;
  assign n8838 = n8837 ^ n8836 ;
  assign n8684 = n8586 ^ n8452 ;
  assign n8685 = n8587 & n8684 ;
  assign n8686 = n8685 ^ n8586 ;
  assign n8839 = n8838 ^ n8686 ;
  assign n8840 = n8839 ^ x26 ;
  assign n8683 = x97 & n2032 ;
  assign n8841 = n8840 ^ n8683 ;
  assign n8682 = x99 & n2028 ;
  assign n8842 = n8841 ^ n8682 ;
  assign n8681 = n2029 & n3851 ;
  assign n8843 = n8842 ^ n8681 ;
  assign n8845 = n8844 ^ n8843 ;
  assign n8849 = n8848 ^ n8845 ;
  assign n8850 = n8849 ^ x23 ;
  assign n8680 = x100 & n1665 ;
  assign n8851 = n8850 ^ n8680 ;
  assign n8679 = x102 & n1668 ;
  assign n8852 = n8851 ^ n8679 ;
  assign n8678 = n1669 & n4425 ;
  assign n8853 = n8852 ^ n8678 ;
  assign n8855 = n8854 ^ n8853 ;
  assign n8859 = n8858 ^ n8855 ;
  assign n8860 = n8859 ^ x20 ;
  assign n8677 = x103 & n1340 ;
  assign n8861 = n8860 ^ n8677 ;
  assign n8676 = x105 & n1343 ;
  assign n8862 = n8861 ^ n8676 ;
  assign n8675 = n1344 & ~n5034 ;
  assign n8863 = n8862 ^ n8675 ;
  assign n8865 = n8864 ^ n8863 ;
  assign n8672 = n8611 ^ n8602 ;
  assign n8673 = ~n8608 & n8672 ;
  assign n8674 = n8673 ^ n8611 ;
  assign n8866 = n8865 ^ n8674 ;
  assign n8867 = n8866 ^ x17 ;
  assign n8671 = x106 & n1060 ;
  assign n8868 = n8867 ^ n8671 ;
  assign n8670 = x108 & n1063 ;
  assign n8869 = n8868 ^ n8670 ;
  assign n8669 = n1064 & n5687 ;
  assign n8870 = n8869 ^ n8669 ;
  assign n8872 = n8871 ^ n8870 ;
  assign n8876 = n8875 ^ n8872 ;
  assign n8877 = n8876 ^ x14 ;
  assign n8668 = x109 & n884 ;
  assign n8878 = n8877 ^ n8668 ;
  assign n8667 = x111 & n789 ;
  assign n8879 = n8878 ^ n8667 ;
  assign n8666 = n790 & ~n6370 ;
  assign n8880 = n8879 ^ n8666 ;
  assign n8882 = n8881 ^ n8880 ;
  assign n8886 = n8885 ^ n8882 ;
  assign n8887 = n8886 ^ x11 ;
  assign n8665 = x112 & n650 ;
  assign n8888 = n8887 ^ n8665 ;
  assign n8664 = x114 & ~n578 ;
  assign n8889 = n8888 ^ n8664 ;
  assign n8663 = ~n579 & ~n7108 ;
  assign n8890 = n8889 ^ n8663 ;
  assign n8892 = n8891 ^ n8890 ;
  assign n8660 = n8635 ^ n8626 ;
  assign n8661 = ~n8632 & n8660 ;
  assign n8662 = n8661 ^ n8635 ;
  assign n8893 = n8892 ^ n8662 ;
  assign n8894 = n8893 ^ x8 ;
  assign n8659 = x115 & n456 ;
  assign n8895 = n8894 ^ n8659 ;
  assign n8658 = x117 & n384 ;
  assign n8896 = n8895 ^ n8658 ;
  assign n8657 = n385 & ~n7860 ;
  assign n8897 = n8896 ^ n8657 ;
  assign n8899 = n8898 ^ n8897 ;
  assign n8903 = n8902 ^ n8899 ;
  assign n8933 = n8932 ^ n8903 ;
  assign n8653 = n8651 ^ n8403 ;
  assign n8655 = n8654 ^ n8653 ;
  assign n8656 = ~n8413 & ~n8655 ;
  assign n8934 = n8933 ^ n8656 ;
  assign n8937 = n8936 ^ n8934 ;
  assign n9227 = x117 & n391 ;
  assign n9219 = n8886 ^ n8662 ;
  assign n9220 = n8892 & n9219 ;
  assign n9221 = n9220 ^ n8886 ;
  assign n9217 = x114 & n584 ;
  assign n9210 = x111 & n795 ;
  assign n9203 = x108 & n1068 ;
  assign n9195 = n8859 ^ n8674 ;
  assign n9196 = n8865 & n9195 ;
  assign n9197 = n9196 ^ n8859 ;
  assign n9193 = x105 & n1348 ;
  assign n9186 = x102 & n1673 ;
  assign n9179 = x99 & n2025 ;
  assign n9171 = n8829 ^ n8686 ;
  assign n9172 = n8838 & n9171 ;
  assign n9173 = n9172 ^ n8829 ;
  assign n9165 = x95 & n2593 ;
  assign n9164 = x97 & n2428 ;
  assign n9166 = n9165 ^ n9164 ;
  assign n9167 = n9166 ^ x29 ;
  assign n9163 = n2429 & n3501 ;
  assign n9168 = n9167 ^ n9163 ;
  assign n9162 = x96 & n2435 ;
  assign n9169 = n9168 ^ n9162 ;
  assign n9158 = n8822 ^ n8689 ;
  assign n9159 = n8828 & n9158 ;
  assign n9160 = n9159 ^ n8822 ;
  assign n9156 = x93 & n2899 ;
  assign n9149 = x90 & n3395 ;
  assign n9141 = n8805 ^ n8698 ;
  assign n9142 = n8811 & n9141 ;
  assign n9143 = n9142 ^ n8805 ;
  assign n9139 = x87 & n3940 ;
  assign n9132 = x84 & n4475 ;
  assign n9125 = x81 & n5121 ;
  assign n9118 = x78 & n5755 ;
  assign n9111 = x75 & n6449 ;
  assign n9103 = n8779 ^ n8739 ;
  assign n9104 = n8785 & n9103 ;
  assign n9105 = n9104 ^ n8779 ;
  assign n9101 = x72 & n7191 ;
  assign n9093 = n8778 ^ n8765 ;
  assign n9094 = n8770 & n9093 ;
  assign n9095 = n9094 ^ n8765 ;
  assign n9091 = x69 & n7947 ;
  assign n9081 = x65 & n8750 ;
  assign n9080 = x66 & n8743 ;
  assign n9082 = n9081 ^ n9080 ;
  assign n9083 = n9082 ^ x59 ;
  assign n9077 = ~n155 & ~n8745 ;
  assign n9078 = n9077 ^ n295 ;
  assign n9079 = n8234 & ~n9078 ;
  assign n9084 = n9083 ^ n9079 ;
  assign n9069 = x60 ^ x59 ;
  assign n9070 = x64 & n9069 ;
  assign n9071 = ~n8761 & n8763 ;
  assign n9073 = ~n9070 & ~n9071 ;
  assign n9085 = n9084 ^ n9073 ;
  assign n9072 = n9071 ^ n9070 ;
  assign n9074 = n9073 ^ n9072 ;
  assign n9086 = n9085 ^ n9074 ;
  assign n9087 = n9086 ^ x56 ;
  assign n9068 = x68 & n7954 ;
  assign n9088 = n9087 ^ n9068 ;
  assign n9067 = x70 & n7950 ;
  assign n9089 = n9088 ^ n9067 ;
  assign n9066 = ~n443 & n7951 ;
  assign n9090 = n9089 ^ n9066 ;
  assign n9092 = n9091 ^ n9090 ;
  assign n9096 = n9095 ^ n9092 ;
  assign n9097 = n9096 ^ x53 ;
  assign n9065 = x71 & n7183 ;
  assign n9098 = n9097 ^ n9065 ;
  assign n9064 = x73 & n7186 ;
  assign n9099 = n9098 ^ n9064 ;
  assign n9063 = n636 & n7187 ;
  assign n9100 = n9099 ^ n9063 ;
  assign n9102 = n9101 ^ n9100 ;
  assign n9106 = n9105 ^ n9102 ;
  assign n9107 = n9106 ^ x50 ;
  assign n9062 = x74 & n6687 ;
  assign n9108 = n9107 ^ n9062 ;
  assign n9061 = x76 & n6444 ;
  assign n9109 = n9108 ^ n9061 ;
  assign n9060 = ~n863 & n6445 ;
  assign n9110 = n9109 ^ n9060 ;
  assign n9112 = n9111 ^ n9110 ;
  assign n9057 = n8786 ^ n8731 ;
  assign n9058 = n8736 & n9057 ;
  assign n9059 = n9058 ^ n8731 ;
  assign n9113 = n9112 ^ n9059 ;
  assign n9114 = n9113 ^ x47 ;
  assign n9056 = x77 & n5981 ;
  assign n9115 = n9114 ^ n9056 ;
  assign n9055 = x79 & n5748 ;
  assign n9116 = n9115 ^ n9055 ;
  assign n9054 = n1123 & n5749 ;
  assign n9117 = n9116 ^ n9054 ;
  assign n9119 = n9118 ^ n9117 ;
  assign n9051 = n8787 ^ n8718 ;
  assign n9052 = n8723 & n9051 ;
  assign n9053 = n9052 ^ n8718 ;
  assign n9120 = n9119 ^ n9053 ;
  assign n9121 = n9120 ^ x44 ;
  assign n9050 = x80 & n5113 ;
  assign n9122 = n9121 ^ n9050 ;
  assign n9049 = x82 & n5116 ;
  assign n9123 = n9122 ^ n9049 ;
  assign n9048 = n1422 & n5117 ;
  assign n9124 = n9123 ^ n9048 ;
  assign n9126 = n9125 ^ n9124 ;
  assign n9045 = n8788 ^ n8707 ;
  assign n9046 = n8794 & n9045 ;
  assign n9047 = n9046 ^ n8788 ;
  assign n9127 = n9126 ^ n9047 ;
  assign n9128 = n9127 ^ x41 ;
  assign n9044 = x83 & n4482 ;
  assign n9129 = n9128 ^ n9044 ;
  assign n9043 = x85 & n4478 ;
  assign n9130 = n9129 ^ n9043 ;
  assign n9042 = n1748 & n4479 ;
  assign n9131 = n9130 ^ n9042 ;
  assign n9133 = n9132 ^ n9131 ;
  assign n9039 = n8804 ^ n8795 ;
  assign n9040 = ~n8801 & n9039 ;
  assign n9041 = n9040 ^ n8804 ;
  assign n9134 = n9133 ^ n9041 ;
  assign n9135 = n9134 ^ x38 ;
  assign n9038 = x86 & n3932 ;
  assign n9136 = n9135 ^ n9038 ;
  assign n9037 = x88 & n3935 ;
  assign n9137 = n9136 ^ n9037 ;
  assign n9036 = n2131 & n3936 ;
  assign n9138 = n9137 ^ n9036 ;
  assign n9140 = n9139 ^ n9138 ;
  assign n9144 = n9143 ^ n9140 ;
  assign n9145 = n9144 ^ x35 ;
  assign n9035 = x89 & n3387 ;
  assign n9146 = n9145 ^ n9035 ;
  assign n9034 = x91 & n3390 ;
  assign n9147 = n9146 ^ n9034 ;
  assign n9033 = n2548 & n3391 ;
  assign n9148 = n9147 ^ n9033 ;
  assign n9150 = n9149 ^ n9148 ;
  assign n9030 = n8821 ^ n8812 ;
  assign n9031 = ~n8818 & n9030 ;
  assign n9032 = n9031 ^ n8821 ;
  assign n9151 = n9150 ^ n9032 ;
  assign n9152 = n9151 ^ x32 ;
  assign n9029 = x92 & n2890 ;
  assign n9153 = n9152 ^ n9029 ;
  assign n9028 = x94 & n2893 ;
  assign n9154 = n9153 ^ n9028 ;
  assign n9027 = n2894 & n3010 ;
  assign n9155 = n9154 ^ n9027 ;
  assign n9157 = n9156 ^ n9155 ;
  assign n9161 = n9160 ^ n9157 ;
  assign n9170 = n9169 ^ n9161 ;
  assign n9174 = n9173 ^ n9170 ;
  assign n9175 = n9174 ^ x26 ;
  assign n9026 = x98 & n2032 ;
  assign n9176 = n9175 ^ n9026 ;
  assign n9025 = x100 & n2028 ;
  assign n9177 = n9176 ^ n9025 ;
  assign n9024 = n2029 & n4048 ;
  assign n9178 = n9177 ^ n9024 ;
  assign n9180 = n9179 ^ n9178 ;
  assign n9021 = n8848 ^ n8839 ;
  assign n9022 = ~n8845 & n9021 ;
  assign n9023 = n9022 ^ n8848 ;
  assign n9181 = n9180 ^ n9023 ;
  assign n9182 = n9181 ^ x23 ;
  assign n9020 = x101 & n1665 ;
  assign n9183 = n9182 ^ n9020 ;
  assign n9019 = x103 & n1668 ;
  assign n9184 = n9183 ^ n9019 ;
  assign n9018 = n1669 & ~n4624 ;
  assign n9185 = n9184 ^ n9018 ;
  assign n9187 = n9186 ^ n9185 ;
  assign n9015 = n8858 ^ n8849 ;
  assign n9016 = ~n8855 & n9015 ;
  assign n9017 = n9016 ^ n8858 ;
  assign n9188 = n9187 ^ n9017 ;
  assign n9189 = n9188 ^ x20 ;
  assign n9014 = x104 & n1340 ;
  assign n9190 = n9189 ^ n9014 ;
  assign n9013 = x106 & n1343 ;
  assign n9191 = n9190 ^ n9013 ;
  assign n9012 = n1344 & ~n5257 ;
  assign n9192 = n9191 ^ n9012 ;
  assign n9194 = n9193 ^ n9192 ;
  assign n9198 = n9197 ^ n9194 ;
  assign n9199 = n9198 ^ x17 ;
  assign n9011 = x107 & n1060 ;
  assign n9200 = n9199 ^ n9011 ;
  assign n9010 = x109 & n1063 ;
  assign n9201 = n9200 ^ n9010 ;
  assign n9009 = n1064 & n5912 ;
  assign n9202 = n9201 ^ n9009 ;
  assign n9204 = n9203 ^ n9202 ;
  assign n9006 = n8875 ^ n8866 ;
  assign n9007 = ~n8872 & n9006 ;
  assign n9008 = n9007 ^ n8875 ;
  assign n9205 = n9204 ^ n9008 ;
  assign n9206 = n9205 ^ x14 ;
  assign n9005 = x110 & n884 ;
  assign n9207 = n9206 ^ n9005 ;
  assign n9004 = x112 & n789 ;
  assign n9208 = n9207 ^ n9004 ;
  assign n9003 = n790 & ~n6616 ;
  assign n9209 = n9208 ^ n9003 ;
  assign n9211 = n9210 ^ n9209 ;
  assign n9000 = n8885 ^ n8876 ;
  assign n9001 = ~n8882 & n9000 ;
  assign n9002 = n9001 ^ n8885 ;
  assign n9212 = n9211 ^ n9002 ;
  assign n9213 = n9212 ^ x11 ;
  assign n8999 = x113 & n650 ;
  assign n9214 = n9213 ^ n8999 ;
  assign n8998 = x115 & ~n578 ;
  assign n9215 = n9214 ^ n8998 ;
  assign n8997 = ~n579 & ~n7353 ;
  assign n9216 = n9215 ^ n8997 ;
  assign n9218 = n9217 ^ n9216 ;
  assign n9222 = n9221 ^ n9218 ;
  assign n9223 = n9222 ^ x8 ;
  assign n8996 = x116 & n456 ;
  assign n9224 = n9223 ^ n8996 ;
  assign n8995 = x118 & n384 ;
  assign n9225 = n9224 ^ n8995 ;
  assign n8994 = n385 & ~n8140 ;
  assign n9226 = n9225 ^ n8994 ;
  assign n9228 = n9227 ^ n9226 ;
  assign n8991 = n8902 ^ n8893 ;
  assign n8992 = ~n8899 & n8991 ;
  assign n8993 = n8992 ^ n8902 ;
  assign n9229 = n9228 ^ n8993 ;
  assign n8988 = n8926 ^ n8903 ;
  assign n8989 = n8932 & n8988 ;
  assign n8990 = n8989 ^ n8926 ;
  assign n9230 = n9229 ^ n8990 ;
  assign n8982 = x119 & n238 ;
  assign n8981 = x121 & n234 ;
  assign n8983 = n8982 ^ n8981 ;
  assign n8984 = n8983 ^ x5 ;
  assign n8979 = n8122 ^ x121 ;
  assign n8980 = n235 & n8979 ;
  assign n8985 = n8984 ^ n8980 ;
  assign n8978 = x120 & n231 ;
  assign n8986 = n8985 ^ n8978 ;
  assign n8972 = x2 & x122 ;
  assign n8973 = n8972 ^ x123 ;
  assign n8974 = ~x1 & n8973 ;
  assign n8961 = x123 ^ x122 ;
  assign n8962 = n8910 & n8961 ;
  assign n8964 = x124 ^ x1 ;
  assign n8963 = x124 ^ x2 ;
  assign n8965 = n8964 ^ n8963 ;
  assign n8966 = ~n8962 & n8965 ;
  assign n8967 = n8966 ^ n8964 ;
  assign n8969 = n8967 ^ n8911 ;
  assign n8975 = n8974 ^ n8969 ;
  assign n8976 = ~x0 & n8975 ;
  assign n8977 = n8976 ^ n8967 ;
  assign n8987 = n8986 ^ n8977 ;
  assign n9231 = n9230 ^ n8987 ;
  assign n8938 = n8403 & n8412 ;
  assign n8939 = n8938 ^ n8413 ;
  assign n8940 = n8643 & ~n8939 ;
  assign n8941 = n8647 & ~n8940 ;
  assign n8942 = ~n8643 & n8938 ;
  assign n8943 = n8942 ^ n8644 ;
  assign n8944 = n8941 & ~n8943 ;
  assign n8945 = n8944 ^ n8940 ;
  assign n8946 = ~n8647 & n8942 ;
  assign n8947 = n8933 & ~n8946 ;
  assign n8948 = ~n8945 & n8947 ;
  assign n8950 = n8948 ^ n8651 ;
  assign n8952 = n8933 ^ n8647 ;
  assign n8951 = n8933 ^ n8643 ;
  assign n8953 = n8952 ^ n8951 ;
  assign n8954 = n8933 ^ n8412 ;
  assign n8955 = n8954 ^ n8951 ;
  assign n8956 = n8953 & ~n8955 ;
  assign n8957 = n8956 ^ n8951 ;
  assign n8958 = n8648 & ~n8957 ;
  assign n8959 = ~n8950 & n8958 ;
  assign n8949 = n8948 ^ n8946 ;
  assign n8960 = n8959 ^ n8949 ;
  assign n9232 = n9231 ^ n8960 ;
  assign n9526 = n9222 ^ n8993 ;
  assign n9527 = n9228 & n9526 ;
  assign n9528 = n9527 ^ n9222 ;
  assign n9522 = x115 & n584 ;
  assign n9514 = n9205 ^ n9002 ;
  assign n9515 = n9211 & n9514 ;
  assign n9516 = n9515 ^ n9205 ;
  assign n9512 = x112 & n795 ;
  assign n9504 = n9198 ^ n9008 ;
  assign n9505 = n9204 & n9504 ;
  assign n9506 = n9505 ^ n9198 ;
  assign n9502 = x109 & n1068 ;
  assign n9495 = x106 & n1348 ;
  assign n9487 = n9181 ^ n9017 ;
  assign n9488 = n9187 & n9487 ;
  assign n9489 = n9488 ^ n9181 ;
  assign n9485 = x103 & n1673 ;
  assign n9477 = n9174 ^ n9023 ;
  assign n9478 = n9180 & n9477 ;
  assign n9479 = n9478 ^ n9174 ;
  assign n9475 = x100 & n2025 ;
  assign n9468 = x97 & n2435 ;
  assign n9466 = n2429 & n3673 ;
  assign n9462 = x96 & n2593 ;
  assign n9461 = x98 & n2428 ;
  assign n9463 = n9462 ^ n9461 ;
  assign n9464 = n9463 ^ x29 ;
  assign n9458 = x94 & n2899 ;
  assign n9450 = n9144 ^ n9032 ;
  assign n9451 = n9150 & n9450 ;
  assign n9452 = n9451 ^ n9144 ;
  assign n9448 = x91 & n3395 ;
  assign n9441 = x88 & n3940 ;
  assign n9433 = n9127 ^ n9041 ;
  assign n9434 = n9133 & n9433 ;
  assign n9435 = n9434 ^ n9127 ;
  assign n9431 = x85 & n4475 ;
  assign n9424 = x82 & n5121 ;
  assign n9417 = x79 & n5755 ;
  assign n9409 = x73 & n7191 ;
  assign n9398 = x69 & n7954 ;
  assign n9397 = x71 & n7950 ;
  assign n9399 = n9398 ^ n9397 ;
  assign n9400 = n9399 ^ x56 ;
  assign n9396 = ~n495 & n7951 ;
  assign n9401 = n9400 ^ n9396 ;
  assign n9395 = x70 & n7947 ;
  assign n9402 = n9401 ^ n9395 ;
  assign n9392 = ~n9073 & n9084 ;
  assign n9389 = x65 ^ x60 ;
  assign n9390 = n9069 & ~n9389 ;
  assign n9385 = x59 & x60 ;
  assign n9386 = n9385 ^ x61 ;
  assign n9387 = ~x64 & n9386 ;
  assign n9381 = x61 ^ x59 ;
  assign n9388 = n9387 ^ n9381 ;
  assign n9391 = n9390 ^ n9388 ;
  assign n9393 = n9392 ^ n9391 ;
  assign n9377 = ~n351 & n8747 ;
  assign n9376 = x67 & n8743 ;
  assign n9378 = n9377 ^ n9376 ;
  assign n9374 = x66 & n8750 ;
  assign n9373 = x68 & n8746 ;
  assign n9375 = n9374 ^ n9373 ;
  assign n9379 = n9378 ^ n9375 ;
  assign n9380 = n9379 ^ x59 ;
  assign n9394 = n9393 ^ n9380 ;
  assign n9403 = n9402 ^ n9394 ;
  assign n9370 = n9095 ^ n9086 ;
  assign n9371 = ~n9092 & n9370 ;
  assign n9372 = n9371 ^ n9095 ;
  assign n9404 = n9403 ^ n9372 ;
  assign n9405 = n9404 ^ x53 ;
  assign n9369 = x72 & n7183 ;
  assign n9406 = n9405 ^ n9369 ;
  assign n9368 = x74 & n7186 ;
  assign n9407 = n9406 ^ n9368 ;
  assign n9367 = n708 & n7187 ;
  assign n9408 = n9407 ^ n9367 ;
  assign n9410 = n9409 ^ n9408 ;
  assign n9364 = n9105 ^ n9096 ;
  assign n9365 = ~n9102 & n9364 ;
  assign n9366 = n9365 ^ n9105 ;
  assign n9411 = n9410 ^ n9366 ;
  assign n9354 = x75 & n6687 ;
  assign n9353 = x77 & n6444 ;
  assign n9355 = n9354 ^ n9353 ;
  assign n9356 = n9355 ^ x50 ;
  assign n9352 = ~n943 & n6445 ;
  assign n9357 = n9356 ^ n9352 ;
  assign n9351 = x76 & n6449 ;
  assign n9358 = n9357 ^ n9351 ;
  assign n9359 = n9358 ^ n9106 ;
  assign n9360 = n9359 ^ n9059 ;
  assign n9361 = n9360 ^ n9358 ;
  assign n9362 = n9112 & n9361 ;
  assign n9363 = n9362 ^ n9359 ;
  assign n9412 = n9411 ^ n9363 ;
  assign n9413 = n9412 ^ x47 ;
  assign n9350 = x78 & n5981 ;
  assign n9414 = n9413 ^ n9350 ;
  assign n9349 = x80 & n5748 ;
  assign n9415 = n9414 ^ n9349 ;
  assign n9348 = n1217 & n5749 ;
  assign n9416 = n9415 ^ n9348 ;
  assign n9418 = n9417 ^ n9416 ;
  assign n9345 = n9113 ^ n9053 ;
  assign n9346 = n9119 & n9345 ;
  assign n9347 = n9346 ^ n9113 ;
  assign n9419 = n9418 ^ n9347 ;
  assign n9420 = n9419 ^ x44 ;
  assign n9344 = x81 & n5113 ;
  assign n9421 = n9420 ^ n9344 ;
  assign n9343 = x83 & n5116 ;
  assign n9422 = n9421 ^ n9343 ;
  assign n9342 = n1517 & n5117 ;
  assign n9423 = n9422 ^ n9342 ;
  assign n9425 = n9424 ^ n9423 ;
  assign n9339 = n9120 ^ n9047 ;
  assign n9340 = n9126 & n9339 ;
  assign n9341 = n9340 ^ n9120 ;
  assign n9426 = n9425 ^ n9341 ;
  assign n9427 = n9426 ^ x41 ;
  assign n9338 = x84 & n4482 ;
  assign n9428 = n9427 ^ n9338 ;
  assign n9337 = x86 & n4478 ;
  assign n9429 = n9428 ^ n9337 ;
  assign n9336 = n1868 & n4479 ;
  assign n9430 = n9429 ^ n9336 ;
  assign n9432 = n9431 ^ n9430 ;
  assign n9436 = n9435 ^ n9432 ;
  assign n9437 = n9436 ^ x38 ;
  assign n9335 = x87 & n3932 ;
  assign n9438 = n9437 ^ n9335 ;
  assign n9334 = x89 & n3935 ;
  assign n9439 = n9438 ^ n9334 ;
  assign n9333 = n2255 & n3936 ;
  assign n9440 = n9439 ^ n9333 ;
  assign n9442 = n9441 ^ n9440 ;
  assign n9330 = n9143 ^ n9134 ;
  assign n9331 = ~n9140 & n9330 ;
  assign n9332 = n9331 ^ n9143 ;
  assign n9443 = n9442 ^ n9332 ;
  assign n9444 = n9443 ^ x35 ;
  assign n9329 = x90 & n3387 ;
  assign n9445 = n9444 ^ n9329 ;
  assign n9328 = x92 & n3390 ;
  assign n9446 = n9445 ^ n9328 ;
  assign n9327 = n2696 & n3391 ;
  assign n9447 = n9446 ^ n9327 ;
  assign n9449 = n9448 ^ n9447 ;
  assign n9453 = n9452 ^ n9449 ;
  assign n9454 = n9453 ^ x32 ;
  assign n9326 = x93 & n2890 ;
  assign n9455 = n9454 ^ n9326 ;
  assign n9325 = x95 & n2893 ;
  assign n9456 = n9455 ^ n9325 ;
  assign n9324 = n2894 & n3166 ;
  assign n9457 = n9456 ^ n9324 ;
  assign n9459 = n9458 ^ n9457 ;
  assign n9321 = n9160 ^ n9151 ;
  assign n9322 = ~n9157 & n9321 ;
  assign n9323 = n9322 ^ n9160 ;
  assign n9460 = n9459 ^ n9323 ;
  assign n9465 = n9464 ^ n9460 ;
  assign n9467 = n9466 ^ n9465 ;
  assign n9469 = n9468 ^ n9467 ;
  assign n9318 = n9173 ^ n9169 ;
  assign n9319 = ~n9170 & n9318 ;
  assign n9320 = n9319 ^ n9173 ;
  assign n9470 = n9469 ^ n9320 ;
  assign n9471 = n9470 ^ x26 ;
  assign n9317 = x99 & n2032 ;
  assign n9472 = n9471 ^ n9317 ;
  assign n9316 = x101 & n2028 ;
  assign n9473 = n9472 ^ n9316 ;
  assign n9315 = n2029 & n4223 ;
  assign n9474 = n9473 ^ n9315 ;
  assign n9476 = n9475 ^ n9474 ;
  assign n9480 = n9479 ^ n9476 ;
  assign n9481 = n9480 ^ x23 ;
  assign n9314 = x102 & n1665 ;
  assign n9482 = n9481 ^ n9314 ;
  assign n9313 = x104 & n1668 ;
  assign n9483 = n9482 ^ n9313 ;
  assign n9312 = n1669 & ~n4830 ;
  assign n9484 = n9483 ^ n9312 ;
  assign n9486 = n9485 ^ n9484 ;
  assign n9490 = n9489 ^ n9486 ;
  assign n9491 = n9490 ^ x20 ;
  assign n9311 = x105 & n1340 ;
  assign n9492 = n9491 ^ n9311 ;
  assign n9310 = x107 & n1343 ;
  assign n9493 = n9492 ^ n9310 ;
  assign n9309 = n1344 & ~n5459 ;
  assign n9494 = n9493 ^ n9309 ;
  assign n9496 = n9495 ^ n9494 ;
  assign n9306 = n9197 ^ n9188 ;
  assign n9307 = ~n9194 & n9306 ;
  assign n9308 = n9307 ^ n9197 ;
  assign n9497 = n9496 ^ n9308 ;
  assign n9498 = n9497 ^ x17 ;
  assign n9305 = x108 & n1060 ;
  assign n9499 = n9498 ^ n9305 ;
  assign n9304 = x110 & n1063 ;
  assign n9500 = n9499 ^ n9304 ;
  assign n9303 = n1064 & n6145 ;
  assign n9501 = n9500 ^ n9303 ;
  assign n9503 = n9502 ^ n9501 ;
  assign n9507 = n9506 ^ n9503 ;
  assign n9508 = n9507 ^ x14 ;
  assign n9302 = x111 & n884 ;
  assign n9509 = n9508 ^ n9302 ;
  assign n9301 = x113 & n789 ;
  assign n9510 = n9509 ^ n9301 ;
  assign n9300 = n790 & ~n6849 ;
  assign n9511 = n9510 ^ n9300 ;
  assign n9513 = n9512 ^ n9511 ;
  assign n9517 = n9516 ^ n9513 ;
  assign n9518 = n9517 ^ x11 ;
  assign n9299 = x114 & n650 ;
  assign n9519 = n9518 ^ n9299 ;
  assign n9298 = x116 & ~n578 ;
  assign n9520 = n9519 ^ n9298 ;
  assign n9297 = ~n579 & ~n7604 ;
  assign n9521 = n9520 ^ n9297 ;
  assign n9523 = n9522 ^ n9521 ;
  assign n9294 = n9221 ^ n9212 ;
  assign n9295 = ~n9218 & n9294 ;
  assign n9296 = n9295 ^ n9221 ;
  assign n9524 = n9523 ^ n9296 ;
  assign n9287 = x2 & x123 ;
  assign n9288 = n9287 ^ x124 ;
  assign n9289 = ~x1 & n9288 ;
  assign n9270 = ~x124 & n8909 ;
  assign n9271 = ~x123 & x124 ;
  assign n9272 = n8908 & n9271 ;
  assign n9273 = n9272 ^ x123 ;
  assign n9274 = n9270 & n9273 ;
  assign n9275 = n9274 ^ n9273 ;
  assign n9276 = n9275 ^ x124 ;
  assign n9277 = x125 ^ x1 ;
  assign n9278 = n9277 ^ x2 ;
  assign n9279 = n9278 ^ x125 ;
  assign n9280 = ~n9276 & n9279 ;
  assign n9281 = n9280 ^ n9277 ;
  assign n9284 = n9281 ^ n8963 ;
  assign n9290 = n9289 ^ n9284 ;
  assign n9291 = ~x0 & n9290 ;
  assign n9292 = n9291 ^ n9281 ;
  assign n9264 = x120 & n238 ;
  assign n9263 = x122 & n234 ;
  assign n9265 = n9264 ^ n9263 ;
  assign n9266 = n9265 ^ x5 ;
  assign n9261 = n8387 ^ x122 ;
  assign n9262 = n235 & ~n9261 ;
  assign n9267 = n9266 ^ n9262 ;
  assign n9260 = x121 & n231 ;
  assign n9268 = n9267 ^ n9260 ;
  assign n9255 = x117 & n456 ;
  assign n9254 = x119 & n384 ;
  assign n9256 = n9255 ^ n9254 ;
  assign n9257 = n9256 ^ x8 ;
  assign n9253 = n385 & n8405 ;
  assign n9258 = n9257 ^ n9253 ;
  assign n9252 = x118 & n391 ;
  assign n9259 = n9258 ^ n9252 ;
  assign n9269 = n9268 ^ n9259 ;
  assign n9293 = n9292 ^ n9269 ;
  assign n9525 = n9524 ^ n9293 ;
  assign n9529 = n9528 ^ n9525 ;
  assign n9234 = n8977 & n8986 ;
  assign n9233 = ~n8990 & ~n9229 ;
  assign n9237 = n9233 ^ n9230 ;
  assign n9238 = n9234 & ~n9237 ;
  assign n9235 = n9234 ^ n8987 ;
  assign n9236 = n9233 & ~n9235 ;
  assign n9239 = n9238 ^ n9236 ;
  assign n9240 = n9235 ^ n9229 ;
  assign n9241 = n9235 ^ n8990 ;
  assign n9242 = n9240 & ~n9241 ;
  assign n9243 = n9242 ^ n9229 ;
  assign n9244 = ~n9234 & ~n9243 ;
  assign n9245 = n9244 ^ n8960 ;
  assign n9246 = n9245 ^ n9244 ;
  assign n9247 = n9244 ^ n9231 ;
  assign n9248 = n9247 ^ n9244 ;
  assign n9249 = n9246 & n9248 ;
  assign n9250 = n9249 ^ n9244 ;
  assign n9251 = ~n9239 & ~n9250 ;
  assign n9530 = n9529 ^ n9251 ;
  assign n9830 = n9239 ^ n9231 ;
  assign n9831 = n9830 ^ n9244 ;
  assign n9829 = ~n9236 & n9529 ;
  assign n9832 = n9831 ^ n9829 ;
  assign n9833 = ~n8960 & n9832 ;
  assign n9834 = n9529 ^ n9237 ;
  assign n9835 = n9834 ^ n9234 ;
  assign n9836 = n9833 & ~n9835 ;
  assign n9837 = n9836 ^ n9832 ;
  assign n9838 = n9243 & n9529 ;
  assign n9839 = ~n9837 & n9838 ;
  assign n9840 = n9839 ^ n9837 ;
  assign n9532 = n9524 ^ n9259 ;
  assign n9531 = n9528 ^ n9268 ;
  assign n9533 = n9532 ^ n9531 ;
  assign n9818 = x119 & n391 ;
  assign n9815 = x120 & n384 ;
  assign n9813 = x118 & n456 ;
  assign n9807 = x121 & n238 ;
  assign n9806 = x123 & n234 ;
  assign n9808 = n9807 ^ n9806 ;
  assign n9809 = n9808 ^ x5 ;
  assign n9804 = n8910 ^ x123 ;
  assign n9805 = n235 & ~n9804 ;
  assign n9810 = n9809 ^ n9805 ;
  assign n9803 = x122 & n231 ;
  assign n9811 = n9810 ^ n9803 ;
  assign n9812 = n9811 ^ x8 ;
  assign n9814 = n9813 ^ n9812 ;
  assign n9816 = n9815 ^ n9814 ;
  assign n9802 = n385 & n8904 ;
  assign n9817 = n9816 ^ n9802 ;
  assign n9819 = n9818 ^ n9817 ;
  assign n9798 = n9517 ^ n9296 ;
  assign n9799 = n9523 & n9798 ;
  assign n9800 = n9799 ^ n9517 ;
  assign n9796 = x116 & n584 ;
  assign n9789 = x113 & n795 ;
  assign n9782 = x110 & n1068 ;
  assign n9774 = n9490 ^ n9308 ;
  assign n9775 = n9496 & n9774 ;
  assign n9776 = n9775 ^ n9490 ;
  assign n9772 = x107 & n1348 ;
  assign n9765 = x104 & n1673 ;
  assign n9758 = x101 & n2025 ;
  assign n9750 = n9460 ^ n9320 ;
  assign n9751 = n9469 & n9750 ;
  assign n9752 = n9751 ^ n9460 ;
  assign n9744 = x97 & n2593 ;
  assign n9743 = x99 & n2428 ;
  assign n9745 = n9744 ^ n9743 ;
  assign n9746 = n9745 ^ x29 ;
  assign n9742 = n2429 & n3851 ;
  assign n9747 = n9746 ^ n9742 ;
  assign n9741 = x98 & n2435 ;
  assign n9748 = n9747 ^ n9741 ;
  assign n9737 = n9453 ^ n9323 ;
  assign n9738 = n9459 & n9737 ;
  assign n9739 = n9738 ^ n9453 ;
  assign n9735 = x95 & n2899 ;
  assign n9728 = x92 & n3395 ;
  assign n9720 = n9436 ^ n9332 ;
  assign n9721 = n9442 & n9720 ;
  assign n9722 = n9721 ^ n9436 ;
  assign n9718 = x89 & n3940 ;
  assign n9711 = x86 & n4475 ;
  assign n9704 = x83 & n5121 ;
  assign n9696 = n9412 ^ n9347 ;
  assign n9697 = n9418 & n9696 ;
  assign n9698 = n9697 ^ n9412 ;
  assign n9689 = n9402 ^ n9372 ;
  assign n9690 = n9403 & n9689 ;
  assign n9691 = n9690 ^ n9402 ;
  assign n9687 = x71 & n7947 ;
  assign n9680 = n9391 ^ n9380 ;
  assign n9681 = ~n9393 & n9680 ;
  assign n9675 = ~n376 & n8747 ;
  assign n9674 = x68 & n8743 ;
  assign n9676 = n9675 ^ n9674 ;
  assign n9672 = x67 & n8750 ;
  assign n9671 = x69 & n8746 ;
  assign n9673 = n9672 ^ n9671 ;
  assign n9677 = n9676 ^ n9673 ;
  assign n9667 = ~n9070 & ~n9391 ;
  assign n9668 = x62 & n9667 ;
  assign n9669 = n9668 ^ x62 ;
  assign n9664 = x66 & n9069 ;
  assign n9650 = x62 ^ x61 ;
  assign n9651 = n9069 & ~n9650 ;
  assign n9652 = n9651 ^ n9069 ;
  assign n9660 = x65 & n9652 ;
  assign n9653 = x62 ^ x60 ;
  assign n9654 = ~n9069 & n9653 ;
  assign n9655 = n9650 & n9654 ;
  assign n9661 = n9660 ^ n9655 ;
  assign n9662 = ~x64 & n9661 ;
  assign n9663 = n9662 ^ n9655 ;
  assign n9665 = n9664 ^ n9663 ;
  assign n9383 = x61 ^ x60 ;
  assign n9648 = ~n9069 & n9383 ;
  assign n9649 = x65 & n9648 ;
  assign n9666 = n9665 ^ n9649 ;
  assign n9670 = n9669 ^ n9666 ;
  assign n9678 = n9677 ^ n9670 ;
  assign n9679 = n9678 ^ n9379 ;
  assign n9682 = n9681 ^ n9679 ;
  assign n9683 = n9682 ^ x56 ;
  assign n9647 = x70 & n7954 ;
  assign n9684 = n9683 ^ n9647 ;
  assign n9646 = x72 & n7950 ;
  assign n9685 = n9684 ^ n9646 ;
  assign n9645 = n565 & n7951 ;
  assign n9686 = n9685 ^ n9645 ;
  assign n9688 = n9687 ^ n9686 ;
  assign n9692 = n9691 ^ n9688 ;
  assign n9642 = n9404 ^ n9366 ;
  assign n9643 = n9410 & n9642 ;
  assign n9635 = x73 & n7183 ;
  assign n9634 = x75 & n7186 ;
  assign n9636 = n9635 ^ n9634 ;
  assign n9637 = n9636 ^ x53 ;
  assign n9633 = ~n778 & n7187 ;
  assign n9638 = n9637 ^ n9633 ;
  assign n9632 = x74 & n7191 ;
  assign n9639 = n9638 ^ n9632 ;
  assign n9640 = n9639 ^ n9404 ;
  assign n9644 = n9643 ^ n9640 ;
  assign n9693 = n9692 ^ n9644 ;
  assign n9626 = x79 & n5981 ;
  assign n9625 = x81 & n5748 ;
  assign n9627 = n9626 ^ n9625 ;
  assign n9628 = n9627 ^ x47 ;
  assign n9624 = n1310 & n5749 ;
  assign n9629 = n9628 ^ n9624 ;
  assign n9623 = x80 & n5755 ;
  assign n9630 = n9629 ^ n9623 ;
  assign n9618 = x76 & n6687 ;
  assign n9617 = x78 & n6444 ;
  assign n9619 = n9618 ^ n9617 ;
  assign n9620 = n9619 ^ x50 ;
  assign n9616 = ~n1036 & n6445 ;
  assign n9621 = n9620 ^ n9616 ;
  assign n9615 = x77 & n6449 ;
  assign n9622 = n9621 ^ n9615 ;
  assign n9631 = n9630 ^ n9622 ;
  assign n9694 = n9693 ^ n9631 ;
  assign n9612 = n9411 ^ n9358 ;
  assign n9613 = n9363 & n9612 ;
  assign n9614 = n9613 ^ n9358 ;
  assign n9695 = n9694 ^ n9614 ;
  assign n9699 = n9698 ^ n9695 ;
  assign n9700 = n9699 ^ x44 ;
  assign n9611 = x82 & n5113 ;
  assign n9701 = n9700 ^ n9611 ;
  assign n9610 = x84 & n5116 ;
  assign n9702 = n9701 ^ n9610 ;
  assign n9609 = n1635 & n5117 ;
  assign n9703 = n9702 ^ n9609 ;
  assign n9705 = n9704 ^ n9703 ;
  assign n9606 = n9419 ^ n9341 ;
  assign n9607 = n9425 & n9606 ;
  assign n9608 = n9607 ^ n9419 ;
  assign n9706 = n9705 ^ n9608 ;
  assign n9707 = n9706 ^ x41 ;
  assign n9605 = x85 & n4482 ;
  assign n9708 = n9707 ^ n9605 ;
  assign n9604 = x87 & n4478 ;
  assign n9709 = n9708 ^ n9604 ;
  assign n9603 = n1987 & n4479 ;
  assign n9710 = n9709 ^ n9603 ;
  assign n9712 = n9711 ^ n9710 ;
  assign n9600 = n9435 ^ n9426 ;
  assign n9601 = ~n9432 & n9600 ;
  assign n9602 = n9601 ^ n9435 ;
  assign n9713 = n9712 ^ n9602 ;
  assign n9714 = n9713 ^ x38 ;
  assign n9599 = x88 & n3932 ;
  assign n9715 = n9714 ^ n9599 ;
  assign n9598 = x90 & n3935 ;
  assign n9716 = n9715 ^ n9598 ;
  assign n9597 = n2398 & n3936 ;
  assign n9717 = n9716 ^ n9597 ;
  assign n9719 = n9718 ^ n9717 ;
  assign n9723 = n9722 ^ n9719 ;
  assign n9724 = n9723 ^ x35 ;
  assign n9596 = x91 & n3387 ;
  assign n9725 = n9724 ^ n9596 ;
  assign n9595 = x93 & n3390 ;
  assign n9726 = n9725 ^ n9595 ;
  assign n9594 = n2842 & n3391 ;
  assign n9727 = n9726 ^ n9594 ;
  assign n9729 = n9728 ^ n9727 ;
  assign n9591 = n9452 ^ n9443 ;
  assign n9592 = ~n9449 & n9591 ;
  assign n9593 = n9592 ^ n9452 ;
  assign n9730 = n9729 ^ n9593 ;
  assign n9731 = n9730 ^ x32 ;
  assign n9590 = x94 & n2890 ;
  assign n9732 = n9731 ^ n9590 ;
  assign n9589 = x96 & n2893 ;
  assign n9733 = n9732 ^ n9589 ;
  assign n9588 = n2894 & n3336 ;
  assign n9734 = n9733 ^ n9588 ;
  assign n9736 = n9735 ^ n9734 ;
  assign n9740 = n9739 ^ n9736 ;
  assign n9749 = n9748 ^ n9740 ;
  assign n9753 = n9752 ^ n9749 ;
  assign n9754 = n9753 ^ x26 ;
  assign n9587 = x100 & n2032 ;
  assign n9755 = n9754 ^ n9587 ;
  assign n9586 = x102 & n2028 ;
  assign n9756 = n9755 ^ n9586 ;
  assign n9585 = n2029 & n4425 ;
  assign n9757 = n9756 ^ n9585 ;
  assign n9759 = n9758 ^ n9757 ;
  assign n9582 = n9479 ^ n9470 ;
  assign n9583 = ~n9476 & n9582 ;
  assign n9584 = n9583 ^ n9479 ;
  assign n9760 = n9759 ^ n9584 ;
  assign n9761 = n9760 ^ x23 ;
  assign n9581 = x103 & n1665 ;
  assign n9762 = n9761 ^ n9581 ;
  assign n9580 = x105 & n1668 ;
  assign n9763 = n9762 ^ n9580 ;
  assign n9579 = n1669 & ~n5034 ;
  assign n9764 = n9763 ^ n9579 ;
  assign n9766 = n9765 ^ n9764 ;
  assign n9576 = n9489 ^ n9480 ;
  assign n9577 = ~n9486 & n9576 ;
  assign n9578 = n9577 ^ n9489 ;
  assign n9767 = n9766 ^ n9578 ;
  assign n9768 = n9767 ^ x20 ;
  assign n9575 = x106 & n1340 ;
  assign n9769 = n9768 ^ n9575 ;
  assign n9574 = x108 & n1343 ;
  assign n9770 = n9769 ^ n9574 ;
  assign n9573 = n1344 & n5687 ;
  assign n9771 = n9770 ^ n9573 ;
  assign n9773 = n9772 ^ n9771 ;
  assign n9777 = n9776 ^ n9773 ;
  assign n9778 = n9777 ^ x17 ;
  assign n9572 = x109 & n1060 ;
  assign n9779 = n9778 ^ n9572 ;
  assign n9571 = x111 & n1063 ;
  assign n9780 = n9779 ^ n9571 ;
  assign n9570 = n1064 & ~n6370 ;
  assign n9781 = n9780 ^ n9570 ;
  assign n9783 = n9782 ^ n9781 ;
  assign n9567 = n9506 ^ n9497 ;
  assign n9568 = ~n9503 & n9567 ;
  assign n9569 = n9568 ^ n9506 ;
  assign n9784 = n9783 ^ n9569 ;
  assign n9785 = n9784 ^ x14 ;
  assign n9566 = x112 & n884 ;
  assign n9786 = n9785 ^ n9566 ;
  assign n9565 = x114 & n789 ;
  assign n9787 = n9786 ^ n9565 ;
  assign n9564 = n790 & ~n7108 ;
  assign n9788 = n9787 ^ n9564 ;
  assign n9790 = n9789 ^ n9788 ;
  assign n9561 = n9516 ^ n9507 ;
  assign n9562 = ~n9513 & n9561 ;
  assign n9563 = n9562 ^ n9516 ;
  assign n9791 = n9790 ^ n9563 ;
  assign n9792 = n9791 ^ x11 ;
  assign n9560 = x115 & n650 ;
  assign n9793 = n9792 ^ n9560 ;
  assign n9559 = x117 & ~n578 ;
  assign n9794 = n9793 ^ n9559 ;
  assign n9558 = ~n579 & ~n7860 ;
  assign n9795 = n9794 ^ n9558 ;
  assign n9797 = n9796 ^ n9795 ;
  assign n9801 = n9800 ^ n9797 ;
  assign n9820 = n9819 ^ n9801 ;
  assign n9539 = ~x124 & x125 ;
  assign n9542 = ~n9275 & n9539 ;
  assign n9537 = x125 ^ x124 ;
  assign n9540 = n9539 ^ n9537 ;
  assign n9541 = n9273 & n9540 ;
  assign n9543 = n9542 ^ n9541 ;
  assign n9545 = x126 ^ x1 ;
  assign n9544 = x126 ^ x2 ;
  assign n9546 = n9545 ^ n9544 ;
  assign n9547 = ~n9543 & n9546 ;
  assign n9548 = n9547 ^ n9545 ;
  assign n9821 = n9820 ^ n9548 ;
  assign n9553 = x2 & x124 ;
  assign n9554 = n9553 ^ x125 ;
  assign n9555 = ~n259 & n9554 ;
  assign n9549 = x125 ^ x2 ;
  assign n9550 = n9549 ^ n9548 ;
  assign n9556 = n9555 ^ n9550 ;
  assign n9557 = ~x0 & n9556 ;
  assign n9822 = n9821 ^ n9557 ;
  assign n9534 = n9528 ^ n9524 ;
  assign n9535 = ~n9532 & n9534 ;
  assign n9536 = n9535 ^ n9528 ;
  assign n9823 = n9822 ^ n9536 ;
  assign n9824 = n9823 ^ n9292 ;
  assign n9825 = n9824 ^ n9268 ;
  assign n9826 = n9825 ^ n9823 ;
  assign n9827 = ~n9533 & n9826 ;
  assign n9828 = n9827 ^ n9824 ;
  assign n9841 = n9840 ^ n9828 ;
  assign n10136 = n9820 ^ n9536 ;
  assign n10137 = n9822 & n10136 ;
  assign n10138 = n10137 ^ n9820 ;
  assign n10131 = x120 & n391 ;
  assign n10128 = x121 & n384 ;
  assign n10126 = x119 & n456 ;
  assign n10120 = x122 & n238 ;
  assign n10119 = x124 & n234 ;
  assign n10121 = n10120 ^ n10119 ;
  assign n10122 = n10121 ^ x5 ;
  assign n10117 = n8962 ^ x124 ;
  assign n10118 = n235 & n10117 ;
  assign n10123 = n10122 ^ n10118 ;
  assign n10116 = x123 & n231 ;
  assign n10124 = n10123 ^ n10116 ;
  assign n10125 = n10124 ^ x8 ;
  assign n10127 = n10126 ^ n10125 ;
  assign n10129 = n10128 ^ n10127 ;
  assign n10115 = n385 & n8979 ;
  assign n10130 = n10129 ^ n10115 ;
  assign n10132 = n10131 ^ n10130 ;
  assign n10112 = x117 & n584 ;
  assign n10104 = n9784 ^ n9563 ;
  assign n10105 = n9790 & n10104 ;
  assign n10106 = n10105 ^ n9784 ;
  assign n10102 = x114 & n795 ;
  assign n10094 = n9777 ^ n9569 ;
  assign n10095 = n9783 & n10094 ;
  assign n10096 = n10095 ^ n9777 ;
  assign n10092 = x111 & n1068 ;
  assign n10085 = x108 & n1348 ;
  assign n10077 = n9760 ^ n9578 ;
  assign n10078 = n9766 & n10077 ;
  assign n10079 = n10078 ^ n9760 ;
  assign n10075 = x105 & n1673 ;
  assign n10067 = n9753 ^ n9584 ;
  assign n10068 = n9759 & n10067 ;
  assign n10069 = n10068 ^ n9753 ;
  assign n10065 = x102 & n2025 ;
  assign n10058 = x99 & n2435 ;
  assign n10051 = x96 & n2899 ;
  assign n10043 = n9723 ^ n9593 ;
  assign n10044 = n9729 & n10043 ;
  assign n10045 = n10044 ^ n9723 ;
  assign n10041 = x93 & n3395 ;
  assign n10034 = x90 & n3940 ;
  assign n10026 = n9706 ^ n9602 ;
  assign n10027 = n9712 & n10026 ;
  assign n10028 = n10027 ^ n9706 ;
  assign n10024 = x87 & n4475 ;
  assign n10017 = x84 & n5121 ;
  assign n10010 = x81 & n5755 ;
  assign n10000 = x77 & n6687 ;
  assign n9999 = x79 & n6444 ;
  assign n10001 = n10000 ^ n9999 ;
  assign n10002 = n10001 ^ x50 ;
  assign n9998 = n1123 & n6445 ;
  assign n10003 = n10002 ^ n9998 ;
  assign n9997 = x78 & n6449 ;
  assign n10004 = n10003 ^ n9997 ;
  assign n9993 = x75 & n7191 ;
  assign n9976 = n9380 & ~n9679 ;
  assign n9977 = n9391 & n9392 ;
  assign n9978 = n9977 ^ n9393 ;
  assign n9979 = n9977 ^ n9670 ;
  assign n9980 = n9677 ^ x59 ;
  assign n9981 = n9980 ^ n9977 ;
  assign n9982 = n9979 & ~n9981 ;
  assign n9983 = n9982 ^ n9670 ;
  assign n9984 = n9978 & ~n9983 ;
  assign n9985 = n9976 & n9984 ;
  assign n9986 = n9985 ^ n9983 ;
  assign n9974 = x69 & n8743 ;
  assign n9964 = x65 & n9655 ;
  assign n9963 = x66 & n9648 ;
  assign n9965 = n9964 ^ n9963 ;
  assign n9960 = ~n155 & n9650 ;
  assign n9961 = n9960 ^ x67 ;
  assign n9962 = n9069 & n9961 ;
  assign n9966 = n9965 ^ n9962 ;
  assign n9967 = n9966 ^ x62 ;
  assign n9956 = x63 ^ x62 ;
  assign n9957 = x64 & n9956 ;
  assign n9968 = n9967 ^ n9957 ;
  assign n9955 = ~n9666 & n9668 ;
  assign n9969 = n9968 ^ n9955 ;
  assign n9970 = n9969 ^ x59 ;
  assign n9954 = x68 & n8750 ;
  assign n9971 = n9970 ^ n9954 ;
  assign n9953 = x70 & n8746 ;
  assign n9972 = n9971 ^ n9953 ;
  assign n9952 = ~n443 & n8747 ;
  assign n9973 = n9972 ^ n9952 ;
  assign n9975 = n9974 ^ n9973 ;
  assign n9987 = n9986 ^ n9975 ;
  assign n9942 = x71 & n7954 ;
  assign n9941 = x73 & n7950 ;
  assign n9943 = n9942 ^ n9941 ;
  assign n9944 = n9943 ^ x56 ;
  assign n9940 = n636 & n7951 ;
  assign n9945 = n9944 ^ n9940 ;
  assign n9939 = x72 & n7947 ;
  assign n9946 = n9945 ^ n9939 ;
  assign n9947 = n9946 ^ n9691 ;
  assign n9948 = n9947 ^ n9682 ;
  assign n9949 = n9948 ^ n9946 ;
  assign n9950 = ~n9688 & n9949 ;
  assign n9951 = n9950 ^ n9947 ;
  assign n9988 = n9987 ^ n9951 ;
  assign n9989 = n9988 ^ x53 ;
  assign n9938 = x74 & n7183 ;
  assign n9990 = n9989 ^ n9938 ;
  assign n9937 = x76 & n7186 ;
  assign n9991 = n9990 ^ n9937 ;
  assign n9936 = ~n863 & n7187 ;
  assign n9992 = n9991 ^ n9936 ;
  assign n9994 = n9993 ^ n9992 ;
  assign n9933 = n9692 ^ n9639 ;
  assign n9934 = n9644 & n9933 ;
  assign n9935 = n9934 ^ n9639 ;
  assign n9995 = n9994 ^ n9935 ;
  assign n9929 = n9693 ^ n9622 ;
  assign n9930 = n9622 ^ n9614 ;
  assign n9931 = n9929 & ~n9930 ;
  assign n9932 = n9931 ^ n9693 ;
  assign n9996 = n9995 ^ n9932 ;
  assign n10005 = n10004 ^ n9996 ;
  assign n10006 = n10005 ^ x47 ;
  assign n9928 = x80 & n5981 ;
  assign n10007 = n10006 ^ n9928 ;
  assign n9927 = x82 & n5748 ;
  assign n10008 = n10007 ^ n9927 ;
  assign n9926 = n1422 & n5749 ;
  assign n10009 = n10008 ^ n9926 ;
  assign n10011 = n10010 ^ n10009 ;
  assign n9923 = n9698 ^ n9630 ;
  assign n9924 = ~n9695 & n9923 ;
  assign n9925 = n9924 ^ n9698 ;
  assign n10012 = n10011 ^ n9925 ;
  assign n10013 = n10012 ^ x44 ;
  assign n9922 = x83 & n5113 ;
  assign n10014 = n10013 ^ n9922 ;
  assign n9921 = x85 & n5116 ;
  assign n10015 = n10014 ^ n9921 ;
  assign n9920 = n1748 & n5117 ;
  assign n10016 = n10015 ^ n9920 ;
  assign n10018 = n10017 ^ n10016 ;
  assign n9917 = n9699 ^ n9608 ;
  assign n9918 = n9705 & n9917 ;
  assign n9919 = n9918 ^ n9699 ;
  assign n10019 = n10018 ^ n9919 ;
  assign n10020 = n10019 ^ x41 ;
  assign n9916 = x86 & n4482 ;
  assign n10021 = n10020 ^ n9916 ;
  assign n9915 = x88 & n4478 ;
  assign n10022 = n10021 ^ n9915 ;
  assign n9914 = n2131 & n4479 ;
  assign n10023 = n10022 ^ n9914 ;
  assign n10025 = n10024 ^ n10023 ;
  assign n10029 = n10028 ^ n10025 ;
  assign n10030 = n10029 ^ x38 ;
  assign n9913 = x89 & n3932 ;
  assign n10031 = n10030 ^ n9913 ;
  assign n9912 = x91 & n3935 ;
  assign n10032 = n10031 ^ n9912 ;
  assign n9911 = n2548 & n3936 ;
  assign n10033 = n10032 ^ n9911 ;
  assign n10035 = n10034 ^ n10033 ;
  assign n9908 = n9722 ^ n9713 ;
  assign n9909 = ~n9719 & n9908 ;
  assign n9910 = n9909 ^ n9722 ;
  assign n10036 = n10035 ^ n9910 ;
  assign n10037 = n10036 ^ x35 ;
  assign n9907 = x92 & n3387 ;
  assign n10038 = n10037 ^ n9907 ;
  assign n9906 = x94 & n3390 ;
  assign n10039 = n10038 ^ n9906 ;
  assign n9905 = n3010 & n3391 ;
  assign n10040 = n10039 ^ n9905 ;
  assign n10042 = n10041 ^ n10040 ;
  assign n10046 = n10045 ^ n10042 ;
  assign n10047 = n10046 ^ x32 ;
  assign n9904 = x95 & n2890 ;
  assign n10048 = n10047 ^ n9904 ;
  assign n9903 = x97 & n2893 ;
  assign n10049 = n10048 ^ n9903 ;
  assign n9902 = n2894 & n3501 ;
  assign n10050 = n10049 ^ n9902 ;
  assign n10052 = n10051 ^ n10050 ;
  assign n9899 = n9739 ^ n9730 ;
  assign n9900 = ~n9736 & n9899 ;
  assign n9901 = n9900 ^ n9739 ;
  assign n10053 = n10052 ^ n9901 ;
  assign n10054 = n10053 ^ x29 ;
  assign n9898 = x98 & n2593 ;
  assign n10055 = n10054 ^ n9898 ;
  assign n9897 = x100 & n2428 ;
  assign n10056 = n10055 ^ n9897 ;
  assign n9896 = n2429 & n4048 ;
  assign n10057 = n10056 ^ n9896 ;
  assign n10059 = n10058 ^ n10057 ;
  assign n9893 = n9752 ^ n9748 ;
  assign n9894 = ~n9749 & n9893 ;
  assign n9895 = n9894 ^ n9752 ;
  assign n10060 = n10059 ^ n9895 ;
  assign n10061 = n10060 ^ x26 ;
  assign n9892 = x101 & n2032 ;
  assign n10062 = n10061 ^ n9892 ;
  assign n9891 = x103 & n2028 ;
  assign n10063 = n10062 ^ n9891 ;
  assign n9890 = n2029 & ~n4624 ;
  assign n10064 = n10063 ^ n9890 ;
  assign n10066 = n10065 ^ n10064 ;
  assign n10070 = n10069 ^ n10066 ;
  assign n10071 = n10070 ^ x23 ;
  assign n9889 = x104 & n1665 ;
  assign n10072 = n10071 ^ n9889 ;
  assign n9888 = x106 & n1668 ;
  assign n10073 = n10072 ^ n9888 ;
  assign n9887 = n1669 & ~n5257 ;
  assign n10074 = n10073 ^ n9887 ;
  assign n10076 = n10075 ^ n10074 ;
  assign n10080 = n10079 ^ n10076 ;
  assign n10081 = n10080 ^ x20 ;
  assign n9886 = x107 & n1340 ;
  assign n10082 = n10081 ^ n9886 ;
  assign n9885 = x109 & n1343 ;
  assign n10083 = n10082 ^ n9885 ;
  assign n9884 = n1344 & n5912 ;
  assign n10084 = n10083 ^ n9884 ;
  assign n10086 = n10085 ^ n10084 ;
  assign n9881 = n9776 ^ n9767 ;
  assign n9882 = ~n9773 & n9881 ;
  assign n9883 = n9882 ^ n9776 ;
  assign n10087 = n10086 ^ n9883 ;
  assign n10088 = n10087 ^ x17 ;
  assign n9880 = x110 & n1060 ;
  assign n10089 = n10088 ^ n9880 ;
  assign n9879 = x112 & n1063 ;
  assign n10090 = n10089 ^ n9879 ;
  assign n9878 = n1064 & ~n6616 ;
  assign n10091 = n10090 ^ n9878 ;
  assign n10093 = n10092 ^ n10091 ;
  assign n10097 = n10096 ^ n10093 ;
  assign n10098 = n10097 ^ x14 ;
  assign n9877 = x113 & n884 ;
  assign n10099 = n10098 ^ n9877 ;
  assign n9876 = x115 & n789 ;
  assign n10100 = n10099 ^ n9876 ;
  assign n9875 = n790 & ~n7353 ;
  assign n10101 = n10100 ^ n9875 ;
  assign n10103 = n10102 ^ n10101 ;
  assign n10107 = n10106 ^ n10103 ;
  assign n10108 = n10107 ^ x11 ;
  assign n9874 = x116 & n650 ;
  assign n10109 = n10108 ^ n9874 ;
  assign n9873 = x118 & ~n578 ;
  assign n10110 = n10109 ^ n9873 ;
  assign n9872 = ~n579 & ~n8140 ;
  assign n10111 = n10110 ^ n9872 ;
  assign n10113 = n10112 ^ n10111 ;
  assign n9869 = n9800 ^ n9791 ;
  assign n9870 = ~n9797 & n9869 ;
  assign n9871 = n9870 ^ n9800 ;
  assign n10114 = n10113 ^ n9871 ;
  assign n10133 = n10132 ^ n10114 ;
  assign n9863 = x2 & x125 ;
  assign n9864 = n9863 ^ x126 ;
  assign n9865 = ~x1 & n9864 ;
  assign n9849 = x125 & ~x126 ;
  assign n9852 = ~n9542 & n9849 ;
  assign n9848 = x126 ^ x125 ;
  assign n9850 = n9849 ^ n9848 ;
  assign n9851 = ~n9541 & n9850 ;
  assign n9853 = n9852 ^ n9851 ;
  assign n9855 = x127 ^ x1 ;
  assign n9854 = x127 ^ x2 ;
  assign n9856 = n9855 ^ n9854 ;
  assign n9857 = ~n9853 & n9856 ;
  assign n9858 = n9857 ^ n9855 ;
  assign n9860 = n9858 ^ n9544 ;
  assign n9866 = n9865 ^ n9860 ;
  assign n9867 = ~x0 & n9866 ;
  assign n9868 = n9867 ^ n9858 ;
  assign n10134 = n10133 ^ n9868 ;
  assign n9845 = n9811 ^ n9801 ;
  assign n9846 = n9819 & n9845 ;
  assign n9847 = n9846 ^ n9811 ;
  assign n10135 = n10134 ^ n9847 ;
  assign n10139 = n10138 ^ n10135 ;
  assign n9842 = n9840 ^ n9823 ;
  assign n9843 = ~n9828 & n9842 ;
  assign n9844 = n9843 ^ n9840 ;
  assign n10140 = n10139 ^ n9844 ;
  assign n10440 = n10138 ^ n9844 ;
  assign n10441 = n10139 & n10440 ;
  assign n10442 = n10441 ^ n10138 ;
  assign n10430 = x121 & n391 ;
  assign n10427 = x122 & n384 ;
  assign n10425 = x120 & n456 ;
  assign n10419 = x123 & n238 ;
  assign n10418 = x125 & n234 ;
  assign n10420 = n10419 ^ n10418 ;
  assign n10421 = n10420 ^ x5 ;
  assign n10416 = n9537 ^ n9275 ;
  assign n10417 = n235 & n10416 ;
  assign n10422 = n10421 ^ n10417 ;
  assign n10415 = x124 & n231 ;
  assign n10423 = n10422 ^ n10415 ;
  assign n10424 = n10423 ^ x8 ;
  assign n10426 = n10425 ^ n10424 ;
  assign n10428 = n10427 ^ n10426 ;
  assign n10414 = n385 & ~n9261 ;
  assign n10429 = n10428 ^ n10414 ;
  assign n10431 = n10430 ^ n10429 ;
  assign n10410 = n10107 ^ n9871 ;
  assign n10411 = n10113 & n10410 ;
  assign n10412 = n10411 ^ n10107 ;
  assign n10408 = x118 & n584 ;
  assign n10401 = x115 & n795 ;
  assign n10394 = x112 & n1068 ;
  assign n10386 = n10080 ^ n9883 ;
  assign n10387 = n10086 & n10386 ;
  assign n10388 = n10387 ^ n10080 ;
  assign n10384 = x109 & n1348 ;
  assign n10377 = x106 & n1673 ;
  assign n10370 = x103 & n2025 ;
  assign n10362 = n10053 ^ n9895 ;
  assign n10363 = n10059 & n10362 ;
  assign n10364 = n10363 ^ n10053 ;
  assign n10360 = x100 & n2435 ;
  assign n10352 = n10046 ^ n9901 ;
  assign n10353 = n10052 & n10352 ;
  assign n10354 = n10353 ^ n10046 ;
  assign n10350 = x97 & n2899 ;
  assign n10343 = x94 & n3395 ;
  assign n10335 = n10029 ^ n9910 ;
  assign n10336 = n10035 & n10335 ;
  assign n10337 = n10336 ^ n10029 ;
  assign n10333 = x91 & n3940 ;
  assign n10326 = x88 & n4475 ;
  assign n10319 = x85 & n5121 ;
  assign n10311 = n10005 ^ n9925 ;
  assign n10312 = n10011 & n10311 ;
  assign n10313 = n10312 ^ n10005 ;
  assign n10309 = x82 & n5755 ;
  assign n10302 = x79 & n6449 ;
  assign n10294 = x73 & n7947 ;
  assign n10287 = x70 & n8743 ;
  assign n10278 = ~x63 & x64 ;
  assign n337 = x65 ^ x64 ;
  assign n10279 = n10278 ^ n337 ;
  assign n10280 = ~n9956 & n10279 ;
  assign n10268 = x66 & n9655 ;
  assign n10267 = x68 & n9651 ;
  assign n10269 = n10268 ^ n10267 ;
  assign n10270 = n10269 ^ x62 ;
  assign n10266 = ~n351 & n9652 ;
  assign n10271 = n10270 ^ n10266 ;
  assign n10265 = x67 & n9648 ;
  assign n10272 = n10271 ^ n10265 ;
  assign n10273 = n10272 ^ x65 ;
  assign n10281 = n10280 ^ n10273 ;
  assign n10257 = x62 & n9957 ;
  assign n10258 = n9957 ^ n9955 ;
  assign n10259 = ~n10257 & ~n10258 ;
  assign n10260 = n9966 ^ n9957 ;
  assign n10261 = n10260 ^ n10257 ;
  assign n10262 = n10261 ^ n9957 ;
  assign n10263 = n10259 & ~n10262 ;
  assign n10264 = n10263 ^ n10261 ;
  assign n10282 = n10281 ^ n10264 ;
  assign n10283 = n10282 ^ x59 ;
  assign n10256 = x69 & n8750 ;
  assign n10284 = n10283 ^ n10256 ;
  assign n10255 = x71 & n8746 ;
  assign n10285 = n10284 ^ n10255 ;
  assign n10254 = ~n495 & n8747 ;
  assign n10286 = n10285 ^ n10254 ;
  assign n10288 = n10287 ^ n10286 ;
  assign n10251 = n9986 ^ n9969 ;
  assign n10252 = ~n9975 & n10251 ;
  assign n10253 = n10252 ^ n9986 ;
  assign n10289 = n10288 ^ n10253 ;
  assign n10290 = n10289 ^ x56 ;
  assign n10250 = x72 & n7954 ;
  assign n10291 = n10290 ^ n10250 ;
  assign n10249 = x74 & n7950 ;
  assign n10292 = n10291 ^ n10249 ;
  assign n10248 = n708 & n7951 ;
  assign n10293 = n10292 ^ n10248 ;
  assign n10295 = n10294 ^ n10293 ;
  assign n10245 = n9987 ^ n9946 ;
  assign n10246 = n9951 & n10245 ;
  assign n10247 = n10246 ^ n9946 ;
  assign n10296 = n10295 ^ n10247 ;
  assign n10235 = x75 & n7183 ;
  assign n10234 = x77 & n7186 ;
  assign n10236 = n10235 ^ n10234 ;
  assign n10237 = n10236 ^ x53 ;
  assign n10233 = ~n943 & n7187 ;
  assign n10238 = n10237 ^ n10233 ;
  assign n10232 = x76 & n7191 ;
  assign n10239 = n10238 ^ n10232 ;
  assign n10240 = n10239 ^ n9988 ;
  assign n10241 = n10240 ^ n9935 ;
  assign n10242 = n10241 ^ n10239 ;
  assign n10243 = n9994 & n10242 ;
  assign n10244 = n10243 ^ n10240 ;
  assign n10297 = n10296 ^ n10244 ;
  assign n10298 = n10297 ^ x50 ;
  assign n10231 = x78 & n6687 ;
  assign n10299 = n10298 ^ n10231 ;
  assign n10230 = x80 & n6444 ;
  assign n10300 = n10299 ^ n10230 ;
  assign n10229 = n1217 & n6445 ;
  assign n10301 = n10300 ^ n10229 ;
  assign n10303 = n10302 ^ n10301 ;
  assign n10226 = n10004 ^ n9932 ;
  assign n10227 = ~n9996 & n10226 ;
  assign n10228 = n10227 ^ n10004 ;
  assign n10304 = n10303 ^ n10228 ;
  assign n10305 = n10304 ^ x47 ;
  assign n10225 = x81 & n5981 ;
  assign n10306 = n10305 ^ n10225 ;
  assign n10224 = x83 & n5748 ;
  assign n10307 = n10306 ^ n10224 ;
  assign n10223 = n1517 & n5749 ;
  assign n10308 = n10307 ^ n10223 ;
  assign n10310 = n10309 ^ n10308 ;
  assign n10314 = n10313 ^ n10310 ;
  assign n10315 = n10314 ^ x44 ;
  assign n10222 = x84 & n5113 ;
  assign n10316 = n10315 ^ n10222 ;
  assign n10221 = x86 & n5116 ;
  assign n10317 = n10316 ^ n10221 ;
  assign n10220 = n1868 & n5117 ;
  assign n10318 = n10317 ^ n10220 ;
  assign n10320 = n10319 ^ n10318 ;
  assign n10217 = n10012 ^ n9919 ;
  assign n10218 = n10018 & n10217 ;
  assign n10219 = n10218 ^ n10012 ;
  assign n10321 = n10320 ^ n10219 ;
  assign n10322 = n10321 ^ x41 ;
  assign n10216 = x87 & n4482 ;
  assign n10323 = n10322 ^ n10216 ;
  assign n10215 = x89 & n4478 ;
  assign n10324 = n10323 ^ n10215 ;
  assign n10214 = n2255 & n4479 ;
  assign n10325 = n10324 ^ n10214 ;
  assign n10327 = n10326 ^ n10325 ;
  assign n10211 = n10028 ^ n10019 ;
  assign n10212 = ~n10025 & n10211 ;
  assign n10213 = n10212 ^ n10028 ;
  assign n10328 = n10327 ^ n10213 ;
  assign n10329 = n10328 ^ x38 ;
  assign n10210 = x90 & n3932 ;
  assign n10330 = n10329 ^ n10210 ;
  assign n10209 = x92 & n3935 ;
  assign n10331 = n10330 ^ n10209 ;
  assign n10208 = n2696 & n3936 ;
  assign n10332 = n10331 ^ n10208 ;
  assign n10334 = n10333 ^ n10332 ;
  assign n10338 = n10337 ^ n10334 ;
  assign n10339 = n10338 ^ x35 ;
  assign n10207 = x93 & n3387 ;
  assign n10340 = n10339 ^ n10207 ;
  assign n10206 = x95 & n3390 ;
  assign n10341 = n10340 ^ n10206 ;
  assign n10205 = n3166 & n3391 ;
  assign n10342 = n10341 ^ n10205 ;
  assign n10344 = n10343 ^ n10342 ;
  assign n10202 = n10045 ^ n10036 ;
  assign n10203 = ~n10042 & n10202 ;
  assign n10204 = n10203 ^ n10045 ;
  assign n10345 = n10344 ^ n10204 ;
  assign n10346 = n10345 ^ x32 ;
  assign n10201 = x96 & n2890 ;
  assign n10347 = n10346 ^ n10201 ;
  assign n10200 = x98 & n2893 ;
  assign n10348 = n10347 ^ n10200 ;
  assign n10199 = n2894 & n3673 ;
  assign n10349 = n10348 ^ n10199 ;
  assign n10351 = n10350 ^ n10349 ;
  assign n10355 = n10354 ^ n10351 ;
  assign n10356 = n10355 ^ x29 ;
  assign n10198 = x99 & n2593 ;
  assign n10357 = n10356 ^ n10198 ;
  assign n10197 = x101 & n2428 ;
  assign n10358 = n10357 ^ n10197 ;
  assign n10196 = n2429 & n4223 ;
  assign n10359 = n10358 ^ n10196 ;
  assign n10361 = n10360 ^ n10359 ;
  assign n10365 = n10364 ^ n10361 ;
  assign n10366 = n10365 ^ x26 ;
  assign n10195 = x102 & n2032 ;
  assign n10367 = n10366 ^ n10195 ;
  assign n10194 = x104 & n2028 ;
  assign n10368 = n10367 ^ n10194 ;
  assign n10193 = n2029 & ~n4830 ;
  assign n10369 = n10368 ^ n10193 ;
  assign n10371 = n10370 ^ n10369 ;
  assign n10190 = n10069 ^ n10060 ;
  assign n10191 = ~n10066 & n10190 ;
  assign n10192 = n10191 ^ n10069 ;
  assign n10372 = n10371 ^ n10192 ;
  assign n10373 = n10372 ^ x23 ;
  assign n10189 = x105 & n1665 ;
  assign n10374 = n10373 ^ n10189 ;
  assign n10188 = x107 & n1668 ;
  assign n10375 = n10374 ^ n10188 ;
  assign n10187 = n1669 & ~n5459 ;
  assign n10376 = n10375 ^ n10187 ;
  assign n10378 = n10377 ^ n10376 ;
  assign n10184 = n10079 ^ n10070 ;
  assign n10185 = ~n10076 & n10184 ;
  assign n10186 = n10185 ^ n10079 ;
  assign n10379 = n10378 ^ n10186 ;
  assign n10380 = n10379 ^ x20 ;
  assign n10183 = x108 & n1340 ;
  assign n10381 = n10380 ^ n10183 ;
  assign n10182 = x110 & n1343 ;
  assign n10382 = n10381 ^ n10182 ;
  assign n10181 = n1344 & n6145 ;
  assign n10383 = n10382 ^ n10181 ;
  assign n10385 = n10384 ^ n10383 ;
  assign n10389 = n10388 ^ n10385 ;
  assign n10390 = n10389 ^ x17 ;
  assign n10180 = x111 & n1060 ;
  assign n10391 = n10390 ^ n10180 ;
  assign n10179 = x113 & n1063 ;
  assign n10392 = n10391 ^ n10179 ;
  assign n10178 = n1064 & ~n6849 ;
  assign n10393 = n10392 ^ n10178 ;
  assign n10395 = n10394 ^ n10393 ;
  assign n10175 = n10096 ^ n10087 ;
  assign n10176 = ~n10093 & n10175 ;
  assign n10177 = n10176 ^ n10096 ;
  assign n10396 = n10395 ^ n10177 ;
  assign n10397 = n10396 ^ x14 ;
  assign n10174 = x114 & n884 ;
  assign n10398 = n10397 ^ n10174 ;
  assign n10173 = x116 & n789 ;
  assign n10399 = n10398 ^ n10173 ;
  assign n10172 = n790 & ~n7604 ;
  assign n10400 = n10399 ^ n10172 ;
  assign n10402 = n10401 ^ n10400 ;
  assign n10169 = n10106 ^ n10097 ;
  assign n10170 = ~n10103 & n10169 ;
  assign n10171 = n10170 ^ n10106 ;
  assign n10403 = n10402 ^ n10171 ;
  assign n10404 = n10403 ^ x11 ;
  assign n10168 = x117 & n650 ;
  assign n10405 = n10404 ^ n10168 ;
  assign n10167 = x119 & ~n578 ;
  assign n10406 = n10405 ^ n10167 ;
  assign n10166 = ~n579 & n8405 ;
  assign n10407 = n10406 ^ n10166 ;
  assign n10409 = n10408 ^ n10407 ;
  assign n10413 = n10412 ^ n10409 ;
  assign n10432 = n10431 ^ n10413 ;
  assign n10144 = x2 & ~x127 ;
  assign n10151 = ~x126 & x127 ;
  assign n10154 = ~n9852 & n10151 ;
  assign n10146 = x127 ^ x126 ;
  assign n10152 = n10151 ^ n10146 ;
  assign n10153 = ~n9851 & n10152 ;
  assign n10155 = n10154 ^ n10153 ;
  assign n10156 = n10145 & ~n10155 ;
  assign n10157 = n10156 ^ x1 ;
  assign n10148 = ~x2 & ~n10146 ;
  assign n10149 = n10148 ^ x126 ;
  assign n10150 = n10145 & ~n10149 ;
  assign n10158 = n10157 ^ n10150 ;
  assign n10159 = ~x0 & n10158 ;
  assign n10160 = n10159 ^ n10157 ;
  assign n10161 = n10144 & ~n10160 ;
  assign n10163 = ~x1 & x126 ;
  assign n10164 = n10161 & n10163 ;
  assign n10162 = n10161 ^ n10160 ;
  assign n10165 = n10164 ^ n10162 ;
  assign n10433 = n10432 ^ n10165 ;
  assign n10141 = n10124 ^ n10114 ;
  assign n10142 = n10132 & n10141 ;
  assign n10143 = n10142 ^ n10124 ;
  assign n10434 = n10433 ^ n10143 ;
  assign n10435 = n10434 ^ n9868 ;
  assign n10436 = n10435 ^ n10434 ;
  assign n10437 = n10436 ^ n9847 ;
  assign n10438 = n10134 & n10437 ;
  assign n10439 = n10438 ^ n10435 ;
  assign n10443 = n10442 ^ n10439 ;
  assign n10719 = x125 & n231 ;
  assign n10712 = x119 & n584 ;
  assign n10709 = x120 & ~n578 ;
  assign n10707 = x118 & n650 ;
  assign n10701 = x121 & n456 ;
  assign n10700 = x123 & n384 ;
  assign n10702 = n10701 ^ n10700 ;
  assign n10703 = n10702 ^ x8 ;
  assign n10699 = n385 & ~n9804 ;
  assign n10704 = n10703 ^ n10699 ;
  assign n10698 = x122 & n391 ;
  assign n10705 = n10704 ^ n10698 ;
  assign n10706 = n10705 ^ x11 ;
  assign n10708 = n10707 ^ n10706 ;
  assign n10710 = n10709 ^ n10708 ;
  assign n10697 = ~n579 & n8904 ;
  assign n10711 = n10710 ^ n10697 ;
  assign n10713 = n10712 ^ n10711 ;
  assign n10693 = n10396 ^ n10171 ;
  assign n10694 = ~n10402 & ~n10693 ;
  assign n10695 = n10694 ^ n10396 ;
  assign n10691 = x116 & n795 ;
  assign n10683 = n10389 ^ n10177 ;
  assign n10684 = ~n10395 & ~n10683 ;
  assign n10685 = n10684 ^ n10389 ;
  assign n10681 = x113 & n1068 ;
  assign n10674 = x110 & n1348 ;
  assign n10666 = n10372 ^ n10186 ;
  assign n10667 = ~n10378 & ~n10666 ;
  assign n10668 = n10667 ^ n10372 ;
  assign n10664 = x107 & n1673 ;
  assign n10656 = n10365 ^ n10192 ;
  assign n10657 = ~n10371 & ~n10656 ;
  assign n10658 = n10657 ^ n10365 ;
  assign n10654 = x104 & n2025 ;
  assign n10647 = x101 & n2435 ;
  assign n10640 = x98 & n2899 ;
  assign n10632 = n10338 ^ n10204 ;
  assign n10633 = ~n10344 & ~n10632 ;
  assign n10634 = n10633 ^ n10338 ;
  assign n10630 = x95 & n3395 ;
  assign n10623 = x92 & n3940 ;
  assign n10615 = n10321 ^ n10213 ;
  assign n10616 = ~n10327 & ~n10615 ;
  assign n10617 = n10616 ^ n10321 ;
  assign n10613 = x89 & n4475 ;
  assign n10606 = x86 & n5121 ;
  assign n10599 = x83 & n5755 ;
  assign n10592 = x80 & n6449 ;
  assign n10582 = n10282 ^ n10253 ;
  assign n10583 = ~n10288 & ~n10582 ;
  assign n10584 = n10583 ^ n10282 ;
  assign n10580 = x71 & n8743 ;
  assign n10570 = x67 & n9655 ;
  assign n10569 = x69 & n9651 ;
  assign n10571 = n10570 ^ n10569 ;
  assign n10572 = n10571 ^ x62 ;
  assign n10568 = ~n376 & n9652 ;
  assign n10573 = n10572 ^ n10568 ;
  assign n10567 = x68 & n9648 ;
  assign n10574 = n10573 ^ n10567 ;
  assign n10563 = x63 & x65 ;
  assign n10564 = n10563 ^ x66 ;
  assign n10565 = ~n9956 & n10564 ;
  assign n10554 = n10272 ^ n10264 ;
  assign n10555 = n10281 & ~n10554 ;
  assign n10556 = n10555 ^ n10272 ;
  assign n10557 = n10556 ^ x66 ;
  assign n10566 = n10565 ^ n10557 ;
  assign n10575 = n10574 ^ n10566 ;
  assign n10576 = n10575 ^ x59 ;
  assign n10553 = x70 & n8750 ;
  assign n10577 = n10576 ^ n10553 ;
  assign n10552 = x72 & n8746 ;
  assign n10578 = n10577 ^ n10552 ;
  assign n10551 = n565 & n8747 ;
  assign n10579 = n10578 ^ n10551 ;
  assign n10581 = n10580 ^ n10579 ;
  assign n10585 = n10584 ^ n10581 ;
  assign n10541 = x73 & n7954 ;
  assign n10540 = x75 & n7950 ;
  assign n10542 = n10541 ^ n10540 ;
  assign n10543 = n10542 ^ x56 ;
  assign n10539 = ~n778 & n7951 ;
  assign n10544 = n10543 ^ n10539 ;
  assign n10538 = x74 & n7947 ;
  assign n10545 = n10544 ^ n10538 ;
  assign n10546 = n10545 ^ n10289 ;
  assign n10547 = n10546 ^ n10247 ;
  assign n10548 = n10547 ^ n10545 ;
  assign n10549 = ~n10295 & ~n10548 ;
  assign n10550 = n10549 ^ n10546 ;
  assign n10586 = n10585 ^ n10550 ;
  assign n10528 = x76 & n7183 ;
  assign n10527 = x78 & n7186 ;
  assign n10529 = n10528 ^ n10527 ;
  assign n10530 = n10529 ^ x53 ;
  assign n10526 = ~n1036 & n7187 ;
  assign n10531 = n10530 ^ n10526 ;
  assign n10525 = x77 & n7191 ;
  assign n10532 = n10531 ^ n10525 ;
  assign n10534 = n10532 ^ n10239 ;
  assign n10533 = n10532 ^ n10296 ;
  assign n10535 = n10534 ^ n10533 ;
  assign n10536 = n10244 & ~n10535 ;
  assign n10537 = n10536 ^ n10534 ;
  assign n10587 = n10586 ^ n10537 ;
  assign n10588 = n10587 ^ x50 ;
  assign n10524 = x79 & n6687 ;
  assign n10589 = n10588 ^ n10524 ;
  assign n10523 = x81 & n6444 ;
  assign n10590 = n10589 ^ n10523 ;
  assign n10522 = n1310 & n6445 ;
  assign n10591 = n10590 ^ n10522 ;
  assign n10593 = n10592 ^ n10591 ;
  assign n10519 = n10297 ^ n10228 ;
  assign n10520 = ~n10303 & ~n10519 ;
  assign n10521 = n10520 ^ n10297 ;
  assign n10594 = n10593 ^ n10521 ;
  assign n10595 = n10594 ^ x47 ;
  assign n10518 = x82 & n5981 ;
  assign n10596 = n10595 ^ n10518 ;
  assign n10517 = x84 & n5748 ;
  assign n10597 = n10596 ^ n10517 ;
  assign n10516 = n1635 & n5749 ;
  assign n10598 = n10597 ^ n10516 ;
  assign n10600 = n10599 ^ n10598 ;
  assign n10513 = n10313 ^ n10304 ;
  assign n10514 = n10310 & ~n10513 ;
  assign n10515 = n10514 ^ n10313 ;
  assign n10601 = n10600 ^ n10515 ;
  assign n10602 = n10601 ^ x44 ;
  assign n10512 = x85 & n5113 ;
  assign n10603 = n10602 ^ n10512 ;
  assign n10511 = x87 & n5116 ;
  assign n10604 = n10603 ^ n10511 ;
  assign n10510 = n1987 & n5117 ;
  assign n10605 = n10604 ^ n10510 ;
  assign n10607 = n10606 ^ n10605 ;
  assign n10507 = n10314 ^ n10219 ;
  assign n10508 = ~n10320 & ~n10507 ;
  assign n10509 = n10508 ^ n10314 ;
  assign n10608 = n10607 ^ n10509 ;
  assign n10609 = n10608 ^ x41 ;
  assign n10506 = x88 & n4482 ;
  assign n10610 = n10609 ^ n10506 ;
  assign n10505 = x90 & n4478 ;
  assign n10611 = n10610 ^ n10505 ;
  assign n10504 = n2398 & n4479 ;
  assign n10612 = n10611 ^ n10504 ;
  assign n10614 = n10613 ^ n10612 ;
  assign n10618 = n10617 ^ n10614 ;
  assign n10619 = n10618 ^ x38 ;
  assign n10503 = x91 & n3932 ;
  assign n10620 = n10619 ^ n10503 ;
  assign n10502 = x93 & n3935 ;
  assign n10621 = n10620 ^ n10502 ;
  assign n10501 = n2842 & n3936 ;
  assign n10622 = n10621 ^ n10501 ;
  assign n10624 = n10623 ^ n10622 ;
  assign n10498 = n10337 ^ n10328 ;
  assign n10499 = n10334 & ~n10498 ;
  assign n10500 = n10499 ^ n10337 ;
  assign n10625 = n10624 ^ n10500 ;
  assign n10626 = n10625 ^ x35 ;
  assign n10497 = x94 & n3387 ;
  assign n10627 = n10626 ^ n10497 ;
  assign n10496 = x96 & n3390 ;
  assign n10628 = n10627 ^ n10496 ;
  assign n10495 = n3336 & n3391 ;
  assign n10629 = n10628 ^ n10495 ;
  assign n10631 = n10630 ^ n10629 ;
  assign n10635 = n10634 ^ n10631 ;
  assign n10636 = n10635 ^ x32 ;
  assign n10494 = x97 & n2890 ;
  assign n10637 = n10636 ^ n10494 ;
  assign n10493 = x99 & n2893 ;
  assign n10638 = n10637 ^ n10493 ;
  assign n10492 = n2894 & n3851 ;
  assign n10639 = n10638 ^ n10492 ;
  assign n10641 = n10640 ^ n10639 ;
  assign n10489 = n10354 ^ n10345 ;
  assign n10490 = n10351 & ~n10489 ;
  assign n10491 = n10490 ^ n10354 ;
  assign n10642 = n10641 ^ n10491 ;
  assign n10643 = n10642 ^ x29 ;
  assign n10488 = x100 & n2593 ;
  assign n10644 = n10643 ^ n10488 ;
  assign n10487 = x102 & n2428 ;
  assign n10645 = n10644 ^ n10487 ;
  assign n10486 = n2429 & n4425 ;
  assign n10646 = n10645 ^ n10486 ;
  assign n10648 = n10647 ^ n10646 ;
  assign n10483 = n10364 ^ n10355 ;
  assign n10484 = n10361 & ~n10483 ;
  assign n10485 = n10484 ^ n10364 ;
  assign n10649 = n10648 ^ n10485 ;
  assign n10650 = n10649 ^ x26 ;
  assign n10482 = x103 & n2032 ;
  assign n10651 = n10650 ^ n10482 ;
  assign n10481 = x105 & n2028 ;
  assign n10652 = n10651 ^ n10481 ;
  assign n10480 = n2029 & ~n5034 ;
  assign n10653 = n10652 ^ n10480 ;
  assign n10655 = n10654 ^ n10653 ;
  assign n10659 = n10658 ^ n10655 ;
  assign n10660 = n10659 ^ x23 ;
  assign n10479 = x106 & n1665 ;
  assign n10661 = n10660 ^ n10479 ;
  assign n10478 = x108 & n1668 ;
  assign n10662 = n10661 ^ n10478 ;
  assign n10477 = n1669 & n5687 ;
  assign n10663 = n10662 ^ n10477 ;
  assign n10665 = n10664 ^ n10663 ;
  assign n10669 = n10668 ^ n10665 ;
  assign n10670 = n10669 ^ x20 ;
  assign n10476 = x109 & n1340 ;
  assign n10671 = n10670 ^ n10476 ;
  assign n10475 = x111 & n1343 ;
  assign n10672 = n10671 ^ n10475 ;
  assign n10474 = n1344 & ~n6370 ;
  assign n10673 = n10672 ^ n10474 ;
  assign n10675 = n10674 ^ n10673 ;
  assign n10471 = n10388 ^ n10379 ;
  assign n10472 = n10385 & ~n10471 ;
  assign n10473 = n10472 ^ n10388 ;
  assign n10676 = n10675 ^ n10473 ;
  assign n10677 = n10676 ^ x17 ;
  assign n10470 = x112 & n1060 ;
  assign n10678 = n10677 ^ n10470 ;
  assign n10469 = x114 & n1063 ;
  assign n10679 = n10678 ^ n10469 ;
  assign n10468 = n1064 & ~n7108 ;
  assign n10680 = n10679 ^ n10468 ;
  assign n10682 = n10681 ^ n10680 ;
  assign n10686 = n10685 ^ n10682 ;
  assign n10687 = n10686 ^ x14 ;
  assign n10467 = x115 & n884 ;
  assign n10688 = n10687 ^ n10467 ;
  assign n10466 = x117 & n789 ;
  assign n10689 = n10688 ^ n10466 ;
  assign n10465 = n790 & ~n7860 ;
  assign n10690 = n10689 ^ n10465 ;
  assign n10692 = n10691 ^ n10690 ;
  assign n10696 = n10695 ^ n10692 ;
  assign n10714 = n10713 ^ n10696 ;
  assign n10715 = n10714 ^ x5 ;
  assign n10464 = x124 & n238 ;
  assign n10716 = n10715 ^ n10464 ;
  assign n10463 = x126 & n234 ;
  assign n10717 = n10716 ^ n10463 ;
  assign n10461 = n9543 ^ x126 ;
  assign n10462 = n235 & n10461 ;
  assign n10718 = n10717 ^ n10462 ;
  assign n10720 = n10719 ^ n10718 ;
  assign n10458 = n10412 ^ n10403 ;
  assign n10459 = n10409 & ~n10458 ;
  assign n10460 = n10459 ^ n10412 ;
  assign n10721 = n10720 ^ n10460 ;
  assign n10447 = x127 & n10145 ;
  assign n10448 = n10154 ^ x2 ;
  assign n10449 = x0 & ~n10448 ;
  assign n10450 = n10449 ^ x2 ;
  assign n10451 = n10447 & n10450 ;
  assign n10452 = n10451 ^ x2 ;
  assign n10453 = n10452 ^ n10423 ;
  assign n10454 = n10453 ^ n10413 ;
  assign n10455 = n10454 ^ n10452 ;
  assign n10456 = n10431 & ~n10455 ;
  assign n10457 = n10456 ^ n10453 ;
  assign n10722 = n10721 ^ n10457 ;
  assign n10723 = n10722 ^ n10165 ;
  assign n10724 = n10723 ^ n10722 ;
  assign n10725 = n10724 ^ n10143 ;
  assign n10726 = ~n10433 & n10725 ;
  assign n10727 = n10726 ^ n10723 ;
  assign n10444 = n10442 ^ n10434 ;
  assign n10445 = n10439 & ~n10444 ;
  assign n10446 = n10445 ^ n10442 ;
  assign n10728 = n10727 ^ n10446 ;
  assign n11000 = n10722 ^ n10446 ;
  assign n11001 = n10727 & n11000 ;
  assign n11002 = n11001 ^ n10722 ;
  assign n10989 = x125 & n238 ;
  assign n10988 = x127 & n234 ;
  assign n10990 = n10989 ^ n10988 ;
  assign n10991 = n10990 ^ x5 ;
  assign n10986 = n9853 ^ x127 ;
  assign n10987 = n235 & n10986 ;
  assign n10992 = n10991 ^ n10987 ;
  assign n10985 = x126 & n231 ;
  assign n10993 = n10992 ^ n10985 ;
  assign n10974 = x122 & n456 ;
  assign n10973 = x124 & n384 ;
  assign n10975 = n10974 ^ n10973 ;
  assign n10976 = n10975 ^ x8 ;
  assign n10972 = n385 & n10117 ;
  assign n10977 = n10976 ^ n10972 ;
  assign n10971 = x123 & n391 ;
  assign n10978 = n10977 ^ n10971 ;
  assign n10963 = x120 & n584 ;
  assign n10956 = x117 & n795 ;
  assign n10948 = n10669 ^ n10473 ;
  assign n10949 = n10675 & n10948 ;
  assign n10950 = n10949 ^ n10669 ;
  assign n10946 = x114 & n1068 ;
  assign n10939 = x111 & n1348 ;
  assign n10932 = x108 & n1673 ;
  assign n10924 = n10642 ^ n10485 ;
  assign n10925 = n10648 & n10924 ;
  assign n10926 = n10925 ^ n10642 ;
  assign n10922 = x105 & n2025 ;
  assign n10914 = n10635 ^ n10491 ;
  assign n10915 = n10641 & n10914 ;
  assign n10916 = n10915 ^ n10635 ;
  assign n10912 = x102 & n2435 ;
  assign n10905 = x99 & n2899 ;
  assign n10897 = n10618 ^ n10500 ;
  assign n10898 = ~n10624 & ~n10897 ;
  assign n10899 = n10898 ^ n10618 ;
  assign n10895 = x96 & n3395 ;
  assign n10888 = x93 & n3940 ;
  assign n10881 = x90 & n4475 ;
  assign n10873 = n10594 ^ n10515 ;
  assign n10874 = ~n10600 & ~n10873 ;
  assign n10875 = n10874 ^ n10594 ;
  assign n10871 = x87 & n5121 ;
  assign n10863 = n10587 ^ n10521 ;
  assign n10864 = n10593 & ~n10863 ;
  assign n10865 = n10864 ^ n10587 ;
  assign n10861 = x84 & n5755 ;
  assign n10854 = x81 & n6449 ;
  assign n10847 = x78 & n7191 ;
  assign n10840 = x75 & n7947 ;
  assign n10828 = x71 & n8750 ;
  assign n10827 = x73 & n8746 ;
  assign n10829 = n10828 ^ n10827 ;
  assign n10830 = n10829 ^ x59 ;
  assign n10826 = n636 & n8747 ;
  assign n10831 = n10830 ^ n10826 ;
  assign n10825 = x72 & n8743 ;
  assign n10832 = n10831 ^ n10825 ;
  assign n10821 = ~n443 & n9652 ;
  assign n10820 = x69 & n9648 ;
  assign n10822 = n10821 ^ n10820 ;
  assign n10818 = x68 & n9655 ;
  assign n10817 = x70 & n9651 ;
  assign n10819 = n10818 ^ n10817 ;
  assign n10823 = n10822 ^ n10819 ;
  assign n10815 = x63 & x67 ;
  assign n10816 = n10815 ^ x2 ;
  assign n10824 = n10823 ^ n10816 ;
  assign n10833 = n10832 ^ n10824 ;
  assign n10812 = x63 & x66 ;
  assign n10813 = n10812 ^ x67 ;
  assign n10814 = x62 & ~n10813 ;
  assign n10834 = n10833 ^ n10814 ;
  assign n10807 = n10574 ^ n10556 ;
  assign n10808 = ~n10566 & n10807 ;
  assign n10809 = n10808 ^ n10574 ;
  assign n10835 = n10834 ^ n10809 ;
  assign n10836 = n10835 ^ x56 ;
  assign n10806 = x74 & n7954 ;
  assign n10837 = n10836 ^ n10806 ;
  assign n10805 = x76 & n7950 ;
  assign n10838 = n10837 ^ n10805 ;
  assign n10804 = ~n863 & n7951 ;
  assign n10839 = n10838 ^ n10804 ;
  assign n10841 = n10840 ^ n10839 ;
  assign n10801 = n10584 ^ n10575 ;
  assign n10802 = ~n10581 & ~n10801 ;
  assign n10803 = n10802 ^ n10584 ;
  assign n10842 = n10841 ^ n10803 ;
  assign n10843 = n10842 ^ x53 ;
  assign n10800 = x77 & n7183 ;
  assign n10844 = n10843 ^ n10800 ;
  assign n10799 = x79 & n7186 ;
  assign n10845 = n10844 ^ n10799 ;
  assign n10798 = n1123 & n7187 ;
  assign n10846 = n10845 ^ n10798 ;
  assign n10848 = n10847 ^ n10846 ;
  assign n10795 = n10585 ^ n10545 ;
  assign n10796 = ~n10550 & ~n10795 ;
  assign n10797 = n10796 ^ n10545 ;
  assign n10849 = n10848 ^ n10797 ;
  assign n10850 = n10849 ^ x50 ;
  assign n10794 = x80 & n6687 ;
  assign n10851 = n10850 ^ n10794 ;
  assign n10793 = x82 & n6444 ;
  assign n10852 = n10851 ^ n10793 ;
  assign n10792 = n1422 & n6445 ;
  assign n10853 = n10852 ^ n10792 ;
  assign n10855 = n10854 ^ n10853 ;
  assign n10789 = n10586 ^ n10532 ;
  assign n10790 = n10537 & n10789 ;
  assign n10791 = n10790 ^ n10532 ;
  assign n10856 = n10855 ^ n10791 ;
  assign n10857 = n10856 ^ x47 ;
  assign n10788 = x83 & n5981 ;
  assign n10858 = n10857 ^ n10788 ;
  assign n10787 = x85 & n5748 ;
  assign n10859 = n10858 ^ n10787 ;
  assign n10786 = n1748 & n5749 ;
  assign n10860 = n10859 ^ n10786 ;
  assign n10862 = n10861 ^ n10860 ;
  assign n10866 = n10865 ^ n10862 ;
  assign n10867 = n10866 ^ x44 ;
  assign n10785 = x86 & n5113 ;
  assign n10868 = n10867 ^ n10785 ;
  assign n10784 = x88 & n5116 ;
  assign n10869 = n10868 ^ n10784 ;
  assign n10783 = n2131 & n5117 ;
  assign n10870 = n10869 ^ n10783 ;
  assign n10872 = n10871 ^ n10870 ;
  assign n10876 = n10875 ^ n10872 ;
  assign n10877 = n10876 ^ x41 ;
  assign n10782 = x89 & n4482 ;
  assign n10878 = n10877 ^ n10782 ;
  assign n10781 = x91 & n4478 ;
  assign n10879 = n10878 ^ n10781 ;
  assign n10780 = n2548 & n4479 ;
  assign n10880 = n10879 ^ n10780 ;
  assign n10882 = n10881 ^ n10880 ;
  assign n10777 = n10601 ^ n10509 ;
  assign n10778 = ~n10607 & n10777 ;
  assign n10779 = n10778 ^ n10601 ;
  assign n10883 = n10882 ^ n10779 ;
  assign n10884 = n10883 ^ x38 ;
  assign n10776 = x92 & n3932 ;
  assign n10885 = n10884 ^ n10776 ;
  assign n10775 = x94 & n3935 ;
  assign n10886 = n10885 ^ n10775 ;
  assign n10774 = n3010 & n3936 ;
  assign n10887 = n10886 ^ n10774 ;
  assign n10889 = n10888 ^ n10887 ;
  assign n10771 = n10617 ^ n10608 ;
  assign n10772 = ~n10614 & ~n10771 ;
  assign n10773 = n10772 ^ n10617 ;
  assign n10890 = n10889 ^ n10773 ;
  assign n10891 = n10890 ^ x35 ;
  assign n10770 = x95 & n3387 ;
  assign n10892 = n10891 ^ n10770 ;
  assign n10769 = x97 & n3390 ;
  assign n10893 = n10892 ^ n10769 ;
  assign n10768 = n3391 & n3501 ;
  assign n10894 = n10893 ^ n10768 ;
  assign n10896 = n10895 ^ n10894 ;
  assign n10900 = n10899 ^ n10896 ;
  assign n10901 = n10900 ^ x32 ;
  assign n10767 = x98 & n2890 ;
  assign n10902 = n10901 ^ n10767 ;
  assign n10766 = x100 & n2893 ;
  assign n10903 = n10902 ^ n10766 ;
  assign n10765 = n2894 & n4048 ;
  assign n10904 = n10903 ^ n10765 ;
  assign n10906 = n10905 ^ n10904 ;
  assign n10762 = n10634 ^ n10625 ;
  assign n10763 = n10631 & n10762 ;
  assign n10764 = n10763 ^ n10634 ;
  assign n10907 = n10906 ^ n10764 ;
  assign n10908 = n10907 ^ x29 ;
  assign n10761 = x101 & n2593 ;
  assign n10909 = n10908 ^ n10761 ;
  assign n10760 = x103 & n2428 ;
  assign n10910 = n10909 ^ n10760 ;
  assign n10759 = n2429 & ~n4624 ;
  assign n10911 = n10910 ^ n10759 ;
  assign n10913 = n10912 ^ n10911 ;
  assign n10917 = n10916 ^ n10913 ;
  assign n10918 = n10917 ^ x26 ;
  assign n10758 = x104 & n2032 ;
  assign n10919 = n10918 ^ n10758 ;
  assign n10757 = x106 & n2028 ;
  assign n10920 = n10919 ^ n10757 ;
  assign n10756 = n2029 & ~n5257 ;
  assign n10921 = n10920 ^ n10756 ;
  assign n10923 = n10922 ^ n10921 ;
  assign n10927 = n10926 ^ n10923 ;
  assign n10928 = n10927 ^ x23 ;
  assign n10755 = x107 & n1665 ;
  assign n10929 = n10928 ^ n10755 ;
  assign n10754 = x109 & n1668 ;
  assign n10930 = n10929 ^ n10754 ;
  assign n10753 = n1669 & n5912 ;
  assign n10931 = n10930 ^ n10753 ;
  assign n10933 = n10932 ^ n10931 ;
  assign n10750 = n10658 ^ n10649 ;
  assign n10751 = ~n10655 & ~n10750 ;
  assign n10752 = n10751 ^ n10658 ;
  assign n10934 = n10933 ^ n10752 ;
  assign n10935 = n10934 ^ x20 ;
  assign n10749 = x110 & n1340 ;
  assign n10936 = n10935 ^ n10749 ;
  assign n10748 = x112 & n1343 ;
  assign n10937 = n10936 ^ n10748 ;
  assign n10747 = n1344 & ~n6616 ;
  assign n10938 = n10937 ^ n10747 ;
  assign n10940 = n10939 ^ n10938 ;
  assign n10744 = n10668 ^ n10659 ;
  assign n10745 = n10665 & n10744 ;
  assign n10746 = n10745 ^ n10668 ;
  assign n10941 = n10940 ^ n10746 ;
  assign n10942 = n10941 ^ x17 ;
  assign n10743 = x113 & n1060 ;
  assign n10943 = n10942 ^ n10743 ;
  assign n10742 = x115 & n1063 ;
  assign n10944 = n10943 ^ n10742 ;
  assign n10741 = n1064 & ~n7353 ;
  assign n10945 = n10944 ^ n10741 ;
  assign n10947 = n10946 ^ n10945 ;
  assign n10951 = n10950 ^ n10947 ;
  assign n10952 = n10951 ^ x14 ;
  assign n10740 = x116 & n884 ;
  assign n10953 = n10952 ^ n10740 ;
  assign n10739 = x118 & n789 ;
  assign n10954 = n10953 ^ n10739 ;
  assign n10738 = n790 & ~n8140 ;
  assign n10955 = n10954 ^ n10738 ;
  assign n10957 = n10956 ^ n10955 ;
  assign n10735 = n10685 ^ n10676 ;
  assign n10736 = ~n10682 & ~n10735 ;
  assign n10737 = n10736 ^ n10685 ;
  assign n10958 = n10957 ^ n10737 ;
  assign n10959 = n10958 ^ x11 ;
  assign n10734 = x119 & n650 ;
  assign n10960 = n10959 ^ n10734 ;
  assign n10733 = x121 & ~n578 ;
  assign n10961 = n10960 ^ n10733 ;
  assign n10732 = ~n579 & n8979 ;
  assign n10962 = n10961 ^ n10732 ;
  assign n10964 = n10963 ^ n10962 ;
  assign n10729 = n10695 ^ n10686 ;
  assign n10730 = n10692 & n10729 ;
  assign n10731 = n10730 ^ n10695 ;
  assign n10965 = n10964 ^ n10731 ;
  assign n10966 = n10965 ^ n10705 ;
  assign n10967 = n10966 ^ n10696 ;
  assign n10968 = n10967 ^ n10965 ;
  assign n10969 = n10713 & n10968 ;
  assign n10970 = n10969 ^ n10966 ;
  assign n10979 = n10978 ^ n10970 ;
  assign n10980 = n10979 ^ n10714 ;
  assign n10981 = n10980 ^ n10979 ;
  assign n10982 = n10981 ^ n10460 ;
  assign n10983 = n10720 & n10982 ;
  assign n10984 = n10983 ^ n10980 ;
  assign n10994 = n10993 ^ n10984 ;
  assign n10996 = n10994 ^ n10721 ;
  assign n10995 = n10994 ^ n10452 ;
  assign n10997 = n10996 ^ n10995 ;
  assign n10998 = ~n10457 & n10997 ;
  assign n10999 = n10998 ^ n10996 ;
  assign n11003 = n11002 ^ n10999 ;
  assign n11269 = n10993 ^ n10979 ;
  assign n11270 = n10984 & n11269 ;
  assign n11271 = n11270 ^ n10979 ;
  assign n11265 = n10978 ^ n10965 ;
  assign n11266 = n10970 & n11265 ;
  assign n11267 = n11266 ^ n10965 ;
  assign n11263 = x127 & n231 ;
  assign n11256 = n10958 ^ n10731 ;
  assign n11257 = ~n10964 & n11256 ;
  assign n11258 = n11257 ^ n10958 ;
  assign n11254 = x124 & n391 ;
  assign n11246 = n10951 ^ n10737 ;
  assign n11247 = n10957 & ~n11246 ;
  assign n11248 = n11247 ^ n10951 ;
  assign n11244 = x121 & n584 ;
  assign n11237 = x118 & n795 ;
  assign n11229 = n10934 ^ n10746 ;
  assign n11230 = ~n10940 & n11229 ;
  assign n11231 = n11230 ^ n10934 ;
  assign n11227 = x115 & n1068 ;
  assign n11219 = n10927 ^ n10752 ;
  assign n11220 = n10933 & ~n11219 ;
  assign n11221 = n11220 ^ n10927 ;
  assign n11217 = x112 & n1348 ;
  assign n11210 = x109 & n1673 ;
  assign n11203 = x106 & n2025 ;
  assign n11195 = n10900 ^ n10764 ;
  assign n11196 = ~n10906 & n11195 ;
  assign n11197 = n11196 ^ n10900 ;
  assign n11193 = x103 & n2435 ;
  assign n11186 = x100 & n2899 ;
  assign n11178 = n10883 ^ n10773 ;
  assign n11179 = ~n10889 & n11178 ;
  assign n11180 = n11179 ^ n10883 ;
  assign n11176 = x97 & n3395 ;
  assign n11169 = x94 & n3940 ;
  assign n11162 = x91 & n4475 ;
  assign n11155 = x88 & n5121 ;
  assign n11148 = x85 & n5755 ;
  assign n11139 = n10835 ^ n10803 ;
  assign n11140 = n10841 & ~n11139 ;
  assign n11141 = n11140 ^ n10835 ;
  assign n11133 = x78 & n7183 ;
  assign n11132 = x80 & n7186 ;
  assign n11134 = n11133 ^ n11132 ;
  assign n11135 = n11134 ^ x53 ;
  assign n11131 = n1217 & n7187 ;
  assign n11136 = n11135 ^ n11131 ;
  assign n11130 = x79 & n7191 ;
  assign n11137 = n11136 ^ n11130 ;
  assign n11123 = x75 & n7954 ;
  assign n11122 = x77 & n7950 ;
  assign n11124 = n11123 ^ n11122 ;
  assign n11125 = n11124 ^ x56 ;
  assign n11121 = ~n943 & n7951 ;
  assign n11126 = n11125 ^ n11121 ;
  assign n11120 = x76 & n7947 ;
  assign n11127 = n11126 ^ n11120 ;
  assign n11114 = x63 & x68 ;
  assign n11115 = n11114 ^ x2 ;
  assign n11111 = ~n495 & n9652 ;
  assign n11110 = x70 & n9648 ;
  assign n11112 = n11111 ^ n11110 ;
  assign n11108 = x69 & n9655 ;
  assign n11107 = x71 & n9651 ;
  assign n11109 = n11108 ^ n11107 ;
  assign n11113 = n11112 ^ n11109 ;
  assign n11116 = n11115 ^ n11113 ;
  assign n11101 = x62 ^ x2 ;
  assign n11102 = n11101 ^ n10823 ;
  assign n11103 = n10823 ^ n10815 ;
  assign n11104 = n11103 ^ n10814 ;
  assign n11105 = n11102 & ~n11104 ;
  assign n11106 = n11105 ^ x2 ;
  assign n11117 = n11116 ^ n11106 ;
  assign n11099 = n10815 ^ x68 ;
  assign n11100 = x62 & ~n11099 ;
  assign n11118 = n11117 ^ n11100 ;
  assign n11094 = x72 & n8750 ;
  assign n11093 = x74 & n8746 ;
  assign n11095 = n11094 ^ n11093 ;
  assign n11096 = n11095 ^ x59 ;
  assign n11092 = n708 & n8747 ;
  assign n11097 = n11096 ^ n11092 ;
  assign n11091 = x73 & n8743 ;
  assign n11098 = n11097 ^ n11091 ;
  assign n11119 = n11118 ^ n11098 ;
  assign n11128 = n11127 ^ n11119 ;
  assign n11088 = n10832 ^ n10809 ;
  assign n11089 = n10834 & n11088 ;
  assign n11090 = n11089 ^ n10832 ;
  assign n11129 = n11128 ^ n11090 ;
  assign n11138 = n11137 ^ n11129 ;
  assign n11142 = n11141 ^ n11138 ;
  assign n11078 = x81 & n6687 ;
  assign n11077 = x83 & n6444 ;
  assign n11079 = n11078 ^ n11077 ;
  assign n11080 = n11079 ^ x50 ;
  assign n11076 = n1517 & n6445 ;
  assign n11081 = n11080 ^ n11076 ;
  assign n11075 = x82 & n6449 ;
  assign n11082 = n11081 ^ n11075 ;
  assign n11083 = n11082 ^ n10842 ;
  assign n11084 = n11083 ^ n10797 ;
  assign n11085 = n11084 ^ n11082 ;
  assign n11086 = ~n10848 & ~n11085 ;
  assign n11087 = n11086 ^ n11083 ;
  assign n11143 = n11142 ^ n11087 ;
  assign n11144 = n11143 ^ x47 ;
  assign n11074 = x84 & n5981 ;
  assign n11145 = n11144 ^ n11074 ;
  assign n11073 = x86 & n5748 ;
  assign n11146 = n11145 ^ n11073 ;
  assign n11072 = n1868 & n5749 ;
  assign n11147 = n11146 ^ n11072 ;
  assign n11149 = n11148 ^ n11147 ;
  assign n11069 = n10849 ^ n10791 ;
  assign n11070 = ~n10855 & ~n11069 ;
  assign n11071 = n11070 ^ n10849 ;
  assign n11150 = n11149 ^ n11071 ;
  assign n11151 = n11150 ^ x44 ;
  assign n11068 = x87 & n5113 ;
  assign n11152 = n11151 ^ n11068 ;
  assign n11067 = x89 & n5116 ;
  assign n11153 = n11152 ^ n11067 ;
  assign n11066 = n2255 & n5117 ;
  assign n11154 = n11153 ^ n11066 ;
  assign n11156 = n11155 ^ n11154 ;
  assign n11063 = n10865 ^ n10856 ;
  assign n11064 = n10862 & ~n11063 ;
  assign n11065 = n11064 ^ n10865 ;
  assign n11157 = n11156 ^ n11065 ;
  assign n11158 = n11157 ^ x41 ;
  assign n11062 = x90 & n4482 ;
  assign n11159 = n11158 ^ n11062 ;
  assign n11061 = x92 & n4478 ;
  assign n11160 = n11159 ^ n11061 ;
  assign n11060 = n2696 & n4479 ;
  assign n11161 = n11160 ^ n11060 ;
  assign n11163 = n11162 ^ n11161 ;
  assign n11057 = n10875 ^ n10866 ;
  assign n11058 = n10872 & n11057 ;
  assign n11059 = n11058 ^ n10875 ;
  assign n11164 = n11163 ^ n11059 ;
  assign n11165 = n11164 ^ x38 ;
  assign n11056 = x93 & n3932 ;
  assign n11166 = n11165 ^ n11056 ;
  assign n11055 = x95 & n3935 ;
  assign n11167 = n11166 ^ n11055 ;
  assign n11054 = n3166 & n3936 ;
  assign n11168 = n11167 ^ n11054 ;
  assign n11170 = n11169 ^ n11168 ;
  assign n11051 = n10876 ^ n10779 ;
  assign n11052 = n10882 & ~n11051 ;
  assign n11053 = n11052 ^ n10876 ;
  assign n11171 = n11170 ^ n11053 ;
  assign n11172 = n11171 ^ x35 ;
  assign n11050 = x96 & n3387 ;
  assign n11173 = n11172 ^ n11050 ;
  assign n11049 = x98 & n3390 ;
  assign n11174 = n11173 ^ n11049 ;
  assign n11048 = n3391 & n3673 ;
  assign n11175 = n11174 ^ n11048 ;
  assign n11177 = n11176 ^ n11175 ;
  assign n11181 = n11180 ^ n11177 ;
  assign n11182 = n11181 ^ x32 ;
  assign n11047 = x99 & n2890 ;
  assign n11183 = n11182 ^ n11047 ;
  assign n11046 = x101 & n2893 ;
  assign n11184 = n11183 ^ n11046 ;
  assign n11045 = n2894 & n4223 ;
  assign n11185 = n11184 ^ n11045 ;
  assign n11187 = n11186 ^ n11185 ;
  assign n11042 = n10899 ^ n10890 ;
  assign n11043 = ~n10896 & ~n11042 ;
  assign n11044 = n11043 ^ n10899 ;
  assign n11188 = n11187 ^ n11044 ;
  assign n11189 = n11188 ^ x29 ;
  assign n11041 = x102 & n2593 ;
  assign n11190 = n11189 ^ n11041 ;
  assign n11040 = x104 & n2428 ;
  assign n11191 = n11190 ^ n11040 ;
  assign n11039 = n2429 & ~n4830 ;
  assign n11192 = n11191 ^ n11039 ;
  assign n11194 = n11193 ^ n11192 ;
  assign n11198 = n11197 ^ n11194 ;
  assign n11199 = n11198 ^ x26 ;
  assign n11038 = x105 & n2032 ;
  assign n11200 = n11199 ^ n11038 ;
  assign n11037 = x107 & n2028 ;
  assign n11201 = n11200 ^ n11037 ;
  assign n11036 = n2029 & ~n5459 ;
  assign n11202 = n11201 ^ n11036 ;
  assign n11204 = n11203 ^ n11202 ;
  assign n11033 = n10916 ^ n10907 ;
  assign n11034 = ~n10913 & n11033 ;
  assign n11035 = n11034 ^ n10916 ;
  assign n11205 = n11204 ^ n11035 ;
  assign n11206 = n11205 ^ x23 ;
  assign n11032 = x108 & n1665 ;
  assign n11207 = n11206 ^ n11032 ;
  assign n11031 = x110 & n1668 ;
  assign n11208 = n11207 ^ n11031 ;
  assign n11030 = n1669 & n6145 ;
  assign n11209 = n11208 ^ n11030 ;
  assign n11211 = n11210 ^ n11209 ;
  assign n11027 = n10926 ^ n10917 ;
  assign n11028 = ~n10923 & n11027 ;
  assign n11029 = n11028 ^ n10926 ;
  assign n11212 = n11211 ^ n11029 ;
  assign n11213 = n11212 ^ x20 ;
  assign n11026 = x111 & n1340 ;
  assign n11214 = n11213 ^ n11026 ;
  assign n11025 = x113 & n1343 ;
  assign n11215 = n11214 ^ n11025 ;
  assign n11024 = n1344 & ~n6849 ;
  assign n11216 = n11215 ^ n11024 ;
  assign n11218 = n11217 ^ n11216 ;
  assign n11222 = n11221 ^ n11218 ;
  assign n11223 = n11222 ^ x17 ;
  assign n11023 = x114 & n1060 ;
  assign n11224 = n11223 ^ n11023 ;
  assign n11022 = x116 & n1063 ;
  assign n11225 = n11224 ^ n11022 ;
  assign n11021 = n1064 & ~n7604 ;
  assign n11226 = n11225 ^ n11021 ;
  assign n11228 = n11227 ^ n11226 ;
  assign n11232 = n11231 ^ n11228 ;
  assign n11233 = n11232 ^ x14 ;
  assign n11020 = x117 & n884 ;
  assign n11234 = n11233 ^ n11020 ;
  assign n11019 = x119 & n789 ;
  assign n11235 = n11234 ^ n11019 ;
  assign n11018 = n790 & n8405 ;
  assign n11236 = n11235 ^ n11018 ;
  assign n11238 = n11237 ^ n11236 ;
  assign n11015 = n10950 ^ n10941 ;
  assign n11016 = ~n10947 & n11015 ;
  assign n11017 = n11016 ^ n10950 ;
  assign n11239 = n11238 ^ n11017 ;
  assign n11240 = n11239 ^ x11 ;
  assign n11014 = x120 & n650 ;
  assign n11241 = n11240 ^ n11014 ;
  assign n11013 = x122 & ~n578 ;
  assign n11242 = n11241 ^ n11013 ;
  assign n11012 = ~n579 & ~n9261 ;
  assign n11243 = n11242 ^ n11012 ;
  assign n11245 = n11244 ^ n11243 ;
  assign n11249 = n11248 ^ n11245 ;
  assign n11250 = n11249 ^ x8 ;
  assign n11011 = x123 & n456 ;
  assign n11251 = n11250 ^ n11011 ;
  assign n11010 = x125 & n384 ;
  assign n11252 = n11251 ^ n11010 ;
  assign n11009 = n385 & n10416 ;
  assign n11253 = n11252 ^ n11009 ;
  assign n11255 = n11254 ^ n11253 ;
  assign n11259 = n11258 ^ n11255 ;
  assign n11260 = n11259 ^ x5 ;
  assign n11008 = x126 & n238 ;
  assign n11261 = n11260 ^ n11008 ;
  assign n11007 = n235 & n10155 ;
  assign n11262 = n11261 ^ n11007 ;
  assign n11264 = n11263 ^ n11262 ;
  assign n11268 = n11267 ^ n11264 ;
  assign n11272 = n11271 ^ n11268 ;
  assign n11004 = n11002 ^ n10994 ;
  assign n11005 = ~n10999 & n11004 ;
  assign n11006 = n11005 ^ n11002 ;
  assign n11273 = n11272 ^ n11006 ;
  assign n11541 = x125 & n391 ;
  assign n11533 = n11232 ^ n11017 ;
  assign n11534 = ~n11238 & ~n11533 ;
  assign n11535 = n11534 ^ n11232 ;
  assign n11531 = x122 & n584 ;
  assign n11524 = x119 & n795 ;
  assign n11517 = x116 & n1068 ;
  assign n11509 = n11205 ^ n11029 ;
  assign n11510 = n11211 & n11509 ;
  assign n11511 = n11510 ^ n11205 ;
  assign n11507 = x113 & n1348 ;
  assign n11499 = n11198 ^ n11035 ;
  assign n11500 = n11204 & n11499 ;
  assign n11501 = n11500 ^ n11198 ;
  assign n11497 = x110 & n1673 ;
  assign n11490 = x107 & n2025 ;
  assign n11482 = n11181 ^ n11044 ;
  assign n11483 = n11187 & ~n11482 ;
  assign n11484 = n11483 ^ n11181 ;
  assign n11480 = x104 & n2435 ;
  assign n11473 = x101 & n2899 ;
  assign n11466 = x98 & n3395 ;
  assign n11458 = n11157 ^ n11059 ;
  assign n11459 = n11163 & ~n11458 ;
  assign n11460 = n11459 ^ n11157 ;
  assign n11456 = x95 & n3940 ;
  assign n11448 = n11150 ^ n11065 ;
  assign n11449 = n11156 & n11448 ;
  assign n11450 = n11449 ^ n11150 ;
  assign n11446 = x92 & n4475 ;
  assign n11438 = n11143 ^ n11071 ;
  assign n11439 = ~n11149 & n11438 ;
  assign n11440 = n11439 ^ n11143 ;
  assign n11436 = x89 & n5121 ;
  assign n11426 = x85 & n5981 ;
  assign n11425 = x87 & n5748 ;
  assign n11427 = n11426 ^ n11425 ;
  assign n11428 = n11427 ^ x47 ;
  assign n11424 = n1987 & n5749 ;
  assign n11429 = n11428 ^ n11424 ;
  assign n11423 = x86 & n5755 ;
  assign n11430 = n11429 ^ n11423 ;
  assign n11411 = x82 & n6687 ;
  assign n11410 = x84 & n6444 ;
  assign n11412 = n11411 ^ n11410 ;
  assign n11413 = n11412 ^ x50 ;
  assign n11409 = n1635 & n6445 ;
  assign n11414 = n11413 ^ n11409 ;
  assign n11408 = x83 & n6449 ;
  assign n11415 = n11414 ^ n11408 ;
  assign n11405 = x80 & n7191 ;
  assign n11403 = n1310 & n7187 ;
  assign n11399 = x79 & n7183 ;
  assign n11398 = x81 & n7186 ;
  assign n11400 = n11399 ^ n11398 ;
  assign n11401 = n11400 ^ x53 ;
  assign n11393 = n11114 ^ x69 ;
  assign n11394 = x62 & ~n11393 ;
  assign n11391 = x63 & x69 ;
  assign n11387 = n565 & n9652 ;
  assign n11386 = x71 & n9648 ;
  assign n11388 = n11387 ^ n11386 ;
  assign n11384 = x70 & n9655 ;
  assign n11383 = x72 & n9651 ;
  assign n11385 = n11384 ^ n11383 ;
  assign n11389 = n11388 ^ n11385 ;
  assign n11390 = n11389 ^ x2 ;
  assign n11392 = n11391 ^ n11390 ;
  assign n11395 = n11394 ^ n11392 ;
  assign n11378 = n11113 ^ n11101 ;
  assign n11379 = n11114 ^ n11113 ;
  assign n11380 = n11379 ^ n11100 ;
  assign n11381 = n11378 & ~n11380 ;
  assign n11372 = x73 & n8750 ;
  assign n11371 = x75 & n8746 ;
  assign n11373 = n11372 ^ n11371 ;
  assign n11374 = n11373 ^ x59 ;
  assign n11370 = ~n778 & n8747 ;
  assign n11375 = n11374 ^ n11370 ;
  assign n11369 = x74 & n8743 ;
  assign n11376 = n11375 ^ n11369 ;
  assign n11377 = n11376 ^ x2 ;
  assign n11382 = n11381 ^ n11377 ;
  assign n11396 = n11395 ^ n11382 ;
  assign n11366 = ~n1036 & n7951 ;
  assign n11364 = x76 & n7954 ;
  assign n11360 = n11106 ^ n11098 ;
  assign n11361 = ~n11118 & n11360 ;
  assign n11362 = n11361 ^ n11098 ;
  assign n11358 = x78 & n7950 ;
  assign n11359 = n11358 ^ x56 ;
  assign n11363 = n11362 ^ n11359 ;
  assign n11365 = n11364 ^ n11363 ;
  assign n11367 = n11366 ^ n11365 ;
  assign n11357 = x77 & n7947 ;
  assign n11368 = n11367 ^ n11357 ;
  assign n11397 = n11396 ^ n11368 ;
  assign n11402 = n11401 ^ n11397 ;
  assign n11404 = n11403 ^ n11402 ;
  assign n11406 = n11405 ^ n11404 ;
  assign n11354 = n11127 ^ n11090 ;
  assign n11355 = n11128 & n11354 ;
  assign n11356 = n11355 ^ n11127 ;
  assign n11407 = n11406 ^ n11356 ;
  assign n11416 = n11415 ^ n11407 ;
  assign n11351 = n11141 ^ n11137 ;
  assign n11352 = ~n11138 & n11351 ;
  assign n11353 = n11352 ^ n11141 ;
  assign n11417 = n11416 ^ n11353 ;
  assign n11419 = n11417 ^ n11082 ;
  assign n11418 = n11417 ^ n11142 ;
  assign n11420 = n11419 ^ n11418 ;
  assign n11421 = ~n11087 & n11420 ;
  assign n11422 = n11421 ^ n11419 ;
  assign n11431 = n11430 ^ n11422 ;
  assign n11432 = n11431 ^ x44 ;
  assign n11350 = x88 & n5113 ;
  assign n11433 = n11432 ^ n11350 ;
  assign n11349 = x90 & n5116 ;
  assign n11434 = n11433 ^ n11349 ;
  assign n11348 = n2398 & n5117 ;
  assign n11435 = n11434 ^ n11348 ;
  assign n11437 = n11436 ^ n11435 ;
  assign n11441 = n11440 ^ n11437 ;
  assign n11442 = n11441 ^ x41 ;
  assign n11347 = x91 & n4482 ;
  assign n11443 = n11442 ^ n11347 ;
  assign n11346 = x93 & n4478 ;
  assign n11444 = n11443 ^ n11346 ;
  assign n11345 = n2842 & n4479 ;
  assign n11445 = n11444 ^ n11345 ;
  assign n11447 = n11446 ^ n11445 ;
  assign n11451 = n11450 ^ n11447 ;
  assign n11452 = n11451 ^ x38 ;
  assign n11344 = x94 & n3932 ;
  assign n11453 = n11452 ^ n11344 ;
  assign n11343 = x96 & n3935 ;
  assign n11454 = n11453 ^ n11343 ;
  assign n11342 = n3336 & n3936 ;
  assign n11455 = n11454 ^ n11342 ;
  assign n11457 = n11456 ^ n11455 ;
  assign n11461 = n11460 ^ n11457 ;
  assign n11462 = n11461 ^ x35 ;
  assign n11341 = x97 & n3387 ;
  assign n11463 = n11462 ^ n11341 ;
  assign n11340 = x99 & n3390 ;
  assign n11464 = n11463 ^ n11340 ;
  assign n11339 = n3391 & n3851 ;
  assign n11465 = n11464 ^ n11339 ;
  assign n11467 = n11466 ^ n11465 ;
  assign n11336 = n11164 ^ n11053 ;
  assign n11337 = ~n11170 & ~n11336 ;
  assign n11338 = n11337 ^ n11164 ;
  assign n11468 = n11467 ^ n11338 ;
  assign n11469 = n11468 ^ x32 ;
  assign n11335 = x100 & n2890 ;
  assign n11470 = n11469 ^ n11335 ;
  assign n11334 = x102 & n2893 ;
  assign n11471 = n11470 ^ n11334 ;
  assign n11333 = n2894 & n4425 ;
  assign n11472 = n11471 ^ n11333 ;
  assign n11474 = n11473 ^ n11472 ;
  assign n11330 = n11180 ^ n11171 ;
  assign n11331 = n11177 & n11330 ;
  assign n11332 = n11331 ^ n11180 ;
  assign n11475 = n11474 ^ n11332 ;
  assign n11476 = n11475 ^ x29 ;
  assign n11329 = x103 & n2593 ;
  assign n11477 = n11476 ^ n11329 ;
  assign n11328 = x105 & n2428 ;
  assign n11478 = n11477 ^ n11328 ;
  assign n11327 = n2429 & ~n5034 ;
  assign n11479 = n11478 ^ n11327 ;
  assign n11481 = n11480 ^ n11479 ;
  assign n11485 = n11484 ^ n11481 ;
  assign n11486 = n11485 ^ x26 ;
  assign n11326 = x106 & n2032 ;
  assign n11487 = n11486 ^ n11326 ;
  assign n11325 = x108 & n2028 ;
  assign n11488 = n11487 ^ n11325 ;
  assign n11324 = n2029 & n5687 ;
  assign n11489 = n11488 ^ n11324 ;
  assign n11491 = n11490 ^ n11489 ;
  assign n11321 = n11197 ^ n11188 ;
  assign n11322 = n11194 & n11321 ;
  assign n11323 = n11322 ^ n11197 ;
  assign n11492 = n11491 ^ n11323 ;
  assign n11493 = n11492 ^ x23 ;
  assign n11320 = x109 & n1665 ;
  assign n11494 = n11493 ^ n11320 ;
  assign n11319 = x111 & n1668 ;
  assign n11495 = n11494 ^ n11319 ;
  assign n11318 = n1669 & ~n6370 ;
  assign n11496 = n11495 ^ n11318 ;
  assign n11498 = n11497 ^ n11496 ;
  assign n11502 = n11501 ^ n11498 ;
  assign n11503 = n11502 ^ x20 ;
  assign n11317 = x112 & n1340 ;
  assign n11504 = n11503 ^ n11317 ;
  assign n11316 = x114 & n1343 ;
  assign n11505 = n11504 ^ n11316 ;
  assign n11315 = n1344 & ~n7108 ;
  assign n11506 = n11505 ^ n11315 ;
  assign n11508 = n11507 ^ n11506 ;
  assign n11512 = n11511 ^ n11508 ;
  assign n11513 = n11512 ^ x17 ;
  assign n11314 = x115 & n1060 ;
  assign n11514 = n11513 ^ n11314 ;
  assign n11313 = x117 & n1063 ;
  assign n11515 = n11514 ^ n11313 ;
  assign n11312 = n1064 & ~n7860 ;
  assign n11516 = n11515 ^ n11312 ;
  assign n11518 = n11517 ^ n11516 ;
  assign n11309 = n11221 ^ n11212 ;
  assign n11310 = ~n11218 & n11309 ;
  assign n11311 = n11310 ^ n11221 ;
  assign n11519 = n11518 ^ n11311 ;
  assign n11520 = n11519 ^ x14 ;
  assign n11308 = x118 & n884 ;
  assign n11521 = n11520 ^ n11308 ;
  assign n11307 = x120 & n789 ;
  assign n11522 = n11521 ^ n11307 ;
  assign n11306 = n790 & n8904 ;
  assign n11523 = n11522 ^ n11306 ;
  assign n11525 = n11524 ^ n11523 ;
  assign n11303 = n11231 ^ n11222 ;
  assign n11304 = ~n11228 & ~n11303 ;
  assign n11305 = n11304 ^ n11231 ;
  assign n11526 = n11525 ^ n11305 ;
  assign n11527 = n11526 ^ x11 ;
  assign n11302 = x121 & n650 ;
  assign n11528 = n11527 ^ n11302 ;
  assign n11301 = x123 & ~n578 ;
  assign n11529 = n11528 ^ n11301 ;
  assign n11300 = ~n579 & ~n9804 ;
  assign n11530 = n11529 ^ n11300 ;
  assign n11532 = n11531 ^ n11530 ;
  assign n11536 = n11535 ^ n11532 ;
  assign n11537 = n11536 ^ x8 ;
  assign n11299 = x124 & n456 ;
  assign n11538 = n11537 ^ n11299 ;
  assign n11298 = x126 & n384 ;
  assign n11539 = n11538 ^ n11298 ;
  assign n11297 = n385 & n10461 ;
  assign n11540 = n11539 ^ n11297 ;
  assign n11542 = n11541 ^ n11540 ;
  assign n11294 = n11248 ^ n11239 ;
  assign n11295 = n11245 & ~n11294 ;
  assign n11296 = n11295 ^ n11248 ;
  assign n11543 = n11542 ^ n11296 ;
  assign n11283 = x127 & n237 ;
  assign n11284 = n11283 ^ n233 ;
  assign n11285 = n10154 ^ x127 ;
  assign n11290 = n202 & n11285 ;
  assign n11291 = n11290 ^ n11283 ;
  assign n11292 = n11284 & ~n11291 ;
  assign n11293 = n11292 ^ x4 ;
  assign n11544 = n11543 ^ n11293 ;
  assign n11280 = n11258 ^ n11249 ;
  assign n11281 = n11255 & n11280 ;
  assign n11282 = n11281 ^ n11258 ;
  assign n11545 = n11544 ^ n11282 ;
  assign n11277 = n11267 ^ n11259 ;
  assign n11278 = ~n11264 & n11277 ;
  assign n11279 = n11278 ^ n11267 ;
  assign n11546 = n11545 ^ n11279 ;
  assign n11274 = n11271 ^ n11006 ;
  assign n11275 = n11272 & n11274 ;
  assign n11276 = n11275 ^ n11271 ;
  assign n11547 = n11546 ^ n11276 ;
  assign n11551 = n11293 ^ n11282 ;
  assign n11809 = n11536 ^ n11296 ;
  assign n11810 = n11542 & n11809 ;
  assign n11811 = n11810 ^ n11536 ;
  assign n11807 = x126 & n391 ;
  assign n11800 = x123 & n584 ;
  assign n11792 = n11519 ^ n11305 ;
  assign n11793 = n11525 & ~n11792 ;
  assign n11794 = n11793 ^ n11519 ;
  assign n11790 = x120 & n795 ;
  assign n11782 = n11512 ^ n11311 ;
  assign n11783 = n11518 & n11782 ;
  assign n11784 = n11783 ^ n11512 ;
  assign n11780 = x117 & n1068 ;
  assign n11773 = x114 & n1348 ;
  assign n11766 = x111 & n1673 ;
  assign n11758 = n11485 ^ n11323 ;
  assign n11759 = ~n11491 & n11758 ;
  assign n11760 = n11759 ^ n11485 ;
  assign n11756 = x108 & n2025 ;
  assign n11749 = x105 & n2435 ;
  assign n11741 = n11468 ^ n11332 ;
  assign n11742 = n11474 & ~n11741 ;
  assign n11743 = n11742 ^ n11468 ;
  assign n11739 = x102 & n2899 ;
  assign n11732 = x99 & n3395 ;
  assign n11725 = x96 & n3940 ;
  assign n11718 = x93 & n4475 ;
  assign n11711 = x90 & n5121 ;
  assign n11701 = x86 & n5981 ;
  assign n11700 = x88 & n5748 ;
  assign n11702 = n11701 ^ n11700 ;
  assign n11703 = n11702 ^ x47 ;
  assign n11699 = n2131 & n5749 ;
  assign n11704 = n11703 ^ n11699 ;
  assign n11698 = x87 & n5755 ;
  assign n11705 = n11704 ^ n11698 ;
  assign n11689 = n11415 ^ n11353 ;
  assign n11690 = n11416 & n11689 ;
  assign n11691 = n11690 ^ n11415 ;
  assign n11687 = x84 & n6449 ;
  assign n11679 = n11397 ^ n11356 ;
  assign n11680 = n11406 & n11679 ;
  assign n11681 = n11680 ^ n11397 ;
  assign n11673 = x80 & n7183 ;
  assign n11672 = x82 & n7186 ;
  assign n11674 = n11673 ^ n11672 ;
  assign n11675 = n11674 ^ x53 ;
  assign n11671 = n1422 & n7187 ;
  assign n11676 = n11675 ^ n11671 ;
  assign n11670 = x81 & n7191 ;
  assign n11677 = n11676 ^ n11670 ;
  assign n11666 = x75 & n8743 ;
  assign n11656 = x71 & n9655 ;
  assign n11655 = x73 & n9651 ;
  assign n11657 = n11656 ^ n11655 ;
  assign n11658 = n11657 ^ x62 ;
  assign n11654 = n636 & n9652 ;
  assign n11659 = n11658 ^ n11654 ;
  assign n11653 = x72 & n9648 ;
  assign n11660 = n11659 ^ n11653 ;
  assign n11647 = n11389 ^ n11101 ;
  assign n11648 = n11394 ^ n11391 ;
  assign n11649 = n11648 ^ n11389 ;
  assign n11650 = n11647 & ~n11649 ;
  assign n11651 = n11650 ^ x2 ;
  assign n11643 = n11391 ^ x70 ;
  assign n11644 = ~n9956 & n11643 ;
  assign n11645 = n11644 ^ x70 ;
  assign n11642 = x5 ^ x2 ;
  assign n11646 = n11645 ^ n11642 ;
  assign n11652 = n11651 ^ n11646 ;
  assign n11661 = n11660 ^ n11652 ;
  assign n11662 = n11661 ^ x59 ;
  assign n11641 = x74 & n8750 ;
  assign n11663 = n11662 ^ n11641 ;
  assign n11640 = x76 & n8746 ;
  assign n11664 = n11663 ^ n11640 ;
  assign n11639 = ~n863 & n8747 ;
  assign n11665 = n11664 ^ n11639 ;
  assign n11667 = n11666 ^ n11665 ;
  assign n11636 = n11395 ^ n11376 ;
  assign n11637 = n11382 & n11636 ;
  assign n11638 = n11637 ^ n11376 ;
  assign n11668 = n11667 ^ n11638 ;
  assign n11626 = x77 & n7954 ;
  assign n11625 = x79 & n7950 ;
  assign n11627 = n11626 ^ n11625 ;
  assign n11628 = n11627 ^ x56 ;
  assign n11624 = n1123 & n7951 ;
  assign n11629 = n11628 ^ n11624 ;
  assign n11623 = x78 & n7947 ;
  assign n11630 = n11629 ^ n11623 ;
  assign n11631 = n11630 ^ n11396 ;
  assign n11632 = n11631 ^ n11362 ;
  assign n11633 = n11632 ^ n11630 ;
  assign n11634 = ~n11368 & n11633 ;
  assign n11635 = n11634 ^ n11631 ;
  assign n11669 = n11668 ^ n11635 ;
  assign n11678 = n11677 ^ n11669 ;
  assign n11682 = n11681 ^ n11678 ;
  assign n11683 = n11682 ^ x50 ;
  assign n11622 = x83 & n6687 ;
  assign n11684 = n11683 ^ n11622 ;
  assign n11621 = x85 & n6444 ;
  assign n11685 = n11684 ^ n11621 ;
  assign n11620 = n1748 & n6445 ;
  assign n11686 = n11685 ^ n11620 ;
  assign n11688 = n11687 ^ n11686 ;
  assign n11692 = n11691 ^ n11688 ;
  assign n11694 = n11692 ^ n11417 ;
  assign n11693 = n11692 ^ n11430 ;
  assign n11695 = n11694 ^ n11693 ;
  assign n11696 = n11422 & n11695 ;
  assign n11697 = n11696 ^ n11694 ;
  assign n11706 = n11705 ^ n11697 ;
  assign n11707 = n11706 ^ x44 ;
  assign n11619 = x89 & n5113 ;
  assign n11708 = n11707 ^ n11619 ;
  assign n11618 = x91 & n5116 ;
  assign n11709 = n11708 ^ n11618 ;
  assign n11617 = n2548 & n5117 ;
  assign n11710 = n11709 ^ n11617 ;
  assign n11712 = n11711 ^ n11710 ;
  assign n11614 = n11440 ^ n11431 ;
  assign n11615 = ~n11437 & ~n11614 ;
  assign n11616 = n11615 ^ n11440 ;
  assign n11713 = n11712 ^ n11616 ;
  assign n11714 = n11713 ^ x41 ;
  assign n11613 = x92 & n4482 ;
  assign n11715 = n11714 ^ n11613 ;
  assign n11612 = x94 & n4478 ;
  assign n11716 = n11715 ^ n11612 ;
  assign n11611 = n3010 & n4479 ;
  assign n11717 = n11716 ^ n11611 ;
  assign n11719 = n11718 ^ n11717 ;
  assign n11608 = n11450 ^ n11441 ;
  assign n11609 = n11447 & ~n11608 ;
  assign n11610 = n11609 ^ n11450 ;
  assign n11720 = n11719 ^ n11610 ;
  assign n11721 = n11720 ^ x38 ;
  assign n11607 = x95 & n3932 ;
  assign n11722 = n11721 ^ n11607 ;
  assign n11606 = x97 & n3935 ;
  assign n11723 = n11722 ^ n11606 ;
  assign n11605 = n3501 & n3936 ;
  assign n11724 = n11723 ^ n11605 ;
  assign n11726 = n11725 ^ n11724 ;
  assign n11602 = n11460 ^ n11451 ;
  assign n11603 = n11457 & ~n11602 ;
  assign n11604 = n11603 ^ n11460 ;
  assign n11727 = n11726 ^ n11604 ;
  assign n11728 = n11727 ^ x35 ;
  assign n11601 = x98 & n3387 ;
  assign n11729 = n11728 ^ n11601 ;
  assign n11600 = x100 & n3390 ;
  assign n11730 = n11729 ^ n11600 ;
  assign n11599 = n3391 & n4048 ;
  assign n11731 = n11730 ^ n11599 ;
  assign n11733 = n11732 ^ n11731 ;
  assign n11596 = n11461 ^ n11338 ;
  assign n11597 = ~n11467 & n11596 ;
  assign n11598 = n11597 ^ n11461 ;
  assign n11734 = n11733 ^ n11598 ;
  assign n11735 = n11734 ^ x32 ;
  assign n11595 = x101 & n2890 ;
  assign n11736 = n11735 ^ n11595 ;
  assign n11594 = x103 & n2893 ;
  assign n11737 = n11736 ^ n11594 ;
  assign n11593 = n2894 & ~n4624 ;
  assign n11738 = n11737 ^ n11593 ;
  assign n11740 = n11739 ^ n11738 ;
  assign n11744 = n11743 ^ n11740 ;
  assign n11745 = n11744 ^ x29 ;
  assign n11592 = x104 & n2593 ;
  assign n11746 = n11745 ^ n11592 ;
  assign n11591 = x106 & n2428 ;
  assign n11747 = n11746 ^ n11591 ;
  assign n11590 = n2429 & ~n5257 ;
  assign n11748 = n11747 ^ n11590 ;
  assign n11750 = n11749 ^ n11748 ;
  assign n11587 = n11484 ^ n11475 ;
  assign n11588 = n11481 & ~n11587 ;
  assign n11589 = n11588 ^ n11484 ;
  assign n11751 = n11750 ^ n11589 ;
  assign n11752 = n11751 ^ x26 ;
  assign n11586 = x107 & n2032 ;
  assign n11753 = n11752 ^ n11586 ;
  assign n11585 = x109 & n2028 ;
  assign n11754 = n11753 ^ n11585 ;
  assign n11584 = n2029 & n5912 ;
  assign n11755 = n11754 ^ n11584 ;
  assign n11757 = n11756 ^ n11755 ;
  assign n11761 = n11760 ^ n11757 ;
  assign n11762 = n11761 ^ x23 ;
  assign n11583 = x110 & n1665 ;
  assign n11763 = n11762 ^ n11583 ;
  assign n11582 = x112 & n1668 ;
  assign n11764 = n11763 ^ n11582 ;
  assign n11581 = n1669 & ~n6616 ;
  assign n11765 = n11764 ^ n11581 ;
  assign n11767 = n11766 ^ n11765 ;
  assign n11578 = n11501 ^ n11492 ;
  assign n11579 = ~n11498 & n11578 ;
  assign n11580 = n11579 ^ n11501 ;
  assign n11768 = n11767 ^ n11580 ;
  assign n11769 = n11768 ^ x20 ;
  assign n11577 = x113 & n1340 ;
  assign n11770 = n11769 ^ n11577 ;
  assign n11576 = x115 & n1343 ;
  assign n11771 = n11770 ^ n11576 ;
  assign n11575 = n1344 & ~n7353 ;
  assign n11772 = n11771 ^ n11575 ;
  assign n11774 = n11773 ^ n11772 ;
  assign n11572 = n11511 ^ n11502 ;
  assign n11573 = ~n11508 & n11572 ;
  assign n11574 = n11573 ^ n11511 ;
  assign n11775 = n11774 ^ n11574 ;
  assign n11776 = n11775 ^ x17 ;
  assign n11571 = x116 & n1060 ;
  assign n11777 = n11776 ^ n11571 ;
  assign n11570 = x118 & n1063 ;
  assign n11778 = n11777 ^ n11570 ;
  assign n11569 = n1064 & ~n8140 ;
  assign n11779 = n11778 ^ n11569 ;
  assign n11781 = n11780 ^ n11779 ;
  assign n11785 = n11784 ^ n11781 ;
  assign n11786 = n11785 ^ x14 ;
  assign n11568 = x119 & n884 ;
  assign n11787 = n11786 ^ n11568 ;
  assign n11567 = x121 & n789 ;
  assign n11788 = n11787 ^ n11567 ;
  assign n11566 = n790 & n8979 ;
  assign n11789 = n11788 ^ n11566 ;
  assign n11791 = n11790 ^ n11789 ;
  assign n11795 = n11794 ^ n11791 ;
  assign n11796 = n11795 ^ x11 ;
  assign n11565 = x122 & n650 ;
  assign n11797 = n11796 ^ n11565 ;
  assign n11564 = x124 & ~n578 ;
  assign n11798 = n11797 ^ n11564 ;
  assign n11563 = ~n579 & n10117 ;
  assign n11799 = n11798 ^ n11563 ;
  assign n11801 = n11800 ^ n11799 ;
  assign n11560 = n11535 ^ n11526 ;
  assign n11561 = n11532 & n11560 ;
  assign n11562 = n11561 ^ n11535 ;
  assign n11802 = n11801 ^ n11562 ;
  assign n11803 = n11802 ^ x8 ;
  assign n11559 = x125 & n456 ;
  assign n11804 = n11803 ^ n11559 ;
  assign n11558 = x127 & n384 ;
  assign n11805 = n11804 ^ n11558 ;
  assign n11557 = n385 & n10986 ;
  assign n11806 = n11805 ^ n11557 ;
  assign n11808 = n11807 ^ n11806 ;
  assign n11812 = n11811 ^ n11808 ;
  assign n11553 = n11543 ^ n11282 ;
  assign n11813 = n11812 ^ n11553 ;
  assign n11552 = n11279 ^ n11276 ;
  assign n11554 = n11553 ^ n11293 ;
  assign n11555 = n11554 ^ n11279 ;
  assign n11556 = ~n11552 & ~n11555 ;
  assign n11814 = n11813 ^ n11556 ;
  assign n11815 = n11814 ^ n11812 ;
  assign n11816 = n11815 ^ n11556 ;
  assign n11817 = n11816 ^ n11815 ;
  assign n11818 = n11815 ^ n11276 ;
  assign n11819 = n11818 ^ n11815 ;
  assign n11820 = n11817 & n11819 ;
  assign n11821 = n11820 ^ n11815 ;
  assign n11822 = ~n11551 & n11821 ;
  assign n11823 = n11822 ^ n11814 ;
  assign n11548 = ~n11279 & ~n11543 ;
  assign n11549 = ~n11545 & n11548 ;
  assign n11550 = ~n11276 & n11549 ;
  assign n11824 = n11823 ^ n11550 ;
  assign n12079 = n11548 ^ n11276 ;
  assign n12081 = n12079 ^ n11276 ;
  assign n12082 = n12081 ^ n12079 ;
  assign n12083 = n11543 ^ n11279 ;
  assign n12084 = n12083 ^ n12079 ;
  assign n12085 = n12082 & n12084 ;
  assign n12086 = n12085 ^ n12079 ;
  assign n12087 = ~n11812 & ~n12086 ;
  assign n12080 = n12079 ^ n11282 ;
  assign n12088 = n12087 ^ n12080 ;
  assign n12089 = ~n11552 & n12083 ;
  assign n12090 = n12089 ^ n11543 ;
  assign n12092 = n12090 ^ n11293 ;
  assign n12091 = n12090 ^ n11282 ;
  assign n12093 = n12092 ^ n12091 ;
  assign n12094 = ~n12088 & ~n12093 ;
  assign n12095 = n12094 ^ n12092 ;
  assign n12096 = n12090 ^ n11812 ;
  assign n12097 = ~n12095 & n12096 ;
  assign n12098 = n12097 ^ n11812 ;
  assign n12074 = n11795 ^ n11562 ;
  assign n12075 = ~n11801 & n12074 ;
  assign n12076 = n12075 ^ n11795 ;
  assign n12072 = x127 & n391 ;
  assign n12066 = x124 & n584 ;
  assign n12055 = x120 & n884 ;
  assign n12054 = x122 & n789 ;
  assign n12056 = n12055 ^ n12054 ;
  assign n12057 = n12056 ^ x14 ;
  assign n12053 = n790 & ~n9261 ;
  assign n12058 = n12057 ^ n12053 ;
  assign n12052 = x121 & n795 ;
  assign n12059 = n12058 ^ n12052 ;
  assign n12048 = n11768 ^ n11574 ;
  assign n12049 = ~n11774 & ~n12048 ;
  assign n12050 = n12049 ^ n11768 ;
  assign n12046 = x118 & n1068 ;
  assign n12038 = n11761 ^ n11580 ;
  assign n12039 = ~n11767 & ~n12038 ;
  assign n12040 = n12039 ^ n11761 ;
  assign n12036 = x115 & n1348 ;
  assign n12029 = x112 & n1673 ;
  assign n12021 = n11744 ^ n11589 ;
  assign n12022 = n11750 & n12021 ;
  assign n12023 = n12022 ^ n11744 ;
  assign n12019 = x109 & n2025 ;
  assign n12012 = x106 & n2435 ;
  assign n12005 = x103 & n2899 ;
  assign n11997 = n11720 ^ n11604 ;
  assign n11998 = ~n11726 & ~n11997 ;
  assign n11999 = n11998 ^ n11720 ;
  assign n11995 = x100 & n3395 ;
  assign n11987 = n11713 ^ n11610 ;
  assign n11988 = ~n11719 & ~n11987 ;
  assign n11989 = n11988 ^ n11713 ;
  assign n11985 = x97 & n3940 ;
  assign n11977 = n11706 ^ n11616 ;
  assign n11978 = n11712 & ~n11977 ;
  assign n11979 = n11978 ^ n11706 ;
  assign n11975 = x94 & n4475 ;
  assign n11967 = n11705 ^ n11692 ;
  assign n11968 = n11697 & n11967 ;
  assign n11969 = n11968 ^ n11692 ;
  assign n11961 = x90 & n5113 ;
  assign n11960 = x92 & n5116 ;
  assign n11962 = n11961 ^ n11960 ;
  assign n11963 = n11962 ^ x44 ;
  assign n11959 = n2696 & n5117 ;
  assign n11964 = n11963 ^ n11959 ;
  assign n11958 = x91 & n5121 ;
  assign n11965 = n11964 ^ n11958 ;
  assign n11951 = x87 & n5981 ;
  assign n11950 = x89 & n5748 ;
  assign n11952 = n11951 ^ n11950 ;
  assign n11953 = n11952 ^ x47 ;
  assign n11949 = n2255 & n5749 ;
  assign n11954 = n11953 ^ n11949 ;
  assign n11948 = x88 & n5755 ;
  assign n11955 = n11954 ^ n11948 ;
  assign n11941 = x84 & n6687 ;
  assign n11940 = x86 & n6444 ;
  assign n11942 = n11941 ^ n11940 ;
  assign n11943 = n11942 ^ x50 ;
  assign n11939 = n1868 & n6445 ;
  assign n11944 = n11943 ^ n11939 ;
  assign n11938 = x85 & n6449 ;
  assign n11945 = n11944 ^ n11938 ;
  assign n11931 = x81 & n7183 ;
  assign n11930 = x83 & n7186 ;
  assign n11932 = n11931 ^ n11930 ;
  assign n11933 = n11932 ^ x53 ;
  assign n11929 = n1517 & n7187 ;
  assign n11934 = n11933 ^ n11929 ;
  assign n11928 = x82 & n7191 ;
  assign n11935 = n11934 ^ n11928 ;
  assign n11925 = x79 & n7947 ;
  assign n11914 = x75 & n8750 ;
  assign n11913 = x77 & n8746 ;
  assign n11915 = n11914 ^ n11913 ;
  assign n11916 = n11915 ^ x59 ;
  assign n11912 = ~n943 & n8747 ;
  assign n11917 = n11916 ^ n11912 ;
  assign n11911 = x76 & n8743 ;
  assign n11918 = n11917 ^ n11911 ;
  assign n11905 = x72 & n9655 ;
  assign n11904 = x74 & n9651 ;
  assign n11906 = n11905 ^ n11904 ;
  assign n11907 = n11906 ^ x62 ;
  assign n11903 = n708 & n9652 ;
  assign n11908 = n11907 ^ n11903 ;
  assign n11902 = x73 & n9648 ;
  assign n11909 = n11908 ^ n11902 ;
  assign n11897 = n11645 ^ x5 ;
  assign n11898 = n11642 & n11897 ;
  assign n11899 = n11898 ^ x2 ;
  assign n11894 = x62 & ~x63 ;
  assign n11895 = n11894 ^ x62 ;
  assign n11896 = x70 & n11895 ;
  assign n11900 = n11899 ^ n11896 ;
  assign n11893 = x71 & n9956 ;
  assign n11901 = n11900 ^ n11893 ;
  assign n11910 = n11909 ^ n11901 ;
  assign n11919 = n11918 ^ n11910 ;
  assign n11890 = n11660 ^ n11651 ;
  assign n11891 = ~n11652 & n11890 ;
  assign n11892 = n11891 ^ n11660 ;
  assign n11920 = n11919 ^ n11892 ;
  assign n11921 = n11920 ^ x56 ;
  assign n11889 = x78 & n7954 ;
  assign n11922 = n11921 ^ n11889 ;
  assign n11888 = x80 & n7950 ;
  assign n11923 = n11922 ^ n11888 ;
  assign n11887 = n1217 & n7951 ;
  assign n11924 = n11923 ^ n11887 ;
  assign n11926 = n11925 ^ n11924 ;
  assign n11884 = n11661 ^ n11638 ;
  assign n11885 = n11667 & n11884 ;
  assign n11886 = n11885 ^ n11661 ;
  assign n11927 = n11926 ^ n11886 ;
  assign n11936 = n11935 ^ n11927 ;
  assign n11881 = n11668 ^ n11630 ;
  assign n11882 = n11635 & n11881 ;
  assign n11883 = n11882 ^ n11630 ;
  assign n11937 = n11936 ^ n11883 ;
  assign n11946 = n11945 ^ n11937 ;
  assign n11878 = n11681 ^ n11677 ;
  assign n11879 = ~n11678 & n11878 ;
  assign n11880 = n11879 ^ n11681 ;
  assign n11947 = n11946 ^ n11880 ;
  assign n11956 = n11955 ^ n11947 ;
  assign n11875 = n11691 ^ n11682 ;
  assign n11876 = ~n11688 & n11875 ;
  assign n11877 = n11876 ^ n11691 ;
  assign n11957 = n11956 ^ n11877 ;
  assign n11966 = n11965 ^ n11957 ;
  assign n11970 = n11969 ^ n11966 ;
  assign n11971 = n11970 ^ x41 ;
  assign n11874 = x93 & n4482 ;
  assign n11972 = n11971 ^ n11874 ;
  assign n11873 = x95 & n4478 ;
  assign n11973 = n11972 ^ n11873 ;
  assign n11872 = n3166 & n4479 ;
  assign n11974 = n11973 ^ n11872 ;
  assign n11976 = n11975 ^ n11974 ;
  assign n11980 = n11979 ^ n11976 ;
  assign n11981 = n11980 ^ x38 ;
  assign n11871 = x96 & n3932 ;
  assign n11982 = n11981 ^ n11871 ;
  assign n11870 = x98 & n3935 ;
  assign n11983 = n11982 ^ n11870 ;
  assign n11869 = n3673 & n3936 ;
  assign n11984 = n11983 ^ n11869 ;
  assign n11986 = n11985 ^ n11984 ;
  assign n11990 = n11989 ^ n11986 ;
  assign n11991 = n11990 ^ x35 ;
  assign n11868 = x99 & n3387 ;
  assign n11992 = n11991 ^ n11868 ;
  assign n11867 = x101 & n3390 ;
  assign n11993 = n11992 ^ n11867 ;
  assign n11866 = n3391 & n4223 ;
  assign n11994 = n11993 ^ n11866 ;
  assign n11996 = n11995 ^ n11994 ;
  assign n12000 = n11999 ^ n11996 ;
  assign n12001 = n12000 ^ x32 ;
  assign n11865 = x102 & n2890 ;
  assign n12002 = n12001 ^ n11865 ;
  assign n11864 = x104 & n2893 ;
  assign n12003 = n12002 ^ n11864 ;
  assign n11863 = n2894 & ~n4830 ;
  assign n12004 = n12003 ^ n11863 ;
  assign n12006 = n12005 ^ n12004 ;
  assign n11860 = n11727 ^ n11598 ;
  assign n11861 = ~n11733 & n11860 ;
  assign n11862 = n11861 ^ n11727 ;
  assign n12007 = n12006 ^ n11862 ;
  assign n12008 = n12007 ^ x29 ;
  assign n11859 = x105 & n2593 ;
  assign n12009 = n12008 ^ n11859 ;
  assign n11858 = x107 & n2428 ;
  assign n12010 = n12009 ^ n11858 ;
  assign n11857 = n2429 & ~n5459 ;
  assign n12011 = n12010 ^ n11857 ;
  assign n12013 = n12012 ^ n12011 ;
  assign n11854 = n11743 ^ n11734 ;
  assign n11855 = ~n11740 & n11854 ;
  assign n11856 = n11855 ^ n11743 ;
  assign n12014 = n12013 ^ n11856 ;
  assign n12015 = n12014 ^ x26 ;
  assign n11853 = x108 & n2032 ;
  assign n12016 = n12015 ^ n11853 ;
  assign n11852 = x110 & n2028 ;
  assign n12017 = n12016 ^ n11852 ;
  assign n11851 = n2029 & n6145 ;
  assign n12018 = n12017 ^ n11851 ;
  assign n12020 = n12019 ^ n12018 ;
  assign n12024 = n12023 ^ n12020 ;
  assign n12025 = n12024 ^ x23 ;
  assign n11850 = x111 & n1665 ;
  assign n12026 = n12025 ^ n11850 ;
  assign n11849 = x113 & n1668 ;
  assign n12027 = n12026 ^ n11849 ;
  assign n11848 = n1669 & ~n6849 ;
  assign n12028 = n12027 ^ n11848 ;
  assign n12030 = n12029 ^ n12028 ;
  assign n11845 = n11760 ^ n11751 ;
  assign n11846 = ~n11757 & ~n11845 ;
  assign n11847 = n11846 ^ n11760 ;
  assign n12031 = n12030 ^ n11847 ;
  assign n12032 = n12031 ^ x20 ;
  assign n11844 = x114 & n1340 ;
  assign n12033 = n12032 ^ n11844 ;
  assign n11843 = x116 & n1343 ;
  assign n12034 = n12033 ^ n11843 ;
  assign n11842 = n1344 & ~n7604 ;
  assign n12035 = n12034 ^ n11842 ;
  assign n12037 = n12036 ^ n12035 ;
  assign n12041 = n12040 ^ n12037 ;
  assign n12042 = n12041 ^ x17 ;
  assign n11841 = x117 & n1060 ;
  assign n12043 = n12042 ^ n11841 ;
  assign n11840 = x119 & n1063 ;
  assign n12044 = n12043 ^ n11840 ;
  assign n11839 = n1064 & n8405 ;
  assign n12045 = n12044 ^ n11839 ;
  assign n12047 = n12046 ^ n12045 ;
  assign n12051 = n12050 ^ n12047 ;
  assign n12060 = n12059 ^ n12051 ;
  assign n11836 = n11784 ^ n11775 ;
  assign n11837 = n11781 & ~n11836 ;
  assign n11838 = n11837 ^ n11784 ;
  assign n12061 = n12060 ^ n11838 ;
  assign n12062 = n12061 ^ x11 ;
  assign n11835 = x123 & n650 ;
  assign n12063 = n12062 ^ n11835 ;
  assign n11834 = x125 & ~n578 ;
  assign n12064 = n12063 ^ n11834 ;
  assign n11833 = ~n579 & n10416 ;
  assign n12065 = n12064 ^ n11833 ;
  assign n12067 = n12066 ^ n12065 ;
  assign n11830 = n11794 ^ n11785 ;
  assign n11831 = n11791 & ~n11830 ;
  assign n11832 = n11831 ^ n11794 ;
  assign n12068 = n12067 ^ n11832 ;
  assign n12069 = n12068 ^ x8 ;
  assign n11829 = x126 & n456 ;
  assign n12070 = n12069 ^ n11829 ;
  assign n11828 = n385 & n10155 ;
  assign n12071 = n12070 ^ n11828 ;
  assign n12073 = n12072 ^ n12071 ;
  assign n12077 = n12076 ^ n12073 ;
  assign n11825 = n11811 ^ n11802 ;
  assign n11826 = ~n11808 & n11825 ;
  assign n11827 = n11826 ^ n11811 ;
  assign n12078 = n12077 ^ n11827 ;
  assign n12099 = n12098 ^ n12078 ;
  assign n12363 = n12061 ^ n11832 ;
  assign n12364 = n12067 & n12363 ;
  assign n12365 = n12364 ^ n12061 ;
  assign n12347 = n335 ^ x7 ;
  assign n12348 = x127 & n383 ;
  assign n12349 = n12347 & n12348 ;
  assign n12350 = n12349 ^ x8 ;
  assign n12343 = n12059 ^ n11838 ;
  assign n12344 = n12060 & n12343 ;
  assign n12345 = n12344 ^ n12059 ;
  assign n12341 = x125 & n584 ;
  assign n12334 = x122 & n795 ;
  assign n12327 = x119 & n1068 ;
  assign n12319 = n12024 ^ n11847 ;
  assign n12320 = ~n12030 & n12319 ;
  assign n12321 = n12320 ^ n12024 ;
  assign n12317 = x116 & n1348 ;
  assign n12310 = x113 & n1673 ;
  assign n12302 = n12007 ^ n11856 ;
  assign n12303 = ~n12013 & ~n12302 ;
  assign n12304 = n12303 ^ n12007 ;
  assign n12300 = x110 & n2025 ;
  assign n12293 = x107 & n2435 ;
  assign n12286 = x104 & n2899 ;
  assign n12279 = x101 & n3395 ;
  assign n12272 = x98 & n3940 ;
  assign n12261 = x94 & n4482 ;
  assign n12260 = x96 & n4478 ;
  assign n12262 = n12261 ^ n12260 ;
  assign n12263 = n12262 ^ x41 ;
  assign n12259 = n3336 & n4479 ;
  assign n12264 = n12263 ^ n12259 ;
  assign n12258 = x95 & n4475 ;
  assign n12265 = n12264 ^ n12258 ;
  assign n12251 = x91 & n5113 ;
  assign n12250 = x93 & n5116 ;
  assign n12252 = n12251 ^ n12250 ;
  assign n12253 = n12252 ^ x44 ;
  assign n12249 = n2842 & n5117 ;
  assign n12254 = n12253 ^ n12249 ;
  assign n12248 = x92 & n5121 ;
  assign n12255 = n12254 ^ n12248 ;
  assign n12240 = x85 & n6687 ;
  assign n12239 = x87 & n6444 ;
  assign n12241 = n12240 ^ n12239 ;
  assign n12242 = n12241 ^ x50 ;
  assign n12238 = n1987 & n6445 ;
  assign n12243 = n12242 ^ n12238 ;
  assign n12237 = x86 & n6449 ;
  assign n12244 = n12243 ^ n12237 ;
  assign n12230 = x82 & n7183 ;
  assign n12229 = x84 & n7186 ;
  assign n12231 = n12230 ^ n12229 ;
  assign n12232 = n12231 ^ x53 ;
  assign n12228 = n1635 & n7187 ;
  assign n12233 = n12232 ^ n12228 ;
  assign n12227 = x83 & n7191 ;
  assign n12234 = n12233 ^ n12227 ;
  assign n12223 = n11918 ^ n11892 ;
  assign n12224 = n11919 & n12223 ;
  assign n12225 = n12224 ^ n11918 ;
  assign n12217 = x79 & n7954 ;
  assign n12216 = x81 & n7950 ;
  assign n12218 = n12217 ^ n12216 ;
  assign n12219 = n12218 ^ x56 ;
  assign n12215 = n1310 & n7951 ;
  assign n12220 = n12219 ^ n12215 ;
  assign n12214 = x80 & n7947 ;
  assign n12221 = n12220 ^ n12214 ;
  assign n12205 = n9956 ^ x71 ;
  assign n12206 = n11894 ^ x63 ;
  assign n12201 = ~x72 & n9956 ;
  assign n12202 = n12201 ^ n11896 ;
  assign n12207 = n12206 ^ n12202 ;
  assign n12208 = n12205 & n12207 ;
  assign n12209 = n12208 ^ n420 ;
  assign n12203 = x71 & n12202 ;
  assign n12204 = n12203 ^ n11896 ;
  assign n12210 = n12209 ^ n12204 ;
  assign n12211 = n12210 ^ n420 ;
  assign n12198 = n11909 ^ n11899 ;
  assign n12199 = ~n11901 & ~n12198 ;
  assign n12200 = n12199 ^ n11909 ;
  assign n12212 = n12211 ^ n12200 ;
  assign n12195 = ~n1036 & n8747 ;
  assign n12193 = x76 & n8750 ;
  assign n12187 = x73 & n9655 ;
  assign n12186 = x75 & n9651 ;
  assign n12188 = n12187 ^ n12186 ;
  assign n12189 = n12188 ^ x62 ;
  assign n12185 = ~n778 & n9652 ;
  assign n12190 = n12189 ^ n12185 ;
  assign n12184 = x74 & n9648 ;
  assign n12191 = n12190 ^ n12184 ;
  assign n12182 = x78 & n8746 ;
  assign n12183 = n12182 ^ x59 ;
  assign n12192 = n12191 ^ n12183 ;
  assign n12194 = n12193 ^ n12192 ;
  assign n12196 = n12195 ^ n12194 ;
  assign n12181 = x77 & n8743 ;
  assign n12197 = n12196 ^ n12181 ;
  assign n12213 = n12212 ^ n12197 ;
  assign n12222 = n12221 ^ n12213 ;
  assign n12226 = n12225 ^ n12222 ;
  assign n12235 = n12234 ^ n12226 ;
  assign n12178 = n11920 ^ n11886 ;
  assign n12179 = n11926 & n12178 ;
  assign n12180 = n12179 ^ n11920 ;
  assign n12236 = n12235 ^ n12180 ;
  assign n12245 = n12244 ^ n12236 ;
  assign n12175 = n11935 ^ n11883 ;
  assign n12176 = n11936 & n12175 ;
  assign n12177 = n12176 ^ n11935 ;
  assign n12246 = n12245 ^ n12177 ;
  assign n12172 = n2398 & n5749 ;
  assign n12170 = x88 & n5981 ;
  assign n12166 = n11945 ^ n11880 ;
  assign n12167 = n11946 & n12166 ;
  assign n12168 = n12167 ^ n11945 ;
  assign n12164 = x90 & n5748 ;
  assign n12165 = n12164 ^ x47 ;
  assign n12169 = n12168 ^ n12165 ;
  assign n12171 = n12170 ^ n12169 ;
  assign n12173 = n12172 ^ n12171 ;
  assign n12163 = x89 & n5755 ;
  assign n12174 = n12173 ^ n12163 ;
  assign n12247 = n12246 ^ n12174 ;
  assign n12256 = n12255 ^ n12247 ;
  assign n12160 = n11947 ^ n11877 ;
  assign n12161 = n11956 & ~n12160 ;
  assign n12162 = n12161 ^ n11955 ;
  assign n12257 = n12256 ^ n12162 ;
  assign n12266 = n12265 ^ n12257 ;
  assign n12157 = n11969 ^ n11965 ;
  assign n12158 = ~n11966 & n12157 ;
  assign n12159 = n12158 ^ n11969 ;
  assign n12267 = n12266 ^ n12159 ;
  assign n12268 = n12267 ^ x38 ;
  assign n12156 = x97 & n3932 ;
  assign n12269 = n12268 ^ n12156 ;
  assign n12155 = x99 & n3935 ;
  assign n12270 = n12269 ^ n12155 ;
  assign n12154 = n3851 & n3936 ;
  assign n12271 = n12270 ^ n12154 ;
  assign n12273 = n12272 ^ n12271 ;
  assign n12151 = n11979 ^ n11970 ;
  assign n12152 = ~n11976 & n12151 ;
  assign n12153 = n12152 ^ n11979 ;
  assign n12274 = n12273 ^ n12153 ;
  assign n12275 = n12274 ^ x35 ;
  assign n12150 = x100 & n3387 ;
  assign n12276 = n12275 ^ n12150 ;
  assign n12149 = x102 & n3390 ;
  assign n12277 = n12276 ^ n12149 ;
  assign n12148 = n3391 & n4425 ;
  assign n12278 = n12277 ^ n12148 ;
  assign n12280 = n12279 ^ n12278 ;
  assign n12145 = n11989 ^ n11980 ;
  assign n12146 = ~n11986 & ~n12145 ;
  assign n12147 = n12146 ^ n11989 ;
  assign n12281 = n12280 ^ n12147 ;
  assign n12282 = n12281 ^ x32 ;
  assign n12144 = x103 & n2890 ;
  assign n12283 = n12282 ^ n12144 ;
  assign n12143 = x105 & n2893 ;
  assign n12284 = n12283 ^ n12143 ;
  assign n12142 = n2894 & ~n5034 ;
  assign n12285 = n12284 ^ n12142 ;
  assign n12287 = n12286 ^ n12285 ;
  assign n12139 = n11999 ^ n11990 ;
  assign n12140 = n11996 & n12139 ;
  assign n12141 = n12140 ^ n11999 ;
  assign n12288 = n12287 ^ n12141 ;
  assign n12289 = n12288 ^ x29 ;
  assign n12138 = x106 & n2593 ;
  assign n12290 = n12289 ^ n12138 ;
  assign n12137 = x108 & n2428 ;
  assign n12291 = n12290 ^ n12137 ;
  assign n12136 = n2429 & n5687 ;
  assign n12292 = n12291 ^ n12136 ;
  assign n12294 = n12293 ^ n12292 ;
  assign n12133 = n12000 ^ n11862 ;
  assign n12134 = n12006 & ~n12133 ;
  assign n12135 = n12134 ^ n12000 ;
  assign n12295 = n12294 ^ n12135 ;
  assign n12296 = n12295 ^ x26 ;
  assign n12132 = x109 & n2032 ;
  assign n12297 = n12296 ^ n12132 ;
  assign n12131 = x111 & n2028 ;
  assign n12298 = n12297 ^ n12131 ;
  assign n12130 = n2029 & ~n6370 ;
  assign n12299 = n12298 ^ n12130 ;
  assign n12301 = n12300 ^ n12299 ;
  assign n12305 = n12304 ^ n12301 ;
  assign n12306 = n12305 ^ x23 ;
  assign n12129 = x112 & n1665 ;
  assign n12307 = n12306 ^ n12129 ;
  assign n12128 = x114 & n1668 ;
  assign n12308 = n12307 ^ n12128 ;
  assign n12127 = n1669 & ~n7108 ;
  assign n12309 = n12308 ^ n12127 ;
  assign n12311 = n12310 ^ n12309 ;
  assign n12124 = n12023 ^ n12014 ;
  assign n12125 = n12020 & ~n12124 ;
  assign n12126 = n12125 ^ n12023 ;
  assign n12312 = n12311 ^ n12126 ;
  assign n12313 = n12312 ^ x20 ;
  assign n12123 = x115 & n1340 ;
  assign n12314 = n12313 ^ n12123 ;
  assign n12122 = x117 & n1343 ;
  assign n12315 = n12314 ^ n12122 ;
  assign n12121 = n1344 & ~n7860 ;
  assign n12316 = n12315 ^ n12121 ;
  assign n12318 = n12317 ^ n12316 ;
  assign n12322 = n12321 ^ n12318 ;
  assign n12323 = n12322 ^ x17 ;
  assign n12120 = x118 & n1060 ;
  assign n12324 = n12323 ^ n12120 ;
  assign n12119 = x120 & n1063 ;
  assign n12325 = n12324 ^ n12119 ;
  assign n12118 = n1064 & n8904 ;
  assign n12326 = n12325 ^ n12118 ;
  assign n12328 = n12327 ^ n12326 ;
  assign n12115 = n12040 ^ n12031 ;
  assign n12116 = ~n12037 & ~n12115 ;
  assign n12117 = n12116 ^ n12040 ;
  assign n12329 = n12328 ^ n12117 ;
  assign n12330 = n12329 ^ x14 ;
  assign n12114 = x121 & n884 ;
  assign n12331 = n12330 ^ n12114 ;
  assign n12113 = x123 & n789 ;
  assign n12332 = n12331 ^ n12113 ;
  assign n12112 = n790 & ~n9804 ;
  assign n12333 = n12332 ^ n12112 ;
  assign n12335 = n12334 ^ n12333 ;
  assign n12109 = n12050 ^ n12041 ;
  assign n12110 = n12047 & n12109 ;
  assign n12111 = n12110 ^ n12050 ;
  assign n12336 = n12335 ^ n12111 ;
  assign n12337 = n12336 ^ x11 ;
  assign n12108 = x124 & n650 ;
  assign n12338 = n12337 ^ n12108 ;
  assign n12107 = x126 & ~n578 ;
  assign n12339 = n12338 ^ n12107 ;
  assign n12106 = ~n579 & n10461 ;
  assign n12340 = n12339 ^ n12106 ;
  assign n12342 = n12341 ^ n12340 ;
  assign n12346 = n12345 ^ n12342 ;
  assign n12351 = n12350 ^ n12346 ;
  assign n12352 = n12351 ^ n12346 ;
  assign n12356 = ~x7 & ~x127 ;
  assign n12357 = n12356 ^ n383 ;
  assign n12358 = ~n10154 & n12357 ;
  assign n12359 = n12358 ^ x8 ;
  assign n12360 = n336 & ~n12359 ;
  assign n12361 = n12352 & n12360 ;
  assign n12362 = n12361 ^ n12351 ;
  assign n12366 = n12365 ^ n12362 ;
  assign n12103 = n12076 ^ n12068 ;
  assign n12104 = ~n12073 & ~n12103 ;
  assign n12105 = n12104 ^ n12076 ;
  assign n12367 = n12366 ^ n12105 ;
  assign n12100 = n12098 ^ n11827 ;
  assign n12101 = n12078 & n12100 ;
  assign n12102 = n12101 ^ n12098 ;
  assign n12368 = n12367 ^ n12102 ;
  assign n12614 = n12365 ^ n12346 ;
  assign n12615 = n12362 & ~n12614 ;
  assign n12616 = n12615 ^ n12362 ;
  assign n12607 = x125 & n650 ;
  assign n12606 = x127 & ~n578 ;
  assign n12608 = n12607 ^ n12606 ;
  assign n12609 = n12608 ^ x11 ;
  assign n12605 = ~n579 & n10986 ;
  assign n12610 = n12609 ^ n12605 ;
  assign n12604 = x126 & n584 ;
  assign n12611 = n12610 ^ n12604 ;
  assign n12600 = n12329 ^ n12111 ;
  assign n12601 = n12335 & ~n12600 ;
  assign n12602 = n12601 ^ n12329 ;
  assign n12598 = x123 & n795 ;
  assign n12590 = n12322 ^ n12117 ;
  assign n12591 = ~n12328 & n12590 ;
  assign n12592 = n12591 ^ n12322 ;
  assign n12588 = x120 & n1068 ;
  assign n12581 = x117 & n1348 ;
  assign n12573 = n12305 ^ n12126 ;
  assign n12574 = n12311 & n12573 ;
  assign n12575 = n12574 ^ n12305 ;
  assign n12571 = x114 & n1673 ;
  assign n12564 = x111 & n2025 ;
  assign n12557 = x108 & n2435 ;
  assign n12549 = n12281 ^ n12141 ;
  assign n12550 = n12287 & ~n12549 ;
  assign n12551 = n12550 ^ n12281 ;
  assign n12547 = x105 & n2899 ;
  assign n12539 = n12274 ^ n12147 ;
  assign n12540 = ~n12280 & n12539 ;
  assign n12541 = n12540 ^ n12274 ;
  assign n12537 = x102 & n3395 ;
  assign n12529 = n12267 ^ n12153 ;
  assign n12530 = ~n12273 & ~n12529 ;
  assign n12531 = n12530 ^ n12267 ;
  assign n12527 = x99 & n3940 ;
  assign n12519 = n12265 ^ n12159 ;
  assign n12520 = ~n12266 & n12519 ;
  assign n12521 = n12520 ^ n12265 ;
  assign n12513 = x95 & n4482 ;
  assign n12512 = x97 & n4478 ;
  assign n12514 = n12513 ^ n12512 ;
  assign n12515 = n12514 ^ x41 ;
  assign n12511 = n3501 & n4479 ;
  assign n12516 = n12515 ^ n12511 ;
  assign n12510 = x96 & n4475 ;
  assign n12517 = n12516 ^ n12510 ;
  assign n12504 = x92 & n5113 ;
  assign n12503 = x94 & n5116 ;
  assign n12505 = n12504 ^ n12503 ;
  assign n12506 = n12505 ^ x44 ;
  assign n12502 = n3010 & n5117 ;
  assign n12507 = n12506 ^ n12502 ;
  assign n12501 = x93 & n5121 ;
  assign n12508 = n12507 ^ n12501 ;
  assign n12498 = n12247 ^ n12162 ;
  assign n12499 = ~n12256 & ~n12498 ;
  assign n12489 = x89 & n5981 ;
  assign n12488 = x91 & n5748 ;
  assign n12490 = n12489 ^ n12488 ;
  assign n12491 = n12490 ^ x47 ;
  assign n12487 = n2548 & n5749 ;
  assign n12492 = n12491 ^ n12487 ;
  assign n12486 = x90 & n5755 ;
  assign n12493 = n12492 ^ n12486 ;
  assign n12482 = n12244 ^ n12177 ;
  assign n12483 = ~n12245 & n12482 ;
  assign n12484 = n12483 ^ n12244 ;
  assign n12476 = x86 & n6687 ;
  assign n12475 = x88 & n6444 ;
  assign n12477 = n12476 ^ n12475 ;
  assign n12478 = n12477 ^ x50 ;
  assign n12474 = n2131 & n6445 ;
  assign n12479 = n12478 ^ n12474 ;
  assign n12473 = x87 & n6449 ;
  assign n12480 = n12479 ^ n12473 ;
  assign n12469 = n12234 ^ n12180 ;
  assign n12470 = ~n12235 & n12469 ;
  assign n12471 = n12470 ^ n12234 ;
  assign n12467 = x84 & n7191 ;
  assign n12460 = x81 & n7947 ;
  assign n12458 = n1422 & n7951 ;
  assign n12454 = x80 & n7954 ;
  assign n12453 = x82 & n7950 ;
  assign n12455 = n12454 ^ n12453 ;
  assign n12456 = n12455 ^ x56 ;
  assign n12449 = ~n12200 & ~n12211 ;
  assign n12450 = n12449 ^ n12208 ;
  assign n12441 = x74 & n9655 ;
  assign n12440 = x76 & n9651 ;
  assign n12442 = n12441 ^ n12440 ;
  assign n12443 = n12442 ^ x62 ;
  assign n12439 = ~n863 & n9652 ;
  assign n12444 = n12443 ^ n12439 ;
  assign n12438 = x75 & n9648 ;
  assign n12445 = n12444 ^ n12438 ;
  assign n12446 = n12445 ^ x8 ;
  assign n12434 = x73 ^ x71 ;
  assign n12435 = ~n11895 & n12434 ;
  assign n12436 = n12435 ^ n420 ;
  assign n12437 = n12206 & n12436 ;
  assign n12447 = n12446 ^ n12437 ;
  assign n12451 = n12450 ^ n12447 ;
  assign n12424 = x77 & n8750 ;
  assign n12423 = x79 & n8746 ;
  assign n12425 = n12424 ^ n12423 ;
  assign n12426 = n12425 ^ x59 ;
  assign n12422 = n1123 & n8747 ;
  assign n12427 = n12426 ^ n12422 ;
  assign n12421 = x78 & n8743 ;
  assign n12428 = n12427 ^ n12421 ;
  assign n12429 = n12428 ^ n12212 ;
  assign n12430 = n12429 ^ n12191 ;
  assign n12431 = n12430 ^ n12428 ;
  assign n12432 = ~n12197 & ~n12431 ;
  assign n12433 = n12432 ^ n12429 ;
  assign n12452 = n12451 ^ n12433 ;
  assign n12457 = n12456 ^ n12452 ;
  assign n12459 = n12458 ^ n12457 ;
  assign n12461 = n12460 ^ n12459 ;
  assign n12418 = n12225 ^ n12221 ;
  assign n12419 = n12222 & n12418 ;
  assign n12420 = n12419 ^ n12225 ;
  assign n12462 = n12461 ^ n12420 ;
  assign n12463 = n12462 ^ x53 ;
  assign n12417 = x83 & n7183 ;
  assign n12464 = n12463 ^ n12417 ;
  assign n12416 = x85 & n7186 ;
  assign n12465 = n12464 ^ n12416 ;
  assign n12415 = n1748 & n7187 ;
  assign n12466 = n12465 ^ n12415 ;
  assign n12468 = n12467 ^ n12466 ;
  assign n12472 = n12471 ^ n12468 ;
  assign n12481 = n12480 ^ n12472 ;
  assign n12485 = n12484 ^ n12481 ;
  assign n12494 = n12493 ^ n12485 ;
  assign n12412 = n12246 ^ n12168 ;
  assign n12413 = ~n12174 & ~n12412 ;
  assign n12414 = n12413 ^ n12246 ;
  assign n12495 = n12494 ^ n12414 ;
  assign n12496 = n12495 ^ n12247 ;
  assign n12500 = n12499 ^ n12496 ;
  assign n12509 = n12508 ^ n12500 ;
  assign n12518 = n12517 ^ n12509 ;
  assign n12522 = n12521 ^ n12518 ;
  assign n12523 = n12522 ^ x38 ;
  assign n12411 = x98 & n3932 ;
  assign n12524 = n12523 ^ n12411 ;
  assign n12410 = x100 & n3935 ;
  assign n12525 = n12524 ^ n12410 ;
  assign n12409 = n3936 & n4048 ;
  assign n12526 = n12525 ^ n12409 ;
  assign n12528 = n12527 ^ n12526 ;
  assign n12532 = n12531 ^ n12528 ;
  assign n12533 = n12532 ^ x35 ;
  assign n12408 = x101 & n3387 ;
  assign n12534 = n12533 ^ n12408 ;
  assign n12407 = x103 & n3390 ;
  assign n12535 = n12534 ^ n12407 ;
  assign n12406 = n3391 & ~n4624 ;
  assign n12536 = n12535 ^ n12406 ;
  assign n12538 = n12537 ^ n12536 ;
  assign n12542 = n12541 ^ n12538 ;
  assign n12543 = n12542 ^ x32 ;
  assign n12405 = x104 & n2890 ;
  assign n12544 = n12543 ^ n12405 ;
  assign n12404 = x106 & n2893 ;
  assign n12545 = n12544 ^ n12404 ;
  assign n12403 = n2894 & ~n5257 ;
  assign n12546 = n12545 ^ n12403 ;
  assign n12548 = n12547 ^ n12546 ;
  assign n12552 = n12551 ^ n12548 ;
  assign n12553 = n12552 ^ x29 ;
  assign n12402 = x107 & n2593 ;
  assign n12554 = n12553 ^ n12402 ;
  assign n12401 = x109 & n2428 ;
  assign n12555 = n12554 ^ n12401 ;
  assign n12400 = n2429 & n5912 ;
  assign n12556 = n12555 ^ n12400 ;
  assign n12558 = n12557 ^ n12556 ;
  assign n12397 = n12288 ^ n12135 ;
  assign n12398 = ~n12294 & ~n12397 ;
  assign n12399 = n12398 ^ n12288 ;
  assign n12559 = n12558 ^ n12399 ;
  assign n12560 = n12559 ^ x26 ;
  assign n12396 = x110 & n2032 ;
  assign n12561 = n12560 ^ n12396 ;
  assign n12395 = x112 & n2028 ;
  assign n12562 = n12561 ^ n12395 ;
  assign n12394 = n2029 & ~n6616 ;
  assign n12563 = n12562 ^ n12394 ;
  assign n12565 = n12564 ^ n12563 ;
  assign n12391 = n12304 ^ n12295 ;
  assign n12392 = n12301 & n12391 ;
  assign n12393 = n12392 ^ n12304 ;
  assign n12566 = n12565 ^ n12393 ;
  assign n12567 = n12566 ^ x23 ;
  assign n12390 = x113 & n1665 ;
  assign n12568 = n12567 ^ n12390 ;
  assign n12389 = x115 & n1668 ;
  assign n12569 = n12568 ^ n12389 ;
  assign n12388 = n1669 & ~n7353 ;
  assign n12570 = n12569 ^ n12388 ;
  assign n12572 = n12571 ^ n12570 ;
  assign n12576 = n12575 ^ n12572 ;
  assign n12577 = n12576 ^ x20 ;
  assign n12387 = x116 & n1340 ;
  assign n12578 = n12577 ^ n12387 ;
  assign n12386 = x118 & n1343 ;
  assign n12579 = n12578 ^ n12386 ;
  assign n12385 = n1344 & ~n8140 ;
  assign n12580 = n12579 ^ n12385 ;
  assign n12582 = n12581 ^ n12580 ;
  assign n12382 = n12321 ^ n12312 ;
  assign n12383 = ~n12318 & ~n12382 ;
  assign n12384 = n12383 ^ n12321 ;
  assign n12583 = n12582 ^ n12384 ;
  assign n12584 = n12583 ^ x17 ;
  assign n12381 = x119 & n1060 ;
  assign n12585 = n12584 ^ n12381 ;
  assign n12380 = x121 & n1063 ;
  assign n12586 = n12585 ^ n12380 ;
  assign n12379 = n1064 & n8979 ;
  assign n12587 = n12586 ^ n12379 ;
  assign n12589 = n12588 ^ n12587 ;
  assign n12593 = n12592 ^ n12589 ;
  assign n12594 = n12593 ^ x14 ;
  assign n12378 = x122 & n884 ;
  assign n12595 = n12594 ^ n12378 ;
  assign n12377 = x124 & n789 ;
  assign n12596 = n12595 ^ n12377 ;
  assign n12376 = n790 & n10117 ;
  assign n12597 = n12596 ^ n12376 ;
  assign n12599 = n12598 ^ n12597 ;
  assign n12603 = n12602 ^ n12599 ;
  assign n12612 = n12611 ^ n12603 ;
  assign n12373 = n12345 ^ n12336 ;
  assign n12374 = n12342 & ~n12373 ;
  assign n12375 = n12374 ^ n12345 ;
  assign n12613 = n12612 ^ n12375 ;
  assign n12617 = n12616 ^ n12613 ;
  assign n12369 = n12105 ^ n12102 ;
  assign n12370 = n12365 ^ n12105 ;
  assign n12371 = n12370 ^ n12362 ;
  assign n12372 = n12369 & n12371 ;
  assign n12618 = n12617 ^ n12372 ;
  assign n12862 = n12615 ^ n12365 ;
  assign n12863 = ~n12613 & n12862 ;
  assign n12864 = n12613 ^ n12365 ;
  assign n12865 = n12362 & ~n12864 ;
  assign n12866 = n12613 ^ n12346 ;
  assign n12867 = n12865 & n12866 ;
  assign n12868 = n12867 ^ n12613 ;
  assign n12869 = ~n12105 & ~n12868 ;
  assign n12870 = ~n12863 & ~n12869 ;
  assign n12871 = n12862 ^ n12613 ;
  assign n12872 = n12871 ^ n12863 ;
  assign n12873 = n12868 ^ n12105 ;
  assign n12874 = n12873 ^ n12869 ;
  assign n12875 = ~n12872 & n12874 ;
  assign n12876 = n12102 & n12875 ;
  assign n12877 = n12870 & ~n12876 ;
  assign n12858 = n12611 ^ n12375 ;
  assign n12859 = ~n12612 & n12858 ;
  assign n12860 = n12859 ^ n12611 ;
  assign n12855 = x127 & n584 ;
  assign n12849 = x124 & n795 ;
  assign n12841 = n12576 ^ n12384 ;
  assign n12842 = ~n12582 & n12841 ;
  assign n12843 = n12842 ^ n12576 ;
  assign n12839 = x121 & n1068 ;
  assign n12832 = x118 & n1348 ;
  assign n12824 = n12559 ^ n12393 ;
  assign n12825 = n12565 & ~n12824 ;
  assign n12826 = n12825 ^ n12559 ;
  assign n12822 = x115 & n1673 ;
  assign n12815 = x112 & n2025 ;
  assign n12808 = x109 & n2435 ;
  assign n12801 = x106 & n2899 ;
  assign n12794 = x103 & n3395 ;
  assign n12783 = x99 & n3932 ;
  assign n12782 = x101 & n3935 ;
  assign n12784 = n12783 ^ n12782 ;
  assign n12785 = n12784 ^ x38 ;
  assign n12781 = n3936 & n4223 ;
  assign n12786 = n12785 ^ n12781 ;
  assign n12780 = x100 & n3940 ;
  assign n12787 = n12786 ^ n12780 ;
  assign n12777 = x97 & n4475 ;
  assign n12775 = n3673 & n4479 ;
  assign n12771 = x96 & n4482 ;
  assign n12770 = x98 & n4478 ;
  assign n12772 = n12771 ^ n12770 ;
  assign n12773 = n12772 ^ x41 ;
  assign n12767 = x94 & n5121 ;
  assign n12765 = n3166 & n5117 ;
  assign n12761 = x93 & n5113 ;
  assign n12760 = x95 & n5116 ;
  assign n12762 = n12761 ^ n12760 ;
  assign n12763 = n12762 ^ x44 ;
  assign n12753 = x90 & n5981 ;
  assign n12752 = x92 & n5748 ;
  assign n12754 = n12753 ^ n12752 ;
  assign n12755 = n12754 ^ x47 ;
  assign n12751 = n2696 & n5749 ;
  assign n12756 = n12755 ^ n12751 ;
  assign n12750 = x91 & n5755 ;
  assign n12757 = n12756 ^ n12750 ;
  assign n12743 = x87 & n6687 ;
  assign n12742 = x89 & n6444 ;
  assign n12744 = n12743 ^ n12742 ;
  assign n12745 = n12744 ^ x50 ;
  assign n12741 = n2255 & n6445 ;
  assign n12746 = n12745 ^ n12741 ;
  assign n12740 = x88 & n6449 ;
  assign n12747 = n12746 ^ n12740 ;
  assign n12732 = x81 & n7954 ;
  assign n12731 = x83 & n7950 ;
  assign n12733 = n12732 ^ n12731 ;
  assign n12734 = n12733 ^ x56 ;
  assign n12730 = n1517 & n7951 ;
  assign n12735 = n12734 ^ n12730 ;
  assign n12729 = x82 & n7947 ;
  assign n12736 = n12735 ^ n12729 ;
  assign n12722 = x78 & n8750 ;
  assign n12721 = x80 & n8746 ;
  assign n12723 = n12722 ^ n12721 ;
  assign n12724 = n12723 ^ x59 ;
  assign n12720 = n1217 & n8747 ;
  assign n12725 = n12724 ^ n12720 ;
  assign n12719 = x79 & n8743 ;
  assign n12726 = n12725 ^ n12719 ;
  assign n12713 = x75 & n9655 ;
  assign n12712 = x77 & n9651 ;
  assign n12714 = n12713 ^ n12712 ;
  assign n12715 = n12714 ^ x62 ;
  assign n12711 = ~n943 & n9652 ;
  assign n12716 = n12715 ^ n12711 ;
  assign n12710 = x76 & n9648 ;
  assign n12717 = n12716 ^ n12710 ;
  assign n12707 = x73 & n11895 ;
  assign n12706 = x74 & n9956 ;
  assign n12708 = n12707 ^ n12706 ;
  assign n12700 = x72 ^ x8 ;
  assign n12703 = n12436 & ~n12700 ;
  assign n12704 = n12703 ^ x72 ;
  assign n12705 = n12206 & n12704 ;
  assign n12709 = n12708 ^ n12705 ;
  assign n12718 = n12717 ^ n12709 ;
  assign n12727 = n12726 ^ n12718 ;
  assign n12697 = n12450 ^ n12445 ;
  assign n12698 = n12447 & ~n12697 ;
  assign n12699 = n12698 ^ n12450 ;
  assign n12728 = n12727 ^ n12699 ;
  assign n12737 = n12736 ^ n12728 ;
  assign n12694 = n12451 ^ n12428 ;
  assign n12695 = ~n12433 & n12694 ;
  assign n12696 = n12695 ^ n12428 ;
  assign n12738 = n12737 ^ n12696 ;
  assign n12691 = n12452 ^ n12420 ;
  assign n12692 = ~n12461 & ~n12691 ;
  assign n12684 = x84 & n7183 ;
  assign n12683 = x86 & n7186 ;
  assign n12685 = n12684 ^ n12683 ;
  assign n12686 = n12685 ^ x53 ;
  assign n12682 = n1868 & n7187 ;
  assign n12687 = n12686 ^ n12682 ;
  assign n12681 = x85 & n7191 ;
  assign n12688 = n12687 ^ n12681 ;
  assign n12689 = n12688 ^ n12452 ;
  assign n12693 = n12692 ^ n12689 ;
  assign n12739 = n12738 ^ n12693 ;
  assign n12748 = n12747 ^ n12739 ;
  assign n12678 = n12471 ^ n12462 ;
  assign n12679 = n12468 & ~n12678 ;
  assign n12680 = n12679 ^ n12471 ;
  assign n12749 = n12748 ^ n12680 ;
  assign n12758 = n12757 ^ n12749 ;
  assign n12675 = n12484 ^ n12480 ;
  assign n12676 = n12481 & n12675 ;
  assign n12677 = n12676 ^ n12484 ;
  assign n12759 = n12758 ^ n12677 ;
  assign n12764 = n12763 ^ n12759 ;
  assign n12766 = n12765 ^ n12764 ;
  assign n12768 = n12767 ^ n12766 ;
  assign n12672 = n12493 ^ n12414 ;
  assign n12673 = ~n12494 & ~n12672 ;
  assign n12674 = n12673 ^ n12493 ;
  assign n12769 = n12768 ^ n12674 ;
  assign n12774 = n12773 ^ n12769 ;
  assign n12776 = n12775 ^ n12774 ;
  assign n12778 = n12777 ^ n12776 ;
  assign n12669 = n12508 ^ n12495 ;
  assign n12670 = ~n12500 & n12669 ;
  assign n12671 = n12670 ^ n12495 ;
  assign n12779 = n12778 ^ n12671 ;
  assign n12788 = n12787 ^ n12779 ;
  assign n12666 = n12521 ^ n12517 ;
  assign n12667 = n12518 & n12666 ;
  assign n12668 = n12667 ^ n12521 ;
  assign n12789 = n12788 ^ n12668 ;
  assign n12790 = n12789 ^ x35 ;
  assign n12665 = x102 & n3387 ;
  assign n12791 = n12790 ^ n12665 ;
  assign n12664 = x104 & n3390 ;
  assign n12792 = n12791 ^ n12664 ;
  assign n12663 = n3391 & ~n4830 ;
  assign n12793 = n12792 ^ n12663 ;
  assign n12795 = n12794 ^ n12793 ;
  assign n12660 = n12531 ^ n12522 ;
  assign n12661 = n12528 & n12660 ;
  assign n12662 = n12661 ^ n12531 ;
  assign n12796 = n12795 ^ n12662 ;
  assign n12797 = n12796 ^ x32 ;
  assign n12659 = x105 & n2890 ;
  assign n12798 = n12797 ^ n12659 ;
  assign n12658 = x107 & n2893 ;
  assign n12799 = n12798 ^ n12658 ;
  assign n12657 = n2894 & ~n5459 ;
  assign n12800 = n12799 ^ n12657 ;
  assign n12802 = n12801 ^ n12800 ;
  assign n12654 = n12541 ^ n12532 ;
  assign n12655 = ~n12538 & ~n12654 ;
  assign n12656 = n12655 ^ n12541 ;
  assign n12803 = n12802 ^ n12656 ;
  assign n12804 = n12803 ^ x29 ;
  assign n12653 = x108 & n2593 ;
  assign n12805 = n12804 ^ n12653 ;
  assign n12652 = x110 & n2428 ;
  assign n12806 = n12805 ^ n12652 ;
  assign n12651 = n2429 & n6145 ;
  assign n12807 = n12806 ^ n12651 ;
  assign n12809 = n12808 ^ n12807 ;
  assign n12648 = n12551 ^ n12542 ;
  assign n12649 = n12548 & ~n12648 ;
  assign n12650 = n12649 ^ n12551 ;
  assign n12810 = n12809 ^ n12650 ;
  assign n12811 = n12810 ^ x26 ;
  assign n12647 = x111 & n2032 ;
  assign n12812 = n12811 ^ n12647 ;
  assign n12646 = x113 & n2028 ;
  assign n12813 = n12812 ^ n12646 ;
  assign n12645 = n2029 & ~n6849 ;
  assign n12814 = n12813 ^ n12645 ;
  assign n12816 = n12815 ^ n12814 ;
  assign n12642 = n12552 ^ n12399 ;
  assign n12643 = ~n12558 & n12642 ;
  assign n12644 = n12643 ^ n12552 ;
  assign n12817 = n12816 ^ n12644 ;
  assign n12818 = n12817 ^ x23 ;
  assign n12641 = x114 & n1665 ;
  assign n12819 = n12818 ^ n12641 ;
  assign n12640 = x116 & n1668 ;
  assign n12820 = n12819 ^ n12640 ;
  assign n12639 = n1669 & ~n7604 ;
  assign n12821 = n12820 ^ n12639 ;
  assign n12823 = n12822 ^ n12821 ;
  assign n12827 = n12826 ^ n12823 ;
  assign n12828 = n12827 ^ x20 ;
  assign n12638 = x117 & n1340 ;
  assign n12829 = n12828 ^ n12638 ;
  assign n12637 = x119 & n1343 ;
  assign n12830 = n12829 ^ n12637 ;
  assign n12636 = n1344 & n8405 ;
  assign n12831 = n12830 ^ n12636 ;
  assign n12833 = n12832 ^ n12831 ;
  assign n12633 = n12575 ^ n12566 ;
  assign n12634 = n12572 & ~n12633 ;
  assign n12635 = n12634 ^ n12575 ;
  assign n12834 = n12833 ^ n12635 ;
  assign n12835 = n12834 ^ x17 ;
  assign n12632 = x120 & n1060 ;
  assign n12836 = n12835 ^ n12632 ;
  assign n12631 = x122 & n1063 ;
  assign n12837 = n12836 ^ n12631 ;
  assign n12630 = n1064 & ~n9261 ;
  assign n12838 = n12837 ^ n12630 ;
  assign n12840 = n12839 ^ n12838 ;
  assign n12844 = n12843 ^ n12840 ;
  assign n12845 = n12844 ^ x14 ;
  assign n12629 = x123 & n884 ;
  assign n12846 = n12845 ^ n12629 ;
  assign n12628 = x125 & n789 ;
  assign n12847 = n12846 ^ n12628 ;
  assign n12627 = n790 & n10416 ;
  assign n12848 = n12847 ^ n12627 ;
  assign n12850 = n12849 ^ n12848 ;
  assign n12624 = n12592 ^ n12583 ;
  assign n12625 = ~n12589 & ~n12624 ;
  assign n12626 = n12625 ^ n12592 ;
  assign n12851 = n12850 ^ n12626 ;
  assign n12852 = n12851 ^ x11 ;
  assign n12623 = x126 & n650 ;
  assign n12853 = n12852 ^ n12623 ;
  assign n12622 = ~n579 & n10155 ;
  assign n12854 = n12853 ^ n12622 ;
  assign n12856 = n12855 ^ n12854 ;
  assign n12619 = n12602 ^ n12593 ;
  assign n12620 = n12599 & ~n12619 ;
  assign n12621 = n12620 ^ n12602 ;
  assign n12857 = n12856 ^ n12621 ;
  assign n12861 = n12860 ^ n12857 ;
  assign n12878 = n12877 ^ n12861 ;
  assign n13130 = n12851 ^ n12621 ;
  assign n13131 = n12856 & n13130 ;
  assign n13132 = n13131 ^ n12851 ;
  assign n13126 = n12844 ^ n12626 ;
  assign n13127 = ~n12850 & n13126 ;
  assign n13128 = n13127 ^ n12844 ;
  assign n12882 = n514 ^ x10 ;
  assign n12883 = x127 & n12882 ;
  assign n13108 = x125 & n795 ;
  assign n13100 = n12827 ^ n12635 ;
  assign n13101 = n12833 & n13100 ;
  assign n13102 = n13101 ^ n12827 ;
  assign n13098 = x122 & n1068 ;
  assign n13091 = x119 & n1348 ;
  assign n13084 = x116 & n1673 ;
  assign n13076 = n12803 ^ n12650 ;
  assign n13077 = ~n12809 & ~n13076 ;
  assign n13078 = n13077 ^ n12803 ;
  assign n13074 = x113 & n2025 ;
  assign n13066 = n12796 ^ n12656 ;
  assign n13067 = n12802 & ~n13066 ;
  assign n13068 = n13067 ^ n12796 ;
  assign n13064 = x110 & n2435 ;
  assign n13056 = n12789 ^ n12662 ;
  assign n13057 = ~n12795 & n13056 ;
  assign n13058 = n13057 ^ n12789 ;
  assign n13054 = x107 & n2899 ;
  assign n13046 = n12787 ^ n12668 ;
  assign n13047 = ~n12788 & n13046 ;
  assign n13048 = n13047 ^ n12787 ;
  assign n13040 = x103 & n3387 ;
  assign n13039 = x105 & n3390 ;
  assign n13041 = n13040 ^ n13039 ;
  assign n13042 = n13041 ^ x35 ;
  assign n13038 = n3391 & ~n5034 ;
  assign n13043 = n13042 ^ n13038 ;
  assign n13037 = x104 & n3395 ;
  assign n13044 = n13043 ^ n13037 ;
  assign n13031 = x100 & n3932 ;
  assign n13030 = x102 & n3935 ;
  assign n13032 = n13031 ^ n13030 ;
  assign n13033 = n13032 ^ x38 ;
  assign n13029 = n3936 & n4425 ;
  assign n13034 = n13033 ^ n13029 ;
  assign n13028 = x101 & n3940 ;
  assign n13035 = n13034 ^ n13028 ;
  assign n13024 = n12769 ^ n12671 ;
  assign n13025 = ~n12778 & ~n13024 ;
  assign n13026 = n13025 ^ n12769 ;
  assign n13018 = x97 & n4482 ;
  assign n13017 = x99 & n4478 ;
  assign n13019 = n13018 ^ n13017 ;
  assign n13020 = n13019 ^ x41 ;
  assign n13016 = n3851 & n4479 ;
  assign n13021 = n13020 ^ n13016 ;
  assign n13015 = x98 & n4475 ;
  assign n13022 = n13021 ^ n13015 ;
  assign n13007 = x95 & n5121 ;
  assign n13005 = n3336 & n5117 ;
  assign n13001 = x94 & n5113 ;
  assign n13000 = x96 & n5116 ;
  assign n13002 = n13001 ^ n13000 ;
  assign n13003 = n13002 ^ x44 ;
  assign n12996 = n12747 ^ n12680 ;
  assign n12997 = ~n12748 & n12996 ;
  assign n12998 = n12997 ^ n12747 ;
  assign n12990 = x91 & n5981 ;
  assign n12989 = x93 & n5748 ;
  assign n12991 = n12990 ^ n12989 ;
  assign n12992 = n12991 ^ x47 ;
  assign n12988 = n2842 & n5749 ;
  assign n12993 = n12992 ^ n12988 ;
  assign n12987 = x92 & n5755 ;
  assign n12994 = n12993 ^ n12987 ;
  assign n12979 = x85 & n7183 ;
  assign n12978 = x87 & n7186 ;
  assign n12980 = n12979 ^ n12978 ;
  assign n12981 = n12980 ^ x53 ;
  assign n12977 = n1987 & n7187 ;
  assign n12982 = n12981 ^ n12977 ;
  assign n12976 = x86 & n7191 ;
  assign n12983 = n12982 ^ n12976 ;
  assign n12972 = n12726 ^ n12699 ;
  assign n12973 = ~n12727 & ~n12972 ;
  assign n12974 = n12973 ^ n12726 ;
  assign n12966 = x82 & n7954 ;
  assign n12965 = x84 & n7950 ;
  assign n12967 = n12966 ^ n12965 ;
  assign n12968 = n12967 ^ x56 ;
  assign n12964 = n1635 & n7951 ;
  assign n12969 = n12968 ^ n12964 ;
  assign n12963 = x83 & n7947 ;
  assign n12970 = n12969 ^ n12963 ;
  assign n12957 = x79 & n8750 ;
  assign n12956 = x81 & n8746 ;
  assign n12958 = n12957 ^ n12956 ;
  assign n12959 = n12958 ^ x59 ;
  assign n12955 = n1310 & n8747 ;
  assign n12960 = n12959 ^ n12955 ;
  assign n12954 = x80 & n8743 ;
  assign n12961 = n12960 ^ n12954 ;
  assign n12948 = x76 & n9655 ;
  assign n12947 = x78 & n9651 ;
  assign n12949 = n12948 ^ n12947 ;
  assign n12950 = n12949 ^ x62 ;
  assign n12946 = ~n1036 & n9652 ;
  assign n12951 = n12950 ^ n12946 ;
  assign n12945 = x77 & n9648 ;
  assign n12952 = n12951 ^ n12945 ;
  assign n543 = x74 ^ x73 ;
  assign n12940 = x63 & n543 ;
  assign n618 = x75 ^ x74 ;
  assign n12941 = n12940 ^ n618 ;
  assign n12942 = ~n9956 & n12941 ;
  assign n12943 = n12942 ^ n618 ;
  assign n12933 = n12717 ^ n12708 ;
  assign n12934 = n12709 & ~n12933 ;
  assign n12935 = n12934 ^ n12717 ;
  assign n12944 = n12943 ^ n12935 ;
  assign n12953 = n12952 ^ n12944 ;
  assign n12962 = n12961 ^ n12953 ;
  assign n12971 = n12970 ^ n12962 ;
  assign n12975 = n12974 ^ n12971 ;
  assign n12984 = n12983 ^ n12975 ;
  assign n12930 = n12736 ^ n12696 ;
  assign n12931 = n12737 & n12930 ;
  assign n12932 = n12931 ^ n12736 ;
  assign n12985 = n12984 ^ n12932 ;
  assign n12920 = x88 & n6687 ;
  assign n12919 = x90 & n6444 ;
  assign n12921 = n12920 ^ n12919 ;
  assign n12922 = n12921 ^ x50 ;
  assign n12918 = n2398 & n6445 ;
  assign n12923 = n12922 ^ n12918 ;
  assign n12917 = x89 & n6449 ;
  assign n12924 = n12923 ^ n12917 ;
  assign n12926 = n12924 ^ n12688 ;
  assign n12925 = n12924 ^ n12738 ;
  assign n12927 = n12926 ^ n12925 ;
  assign n12928 = ~n12693 & n12927 ;
  assign n12929 = n12928 ^ n12926 ;
  assign n12986 = n12985 ^ n12929 ;
  assign n12995 = n12994 ^ n12986 ;
  assign n12999 = n12998 ^ n12995 ;
  assign n13004 = n13003 ^ n12999 ;
  assign n13006 = n13005 ^ n13004 ;
  assign n13008 = n13007 ^ n13006 ;
  assign n12914 = n12757 ^ n12677 ;
  assign n12915 = ~n12758 & n12914 ;
  assign n12916 = n12915 ^ n12757 ;
  assign n13009 = n13008 ^ n12916 ;
  assign n13010 = n13009 ^ n12759 ;
  assign n13011 = n13010 ^ n12674 ;
  assign n13012 = n13011 ^ n13009 ;
  assign n13013 = ~n12768 & ~n13012 ;
  assign n13014 = n13013 ^ n13010 ;
  assign n13023 = n13022 ^ n13014 ;
  assign n13027 = n13026 ^ n13023 ;
  assign n13036 = n13035 ^ n13027 ;
  assign n13045 = n13044 ^ n13036 ;
  assign n13049 = n13048 ^ n13045 ;
  assign n13050 = n13049 ^ x32 ;
  assign n12913 = x106 & n2890 ;
  assign n13051 = n13050 ^ n12913 ;
  assign n12912 = x108 & n2893 ;
  assign n13052 = n13051 ^ n12912 ;
  assign n12911 = n2894 & n5687 ;
  assign n13053 = n13052 ^ n12911 ;
  assign n13055 = n13054 ^ n13053 ;
  assign n13059 = n13058 ^ n13055 ;
  assign n13060 = n13059 ^ x29 ;
  assign n12910 = x109 & n2593 ;
  assign n13061 = n13060 ^ n12910 ;
  assign n12909 = x111 & n2428 ;
  assign n13062 = n13061 ^ n12909 ;
  assign n12908 = n2429 & ~n6370 ;
  assign n13063 = n13062 ^ n12908 ;
  assign n13065 = n13064 ^ n13063 ;
  assign n13069 = n13068 ^ n13065 ;
  assign n13070 = n13069 ^ x26 ;
  assign n12907 = x112 & n2032 ;
  assign n13071 = n13070 ^ n12907 ;
  assign n12906 = x114 & n2028 ;
  assign n13072 = n13071 ^ n12906 ;
  assign n12905 = n2029 & ~n7108 ;
  assign n13073 = n13072 ^ n12905 ;
  assign n13075 = n13074 ^ n13073 ;
  assign n13079 = n13078 ^ n13075 ;
  assign n13080 = n13079 ^ x23 ;
  assign n12904 = x115 & n1665 ;
  assign n13081 = n13080 ^ n12904 ;
  assign n12903 = x117 & n1668 ;
  assign n13082 = n13081 ^ n12903 ;
  assign n12902 = n1669 & ~n7860 ;
  assign n13083 = n13082 ^ n12902 ;
  assign n13085 = n13084 ^ n13083 ;
  assign n12899 = n12810 ^ n12644 ;
  assign n12900 = ~n12816 & n12899 ;
  assign n12901 = n12900 ^ n12810 ;
  assign n13086 = n13085 ^ n12901 ;
  assign n13087 = n13086 ^ x20 ;
  assign n12898 = x118 & n1340 ;
  assign n13088 = n13087 ^ n12898 ;
  assign n12897 = x120 & n1343 ;
  assign n13089 = n13088 ^ n12897 ;
  assign n12896 = n1344 & n8904 ;
  assign n13090 = n13089 ^ n12896 ;
  assign n13092 = n13091 ^ n13090 ;
  assign n12893 = n12826 ^ n12817 ;
  assign n12894 = ~n12823 & n12893 ;
  assign n12895 = n12894 ^ n12826 ;
  assign n13093 = n13092 ^ n12895 ;
  assign n13094 = n13093 ^ x17 ;
  assign n12892 = x121 & n1060 ;
  assign n13095 = n13094 ^ n12892 ;
  assign n12891 = x123 & n1063 ;
  assign n13096 = n13095 ^ n12891 ;
  assign n12890 = n1064 & ~n9804 ;
  assign n13097 = n13096 ^ n12890 ;
  assign n13099 = n13098 ^ n13097 ;
  assign n13103 = n13102 ^ n13099 ;
  assign n13104 = n13103 ^ x14 ;
  assign n12889 = x124 & n884 ;
  assign n13105 = n13104 ^ n12889 ;
  assign n12888 = x126 & n789 ;
  assign n13106 = n13105 ^ n12888 ;
  assign n12887 = n790 & n10461 ;
  assign n13107 = n13106 ^ n12887 ;
  assign n13109 = n13108 ^ n13107 ;
  assign n12884 = n12843 ^ n12834 ;
  assign n12885 = ~n12840 & ~n12884 ;
  assign n12886 = n12885 ^ n12843 ;
  assign n13110 = n13109 ^ n12886 ;
  assign n13112 = n13110 ^ x11 ;
  assign n13111 = n13110 ^ n514 ;
  assign n13113 = n13112 ^ n13111 ;
  assign n13114 = n12883 & ~n13113 ;
  assign n13115 = n13114 ^ n13112 ;
  assign n13116 = n13115 ^ n13110 ;
  assign n13119 = ~x10 & x127 ;
  assign n13120 = n13119 ^ x11 ;
  assign n13121 = ~n10154 & ~n13120 ;
  assign n13122 = n13121 ^ x11 ;
  assign n13123 = n515 & ~n13122 ;
  assign n13124 = n13116 & n13123 ;
  assign n13125 = n13124 ^ n13115 ;
  assign n13129 = n13128 ^ n13125 ;
  assign n13133 = n13132 ^ n13129 ;
  assign n12879 = n12877 ^ n12860 ;
  assign n12880 = ~n12861 & ~n12879 ;
  assign n12881 = n12880 ^ n12877 ;
  assign n13134 = n13133 ^ n12881 ;
  assign n13375 = n13103 ^ n12886 ;
  assign n13376 = n13109 & ~n13375 ;
  assign n13377 = n13376 ^ n13103 ;
  assign n13373 = x126 & n795 ;
  assign n13366 = x123 & n1068 ;
  assign n13358 = n13086 ^ n12895 ;
  assign n13359 = n13092 & n13358 ;
  assign n13360 = n13359 ^ n13086 ;
  assign n13356 = x120 & n1348 ;
  assign n13349 = x117 & n1673 ;
  assign n13342 = x114 & n2025 ;
  assign n13335 = x111 & n2435 ;
  assign n13328 = x108 & n2899 ;
  assign n13317 = x104 & n3387 ;
  assign n13316 = x106 & n3390 ;
  assign n13318 = n13317 ^ n13316 ;
  assign n13319 = n13318 ^ x35 ;
  assign n13315 = n3391 & ~n5257 ;
  assign n13320 = n13319 ^ n13315 ;
  assign n13314 = x105 & n3395 ;
  assign n13321 = n13320 ^ n13314 ;
  assign n13308 = x101 & n3932 ;
  assign n13307 = x103 & n3935 ;
  assign n13309 = n13308 ^ n13307 ;
  assign n13310 = n13309 ^ x38 ;
  assign n13306 = n3936 & ~n4624 ;
  assign n13311 = n13310 ^ n13306 ;
  assign n13305 = x102 & n3940 ;
  assign n13312 = n13311 ^ n13305 ;
  assign n13296 = n13022 ^ n13009 ;
  assign n13297 = n13014 & ~n13296 ;
  assign n13298 = n13297 ^ n13009 ;
  assign n13290 = x98 & n4482 ;
  assign n13289 = x100 & n4478 ;
  assign n13291 = n13290 ^ n13289 ;
  assign n13292 = n13291 ^ x41 ;
  assign n13288 = n4048 & n4479 ;
  assign n13293 = n13292 ^ n13288 ;
  assign n13287 = x99 & n4475 ;
  assign n13294 = n13293 ^ n13287 ;
  assign n13283 = n12999 ^ n12916 ;
  assign n13284 = ~n13008 & ~n13283 ;
  assign n13285 = n13284 ^ n12999 ;
  assign n13277 = x95 & n5113 ;
  assign n13276 = x97 & n5116 ;
  assign n13278 = n13277 ^ n13276 ;
  assign n13279 = n13278 ^ x44 ;
  assign n13275 = n3501 & n5117 ;
  assign n13280 = n13279 ^ n13275 ;
  assign n13274 = x96 & n5121 ;
  assign n13281 = n13280 ^ n13274 ;
  assign n13266 = x89 & n6687 ;
  assign n13265 = x91 & n6444 ;
  assign n13267 = n13266 ^ n13265 ;
  assign n13268 = n13267 ^ x50 ;
  assign n13264 = n2548 & n6445 ;
  assign n13269 = n13268 ^ n13264 ;
  assign n13263 = x90 & n6449 ;
  assign n13270 = n13269 ^ n13263 ;
  assign n13259 = n12983 ^ n12932 ;
  assign n13260 = ~n12984 & n13259 ;
  assign n13261 = n13260 ^ n12983 ;
  assign n13253 = x86 & n7183 ;
  assign n13252 = x88 & n7186 ;
  assign n13254 = n13253 ^ n13252 ;
  assign n13255 = n13254 ^ x53 ;
  assign n13251 = n2131 & n7187 ;
  assign n13256 = n13255 ^ n13251 ;
  assign n13250 = x87 & n7191 ;
  assign n13257 = n13256 ^ n13250 ;
  assign n13247 = x84 & n7947 ;
  assign n13240 = x81 & n8743 ;
  assign n13229 = x77 & n9655 ;
  assign n13228 = x79 & n9651 ;
  assign n13230 = n13229 ^ n13228 ;
  assign n13231 = n13230 ^ x62 ;
  assign n13227 = n1123 & n9652 ;
  assign n13232 = n13231 ^ n13227 ;
  assign n13226 = x78 & n9648 ;
  assign n13233 = n13232 ^ n13226 ;
  assign n13221 = x63 & x75 ;
  assign n13222 = n13221 ^ x76 ;
  assign n13223 = ~n9956 & n13222 ;
  assign n13215 = n12708 ^ x76 ;
  assign n13224 = n13223 ^ n13215 ;
  assign n13225 = n13224 ^ x11 ;
  assign n13234 = n13233 ^ n13225 ;
  assign n13209 = ~x75 & n12706 ;
  assign n13208 = ~x74 & n12707 ;
  assign n13210 = n13209 ^ n13208 ;
  assign n13211 = ~n12935 & ~n13210 ;
  assign n13212 = n13208 ^ n12943 ;
  assign n13213 = n13211 & ~n13212 ;
  assign n13214 = n13213 ^ n13210 ;
  assign n13235 = n13234 ^ n13214 ;
  assign n13236 = n13235 ^ x59 ;
  assign n13207 = x80 & n8750 ;
  assign n13237 = n13236 ^ n13207 ;
  assign n13206 = x82 & n8746 ;
  assign n13238 = n13237 ^ n13206 ;
  assign n13205 = n1422 & n8747 ;
  assign n13239 = n13238 ^ n13205 ;
  assign n13241 = n13240 ^ n13239 ;
  assign n13202 = n12961 ^ n12952 ;
  assign n13203 = n12953 & n13202 ;
  assign n13204 = n13203 ^ n12961 ;
  assign n13242 = n13241 ^ n13204 ;
  assign n13243 = n13242 ^ x56 ;
  assign n13201 = x83 & n7954 ;
  assign n13244 = n13243 ^ n13201 ;
  assign n13200 = x85 & n7950 ;
  assign n13245 = n13244 ^ n13200 ;
  assign n13199 = n1748 & n7951 ;
  assign n13246 = n13245 ^ n13199 ;
  assign n13248 = n13247 ^ n13246 ;
  assign n13196 = n12974 ^ n12970 ;
  assign n13197 = n12971 & n13196 ;
  assign n13198 = n13197 ^ n12974 ;
  assign n13249 = n13248 ^ n13198 ;
  assign n13258 = n13257 ^ n13249 ;
  assign n13262 = n13261 ^ n13258 ;
  assign n13271 = n13270 ^ n13262 ;
  assign n13193 = n12985 ^ n12924 ;
  assign n13194 = n12929 & ~n13193 ;
  assign n13195 = n13194 ^ n12924 ;
  assign n13272 = n13271 ^ n13195 ;
  assign n13183 = x92 & n5981 ;
  assign n13182 = x94 & n5748 ;
  assign n13184 = n13183 ^ n13182 ;
  assign n13185 = n13184 ^ x47 ;
  assign n13181 = n3010 & n5749 ;
  assign n13186 = n13185 ^ n13181 ;
  assign n13180 = x93 & n5755 ;
  assign n13187 = n13186 ^ n13180 ;
  assign n13188 = n13187 ^ n12998 ;
  assign n13189 = n13188 ^ n12994 ;
  assign n13190 = n13189 ^ n13187 ;
  assign n13191 = n12995 & n13190 ;
  assign n13192 = n13191 ^ n13188 ;
  assign n13273 = n13272 ^ n13192 ;
  assign n13282 = n13281 ^ n13273 ;
  assign n13286 = n13285 ^ n13282 ;
  assign n13295 = n13294 ^ n13286 ;
  assign n13299 = n13298 ^ n13295 ;
  assign n13300 = n13299 ^ n13035 ;
  assign n13301 = n13300 ^ n13026 ;
  assign n13302 = n13301 ^ n13299 ;
  assign n13303 = n13027 & ~n13302 ;
  assign n13304 = n13303 ^ n13300 ;
  assign n13313 = n13312 ^ n13304 ;
  assign n13322 = n13321 ^ n13313 ;
  assign n13177 = n13048 ^ n13044 ;
  assign n13178 = n13045 & n13177 ;
  assign n13179 = n13178 ^ n13048 ;
  assign n13323 = n13322 ^ n13179 ;
  assign n13324 = n13323 ^ x32 ;
  assign n13176 = x107 & n2890 ;
  assign n13325 = n13324 ^ n13176 ;
  assign n13175 = x109 & n2893 ;
  assign n13326 = n13325 ^ n13175 ;
  assign n13174 = n2894 & n5912 ;
  assign n13327 = n13326 ^ n13174 ;
  assign n13329 = n13328 ^ n13327 ;
  assign n13171 = n13058 ^ n13049 ;
  assign n13172 = n13055 & n13171 ;
  assign n13173 = n13172 ^ n13058 ;
  assign n13330 = n13329 ^ n13173 ;
  assign n13331 = n13330 ^ x29 ;
  assign n13170 = x110 & n2593 ;
  assign n13332 = n13331 ^ n13170 ;
  assign n13169 = x112 & n2428 ;
  assign n13333 = n13332 ^ n13169 ;
  assign n13168 = n2429 & ~n6616 ;
  assign n13334 = n13333 ^ n13168 ;
  assign n13336 = n13335 ^ n13334 ;
  assign n13165 = n13068 ^ n13059 ;
  assign n13166 = ~n13065 & n13165 ;
  assign n13167 = n13166 ^ n13068 ;
  assign n13337 = n13336 ^ n13167 ;
  assign n13338 = n13337 ^ x26 ;
  assign n13164 = x113 & n2032 ;
  assign n13339 = n13338 ^ n13164 ;
  assign n13163 = x115 & n2028 ;
  assign n13340 = n13339 ^ n13163 ;
  assign n13162 = n2029 & ~n7353 ;
  assign n13341 = n13340 ^ n13162 ;
  assign n13343 = n13342 ^ n13341 ;
  assign n13159 = n13078 ^ n13069 ;
  assign n13160 = ~n13075 & ~n13159 ;
  assign n13161 = n13160 ^ n13078 ;
  assign n13344 = n13343 ^ n13161 ;
  assign n13345 = n13344 ^ x23 ;
  assign n13158 = x116 & n1665 ;
  assign n13346 = n13345 ^ n13158 ;
  assign n13157 = x118 & n1668 ;
  assign n13347 = n13346 ^ n13157 ;
  assign n13156 = n1669 & ~n8140 ;
  assign n13348 = n13347 ^ n13156 ;
  assign n13350 = n13349 ^ n13348 ;
  assign n13153 = n13079 ^ n12901 ;
  assign n13154 = ~n13085 & n13153 ;
  assign n13155 = n13154 ^ n13079 ;
  assign n13351 = n13350 ^ n13155 ;
  assign n13352 = n13351 ^ x20 ;
  assign n13152 = x119 & n1340 ;
  assign n13353 = n13352 ^ n13152 ;
  assign n13151 = x121 & n1343 ;
  assign n13354 = n13353 ^ n13151 ;
  assign n13150 = n1344 & n8979 ;
  assign n13355 = n13354 ^ n13150 ;
  assign n13357 = n13356 ^ n13355 ;
  assign n13361 = n13360 ^ n13357 ;
  assign n13362 = n13361 ^ x17 ;
  assign n13149 = x122 & n1060 ;
  assign n13363 = n13362 ^ n13149 ;
  assign n13148 = x124 & n1063 ;
  assign n13364 = n13363 ^ n13148 ;
  assign n13147 = n1064 & n10117 ;
  assign n13365 = n13364 ^ n13147 ;
  assign n13367 = n13366 ^ n13365 ;
  assign n13144 = n13102 ^ n13093 ;
  assign n13145 = ~n13099 & n13144 ;
  assign n13146 = n13145 ^ n13102 ;
  assign n13368 = n13367 ^ n13146 ;
  assign n13369 = n13368 ^ x14 ;
  assign n13143 = x125 & n884 ;
  assign n13370 = n13369 ^ n13143 ;
  assign n13142 = x127 & n789 ;
  assign n13371 = n13370 ^ n13142 ;
  assign n13141 = n790 & n10986 ;
  assign n13372 = n13371 ^ n13141 ;
  assign n13374 = n13373 ^ n13372 ;
  assign n13378 = n13377 ^ n13374 ;
  assign n13138 = n13128 ^ n13110 ;
  assign n13139 = n13125 & n13138 ;
  assign n13140 = n13139 ^ n13128 ;
  assign n13379 = n13378 ^ n13140 ;
  assign n13135 = n13132 ^ n12881 ;
  assign n13136 = n13133 & ~n13135 ;
  assign n13137 = n13136 ^ n13132 ;
  assign n13380 = n13379 ^ n13137 ;
  assign n13608 = n13361 ^ n13146 ;
  assign n13609 = ~n13367 & ~n13608 ;
  assign n13610 = n13609 ^ n13361 ;
  assign n13606 = x127 & n795 ;
  assign n13600 = x124 & n1068 ;
  assign n13593 = x121 & n1348 ;
  assign n13585 = n13337 ^ n13161 ;
  assign n13586 = ~n13343 & n13585 ;
  assign n13587 = n13586 ^ n13337 ;
  assign n13583 = x118 & n1673 ;
  assign n13575 = n13330 ^ n13167 ;
  assign n13576 = ~n13336 & ~n13575 ;
  assign n13577 = n13576 ^ n13330 ;
  assign n13573 = x115 & n2025 ;
  assign n13563 = x111 & n2593 ;
  assign n13562 = x113 & n2428 ;
  assign n13564 = n13563 ^ n13562 ;
  assign n13565 = n13564 ^ x29 ;
  assign n13561 = n2429 & ~n6849 ;
  assign n13566 = n13565 ^ n13561 ;
  assign n13560 = x112 & n2435 ;
  assign n13567 = n13566 ^ n13560 ;
  assign n13548 = x108 & n2890 ;
  assign n13547 = x110 & n2893 ;
  assign n13549 = n13548 ^ n13547 ;
  assign n13550 = n13549 ^ x32 ;
  assign n13546 = n2894 & n6145 ;
  assign n13551 = n13550 ^ n13546 ;
  assign n13545 = x109 & n2899 ;
  assign n13552 = n13551 ^ n13545 ;
  assign n13539 = x105 & n3387 ;
  assign n13538 = x107 & n3390 ;
  assign n13540 = n13539 ^ n13538 ;
  assign n13541 = n13540 ^ x35 ;
  assign n13537 = n3391 & ~n5459 ;
  assign n13542 = n13541 ^ n13537 ;
  assign n13536 = x106 & n3395 ;
  assign n13543 = n13542 ^ n13536 ;
  assign n13532 = n13312 ^ n13299 ;
  assign n13533 = n13304 & n13532 ;
  assign n13534 = n13533 ^ n13299 ;
  assign n13526 = x102 & n3932 ;
  assign n13525 = x104 & n3935 ;
  assign n13527 = n13526 ^ n13525 ;
  assign n13528 = n13527 ^ x38 ;
  assign n13524 = n3936 & ~n4830 ;
  assign n13529 = n13528 ^ n13524 ;
  assign n13523 = x103 & n3940 ;
  assign n13530 = n13529 ^ n13523 ;
  assign n13516 = x99 & n4482 ;
  assign n13515 = x101 & n4478 ;
  assign n13517 = n13516 ^ n13515 ;
  assign n13518 = n13517 ^ x41 ;
  assign n13514 = n4223 & n4479 ;
  assign n13519 = n13518 ^ n13514 ;
  assign n13513 = x100 & n4475 ;
  assign n13520 = n13519 ^ n13513 ;
  assign n13509 = x97 & n5121 ;
  assign n13507 = n3673 & n5117 ;
  assign n13503 = x96 & n5113 ;
  assign n13502 = x98 & n5116 ;
  assign n13504 = n13503 ^ n13502 ;
  assign n13505 = n13504 ^ x44 ;
  assign n13495 = x93 & n5981 ;
  assign n13494 = x95 & n5748 ;
  assign n13496 = n13495 ^ n13494 ;
  assign n13497 = n13496 ^ x47 ;
  assign n13493 = n3166 & n5749 ;
  assign n13498 = n13497 ^ n13493 ;
  assign n13492 = x94 & n5755 ;
  assign n13499 = n13498 ^ n13492 ;
  assign n13485 = x90 & n6687 ;
  assign n13484 = x92 & n6444 ;
  assign n13486 = n13485 ^ n13484 ;
  assign n13487 = n13486 ^ x50 ;
  assign n13483 = n2696 & n6445 ;
  assign n13488 = n13487 ^ n13483 ;
  assign n13482 = x91 & n6449 ;
  assign n13489 = n13488 ^ n13482 ;
  assign n13478 = n13242 ^ n13198 ;
  assign n13479 = n13248 & n13478 ;
  assign n13480 = n13479 ^ n13242 ;
  assign n13472 = x87 & n7183 ;
  assign n13471 = x89 & n7186 ;
  assign n13473 = n13472 ^ n13471 ;
  assign n13474 = n13473 ^ x53 ;
  assign n13470 = n2255 & n7187 ;
  assign n13475 = n13474 ^ n13470 ;
  assign n13469 = x88 & n7191 ;
  assign n13476 = n13475 ^ n13469 ;
  assign n13461 = x81 & n8750 ;
  assign n13460 = x83 & n8746 ;
  assign n13462 = n13461 ^ n13460 ;
  assign n13463 = n13462 ^ x59 ;
  assign n13459 = n1517 & n8747 ;
  assign n13464 = n13463 ^ n13459 ;
  assign n13458 = x82 & n8743 ;
  assign n13465 = n13464 ^ n13458 ;
  assign n13452 = x78 & n9655 ;
  assign n13451 = x80 & n9651 ;
  assign n13453 = n13452 ^ n13451 ;
  assign n13454 = n13453 ^ x62 ;
  assign n13450 = n1217 & n9652 ;
  assign n13455 = n13454 ^ n13450 ;
  assign n13449 = x79 & n9648 ;
  assign n13456 = n13455 ^ n13449 ;
  assign n13445 = n12708 ^ x11 ;
  assign n13446 = ~n13224 & ~n13445 ;
  assign n13447 = n13446 ^ x11 ;
  assign n13441 = x63 & x76 ;
  assign n13442 = n13441 ^ x77 ;
  assign n13443 = ~n9956 & n13442 ;
  assign n13444 = n13443 ^ x77 ;
  assign n13448 = n13447 ^ n13444 ;
  assign n13457 = n13456 ^ n13448 ;
  assign n13466 = n13465 ^ n13457 ;
  assign n13438 = n13233 ^ n13214 ;
  assign n13439 = ~n13234 & ~n13438 ;
  assign n13440 = n13439 ^ n13233 ;
  assign n13467 = n13466 ^ n13440 ;
  assign n13435 = n13235 ^ n13204 ;
  assign n13436 = n13241 & n13435 ;
  assign n13428 = x84 & n7954 ;
  assign n13427 = x86 & n7950 ;
  assign n13429 = n13428 ^ n13427 ;
  assign n13430 = n13429 ^ x56 ;
  assign n13426 = n1868 & n7951 ;
  assign n13431 = n13430 ^ n13426 ;
  assign n13425 = x85 & n7947 ;
  assign n13432 = n13431 ^ n13425 ;
  assign n13433 = n13432 ^ n13235 ;
  assign n13437 = n13436 ^ n13433 ;
  assign n13468 = n13467 ^ n13437 ;
  assign n13477 = n13476 ^ n13468 ;
  assign n13481 = n13480 ^ n13477 ;
  assign n13490 = n13489 ^ n13481 ;
  assign n13422 = n13261 ^ n13257 ;
  assign n13423 = ~n13258 & n13422 ;
  assign n13424 = n13423 ^ n13261 ;
  assign n13491 = n13490 ^ n13424 ;
  assign n13500 = n13499 ^ n13491 ;
  assign n13419 = n13270 ^ n13195 ;
  assign n13420 = n13271 & n13419 ;
  assign n13421 = n13420 ^ n13270 ;
  assign n13501 = n13500 ^ n13421 ;
  assign n13506 = n13505 ^ n13501 ;
  assign n13508 = n13507 ^ n13506 ;
  assign n13510 = n13509 ^ n13508 ;
  assign n13416 = n13272 ^ n13187 ;
  assign n13417 = n13192 & n13416 ;
  assign n13418 = n13417 ^ n13187 ;
  assign n13511 = n13510 ^ n13418 ;
  assign n13413 = n13285 ^ n13281 ;
  assign n13414 = ~n13282 & ~n13413 ;
  assign n13415 = n13414 ^ n13285 ;
  assign n13512 = n13511 ^ n13415 ;
  assign n13521 = n13520 ^ n13512 ;
  assign n13410 = n13298 ^ n13294 ;
  assign n13411 = n13295 & ~n13410 ;
  assign n13412 = n13411 ^ n13298 ;
  assign n13522 = n13521 ^ n13412 ;
  assign n13531 = n13530 ^ n13522 ;
  assign n13535 = n13534 ^ n13531 ;
  assign n13544 = n13543 ^ n13535 ;
  assign n13553 = n13552 ^ n13544 ;
  assign n13407 = n13321 ^ n13179 ;
  assign n13408 = n13322 & n13407 ;
  assign n13409 = n13408 ^ n13321 ;
  assign n13554 = n13553 ^ n13409 ;
  assign n13555 = n13554 ^ n13323 ;
  assign n13556 = n13555 ^ n13554 ;
  assign n13557 = n13556 ^ n13173 ;
  assign n13558 = n13329 & ~n13557 ;
  assign n13559 = n13558 ^ n13555 ;
  assign n13568 = n13567 ^ n13559 ;
  assign n13569 = n13568 ^ x26 ;
  assign n13406 = x114 & n2032 ;
  assign n13570 = n13569 ^ n13406 ;
  assign n13405 = x116 & n2028 ;
  assign n13571 = n13570 ^ n13405 ;
  assign n13404 = n2029 & ~n7604 ;
  assign n13572 = n13571 ^ n13404 ;
  assign n13574 = n13573 ^ n13572 ;
  assign n13578 = n13577 ^ n13574 ;
  assign n13579 = n13578 ^ x23 ;
  assign n13403 = x117 & n1665 ;
  assign n13580 = n13579 ^ n13403 ;
  assign n13402 = x119 & n1668 ;
  assign n13581 = n13580 ^ n13402 ;
  assign n13401 = n1669 & n8405 ;
  assign n13582 = n13581 ^ n13401 ;
  assign n13584 = n13583 ^ n13582 ;
  assign n13588 = n13587 ^ n13584 ;
  assign n13589 = n13588 ^ x20 ;
  assign n13400 = x120 & n1340 ;
  assign n13590 = n13589 ^ n13400 ;
  assign n13399 = x122 & n1343 ;
  assign n13591 = n13590 ^ n13399 ;
  assign n13398 = n1344 & ~n9261 ;
  assign n13592 = n13591 ^ n13398 ;
  assign n13594 = n13593 ^ n13592 ;
  assign n13395 = n13344 ^ n13155 ;
  assign n13396 = n13350 & ~n13395 ;
  assign n13397 = n13396 ^ n13344 ;
  assign n13595 = n13594 ^ n13397 ;
  assign n13596 = n13595 ^ x17 ;
  assign n13394 = x123 & n1060 ;
  assign n13597 = n13596 ^ n13394 ;
  assign n13393 = x125 & n1063 ;
  assign n13598 = n13597 ^ n13393 ;
  assign n13392 = n1064 & n10416 ;
  assign n13599 = n13598 ^ n13392 ;
  assign n13601 = n13600 ^ n13599 ;
  assign n13389 = n13360 ^ n13351 ;
  assign n13390 = n13357 & ~n13389 ;
  assign n13391 = n13390 ^ n13360 ;
  assign n13602 = n13601 ^ n13391 ;
  assign n13603 = n13602 ^ x14 ;
  assign n13388 = x126 & n884 ;
  assign n13604 = n13603 ^ n13388 ;
  assign n13387 = n790 & n10155 ;
  assign n13605 = n13604 ^ n13387 ;
  assign n13607 = n13606 ^ n13605 ;
  assign n13611 = n13610 ^ n13607 ;
  assign n13384 = n13377 ^ n13368 ;
  assign n13385 = n13374 & ~n13384 ;
  assign n13386 = n13385 ^ n13377 ;
  assign n13612 = n13611 ^ n13386 ;
  assign n13381 = n13140 ^ n13137 ;
  assign n13382 = ~n13379 & ~n13381 ;
  assign n13383 = n13382 ^ n13137 ;
  assign n13613 = n13612 ^ n13383 ;
  assign n13848 = n13595 ^ n13391 ;
  assign n13849 = n13601 & n13848 ;
  assign n13850 = n13849 ^ n13595 ;
  assign n13841 = x124 & n1060 ;
  assign n13840 = x126 & n1063 ;
  assign n13842 = n13841 ^ n13840 ;
  assign n13843 = n13842 ^ x17 ;
  assign n13839 = n1064 & n10461 ;
  assign n13844 = n13843 ^ n13839 ;
  assign n13838 = x125 & n1068 ;
  assign n13845 = n13844 ^ n13838 ;
  assign n13831 = x121 & n1340 ;
  assign n13830 = x123 & n1343 ;
  assign n13832 = n13831 ^ n13830 ;
  assign n13833 = n13832 ^ x20 ;
  assign n13829 = n1344 & ~n9804 ;
  assign n13834 = n13833 ^ n13829 ;
  assign n13828 = x122 & n1348 ;
  assign n13835 = n13834 ^ n13828 ;
  assign n13824 = x119 & n1673 ;
  assign n13814 = x115 & n2032 ;
  assign n13813 = x117 & n2028 ;
  assign n13815 = n13814 ^ n13813 ;
  assign n13816 = n13815 ^ x26 ;
  assign n13812 = n2029 & ~n7860 ;
  assign n13817 = n13816 ^ n13812 ;
  assign n13811 = x116 & n2025 ;
  assign n13818 = n13817 ^ n13811 ;
  assign n13800 = x112 & n2593 ;
  assign n13799 = x114 & n2428 ;
  assign n13801 = n13800 ^ n13799 ;
  assign n13802 = n13801 ^ x29 ;
  assign n13798 = n2429 & ~n7108 ;
  assign n13803 = n13802 ^ n13798 ;
  assign n13797 = x113 & n2435 ;
  assign n13804 = n13803 ^ n13797 ;
  assign n13786 = x109 & n2890 ;
  assign n13785 = x111 & n2893 ;
  assign n13787 = n13786 ^ n13785 ;
  assign n13788 = n13787 ^ x32 ;
  assign n13784 = n2894 & ~n6370 ;
  assign n13789 = n13788 ^ n13784 ;
  assign n13783 = x110 & n2899 ;
  assign n13790 = n13789 ^ n13783 ;
  assign n13776 = x106 & n3387 ;
  assign n13775 = x108 & n3390 ;
  assign n13777 = n13776 ^ n13775 ;
  assign n13778 = n13777 ^ x35 ;
  assign n13774 = n3391 & n5687 ;
  assign n13779 = n13778 ^ n13774 ;
  assign n13773 = x107 & n3395 ;
  assign n13780 = n13779 ^ n13773 ;
  assign n13762 = x103 & n3932 ;
  assign n13761 = x105 & n3935 ;
  assign n13763 = n13762 ^ n13761 ;
  assign n13764 = n13763 ^ x38 ;
  assign n13760 = n3936 & ~n5034 ;
  assign n13765 = n13764 ^ n13760 ;
  assign n13759 = x104 & n3940 ;
  assign n13766 = n13765 ^ n13759 ;
  assign n13756 = n13520 ^ n13415 ;
  assign n13757 = n13512 & ~n13756 ;
  assign n13748 = x100 & n4482 ;
  assign n13747 = x102 & n4478 ;
  assign n13749 = n13748 ^ n13747 ;
  assign n13750 = n13749 ^ x41 ;
  assign n13746 = n4425 & n4479 ;
  assign n13751 = n13750 ^ n13746 ;
  assign n13745 = x101 & n4475 ;
  assign n13752 = n13751 ^ n13745 ;
  assign n13737 = x98 & n5121 ;
  assign n13735 = n3851 & n5117 ;
  assign n13731 = x97 & n5113 ;
  assign n13730 = x99 & n5116 ;
  assign n13732 = n13731 ^ n13730 ;
  assign n13733 = n13732 ^ x44 ;
  assign n13727 = x95 & n5755 ;
  assign n13725 = n3336 & n5749 ;
  assign n13721 = x94 & n5981 ;
  assign n13720 = x96 & n5748 ;
  assign n13722 = n13721 ^ n13720 ;
  assign n13723 = n13722 ^ x47 ;
  assign n13713 = x91 & n6687 ;
  assign n13712 = x93 & n6444 ;
  assign n13714 = n13713 ^ n13712 ;
  assign n13715 = n13714 ^ x50 ;
  assign n13711 = n2842 & n6445 ;
  assign n13716 = n13715 ^ n13711 ;
  assign n13710 = x92 & n6449 ;
  assign n13717 = n13716 ^ n13710 ;
  assign n13706 = x86 & n7947 ;
  assign n13704 = n1987 & n7951 ;
  assign n13700 = x85 & n7954 ;
  assign n13699 = x87 & n7950 ;
  assign n13701 = n13700 ^ n13699 ;
  assign n13702 = n13701 ^ x56 ;
  assign n13692 = n1310 & n9652 ;
  assign n13691 = x80 & n9648 ;
  assign n13693 = n13692 ^ n13691 ;
  assign n13689 = x79 & n9655 ;
  assign n13688 = x81 & n9651 ;
  assign n13690 = n13689 ^ n13688 ;
  assign n13694 = n13693 ^ n13690 ;
  assign n13687 = n844 ^ x62 ;
  assign n13695 = n13694 ^ n13687 ;
  assign n13684 = n13456 ^ n13447 ;
  assign n13685 = ~n13448 & ~n13684 ;
  assign n13686 = n13685 ^ n13456 ;
  assign n13696 = n13695 ^ n13686 ;
  assign n13681 = x63 & x78 ;
  assign n13679 = x63 & n844 ;
  assign n13678 = n13442 ^ x78 ;
  assign n13680 = n13679 ^ n13678 ;
  assign n13682 = n13681 ^ n13680 ;
  assign n13683 = ~n9956 & n13682 ;
  assign n13697 = n13696 ^ n13683 ;
  assign n13673 = x82 & n8750 ;
  assign n13672 = x84 & n8746 ;
  assign n13674 = n13673 ^ n13672 ;
  assign n13675 = n13674 ^ x59 ;
  assign n13671 = n1635 & n8747 ;
  assign n13676 = n13675 ^ n13671 ;
  assign n13670 = x83 & n8743 ;
  assign n13677 = n13676 ^ n13670 ;
  assign n13698 = n13697 ^ n13677 ;
  assign n13703 = n13702 ^ n13698 ;
  assign n13705 = n13704 ^ n13703 ;
  assign n13707 = n13706 ^ n13705 ;
  assign n13667 = n13465 ^ n13440 ;
  assign n13668 = n13466 & n13667 ;
  assign n13669 = n13668 ^ n13465 ;
  assign n13708 = n13707 ^ n13669 ;
  assign n13657 = x88 & n7183 ;
  assign n13656 = x90 & n7186 ;
  assign n13658 = n13657 ^ n13656 ;
  assign n13659 = n13658 ^ x53 ;
  assign n13655 = n2398 & n7187 ;
  assign n13660 = n13659 ^ n13655 ;
  assign n13654 = x89 & n7191 ;
  assign n13661 = n13660 ^ n13654 ;
  assign n13663 = n13661 ^ n13432 ;
  assign n13662 = n13661 ^ n13467 ;
  assign n13664 = n13663 ^ n13662 ;
  assign n13665 = n13437 & n13664 ;
  assign n13666 = n13665 ^ n13663 ;
  assign n13709 = n13708 ^ n13666 ;
  assign n13718 = n13717 ^ n13709 ;
  assign n13651 = n13480 ^ n13476 ;
  assign n13652 = ~n13477 & n13651 ;
  assign n13653 = n13652 ^ n13480 ;
  assign n13719 = n13718 ^ n13653 ;
  assign n13724 = n13723 ^ n13719 ;
  assign n13726 = n13725 ^ n13724 ;
  assign n13728 = n13727 ^ n13726 ;
  assign n13648 = n13489 ^ n13424 ;
  assign n13649 = n13490 & n13648 ;
  assign n13650 = n13649 ^ n13489 ;
  assign n13729 = n13728 ^ n13650 ;
  assign n13734 = n13733 ^ n13729 ;
  assign n13736 = n13735 ^ n13734 ;
  assign n13738 = n13737 ^ n13736 ;
  assign n13645 = n13499 ^ n13421 ;
  assign n13646 = n13500 & n13645 ;
  assign n13647 = n13646 ^ n13499 ;
  assign n13739 = n13738 ^ n13647 ;
  assign n13740 = n13739 ^ n13501 ;
  assign n13741 = n13740 ^ n13418 ;
  assign n13742 = n13741 ^ n13739 ;
  assign n13743 = n13510 & n13742 ;
  assign n13744 = n13743 ^ n13740 ;
  assign n13753 = n13752 ^ n13744 ;
  assign n13754 = n13753 ^ n13520 ;
  assign n13758 = n13757 ^ n13754 ;
  assign n13767 = n13766 ^ n13758 ;
  assign n13768 = n13767 ^ n13530 ;
  assign n13769 = n13768 ^ n13767 ;
  assign n13770 = n13769 ^ n13412 ;
  assign n13771 = ~n13522 & ~n13770 ;
  assign n13772 = n13771 ^ n13768 ;
  assign n13781 = n13780 ^ n13772 ;
  assign n13642 = n13543 ^ n13534 ;
  assign n13643 = ~n13535 & n13642 ;
  assign n13644 = n13643 ^ n13543 ;
  assign n13782 = n13781 ^ n13644 ;
  assign n13791 = n13790 ^ n13782 ;
  assign n13792 = n13791 ^ n13552 ;
  assign n13793 = n13792 ^ n13791 ;
  assign n13794 = n13793 ^ n13409 ;
  assign n13795 = n13553 & n13794 ;
  assign n13796 = n13795 ^ n13792 ;
  assign n13805 = n13804 ^ n13796 ;
  assign n13807 = n13805 ^ n13554 ;
  assign n13806 = n13805 ^ n13567 ;
  assign n13808 = n13807 ^ n13806 ;
  assign n13809 = n13559 & n13808 ;
  assign n13810 = n13809 ^ n13807 ;
  assign n13819 = n13818 ^ n13810 ;
  assign n13820 = n13819 ^ x23 ;
  assign n13641 = x118 & n1665 ;
  assign n13821 = n13820 ^ n13641 ;
  assign n13640 = x120 & n1668 ;
  assign n13822 = n13821 ^ n13640 ;
  assign n13639 = n1669 & n8904 ;
  assign n13823 = n13822 ^ n13639 ;
  assign n13825 = n13824 ^ n13823 ;
  assign n13636 = n13577 ^ n13568 ;
  assign n13637 = ~n13574 & ~n13636 ;
  assign n13638 = n13637 ^ n13577 ;
  assign n13826 = n13825 ^ n13638 ;
  assign n13633 = n13587 ^ n13578 ;
  assign n13634 = n13584 & n13633 ;
  assign n13635 = n13634 ^ n13587 ;
  assign n13827 = n13826 ^ n13635 ;
  assign n13836 = n13835 ^ n13827 ;
  assign n13630 = n13588 ^ n13397 ;
  assign n13631 = n13594 & n13630 ;
  assign n13632 = n13631 ^ n13588 ;
  assign n13837 = n13836 ^ n13632 ;
  assign n13846 = n13845 ^ n13837 ;
  assign n13620 = x127 & n883 ;
  assign n13621 = n13620 ^ n788 ;
  assign n13626 = n644 & n11285 ;
  assign n13627 = n13626 ^ n13620 ;
  assign n13628 = n13621 & ~n13627 ;
  assign n13629 = n13628 ^ x13 ;
  assign n13847 = n13846 ^ n13629 ;
  assign n13851 = n13850 ^ n13847 ;
  assign n13617 = n13610 ^ n13602 ;
  assign n13618 = ~n13607 & ~n13617 ;
  assign n13619 = n13618 ^ n13610 ;
  assign n13852 = n13851 ^ n13619 ;
  assign n13614 = n13386 ^ n13383 ;
  assign n13615 = n13612 & n13614 ;
  assign n13616 = n13615 ^ n13383 ;
  assign n13853 = n13852 ^ n13616 ;
  assign n14082 = x126 & n1068 ;
  assign n14075 = x123 & n1348 ;
  assign n14067 = n13819 ^ n13638 ;
  assign n14068 = ~n13825 & n14067 ;
  assign n14069 = n14068 ^ n13819 ;
  assign n14065 = x120 & n1673 ;
  assign n14057 = n13818 ^ n13805 ;
  assign n14058 = ~n13810 & ~n14057 ;
  assign n14059 = n14058 ^ n13805 ;
  assign n14051 = x116 & n2032 ;
  assign n14050 = x118 & n2028 ;
  assign n14052 = n14051 ^ n14050 ;
  assign n14053 = n14052 ^ x26 ;
  assign n14049 = n2029 & ~n8140 ;
  assign n14054 = n14053 ^ n14049 ;
  assign n14048 = x117 & n2025 ;
  assign n14055 = n14054 ^ n14048 ;
  assign n14044 = n13804 ^ n13791 ;
  assign n14045 = ~n13796 & ~n14044 ;
  assign n14046 = n14045 ^ n13791 ;
  assign n14038 = x113 & n2593 ;
  assign n14037 = x115 & n2428 ;
  assign n14039 = n14038 ^ n14037 ;
  assign n14040 = n14039 ^ x29 ;
  assign n14036 = n2429 & ~n7353 ;
  assign n14041 = n14040 ^ n14036 ;
  assign n14035 = x114 & n2435 ;
  assign n14042 = n14041 ^ n14035 ;
  assign n14028 = x110 & n2890 ;
  assign n14027 = x112 & n2893 ;
  assign n14029 = n14028 ^ n14027 ;
  assign n14030 = n14029 ^ x32 ;
  assign n14026 = n2894 & ~n6616 ;
  assign n14031 = n14030 ^ n14026 ;
  assign n14025 = x111 & n2899 ;
  assign n14032 = n14031 ^ n14025 ;
  assign n14021 = n13780 ^ n13767 ;
  assign n14022 = ~n13772 & ~n14021 ;
  assign n14023 = n14022 ^ n13767 ;
  assign n14015 = x107 & n3387 ;
  assign n14014 = x109 & n3390 ;
  assign n14016 = n14015 ^ n14014 ;
  assign n14017 = n14016 ^ x35 ;
  assign n14013 = n3391 & n5912 ;
  assign n14018 = n14017 ^ n14013 ;
  assign n14012 = x108 & n3395 ;
  assign n14019 = n14018 ^ n14012 ;
  assign n14008 = n13766 ^ n13753 ;
  assign n14009 = ~n13758 & ~n14008 ;
  assign n14010 = n14009 ^ n13753 ;
  assign n14002 = x104 & n3932 ;
  assign n14001 = x106 & n3935 ;
  assign n14003 = n14002 ^ n14001 ;
  assign n14004 = n14003 ^ x38 ;
  assign n14000 = n3936 & ~n5257 ;
  assign n14005 = n14004 ^ n14000 ;
  assign n13999 = x105 & n3940 ;
  assign n14006 = n14005 ^ n13999 ;
  assign n13996 = x102 & n4475 ;
  assign n13994 = n4479 & ~n4624 ;
  assign n13990 = x101 & n4482 ;
  assign n13989 = x103 & n4478 ;
  assign n13991 = n13990 ^ n13989 ;
  assign n13992 = n13991 ^ x41 ;
  assign n13985 = n13729 ^ n13647 ;
  assign n13986 = ~n13738 & ~n13985 ;
  assign n13987 = n13986 ^ n13729 ;
  assign n13979 = x98 & n5113 ;
  assign n13978 = x100 & n5116 ;
  assign n13980 = n13979 ^ n13978 ;
  assign n13981 = n13980 ^ x44 ;
  assign n13977 = n4048 & n5117 ;
  assign n13982 = n13981 ^ n13977 ;
  assign n13976 = x99 & n5121 ;
  assign n13983 = n13982 ^ n13976 ;
  assign n13972 = n13719 ^ n13650 ;
  assign n13973 = ~n13728 & ~n13972 ;
  assign n13974 = n13973 ^ n13719 ;
  assign n13966 = x95 & n5981 ;
  assign n13965 = x97 & n5748 ;
  assign n13967 = n13966 ^ n13965 ;
  assign n13968 = n13967 ^ x47 ;
  assign n13964 = n3501 & n5749 ;
  assign n13969 = n13968 ^ n13964 ;
  assign n13963 = x96 & n5755 ;
  assign n13970 = n13969 ^ n13963 ;
  assign n13956 = x92 & n6687 ;
  assign n13955 = x94 & n6444 ;
  assign n13957 = n13956 ^ n13955 ;
  assign n13958 = n13957 ^ x50 ;
  assign n13954 = n3010 & n6445 ;
  assign n13959 = n13958 ^ n13954 ;
  assign n13953 = x93 & n6449 ;
  assign n13960 = n13959 ^ n13953 ;
  assign n13946 = x89 & n7183 ;
  assign n13945 = x91 & n7186 ;
  assign n13947 = n13946 ^ n13945 ;
  assign n13948 = n13947 ^ x53 ;
  assign n13944 = n2548 & n7187 ;
  assign n13949 = n13948 ^ n13944 ;
  assign n13943 = x90 & n7191 ;
  assign n13950 = n13949 ^ n13943 ;
  assign n13939 = n13698 ^ n13669 ;
  assign n13940 = ~n13707 & ~n13939 ;
  assign n13941 = n13940 ^ n13698 ;
  assign n13933 = x86 & n7954 ;
  assign n13932 = x88 & n7950 ;
  assign n13934 = n13933 ^ n13932 ;
  assign n13935 = n13934 ^ x56 ;
  assign n13931 = n2131 & n7951 ;
  assign n13936 = n13935 ^ n13931 ;
  assign n13930 = x87 & n7947 ;
  assign n13937 = n13936 ^ n13930 ;
  assign n13923 = x83 & n8750 ;
  assign n13922 = x85 & n8746 ;
  assign n13924 = n13923 ^ n13922 ;
  assign n13925 = n13924 ^ x59 ;
  assign n13921 = n1748 & n8747 ;
  assign n13926 = n13925 ^ n13921 ;
  assign n13920 = x84 & n8743 ;
  assign n13927 = n13926 ^ n13920 ;
  assign n13913 = x80 & n9655 ;
  assign n13912 = x82 & n9651 ;
  assign n13914 = n13913 ^ n13912 ;
  assign n13915 = n13914 ^ x62 ;
  assign n13911 = n1422 & n9652 ;
  assign n13916 = n13915 ^ n13911 ;
  assign n13910 = x81 & n9648 ;
  assign n13917 = n13916 ^ n13910 ;
  assign n13905 = n13681 ^ x79 ;
  assign n13906 = ~n9956 & n13905 ;
  assign n13907 = n13906 ^ x79 ;
  assign n13908 = n13907 ^ x14 ;
  assign n13909 = n13908 ^ n13444 ;
  assign n13918 = n13917 ^ n13909 ;
  assign n13889 = n13694 ^ x78 ;
  assign n13899 = ~n13679 & n13889 ;
  assign n13900 = n13899 ^ x78 ;
  assign n760 = x77 ^ x76 ;
  assign n13895 = n13694 ^ x76 ;
  assign n13896 = ~n760 & n13895 ;
  assign n13897 = n13896 ^ x76 ;
  assign n13898 = x63 & n13897 ;
  assign n13901 = n13900 ^ n13898 ;
  assign n13902 = x62 & ~n13901 ;
  assign n13903 = n13902 ^ n13900 ;
  assign n13892 = ~n844 & ~n13889 ;
  assign n13893 = n13892 ^ x78 ;
  assign n13894 = n11894 & ~n13893 ;
  assign n13904 = n13903 ^ n13894 ;
  assign n13919 = n13918 ^ n13904 ;
  assign n13928 = n13927 ^ n13919 ;
  assign n13886 = n13686 ^ n13677 ;
  assign n13887 = n13697 & n13886 ;
  assign n13888 = n13887 ^ n13677 ;
  assign n13929 = n13928 ^ n13888 ;
  assign n13938 = n13937 ^ n13929 ;
  assign n13942 = n13941 ^ n13938 ;
  assign n13951 = n13950 ^ n13942 ;
  assign n13883 = n13708 ^ n13661 ;
  assign n13884 = n13666 & ~n13883 ;
  assign n13885 = n13884 ^ n13661 ;
  assign n13952 = n13951 ^ n13885 ;
  assign n13961 = n13960 ^ n13952 ;
  assign n13880 = n13709 ^ n13653 ;
  assign n13881 = ~n13718 & n13880 ;
  assign n13882 = n13881 ^ n13717 ;
  assign n13962 = n13961 ^ n13882 ;
  assign n13971 = n13970 ^ n13962 ;
  assign n13975 = n13974 ^ n13971 ;
  assign n13984 = n13983 ^ n13975 ;
  assign n13988 = n13987 ^ n13984 ;
  assign n13993 = n13992 ^ n13988 ;
  assign n13995 = n13994 ^ n13993 ;
  assign n13997 = n13996 ^ n13995 ;
  assign n13877 = n13752 ^ n13739 ;
  assign n13878 = ~n13744 & ~n13877 ;
  assign n13879 = n13878 ^ n13739 ;
  assign n13998 = n13997 ^ n13879 ;
  assign n14007 = n14006 ^ n13998 ;
  assign n14011 = n14010 ^ n14007 ;
  assign n14020 = n14019 ^ n14011 ;
  assign n14024 = n14023 ^ n14020 ;
  assign n14033 = n14032 ^ n14024 ;
  assign n13874 = n13790 ^ n13644 ;
  assign n13875 = n13782 & n13874 ;
  assign n13876 = n13875 ^ n13790 ;
  assign n14034 = n14033 ^ n13876 ;
  assign n14043 = n14042 ^ n14034 ;
  assign n14047 = n14046 ^ n14043 ;
  assign n14056 = n14055 ^ n14047 ;
  assign n14060 = n14059 ^ n14056 ;
  assign n14061 = n14060 ^ x23 ;
  assign n13873 = x119 & n1665 ;
  assign n14062 = n14061 ^ n13873 ;
  assign n13872 = x121 & n1668 ;
  assign n14063 = n14062 ^ n13872 ;
  assign n13871 = n1669 & n8979 ;
  assign n14064 = n14063 ^ n13871 ;
  assign n14066 = n14065 ^ n14064 ;
  assign n14070 = n14069 ^ n14066 ;
  assign n14071 = n14070 ^ x20 ;
  assign n13870 = x122 & n1340 ;
  assign n14072 = n14071 ^ n13870 ;
  assign n13869 = x124 & n1343 ;
  assign n14073 = n14072 ^ n13869 ;
  assign n13868 = n1344 & n10117 ;
  assign n14074 = n14073 ^ n13868 ;
  assign n14076 = n14075 ^ n14074 ;
  assign n13865 = n13835 ^ n13635 ;
  assign n13866 = n13827 & ~n13865 ;
  assign n13867 = n13866 ^ n13835 ;
  assign n14077 = n14076 ^ n13867 ;
  assign n14078 = n14077 ^ x17 ;
  assign n13864 = x125 & n1060 ;
  assign n14079 = n14078 ^ n13864 ;
  assign n13863 = x127 & n1063 ;
  assign n14080 = n14079 ^ n13863 ;
  assign n13862 = n1064 & n10986 ;
  assign n14081 = n14080 ^ n13862 ;
  assign n14083 = n14082 ^ n14081 ;
  assign n13859 = n13845 ^ n13632 ;
  assign n13860 = n13837 & n13859 ;
  assign n13861 = n13860 ^ n13845 ;
  assign n14084 = n14083 ^ n13861 ;
  assign n13858 = ~n13629 & n13846 ;
  assign n14085 = n14084 ^ n13858 ;
  assign n13857 = ~n13619 & n13850 ;
  assign n14086 = n14085 ^ n13857 ;
  assign n13854 = n13850 ^ n13619 ;
  assign n13855 = n13854 ^ n13616 ;
  assign n13856 = n13852 & n13855 ;
  assign n14087 = n14086 ^ n13856 ;
  assign n14308 = n13858 ^ n13847 ;
  assign n14309 = n14084 ^ n13857 ;
  assign n14310 = n14309 ^ n13854 ;
  assign n14311 = ~n14308 & ~n14310 ;
  assign n14312 = n14085 ^ n14084 ;
  assign n14313 = n14309 ^ n14084 ;
  assign n14314 = ~n14312 & n14313 ;
  assign n14315 = n14314 ^ n14084 ;
  assign n14316 = n13616 & n14315 ;
  assign n14317 = n14311 & ~n14316 ;
  assign n14318 = n13850 ^ n13616 ;
  assign n14319 = n13619 ^ n13616 ;
  assign n14320 = n14318 & n14319 ;
  assign n14321 = n14320 ^ n13850 ;
  assign n14322 = ~n13858 & n14084 ;
  assign n14323 = ~n14321 & n14322 ;
  assign n14324 = n14323 ^ n14321 ;
  assign n14325 = ~n14317 & n14324 ;
  assign n14302 = n1064 & n10155 ;
  assign n14301 = x126 & n1060 ;
  assign n14303 = n14302 ^ n14301 ;
  assign n14304 = n14303 ^ x17 ;
  assign n14300 = x127 & n1068 ;
  assign n14305 = n14304 ^ n14300 ;
  assign n14296 = n14070 ^ n13867 ;
  assign n14297 = n14076 & n14296 ;
  assign n14298 = n14297 ^ n14070 ;
  assign n14290 = x123 & n1340 ;
  assign n14289 = x125 & n1343 ;
  assign n14291 = n14290 ^ n14289 ;
  assign n14292 = n14291 ^ x20 ;
  assign n14288 = n1344 & n10416 ;
  assign n14293 = n14292 ^ n14288 ;
  assign n14287 = x124 & n1348 ;
  assign n14294 = n14293 ^ n14287 ;
  assign n14280 = x120 & n1665 ;
  assign n14279 = x122 & n1668 ;
  assign n14281 = n14280 ^ n14279 ;
  assign n14282 = n14281 ^ x23 ;
  assign n14278 = n1669 & ~n9261 ;
  assign n14283 = n14282 ^ n14278 ;
  assign n14277 = x121 & n1673 ;
  assign n14284 = n14283 ^ n14277 ;
  assign n14269 = x117 & n2032 ;
  assign n14268 = x119 & n2028 ;
  assign n14270 = n14269 ^ n14268 ;
  assign n14271 = n14270 ^ x26 ;
  assign n14267 = n2029 & n8405 ;
  assign n14272 = n14271 ^ n14267 ;
  assign n14266 = x118 & n2025 ;
  assign n14273 = n14272 ^ n14266 ;
  assign n14260 = x114 & n2593 ;
  assign n14259 = x116 & n2428 ;
  assign n14261 = n14260 ^ n14259 ;
  assign n14262 = n14261 ^ x29 ;
  assign n14258 = n2429 & ~n7604 ;
  assign n14263 = n14262 ^ n14258 ;
  assign n14257 = x115 & n2435 ;
  assign n14264 = n14263 ^ n14257 ;
  assign n14253 = n14032 ^ n13876 ;
  assign n14254 = ~n14033 & n14253 ;
  assign n14255 = n14254 ^ n14032 ;
  assign n14247 = x111 & n2890 ;
  assign n14246 = x113 & n2893 ;
  assign n14248 = n14247 ^ n14246 ;
  assign n14249 = n14248 ^ x32 ;
  assign n14245 = n2894 & ~n6849 ;
  assign n14250 = n14249 ^ n14245 ;
  assign n14244 = x112 & n2899 ;
  assign n14251 = n14250 ^ n14244 ;
  assign n14232 = x105 & n3932 ;
  assign n14231 = x107 & n3935 ;
  assign n14233 = n14232 ^ n14231 ;
  assign n14234 = n14233 ^ x38 ;
  assign n14230 = n3936 & ~n5459 ;
  assign n14235 = n14234 ^ n14230 ;
  assign n14229 = x106 & n3940 ;
  assign n14236 = n14235 ^ n14229 ;
  assign n14225 = n13988 ^ n13879 ;
  assign n14226 = n13997 & ~n14225 ;
  assign n14227 = n14226 ^ n13988 ;
  assign n14219 = x102 & n4482 ;
  assign n14218 = x104 & n4478 ;
  assign n14220 = n14219 ^ n14218 ;
  assign n14221 = n14220 ^ x41 ;
  assign n14217 = n4479 & ~n4830 ;
  assign n14222 = n14221 ^ n14217 ;
  assign n14216 = x103 & n4475 ;
  assign n14223 = n14222 ^ n14216 ;
  assign n14212 = x100 & n5121 ;
  assign n14210 = n4223 & n5117 ;
  assign n14206 = x99 & n5113 ;
  assign n14205 = x101 & n5116 ;
  assign n14207 = n14206 ^ n14205 ;
  assign n14208 = n14207 ^ x44 ;
  assign n14202 = n13974 ^ n13970 ;
  assign n14203 = ~n13971 & ~n14202 ;
  assign n14204 = n14203 ^ n13974 ;
  assign n14209 = n14208 ^ n14204 ;
  assign n14211 = n14210 ^ n14209 ;
  assign n14213 = n14212 ^ n14211 ;
  assign n14198 = n13960 ^ n13882 ;
  assign n14199 = n13961 & n14198 ;
  assign n14200 = n14199 ^ n13960 ;
  assign n14192 = x96 & n5981 ;
  assign n14191 = x98 & n5748 ;
  assign n14193 = n14192 ^ n14191 ;
  assign n14194 = n14193 ^ x47 ;
  assign n14190 = n3673 & n5749 ;
  assign n14195 = n14194 ^ n14190 ;
  assign n14189 = x97 & n5755 ;
  assign n14196 = n14195 ^ n14189 ;
  assign n14182 = x93 & n6687 ;
  assign n14181 = x95 & n6444 ;
  assign n14183 = n14182 ^ n14181 ;
  assign n14184 = n14183 ^ x50 ;
  assign n14180 = n3166 & n6445 ;
  assign n14185 = n14184 ^ n14180 ;
  assign n14179 = x94 & n6449 ;
  assign n14186 = n14185 ^ n14179 ;
  assign n14173 = n13917 ^ n13904 ;
  assign n14174 = ~n13918 & n14173 ;
  assign n14175 = n14174 ^ n13917 ;
  assign n14167 = ~x63 & n1017 ;
  assign n14168 = n14167 ^ x79 ;
  assign n14144 = x63 & x80 ;
  assign n14170 = n14168 ^ n14144 ;
  assign n14171 = x62 & ~n14170 ;
  assign n14163 = n1517 & n9652 ;
  assign n14162 = x82 & n9648 ;
  assign n14164 = n14163 ^ n14162 ;
  assign n14160 = x81 & n9655 ;
  assign n14159 = x83 & n9651 ;
  assign n14161 = n14160 ^ n14159 ;
  assign n14165 = n14164 ^ n14161 ;
  assign n14153 = x84 & n8750 ;
  assign n14152 = x86 & n8746 ;
  assign n14154 = n14153 ^ n14152 ;
  assign n14155 = n14154 ^ x59 ;
  assign n14151 = n1868 & n8747 ;
  assign n14156 = n14155 ^ n14151 ;
  assign n14150 = x85 & n8743 ;
  assign n14157 = n14156 ^ n14150 ;
  assign n14145 = n13444 ^ x14 ;
  assign n14146 = n13907 ^ n13444 ;
  assign n14147 = ~n14145 & ~n14146 ;
  assign n14148 = n14147 ^ x14 ;
  assign n14149 = n14148 ^ n14144 ;
  assign n14158 = n14157 ^ n14149 ;
  assign n14166 = n14165 ^ n14158 ;
  assign n14172 = n14171 ^ n14166 ;
  assign n14176 = n14175 ^ n14172 ;
  assign n14134 = x87 & n7954 ;
  assign n14133 = x89 & n7950 ;
  assign n14135 = n14134 ^ n14133 ;
  assign n14136 = n14135 ^ x56 ;
  assign n14132 = n2255 & n7951 ;
  assign n14137 = n14136 ^ n14132 ;
  assign n14131 = x88 & n7947 ;
  assign n14138 = n14137 ^ n14131 ;
  assign n14139 = n14138 ^ n13927 ;
  assign n14140 = n14139 ^ n13888 ;
  assign n14141 = n14140 ^ n14138 ;
  assign n14142 = ~n13928 & n14141 ;
  assign n14143 = n14142 ^ n14139 ;
  assign n14177 = n14176 ^ n14143 ;
  assign n14121 = x90 & n7183 ;
  assign n14120 = x92 & n7186 ;
  assign n14122 = n14121 ^ n14120 ;
  assign n14123 = n14122 ^ x53 ;
  assign n14119 = n2696 & n7187 ;
  assign n14124 = n14123 ^ n14119 ;
  assign n14118 = x91 & n7191 ;
  assign n14125 = n14124 ^ n14118 ;
  assign n14126 = n14125 ^ n13941 ;
  assign n14127 = n14126 ^ n13937 ;
  assign n14128 = n14127 ^ n14125 ;
  assign n14129 = n13938 & ~n14128 ;
  assign n14130 = n14129 ^ n14126 ;
  assign n14178 = n14177 ^ n14130 ;
  assign n14187 = n14186 ^ n14178 ;
  assign n14115 = n13950 ^ n13885 ;
  assign n14116 = n13951 & n14115 ;
  assign n14117 = n14116 ^ n13950 ;
  assign n14188 = n14187 ^ n14117 ;
  assign n14197 = n14196 ^ n14188 ;
  assign n14201 = n14200 ^ n14197 ;
  assign n14214 = n14213 ^ n14201 ;
  assign n14112 = n13987 ^ n13983 ;
  assign n14113 = n13984 & ~n14112 ;
  assign n14114 = n14113 ^ n13987 ;
  assign n14215 = n14214 ^ n14114 ;
  assign n14224 = n14223 ^ n14215 ;
  assign n14228 = n14227 ^ n14224 ;
  assign n14237 = n14236 ^ n14228 ;
  assign n14109 = n3391 & n6145 ;
  assign n14107 = x108 & n3387 ;
  assign n14103 = n14010 ^ n14006 ;
  assign n14104 = n14007 & ~n14103 ;
  assign n14105 = n14104 ^ n14010 ;
  assign n14101 = x110 & n3390 ;
  assign n14102 = n14101 ^ x35 ;
  assign n14106 = n14105 ^ n14102 ;
  assign n14108 = n14107 ^ n14106 ;
  assign n14110 = n14109 ^ n14108 ;
  assign n14100 = x109 & n3395 ;
  assign n14111 = n14110 ^ n14100 ;
  assign n14238 = n14237 ^ n14111 ;
  assign n14239 = n14238 ^ n14023 ;
  assign n14240 = n14239 ^ n14019 ;
  assign n14241 = n14240 ^ n14238 ;
  assign n14242 = ~n14020 & ~n14241 ;
  assign n14243 = n14242 ^ n14239 ;
  assign n14252 = n14251 ^ n14243 ;
  assign n14256 = n14255 ^ n14252 ;
  assign n14265 = n14264 ^ n14256 ;
  assign n14274 = n14273 ^ n14265 ;
  assign n14097 = n14046 ^ n14042 ;
  assign n14098 = n14043 & ~n14097 ;
  assign n14099 = n14098 ^ n14046 ;
  assign n14275 = n14274 ^ n14099 ;
  assign n14094 = n14059 ^ n14055 ;
  assign n14095 = ~n14056 & ~n14094 ;
  assign n14096 = n14095 ^ n14059 ;
  assign n14276 = n14275 ^ n14096 ;
  assign n14285 = n14284 ^ n14276 ;
  assign n14091 = n14069 ^ n14060 ;
  assign n14092 = n14066 & n14091 ;
  assign n14093 = n14092 ^ n14069 ;
  assign n14286 = n14285 ^ n14093 ;
  assign n14295 = n14294 ^ n14286 ;
  assign n14299 = n14298 ^ n14295 ;
  assign n14306 = n14305 ^ n14299 ;
  assign n14088 = n14077 ^ n13861 ;
  assign n14089 = n14083 & n14088 ;
  assign n14090 = n14089 ^ n14077 ;
  assign n14307 = n14306 ^ n14090 ;
  assign n14326 = n14325 ^ n14307 ;
  assign n14543 = x127 & n1059 ;
  assign n14544 = n14543 ^ n1057 ;
  assign n14549 = n873 & n11285 ;
  assign n14550 = n14549 ^ n14543 ;
  assign n14551 = n14544 & ~n14550 ;
  assign n14552 = n14551 ^ x16 ;
  assign n14537 = x124 & n1340 ;
  assign n14536 = x126 & n1343 ;
  assign n14538 = n14537 ^ n14536 ;
  assign n14539 = n14538 ^ x20 ;
  assign n14535 = n1344 & n10461 ;
  assign n14540 = n14539 ^ n14535 ;
  assign n14534 = x125 & n1348 ;
  assign n14541 = n14540 ^ n14534 ;
  assign n14527 = x121 & n1665 ;
  assign n14526 = x123 & n1668 ;
  assign n14528 = n14527 ^ n14526 ;
  assign n14529 = n14528 ^ x23 ;
  assign n14525 = n1669 & ~n9804 ;
  assign n14530 = n14529 ^ n14525 ;
  assign n14524 = x122 & n1673 ;
  assign n14531 = n14530 ^ n14524 ;
  assign n14517 = x118 & n2032 ;
  assign n14516 = x120 & n2028 ;
  assign n14518 = n14517 ^ n14516 ;
  assign n14519 = n14518 ^ x26 ;
  assign n14515 = n2029 & n8904 ;
  assign n14520 = n14519 ^ n14515 ;
  assign n14514 = x119 & n2025 ;
  assign n14521 = n14520 ^ n14514 ;
  assign n14503 = x115 & n2593 ;
  assign n14502 = x117 & n2428 ;
  assign n14504 = n14503 ^ n14502 ;
  assign n14505 = n14504 ^ x29 ;
  assign n14501 = n2429 & ~n7860 ;
  assign n14506 = n14505 ^ n14501 ;
  assign n14500 = x116 & n2435 ;
  assign n14507 = n14506 ^ n14500 ;
  assign n14489 = x112 & n2890 ;
  assign n14488 = x114 & n2893 ;
  assign n14490 = n14489 ^ n14488 ;
  assign n14491 = n14490 ^ x32 ;
  assign n14487 = n2894 & ~n7108 ;
  assign n14492 = n14491 ^ n14487 ;
  assign n14486 = x113 & n2899 ;
  assign n14493 = n14492 ^ n14486 ;
  assign n14475 = x109 & n3387 ;
  assign n14474 = x111 & n3390 ;
  assign n14476 = n14475 ^ n14474 ;
  assign n14477 = n14476 ^ x35 ;
  assign n14473 = n3391 & ~n6370 ;
  assign n14478 = n14477 ^ n14473 ;
  assign n14472 = x110 & n3395 ;
  assign n14479 = n14478 ^ n14472 ;
  assign n14465 = x106 & n3932 ;
  assign n14464 = x108 & n3935 ;
  assign n14466 = n14465 ^ n14464 ;
  assign n14467 = n14466 ^ x38 ;
  assign n14463 = n3936 & n5687 ;
  assign n14468 = n14467 ^ n14463 ;
  assign n14462 = x107 & n3940 ;
  assign n14469 = n14468 ^ n14462 ;
  assign n14459 = n14223 ^ n14114 ;
  assign n14460 = n14215 & ~n14459 ;
  assign n14451 = x103 & n4482 ;
  assign n14450 = x105 & n4478 ;
  assign n14452 = n14451 ^ n14450 ;
  assign n14453 = n14452 ^ x41 ;
  assign n14449 = n4479 & ~n5034 ;
  assign n14454 = n14453 ^ n14449 ;
  assign n14448 = x104 & n4475 ;
  assign n14455 = n14454 ^ n14448 ;
  assign n14444 = n14204 ^ n14201 ;
  assign n14445 = n14213 & n14444 ;
  assign n14446 = n14445 ^ n14201 ;
  assign n14441 = x101 & n5121 ;
  assign n14439 = n4425 & n5117 ;
  assign n14435 = x100 & n5113 ;
  assign n14434 = x102 & n5116 ;
  assign n14436 = n14435 ^ n14434 ;
  assign n14437 = n14436 ^ x44 ;
  assign n14429 = n14177 ^ n14125 ;
  assign n14430 = ~n14130 & n14429 ;
  assign n14431 = n14430 ^ n14125 ;
  assign n14427 = x95 & n6449 ;
  assign n14422 = x94 & n6687 ;
  assign n14421 = x96 & n6444 ;
  assign n14423 = n14422 ^ n14421 ;
  assign n14424 = n14423 ^ x50 ;
  assign n14420 = n3336 & n6445 ;
  assign n14425 = n14424 ^ n14420 ;
  assign n14416 = n14176 ^ n14138 ;
  assign n14417 = n14143 & n14416 ;
  assign n14418 = n14417 ^ n14138 ;
  assign n14414 = x92 & n7191 ;
  assign n14409 = x91 & n7183 ;
  assign n14408 = x93 & n7186 ;
  assign n14410 = n14409 ^ n14408 ;
  assign n14411 = n14410 ^ x53 ;
  assign n14407 = n2842 & n7187 ;
  assign n14412 = n14411 ^ n14407 ;
  assign n14401 = x88 & n7954 ;
  assign n14400 = x90 & n7950 ;
  assign n14402 = n14401 ^ n14400 ;
  assign n14403 = n14402 ^ x56 ;
  assign n14399 = n2398 & n7951 ;
  assign n14404 = n14403 ^ n14399 ;
  assign n14398 = x89 & n7947 ;
  assign n14405 = n14404 ^ n14398 ;
  assign n14394 = n14175 ^ n14157 ;
  assign n14395 = n14172 & n14394 ;
  assign n14396 = n14395 ^ n14157 ;
  assign n14381 = n14148 ^ x62 ;
  assign n14382 = n14381 ^ n14165 ;
  assign n14383 = n14168 ^ n14165 ;
  assign n14384 = n14383 ^ n14149 ;
  assign n14387 = n14170 & ~n14384 ;
  assign n14388 = n14387 ^ n14149 ;
  assign n14389 = ~n14382 & n14388 ;
  assign n14390 = n14389 ^ n14148 ;
  assign n14378 = x80 ^ x62 ;
  assign n14379 = n14378 ^ x81 ;
  assign n14375 = n1635 & n9652 ;
  assign n14374 = x83 & n9648 ;
  assign n14376 = n14375 ^ n14374 ;
  assign n14372 = x82 & n9655 ;
  assign n14371 = x84 & n9651 ;
  assign n14373 = n14372 ^ n14371 ;
  assign n14377 = n14376 ^ n14373 ;
  assign n14380 = n14379 ^ n14377 ;
  assign n14391 = n14390 ^ n14380 ;
  assign n14369 = n14168 ^ x81 ;
  assign n14370 = ~n9956 & n14369 ;
  assign n14392 = n14391 ^ n14370 ;
  assign n14364 = x85 & n8750 ;
  assign n14363 = x87 & n8746 ;
  assign n14365 = n14364 ^ n14363 ;
  assign n14366 = n14365 ^ x59 ;
  assign n14362 = n1987 & n8747 ;
  assign n14367 = n14366 ^ n14362 ;
  assign n14361 = x86 & n8743 ;
  assign n14368 = n14367 ^ n14361 ;
  assign n14393 = n14392 ^ n14368 ;
  assign n14397 = n14396 ^ n14393 ;
  assign n14406 = n14405 ^ n14397 ;
  assign n14413 = n14412 ^ n14406 ;
  assign n14415 = n14414 ^ n14413 ;
  assign n14419 = n14418 ^ n14415 ;
  assign n14426 = n14425 ^ n14419 ;
  assign n14428 = n14427 ^ n14426 ;
  assign n14432 = n14431 ^ n14428 ;
  assign n14358 = n3851 & n5749 ;
  assign n14356 = x97 & n5981 ;
  assign n14354 = x99 & n5748 ;
  assign n14350 = n14186 ^ n14117 ;
  assign n14351 = ~n14187 & n14350 ;
  assign n14352 = n14351 ^ n14186 ;
  assign n14353 = n14352 ^ x47 ;
  assign n14355 = n14354 ^ n14353 ;
  assign n14357 = n14356 ^ n14355 ;
  assign n14359 = n14358 ^ n14357 ;
  assign n14349 = x98 & n5755 ;
  assign n14360 = n14359 ^ n14349 ;
  assign n14433 = n14432 ^ n14360 ;
  assign n14438 = n14437 ^ n14433 ;
  assign n14440 = n14439 ^ n14438 ;
  assign n14442 = n14441 ^ n14440 ;
  assign n14346 = n14200 ^ n14196 ;
  assign n14347 = n14197 & n14346 ;
  assign n14348 = n14347 ^ n14200 ;
  assign n14443 = n14442 ^ n14348 ;
  assign n14447 = n14446 ^ n14443 ;
  assign n14456 = n14455 ^ n14447 ;
  assign n14457 = n14456 ^ n14223 ;
  assign n14461 = n14460 ^ n14457 ;
  assign n14470 = n14469 ^ n14461 ;
  assign n14343 = n14236 ^ n14227 ;
  assign n14344 = n14228 & n14343 ;
  assign n14345 = n14344 ^ n14236 ;
  assign n14471 = n14470 ^ n14345 ;
  assign n14480 = n14479 ^ n14471 ;
  assign n14481 = n14480 ^ n14237 ;
  assign n14482 = n14481 ^ n14480 ;
  assign n14483 = n14482 ^ n14105 ;
  assign n14484 = n14111 & n14483 ;
  assign n14485 = n14484 ^ n14481 ;
  assign n14494 = n14493 ^ n14485 ;
  assign n14496 = n14494 ^ n14238 ;
  assign n14495 = n14494 ^ n14251 ;
  assign n14497 = n14496 ^ n14495 ;
  assign n14498 = ~n14243 & n14497 ;
  assign n14499 = n14498 ^ n14496 ;
  assign n14508 = n14507 ^ n14499 ;
  assign n14509 = n14508 ^ n14264 ;
  assign n14510 = n14509 ^ n14255 ;
  assign n14511 = n14510 ^ n14508 ;
  assign n14512 = n14256 & n14511 ;
  assign n14513 = n14512 ^ n14509 ;
  assign n14522 = n14521 ^ n14513 ;
  assign n14340 = n14273 ^ n14099 ;
  assign n14341 = ~n14274 & ~n14340 ;
  assign n14342 = n14341 ^ n14273 ;
  assign n14523 = n14522 ^ n14342 ;
  assign n14532 = n14531 ^ n14523 ;
  assign n14337 = n14284 ^ n14096 ;
  assign n14338 = n14276 & ~n14337 ;
  assign n14339 = n14338 ^ n14284 ;
  assign n14533 = n14532 ^ n14339 ;
  assign n14542 = n14541 ^ n14533 ;
  assign n14553 = n14552 ^ n14542 ;
  assign n14334 = n14294 ^ n14093 ;
  assign n14335 = ~n14286 & ~n14334 ;
  assign n14336 = n14335 ^ n14294 ;
  assign n14554 = n14553 ^ n14336 ;
  assign n14330 = n14325 ^ n14295 ;
  assign n14327 = n14305 ^ n14298 ;
  assign n14331 = n14327 ^ n14295 ;
  assign n14332 = n14331 ^ n14090 ;
  assign n14333 = ~n14330 & n14332 ;
  assign n14555 = n14554 ^ n14333 ;
  assign n14328 = n14298 ^ n14090 ;
  assign n14329 = ~n14327 & ~n14328 ;
  assign n14556 = n14555 ^ n14329 ;
  assign n14788 = n14295 & n14305 ;
  assign n14789 = n14788 ^ n14554 ;
  assign n14790 = n14090 & n14298 ;
  assign n14791 = n14790 ^ n14328 ;
  assign n14792 = n14789 & n14791 ;
  assign n14793 = n14305 ^ n14295 ;
  assign n14794 = n14793 ^ n14789 ;
  assign n14795 = n14794 ^ n14554 ;
  assign n14798 = ~n14790 & ~n14795 ;
  assign n14799 = n14798 ^ n14554 ;
  assign n14800 = ~n14325 & ~n14799 ;
  assign n14801 = n14792 & ~n14800 ;
  assign n14802 = n14325 ^ n14305 ;
  assign n14803 = ~n14793 & n14802 ;
  assign n14804 = n14803 ^ n14325 ;
  assign n14805 = ~n14554 & ~n14790 ;
  assign n14806 = n14804 & n14805 ;
  assign n14807 = n14806 ^ n14804 ;
  assign n14808 = ~n14801 & ~n14807 ;
  assign n14784 = n14552 ^ n14336 ;
  assign n14785 = n14553 & n14784 ;
  assign n14786 = n14785 ^ n14552 ;
  assign n14777 = x125 & n1340 ;
  assign n14776 = x127 & n1343 ;
  assign n14778 = n14777 ^ n14776 ;
  assign n14779 = n14778 ^ x20 ;
  assign n14775 = n1344 & n10986 ;
  assign n14780 = n14779 ^ n14775 ;
  assign n14774 = x126 & n1348 ;
  assign n14781 = n14780 ^ n14774 ;
  assign n14767 = x122 & n1665 ;
  assign n14766 = x124 & n1668 ;
  assign n14768 = n14767 ^ n14766 ;
  assign n14769 = n14768 ^ x23 ;
  assign n14765 = n1669 & n10117 ;
  assign n14770 = n14769 ^ n14765 ;
  assign n14764 = x123 & n1673 ;
  assign n14771 = n14770 ^ n14764 ;
  assign n14758 = x119 & n2032 ;
  assign n14757 = x121 & n2028 ;
  assign n14759 = n14758 ^ n14757 ;
  assign n14760 = n14759 ^ x26 ;
  assign n14756 = n2029 & n8979 ;
  assign n14761 = n14760 ^ n14756 ;
  assign n14755 = x120 & n2025 ;
  assign n14762 = n14761 ^ n14755 ;
  assign n14746 = n14507 ^ n14494 ;
  assign n14747 = n14499 & n14746 ;
  assign n14748 = n14747 ^ n14494 ;
  assign n14740 = x116 & n2593 ;
  assign n14739 = x118 & n2428 ;
  assign n14741 = n14740 ^ n14739 ;
  assign n14742 = n14741 ^ x29 ;
  assign n14738 = n2429 & ~n8140 ;
  assign n14743 = n14742 ^ n14738 ;
  assign n14737 = x117 & n2435 ;
  assign n14744 = n14743 ^ n14737 ;
  assign n14733 = n14493 ^ n14480 ;
  assign n14734 = n14485 & ~n14733 ;
  assign n14735 = n14734 ^ n14480 ;
  assign n14727 = x113 & n2890 ;
  assign n14726 = x115 & n2893 ;
  assign n14728 = n14727 ^ n14726 ;
  assign n14729 = n14728 ^ x32 ;
  assign n14725 = n2894 & ~n7353 ;
  assign n14730 = n14729 ^ n14725 ;
  assign n14724 = x114 & n2899 ;
  assign n14731 = n14730 ^ n14724 ;
  assign n14720 = n14479 ^ n14345 ;
  assign n14721 = n14471 & n14720 ;
  assign n14722 = n14721 ^ n14479 ;
  assign n14718 = x111 & n3395 ;
  assign n14713 = x110 & n3387 ;
  assign n14712 = x112 & n3390 ;
  assign n14714 = n14713 ^ n14712 ;
  assign n14715 = n14714 ^ x35 ;
  assign n14711 = n3391 & ~n6616 ;
  assign n14716 = n14715 ^ n14711 ;
  assign n14707 = n14469 ^ n14456 ;
  assign n14708 = ~n14461 & ~n14707 ;
  assign n14709 = n14708 ^ n14456 ;
  assign n14701 = x107 & n3932 ;
  assign n14700 = x109 & n3935 ;
  assign n14702 = n14701 ^ n14700 ;
  assign n14703 = n14702 ^ x38 ;
  assign n14699 = n3936 & n5912 ;
  assign n14704 = n14703 ^ n14699 ;
  assign n14698 = x108 & n3940 ;
  assign n14705 = n14704 ^ n14698 ;
  assign n14691 = x104 & n4482 ;
  assign n14690 = x106 & n4478 ;
  assign n14692 = n14691 ^ n14690 ;
  assign n14693 = n14692 ^ x41 ;
  assign n14689 = n4479 & ~n5257 ;
  assign n14694 = n14693 ^ n14689 ;
  assign n14688 = x105 & n4475 ;
  assign n14695 = n14694 ^ n14688 ;
  assign n14684 = n14433 ^ n14348 ;
  assign n14685 = n14442 & n14684 ;
  assign n14686 = n14685 ^ n14433 ;
  assign n14678 = x101 & n5113 ;
  assign n14677 = x103 & n5116 ;
  assign n14679 = n14678 ^ n14677 ;
  assign n14680 = n14679 ^ x44 ;
  assign n14676 = ~n4624 & n5117 ;
  assign n14681 = n14680 ^ n14676 ;
  assign n14675 = x102 & n5121 ;
  assign n14682 = n14681 ^ n14675 ;
  assign n14671 = n14432 ^ n14352 ;
  assign n14672 = ~n14360 & n14671 ;
  assign n14673 = n14672 ^ n14432 ;
  assign n14665 = x98 & n5981 ;
  assign n14664 = x100 & n5748 ;
  assign n14666 = n14665 ^ n14664 ;
  assign n14667 = n14666 ^ x47 ;
  assign n14663 = n4048 & n5749 ;
  assign n14668 = n14667 ^ n14663 ;
  assign n14662 = x99 & n5755 ;
  assign n14669 = n14668 ^ n14662 ;
  assign n14655 = x95 & n6687 ;
  assign n14654 = x97 & n6444 ;
  assign n14656 = n14655 ^ n14654 ;
  assign n14657 = n14656 ^ x50 ;
  assign n14653 = n3501 & n6445 ;
  assign n14658 = n14657 ^ n14653 ;
  assign n14652 = x96 & n6449 ;
  assign n14659 = n14658 ^ n14652 ;
  assign n14645 = x92 & n7183 ;
  assign n14644 = x94 & n7186 ;
  assign n14646 = n14645 ^ n14644 ;
  assign n14647 = n14646 ^ x53 ;
  assign n14643 = n3010 & n7187 ;
  assign n14648 = n14647 ^ n14643 ;
  assign n14642 = x93 & n7191 ;
  assign n14649 = n14648 ^ n14642 ;
  assign n14638 = n14405 ^ n14396 ;
  assign n14639 = ~n14397 & n14638 ;
  assign n14640 = n14639 ^ n14405 ;
  assign n14632 = x89 & n7954 ;
  assign n14631 = x91 & n7950 ;
  assign n14633 = n14632 ^ n14631 ;
  assign n14634 = n14633 ^ x56 ;
  assign n14630 = n2548 & n7951 ;
  assign n14635 = n14634 ^ n14630 ;
  assign n14629 = x90 & n7947 ;
  assign n14636 = n14635 ^ n14629 ;
  assign n14601 = ~n1107 & ~n14377 ;
  assign n14616 = n14601 ^ n11894 ;
  assign n14605 = n14377 ^ x80 ;
  assign n14621 = n1017 & ~n14605 ;
  assign n14607 = x81 ^ x79 ;
  assign n14622 = n14621 ^ n14607 ;
  assign n14623 = n14616 & n14622 ;
  assign n14606 = n14377 ^ x62 ;
  assign n14624 = n14623 ^ n14606 ;
  assign n14611 = ~x81 & ~n14377 ;
  assign n14612 = n14611 ^ n14606 ;
  assign n14613 = ~n14607 & ~n14612 ;
  assign n14614 = n14613 ^ n14606 ;
  assign n14615 = n14605 & ~n14614 ;
  assign n14625 = n14624 ^ n14615 ;
  assign n14599 = n14377 ^ x81 ;
  assign n14600 = n14377 ^ n1107 ;
  assign n14602 = n14601 ^ n14600 ;
  assign n14585 = ~x63 & n1107 ;
  assign n14603 = n14602 ^ n14585 ;
  assign n14604 = ~n14599 & ~n14603 ;
  assign n14626 = n14625 ^ n14604 ;
  assign n14592 = x83 & n9655 ;
  assign n14591 = x85 & n9651 ;
  assign n14593 = n14592 ^ n14591 ;
  assign n14594 = n14593 ^ x62 ;
  assign n14590 = n1748 & n9652 ;
  assign n14595 = n14594 ^ n14590 ;
  assign n14589 = x84 & n9648 ;
  assign n14596 = n14595 ^ n14589 ;
  assign n14588 = n1198 ^ x17 ;
  assign n14597 = n14596 ^ n14588 ;
  assign n14584 = n1198 ^ n1107 ;
  assign n14586 = n14585 ^ n14584 ;
  assign n14587 = ~n9956 & n14586 ;
  assign n14598 = n14597 ^ n14587 ;
  assign n14627 = n14626 ^ n14598 ;
  assign n14582 = x87 & n8743 ;
  assign n14580 = n2131 & n8747 ;
  assign n14578 = x86 & n8750 ;
  assign n14574 = n14390 ^ n14368 ;
  assign n14575 = n14392 & ~n14574 ;
  assign n14576 = n14575 ^ n14390 ;
  assign n14572 = x88 & n8746 ;
  assign n14573 = n14572 ^ x59 ;
  assign n14577 = n14576 ^ n14573 ;
  assign n14579 = n14578 ^ n14577 ;
  assign n14581 = n14580 ^ n14579 ;
  assign n14583 = n14582 ^ n14581 ;
  assign n14628 = n14627 ^ n14583 ;
  assign n14637 = n14636 ^ n14628 ;
  assign n14641 = n14640 ^ n14637 ;
  assign n14650 = n14649 ^ n14641 ;
  assign n14569 = n14418 ^ n14406 ;
  assign n14570 = n14415 & n14569 ;
  assign n14571 = n14570 ^ n14406 ;
  assign n14651 = n14650 ^ n14571 ;
  assign n14660 = n14659 ^ n14651 ;
  assign n14566 = n14431 ^ n14419 ;
  assign n14567 = n14428 & n14566 ;
  assign n14568 = n14567 ^ n14419 ;
  assign n14661 = n14660 ^ n14568 ;
  assign n14670 = n14669 ^ n14661 ;
  assign n14674 = n14673 ^ n14670 ;
  assign n14683 = n14682 ^ n14674 ;
  assign n14687 = n14686 ^ n14683 ;
  assign n14696 = n14695 ^ n14687 ;
  assign n14563 = n14455 ^ n14446 ;
  assign n14564 = n14447 & ~n14563 ;
  assign n14565 = n14564 ^ n14455 ;
  assign n14697 = n14696 ^ n14565 ;
  assign n14706 = n14705 ^ n14697 ;
  assign n14710 = n14709 ^ n14706 ;
  assign n14717 = n14716 ^ n14710 ;
  assign n14719 = n14718 ^ n14717 ;
  assign n14723 = n14722 ^ n14719 ;
  assign n14732 = n14731 ^ n14723 ;
  assign n14736 = n14735 ^ n14732 ;
  assign n14745 = n14744 ^ n14736 ;
  assign n14749 = n14748 ^ n14745 ;
  assign n14751 = n14749 ^ n14508 ;
  assign n14750 = n14749 ^ n14521 ;
  assign n14752 = n14751 ^ n14750 ;
  assign n14753 = n14513 & n14752 ;
  assign n14754 = n14753 ^ n14751 ;
  assign n14763 = n14762 ^ n14754 ;
  assign n14772 = n14771 ^ n14763 ;
  assign n14560 = n14531 ^ n14342 ;
  assign n14561 = ~n14523 & n14560 ;
  assign n14562 = n14561 ^ n14531 ;
  assign n14773 = n14772 ^ n14562 ;
  assign n14782 = n14781 ^ n14773 ;
  assign n14557 = n14541 ^ n14339 ;
  assign n14558 = ~n14533 & n14557 ;
  assign n14559 = n14558 ^ n14541 ;
  assign n14783 = n14782 ^ n14559 ;
  assign n14787 = n14786 ^ n14783 ;
  assign n14809 = n14808 ^ n14787 ;
  assign n15021 = n14559 & n14786 ;
  assign n15020 = ~n14773 & ~n14781 ;
  assign n15022 = n15021 ^ n15020 ;
  assign n15015 = n1344 & n10155 ;
  assign n15014 = x126 & n1340 ;
  assign n15016 = n15015 ^ n15014 ;
  assign n15017 = n15016 ^ x20 ;
  assign n15013 = x127 & n1348 ;
  assign n15018 = n15017 ^ n15013 ;
  assign n15006 = x123 & n1665 ;
  assign n15005 = x125 & n1668 ;
  assign n15007 = n15006 ^ n15005 ;
  assign n15008 = n15007 ^ x23 ;
  assign n15004 = n1669 & n10416 ;
  assign n15009 = n15008 ^ n15004 ;
  assign n15003 = x124 & n1673 ;
  assign n15010 = n15009 ^ n15003 ;
  assign n14992 = x120 & n2032 ;
  assign n14991 = x122 & n2028 ;
  assign n14993 = n14992 ^ n14991 ;
  assign n14994 = n14993 ^ x26 ;
  assign n14990 = n2029 & ~n9261 ;
  assign n14995 = n14994 ^ n14990 ;
  assign n14989 = x121 & n2025 ;
  assign n14996 = n14995 ^ n14989 ;
  assign n14981 = x117 & n2593 ;
  assign n14980 = x119 & n2428 ;
  assign n14982 = n14981 ^ n14980 ;
  assign n14983 = n14982 ^ x29 ;
  assign n14979 = n2429 & n8405 ;
  assign n14984 = n14983 ^ n14979 ;
  assign n14978 = x118 & n2435 ;
  assign n14985 = n14984 ^ n14978 ;
  assign n14972 = x114 & n2890 ;
  assign n14971 = x116 & n2893 ;
  assign n14973 = n14972 ^ n14971 ;
  assign n14974 = n14973 ^ x32 ;
  assign n14970 = n2894 & ~n7604 ;
  assign n14975 = n14974 ^ n14970 ;
  assign n14969 = x115 & n2899 ;
  assign n14976 = n14975 ^ n14969 ;
  assign n14962 = x111 & n3387 ;
  assign n14961 = x113 & n3390 ;
  assign n14963 = n14962 ^ n14961 ;
  assign n14964 = n14963 ^ x35 ;
  assign n14960 = n3391 & ~n6849 ;
  assign n14965 = n14964 ^ n14960 ;
  assign n14959 = x112 & n3395 ;
  assign n14966 = n14965 ^ n14959 ;
  assign n14948 = x108 & n3932 ;
  assign n14947 = x110 & n3935 ;
  assign n14949 = n14948 ^ n14947 ;
  assign n14950 = n14949 ^ x38 ;
  assign n14946 = n3936 & n6145 ;
  assign n14951 = n14950 ^ n14946 ;
  assign n14945 = x109 & n3940 ;
  assign n14952 = n14951 ^ n14945 ;
  assign n14934 = x105 & n4482 ;
  assign n14933 = x107 & n4478 ;
  assign n14935 = n14934 ^ n14933 ;
  assign n14936 = n14935 ^ x41 ;
  assign n14932 = n4479 & ~n5459 ;
  assign n14937 = n14936 ^ n14932 ;
  assign n14931 = x106 & n4475 ;
  assign n14938 = n14937 ^ n14931 ;
  assign n14924 = x102 & n5113 ;
  assign n14923 = x104 & n5116 ;
  assign n14925 = n14924 ^ n14923 ;
  assign n14926 = n14925 ^ x44 ;
  assign n14922 = ~n4830 & n5117 ;
  assign n14927 = n14926 ^ n14922 ;
  assign n14921 = x103 & n5121 ;
  assign n14928 = n14927 ^ n14921 ;
  assign n14910 = x99 & n5981 ;
  assign n14909 = x101 & n5748 ;
  assign n14911 = n14910 ^ n14909 ;
  assign n14912 = n14911 ^ x47 ;
  assign n14908 = n4223 & n5749 ;
  assign n14913 = n14912 ^ n14908 ;
  assign n14907 = x100 & n5755 ;
  assign n14914 = n14913 ^ n14907 ;
  assign n14903 = n14659 ^ n14568 ;
  assign n14904 = n14660 & n14903 ;
  assign n14905 = n14904 ^ n14659 ;
  assign n14897 = x96 & n6687 ;
  assign n14896 = x98 & n6444 ;
  assign n14898 = n14897 ^ n14896 ;
  assign n14899 = n14898 ^ x50 ;
  assign n14895 = n3673 & n6445 ;
  assign n14900 = n14899 ^ n14895 ;
  assign n14894 = x97 & n6449 ;
  assign n14901 = n14900 ^ n14894 ;
  assign n14890 = n14649 ^ n14571 ;
  assign n14891 = n14650 & n14890 ;
  assign n14892 = n14891 ^ n14649 ;
  assign n14884 = x93 & n7183 ;
  assign n14883 = x95 & n7186 ;
  assign n14885 = n14884 ^ n14883 ;
  assign n14886 = n14885 ^ x53 ;
  assign n14882 = n3166 & n7187 ;
  assign n14887 = n14886 ^ n14882 ;
  assign n14881 = x94 & n7191 ;
  assign n14888 = n14887 ^ n14881 ;
  assign n14872 = x87 & n8750 ;
  assign n14871 = x89 & n8746 ;
  assign n14873 = n14872 ^ n14871 ;
  assign n14874 = n14873 ^ x59 ;
  assign n14870 = n2255 & n8747 ;
  assign n14875 = n14874 ^ n14870 ;
  assign n14869 = x88 & n8743 ;
  assign n14876 = n14875 ^ n14869 ;
  assign n14863 = x84 & n9655 ;
  assign n14862 = x86 & n9651 ;
  assign n14864 = n14863 ^ n14862 ;
  assign n14865 = n14864 ^ x62 ;
  assign n14861 = n1868 & n9652 ;
  assign n14866 = n14865 ^ n14861 ;
  assign n14860 = x85 & n9648 ;
  assign n14867 = n14866 ^ n14860 ;
  assign n14851 = x81 ^ x17 ;
  assign n14854 = ~n11895 & n14584 ;
  assign n14855 = n14854 ^ n1107 ;
  assign n14856 = ~n14851 & ~n14855 ;
  assign n14857 = n14856 ^ x17 ;
  assign n14858 = n12206 & ~n14857 ;
  assign n14849 = x82 & n11895 ;
  assign n14848 = x83 & n9956 ;
  assign n14850 = n14849 ^ n14848 ;
  assign n14859 = n14858 ^ n14850 ;
  assign n14868 = n14867 ^ n14859 ;
  assign n14877 = n14876 ^ n14868 ;
  assign n14845 = n14626 ^ n14596 ;
  assign n14846 = n14598 & n14845 ;
  assign n14847 = n14846 ^ n14626 ;
  assign n14878 = n14877 ^ n14847 ;
  assign n14835 = x90 & n7954 ;
  assign n14834 = x92 & n7950 ;
  assign n14836 = n14835 ^ n14834 ;
  assign n14837 = n14836 ^ x56 ;
  assign n14833 = n2696 & n7951 ;
  assign n14838 = n14837 ^ n14833 ;
  assign n14832 = x91 & n7947 ;
  assign n14839 = n14838 ^ n14832 ;
  assign n14841 = n14839 ^ n14627 ;
  assign n14840 = n14839 ^ n14576 ;
  assign n14842 = n14841 ^ n14840 ;
  assign n14843 = n14583 & n14842 ;
  assign n14844 = n14843 ^ n14841 ;
  assign n14879 = n14878 ^ n14844 ;
  assign n14829 = n14640 ^ n14636 ;
  assign n14830 = ~n14637 & n14829 ;
  assign n14831 = n14830 ^ n14640 ;
  assign n14880 = n14879 ^ n14831 ;
  assign n14889 = n14888 ^ n14880 ;
  assign n14893 = n14892 ^ n14889 ;
  assign n14902 = n14901 ^ n14893 ;
  assign n14906 = n14905 ^ n14902 ;
  assign n14915 = n14914 ^ n14906 ;
  assign n14916 = n14915 ^ n14673 ;
  assign n14917 = n14916 ^ n14669 ;
  assign n14918 = n14917 ^ n14915 ;
  assign n14919 = ~n14670 & n14918 ;
  assign n14920 = n14919 ^ n14916 ;
  assign n14929 = n14928 ^ n14920 ;
  assign n14826 = n14686 ^ n14682 ;
  assign n14827 = ~n14683 & n14826 ;
  assign n14828 = n14827 ^ n14686 ;
  assign n14930 = n14929 ^ n14828 ;
  assign n14939 = n14938 ^ n14930 ;
  assign n14940 = n14939 ^ n14695 ;
  assign n14941 = n14940 ^ n14565 ;
  assign n14942 = n14941 ^ n14939 ;
  assign n14943 = n14696 & n14942 ;
  assign n14944 = n14943 ^ n14940 ;
  assign n14953 = n14952 ^ n14944 ;
  assign n14954 = n14953 ^ n14709 ;
  assign n14955 = n14954 ^ n14705 ;
  assign n14956 = n14955 ^ n14953 ;
  assign n14957 = ~n14706 & ~n14956 ;
  assign n14958 = n14957 ^ n14954 ;
  assign n14967 = n14966 ^ n14958 ;
  assign n14823 = n14722 ^ n14710 ;
  assign n14824 = ~n14719 & ~n14823 ;
  assign n14825 = n14824 ^ n14710 ;
  assign n14968 = n14967 ^ n14825 ;
  assign n14977 = n14976 ^ n14968 ;
  assign n14986 = n14985 ^ n14977 ;
  assign n14820 = n14735 ^ n14731 ;
  assign n14821 = n14732 & ~n14820 ;
  assign n14822 = n14821 ^ n14735 ;
  assign n14987 = n14986 ^ n14822 ;
  assign n14817 = n14748 ^ n14744 ;
  assign n14818 = ~n14745 & n14817 ;
  assign n14819 = n14818 ^ n14748 ;
  assign n14988 = n14987 ^ n14819 ;
  assign n14997 = n14996 ^ n14988 ;
  assign n14999 = n14997 ^ n14749 ;
  assign n14998 = n14997 ^ n14762 ;
  assign n15000 = n14999 ^ n14998 ;
  assign n15001 = n14754 & n15000 ;
  assign n15002 = n15001 ^ n14999 ;
  assign n15011 = n15010 ^ n15002 ;
  assign n14814 = n14771 ^ n14562 ;
  assign n14815 = n14772 & n14814 ;
  assign n14816 = n14815 ^ n14771 ;
  assign n15012 = n15011 ^ n14816 ;
  assign n15019 = n15018 ^ n15012 ;
  assign n15023 = n15022 ^ n15019 ;
  assign n14810 = n14808 ^ n14782 ;
  assign n14811 = n14786 ^ n14559 ;
  assign n14812 = n14811 ^ n14782 ;
  assign n14813 = ~n14810 & n14812 ;
  assign n15024 = n15023 ^ n14813 ;
  assign n15248 = x124 & n1665 ;
  assign n15247 = x126 & n1668 ;
  assign n15249 = n15248 ^ n15247 ;
  assign n15250 = n15249 ^ x23 ;
  assign n15246 = n1669 & n10461 ;
  assign n15251 = n15250 ^ n15246 ;
  assign n15245 = x125 & n1673 ;
  assign n15252 = n15251 ^ n15245 ;
  assign n15234 = x121 & n2032 ;
  assign n15233 = x123 & n2028 ;
  assign n15235 = n15234 ^ n15233 ;
  assign n15236 = n15235 ^ x26 ;
  assign n15232 = n2029 & ~n9804 ;
  assign n15237 = n15236 ^ n15232 ;
  assign n15231 = x122 & n2025 ;
  assign n15238 = n15237 ^ n15231 ;
  assign n15227 = n14985 ^ n14822 ;
  assign n15228 = n14986 & ~n15227 ;
  assign n15229 = n15228 ^ n14985 ;
  assign n15221 = x118 & n2593 ;
  assign n15220 = x120 & n2428 ;
  assign n15222 = n15221 ^ n15220 ;
  assign n15223 = n15222 ^ x29 ;
  assign n15219 = n2429 & n8904 ;
  assign n15224 = n15223 ^ n15219 ;
  assign n15218 = x119 & n2435 ;
  assign n15225 = n15224 ^ n15218 ;
  assign n15207 = x115 & n2890 ;
  assign n15206 = x117 & n2893 ;
  assign n15208 = n15207 ^ n15206 ;
  assign n15209 = n15208 ^ x32 ;
  assign n15205 = n2894 & ~n7860 ;
  assign n15210 = n15209 ^ n15205 ;
  assign n15204 = x116 & n2899 ;
  assign n15211 = n15210 ^ n15204 ;
  assign n15193 = x112 & n3387 ;
  assign n15192 = x114 & n3390 ;
  assign n15194 = n15193 ^ n15192 ;
  assign n15195 = n15194 ^ x35 ;
  assign n15191 = n3391 & ~n7108 ;
  assign n15196 = n15195 ^ n15191 ;
  assign n15190 = x113 & n3395 ;
  assign n15197 = n15196 ^ n15190 ;
  assign n15179 = x109 & n3932 ;
  assign n15178 = x111 & n3935 ;
  assign n15180 = n15179 ^ n15178 ;
  assign n15181 = n15180 ^ x38 ;
  assign n15177 = n3936 & ~n6370 ;
  assign n15182 = n15181 ^ n15177 ;
  assign n15176 = x110 & n3940 ;
  assign n15183 = n15182 ^ n15176 ;
  assign n15169 = x106 & n4482 ;
  assign n15168 = x108 & n4478 ;
  assign n15170 = n15169 ^ n15168 ;
  assign n15171 = n15170 ^ x41 ;
  assign n15167 = n4479 & n5687 ;
  assign n15172 = n15171 ^ n15167 ;
  assign n15166 = x107 & n4475 ;
  assign n15173 = n15172 ^ n15166 ;
  assign n15162 = n14928 ^ n14915 ;
  assign n15163 = n14920 & n15162 ;
  assign n15164 = n15163 ^ n14915 ;
  assign n15156 = x103 & n5113 ;
  assign n15155 = x105 & n5116 ;
  assign n15157 = n15156 ^ n15155 ;
  assign n15158 = n15157 ^ x44 ;
  assign n15154 = ~n5034 & n5117 ;
  assign n15159 = n15158 ^ n15154 ;
  assign n15153 = x104 & n5121 ;
  assign n15160 = n15159 ^ n15153 ;
  assign n15142 = x100 & n5981 ;
  assign n15141 = x102 & n5748 ;
  assign n15143 = n15142 ^ n15141 ;
  assign n15144 = n15143 ^ x47 ;
  assign n15140 = n4425 & n5749 ;
  assign n15145 = n15144 ^ n15140 ;
  assign n15139 = x101 & n5755 ;
  assign n15146 = n15145 ^ n15139 ;
  assign n15129 = n14878 ^ n14839 ;
  assign n15130 = ~n14844 & ~n15129 ;
  assign n15131 = n15130 ^ n14839 ;
  assign n15127 = x95 & n7191 ;
  assign n15122 = x94 & n7183 ;
  assign n15121 = x96 & n7186 ;
  assign n15123 = n15122 ^ n15121 ;
  assign n15124 = n15123 ^ x53 ;
  assign n15120 = n3336 & n7187 ;
  assign n15125 = n15124 ^ n15120 ;
  assign n15113 = x88 & n8750 ;
  assign n15112 = x90 & n8746 ;
  assign n15114 = n15113 ^ n15112 ;
  assign n15115 = n15114 ^ x59 ;
  assign n15111 = n2398 & n8747 ;
  assign n15116 = n15115 ^ n15111 ;
  assign n15110 = x89 & n8743 ;
  assign n15117 = n15116 ^ n15110 ;
  assign n15103 = x85 & n9655 ;
  assign n15102 = x87 & n9651 ;
  assign n15104 = n15103 ^ n15102 ;
  assign n15105 = n15104 ^ x62 ;
  assign n15101 = n1987 & n9652 ;
  assign n15106 = n15105 ^ n15101 ;
  assign n15100 = x86 & n9648 ;
  assign n15107 = n15106 ^ n15100 ;
  assign n15096 = ~x84 & n9956 ;
  assign n15097 = n15096 ^ n14849 ;
  assign n15098 = n15097 ^ n9956 ;
  assign n15095 = x83 & n12206 ;
  assign n15099 = n15098 ^ n15095 ;
  assign n15108 = n15107 ^ n15099 ;
  assign n15092 = n14867 ^ n14858 ;
  assign n15093 = n14859 & n15092 ;
  assign n15094 = n15093 ^ n14867 ;
  assign n15109 = n15108 ^ n15094 ;
  assign n15118 = n15117 ^ n15109 ;
  assign n15089 = n14876 ^ n14847 ;
  assign n15090 = ~n14877 & n15089 ;
  assign n15082 = x91 & n7954 ;
  assign n15081 = x93 & n7950 ;
  assign n15083 = n15082 ^ n15081 ;
  assign n15084 = n15083 ^ x56 ;
  assign n15080 = n2842 & n7951 ;
  assign n15085 = n15084 ^ n15080 ;
  assign n15079 = x92 & n7947 ;
  assign n15086 = n15085 ^ n15079 ;
  assign n15087 = n15086 ^ n14876 ;
  assign n15091 = n15090 ^ n15087 ;
  assign n15119 = n15118 ^ n15091 ;
  assign n15126 = n15125 ^ n15119 ;
  assign n15128 = n15127 ^ n15126 ;
  assign n15132 = n15131 ^ n15128 ;
  assign n15076 = n3851 & n6445 ;
  assign n15074 = x97 & n6687 ;
  assign n15070 = n14888 ^ n14831 ;
  assign n15071 = ~n14880 & n15070 ;
  assign n15072 = n15071 ^ n14888 ;
  assign n15068 = x99 & n6444 ;
  assign n15069 = n15068 ^ x50 ;
  assign n15073 = n15072 ^ n15069 ;
  assign n15075 = n15074 ^ n15073 ;
  assign n15077 = n15076 ^ n15075 ;
  assign n15067 = x98 & n6449 ;
  assign n15078 = n15077 ^ n15067 ;
  assign n15133 = n15132 ^ n15078 ;
  assign n15134 = n15133 ^ n14901 ;
  assign n15135 = n15134 ^ n14892 ;
  assign n15136 = n15135 ^ n15133 ;
  assign n15137 = ~n14893 & n15136 ;
  assign n15138 = n15137 ^ n15134 ;
  assign n15147 = n15146 ^ n15138 ;
  assign n15148 = n15147 ^ n14914 ;
  assign n15149 = n15148 ^ n14905 ;
  assign n15150 = n15149 ^ n15147 ;
  assign n15151 = ~n14906 & n15150 ;
  assign n15152 = n15151 ^ n15148 ;
  assign n15161 = n15160 ^ n15152 ;
  assign n15165 = n15164 ^ n15161 ;
  assign n15174 = n15173 ^ n15165 ;
  assign n15064 = n14938 ^ n14828 ;
  assign n15065 = ~n14930 & n15064 ;
  assign n15066 = n15065 ^ n14938 ;
  assign n15175 = n15174 ^ n15066 ;
  assign n15184 = n15183 ^ n15175 ;
  assign n15186 = n15184 ^ n14939 ;
  assign n15185 = n15184 ^ n14952 ;
  assign n15187 = n15186 ^ n15185 ;
  assign n15188 = n14944 & n15187 ;
  assign n15189 = n15188 ^ n15186 ;
  assign n15198 = n15197 ^ n15189 ;
  assign n15200 = n15198 ^ n14953 ;
  assign n15199 = n15198 ^ n14966 ;
  assign n15201 = n15200 ^ n15199 ;
  assign n15202 = ~n14958 & n15201 ;
  assign n15203 = n15202 ^ n15200 ;
  assign n15212 = n15211 ^ n15203 ;
  assign n15213 = n15212 ^ n14976 ;
  assign n15214 = n15213 ^ n15212 ;
  assign n15215 = n15214 ^ n14825 ;
  assign n15216 = ~n14968 & ~n15215 ;
  assign n15217 = n15216 ^ n15213 ;
  assign n15226 = n15225 ^ n15217 ;
  assign n15230 = n15229 ^ n15226 ;
  assign n15239 = n15238 ^ n15230 ;
  assign n15240 = n15239 ^ n14996 ;
  assign n15241 = n15240 ^ n15239 ;
  assign n15242 = n15241 ^ n14819 ;
  assign n15243 = n14988 & n15242 ;
  assign n15244 = n15243 ^ n15240 ;
  assign n15253 = n15252 ^ n15244 ;
  assign n15061 = n15018 ^ n14816 ;
  assign n15062 = n15012 & n15061 ;
  assign n15063 = n15062 ^ n15018 ;
  assign n15254 = n15253 ^ n15063 ;
  assign n15057 = n15010 ^ n14997 ;
  assign n15058 = ~n15002 & ~n15057 ;
  assign n15059 = n15058 ^ n14997 ;
  assign n15047 = x127 & n1339 ;
  assign n15048 = n15047 ^ n1337 ;
  assign n15053 = n1143 & n11285 ;
  assign n15054 = n15053 ^ n15047 ;
  assign n15055 = n15048 & ~n15054 ;
  assign n15056 = n15055 ^ x19 ;
  assign n15060 = n15059 ^ n15056 ;
  assign n15255 = n15254 ^ n15060 ;
  assign n15025 = n15020 ^ n15019 ;
  assign n15026 = n14808 ^ n14781 ;
  assign n15027 = ~n14782 & ~n15026 ;
  assign n15028 = n15027 ^ n14808 ;
  assign n15029 = n15021 ^ n14811 ;
  assign n15030 = ~n15019 & n15029 ;
  assign n15031 = n15028 & n15030 ;
  assign n15032 = n15031 ^ n15028 ;
  assign n15033 = ~n15021 & ~n15032 ;
  assign n15034 = n15025 & n15033 ;
  assign n15035 = n15034 ^ n15032 ;
  assign n15036 = n15035 ^ n15032 ;
  assign n15037 = n15019 ^ n14782 ;
  assign n15038 = n15037 ^ n15020 ;
  assign n15039 = n15038 ^ n15019 ;
  assign n15042 = n15029 & ~n15039 ;
  assign n15043 = n15042 ^ n15019 ;
  assign n15044 = ~n14808 & ~n15043 ;
  assign n15045 = n15036 & n15044 ;
  assign n15046 = n15045 ^ n15035 ;
  assign n15256 = n15255 ^ n15046 ;
  assign n15454 = n15056 ^ n15046 ;
  assign n15455 = n15060 & n15454 ;
  assign n15449 = n15252 ^ n15239 ;
  assign n15450 = ~n15244 & ~n15449 ;
  assign n15451 = n15450 ^ n15239 ;
  assign n15443 = x125 & n1665 ;
  assign n15442 = x127 & n1668 ;
  assign n15444 = n15443 ^ n15442 ;
  assign n15445 = n15444 ^ x23 ;
  assign n15441 = n1669 & n10986 ;
  assign n15446 = n15445 ^ n15441 ;
  assign n15440 = x126 & n1673 ;
  assign n15447 = n15446 ^ n15440 ;
  assign n15433 = x122 & n2032 ;
  assign n15432 = x124 & n2028 ;
  assign n15434 = n15433 ^ n15432 ;
  assign n15435 = n15434 ^ x26 ;
  assign n15431 = n2029 & n10117 ;
  assign n15436 = n15435 ^ n15431 ;
  assign n15430 = x123 & n2025 ;
  assign n15437 = n15436 ^ n15430 ;
  assign n15424 = x119 & n2593 ;
  assign n15423 = x121 & n2428 ;
  assign n15425 = n15424 ^ n15423 ;
  assign n15426 = n15425 ^ x29 ;
  assign n15422 = n2429 & n8979 ;
  assign n15427 = n15426 ^ n15422 ;
  assign n15421 = x120 & n2435 ;
  assign n15428 = n15427 ^ n15421 ;
  assign n15417 = n15225 ^ n15212 ;
  assign n15418 = ~n15217 & ~n15417 ;
  assign n15419 = n15418 ^ n15212 ;
  assign n15413 = n15211 ^ n15198 ;
  assign n15414 = ~n15203 & ~n15413 ;
  assign n15415 = n15414 ^ n15198 ;
  assign n15407 = x116 & n2890 ;
  assign n15406 = x118 & n2893 ;
  assign n15408 = n15407 ^ n15406 ;
  assign n15409 = n15408 ^ x32 ;
  assign n15405 = n2894 & ~n8140 ;
  assign n15410 = n15409 ^ n15405 ;
  assign n15404 = x117 & n2899 ;
  assign n15411 = n15410 ^ n15404 ;
  assign n15400 = n15197 ^ n15184 ;
  assign n15401 = ~n15189 & ~n15400 ;
  assign n15402 = n15401 ^ n15184 ;
  assign n15394 = x113 & n3387 ;
  assign n15393 = x115 & n3390 ;
  assign n15395 = n15394 ^ n15393 ;
  assign n15396 = n15395 ^ x35 ;
  assign n15392 = n3391 & ~n7353 ;
  assign n15397 = n15396 ^ n15392 ;
  assign n15391 = x114 & n3395 ;
  assign n15398 = n15397 ^ n15391 ;
  assign n15384 = x110 & n3932 ;
  assign n15383 = x112 & n3935 ;
  assign n15385 = n15384 ^ n15383 ;
  assign n15386 = n15385 ^ x38 ;
  assign n15382 = n3936 & ~n6616 ;
  assign n15387 = n15386 ^ n15382 ;
  assign n15381 = x111 & n3940 ;
  assign n15388 = n15387 ^ n15381 ;
  assign n15377 = n15173 ^ n15164 ;
  assign n15378 = n15165 & n15377 ;
  assign n15379 = n15378 ^ n15173 ;
  assign n15375 = x108 & n4475 ;
  assign n15370 = x107 & n4482 ;
  assign n15369 = x109 & n4478 ;
  assign n15371 = n15370 ^ n15369 ;
  assign n15372 = n15371 ^ x41 ;
  assign n15368 = n4479 & n5912 ;
  assign n15373 = n15372 ^ n15368 ;
  assign n15364 = n15160 ^ n15147 ;
  assign n15365 = ~n15152 & ~n15364 ;
  assign n15366 = n15365 ^ n15147 ;
  assign n15358 = x104 & n5113 ;
  assign n15357 = x106 & n5116 ;
  assign n15359 = n15358 ^ n15357 ;
  assign n15360 = n15359 ^ x44 ;
  assign n15356 = n5117 & ~n5257 ;
  assign n15361 = n15360 ^ n15356 ;
  assign n15355 = x105 & n5121 ;
  assign n15362 = n15361 ^ n15355 ;
  assign n15349 = x101 & n5981 ;
  assign n15348 = x103 & n5748 ;
  assign n15350 = n15349 ^ n15348 ;
  assign n15351 = n15350 ^ x47 ;
  assign n15347 = ~n4624 & n5749 ;
  assign n15352 = n15351 ^ n15347 ;
  assign n15346 = x102 & n5755 ;
  assign n15353 = n15352 ^ n15346 ;
  assign n15333 = x95 & n7183 ;
  assign n15332 = x97 & n7186 ;
  assign n15334 = n15333 ^ n15332 ;
  assign n15335 = n15334 ^ x53 ;
  assign n15331 = n3501 & n7187 ;
  assign n15336 = n15335 ^ n15331 ;
  assign n15330 = x96 & n7191 ;
  assign n15337 = n15336 ^ n15330 ;
  assign n15323 = x92 & n7954 ;
  assign n15322 = x94 & n7950 ;
  assign n15324 = n15323 ^ n15322 ;
  assign n15325 = n15324 ^ x56 ;
  assign n15321 = n3010 & n7951 ;
  assign n15326 = n15325 ^ n15321 ;
  assign n15320 = x93 & n7947 ;
  assign n15327 = n15326 ^ n15320 ;
  assign n15315 = ~n15099 & n15107 ;
  assign n15314 = x83 & n15097 ;
  assign n15316 = n15315 ^ n15314 ;
  assign n15317 = n15316 ^ n14849 ;
  assign n15307 = x86 & n9655 ;
  assign n15306 = x88 & n9651 ;
  assign n15308 = n15307 ^ n15306 ;
  assign n15309 = n15308 ^ x62 ;
  assign n15305 = n2131 & n9652 ;
  assign n15310 = n15309 ^ n15305 ;
  assign n15304 = x87 & n9648 ;
  assign n15311 = n15310 ^ n15304 ;
  assign n15312 = n15311 ^ x20 ;
  assign n15298 = x85 & n11895 ;
  assign n15299 = n15298 ^ n14848 ;
  assign n15300 = n15299 ^ n15095 ;
  assign n15301 = n15300 ^ x85 ;
  assign n15302 = n15301 ^ x84 ;
  assign n15303 = n12206 & n15302 ;
  assign n15313 = n15312 ^ n15303 ;
  assign n15318 = n15317 ^ n15313 ;
  assign n15295 = n15117 ^ n15094 ;
  assign n15296 = n15109 & n15295 ;
  assign n15288 = x89 & n8750 ;
  assign n15287 = x91 & n8746 ;
  assign n15289 = n15288 ^ n15287 ;
  assign n15290 = n15289 ^ x59 ;
  assign n15286 = n2548 & n8747 ;
  assign n15291 = n15290 ^ n15286 ;
  assign n15285 = x90 & n8743 ;
  assign n15292 = n15291 ^ n15285 ;
  assign n15293 = n15292 ^ n15117 ;
  assign n15297 = n15296 ^ n15293 ;
  assign n15319 = n15318 ^ n15297 ;
  assign n15328 = n15327 ^ n15319 ;
  assign n15282 = n15118 ^ n15086 ;
  assign n15283 = n15091 & ~n15282 ;
  assign n15284 = n15283 ^ n15086 ;
  assign n15329 = n15328 ^ n15284 ;
  assign n15338 = n15337 ^ n15329 ;
  assign n15279 = n15131 ^ n15119 ;
  assign n15280 = ~n15128 & ~n15279 ;
  assign n15281 = n15280 ^ n15119 ;
  assign n15339 = n15338 ^ n15281 ;
  assign n15269 = x98 & n6687 ;
  assign n15268 = x100 & n6444 ;
  assign n15270 = n15269 ^ n15268 ;
  assign n15271 = n15270 ^ x50 ;
  assign n15267 = n4048 & n6445 ;
  assign n15272 = n15271 ^ n15267 ;
  assign n15266 = x99 & n6449 ;
  assign n15273 = n15272 ^ n15266 ;
  assign n15274 = n15273 ^ n15132 ;
  assign n15275 = n15274 ^ n15072 ;
  assign n15276 = n15275 ^ n15273 ;
  assign n15277 = ~n15078 & ~n15276 ;
  assign n15278 = n15277 ^ n15274 ;
  assign n15340 = n15339 ^ n15278 ;
  assign n15342 = n15340 ^ n15133 ;
  assign n15341 = n15340 ^ n15146 ;
  assign n15343 = n15342 ^ n15341 ;
  assign n15344 = ~n15138 & ~n15343 ;
  assign n15345 = n15344 ^ n15342 ;
  assign n15354 = n15353 ^ n15345 ;
  assign n15363 = n15362 ^ n15354 ;
  assign n15367 = n15366 ^ n15363 ;
  assign n15374 = n15373 ^ n15367 ;
  assign n15376 = n15375 ^ n15374 ;
  assign n15380 = n15379 ^ n15376 ;
  assign n15389 = n15388 ^ n15380 ;
  assign n15263 = n15183 ^ n15066 ;
  assign n15264 = n15175 & n15263 ;
  assign n15265 = n15264 ^ n15183 ;
  assign n15390 = n15389 ^ n15265 ;
  assign n15399 = n15398 ^ n15390 ;
  assign n15403 = n15402 ^ n15399 ;
  assign n15412 = n15411 ^ n15403 ;
  assign n15416 = n15415 ^ n15412 ;
  assign n15420 = n15419 ^ n15416 ;
  assign n15429 = n15428 ^ n15420 ;
  assign n15438 = n15437 ^ n15429 ;
  assign n15260 = n15238 ^ n15229 ;
  assign n15261 = n15230 & n15260 ;
  assign n15262 = n15261 ^ n15238 ;
  assign n15439 = n15438 ^ n15262 ;
  assign n15448 = n15447 ^ n15439 ;
  assign n15452 = n15451 ^ n15448 ;
  assign n15257 = n15063 ^ n15060 ;
  assign n15258 = n15257 ^ n15046 ;
  assign n15259 = n15254 & n15258 ;
  assign n15453 = n15452 ^ n15259 ;
  assign n15456 = n15455 ^ n15453 ;
  assign n15680 = n1669 & n10155 ;
  assign n15679 = x126 & n1665 ;
  assign n15681 = n15680 ^ n15679 ;
  assign n15682 = n15681 ^ x23 ;
  assign n15678 = x127 & n1673 ;
  assign n15683 = n15682 ^ n15678 ;
  assign n15671 = x123 & n2032 ;
  assign n15670 = x125 & n2028 ;
  assign n15672 = n15671 ^ n15670 ;
  assign n15673 = n15672 ^ x26 ;
  assign n15669 = n2029 & n10416 ;
  assign n15674 = n15673 ^ n15669 ;
  assign n15668 = x124 & n2025 ;
  assign n15675 = n15674 ^ n15668 ;
  assign n15657 = x120 & n2593 ;
  assign n15656 = x122 & n2428 ;
  assign n15658 = n15657 ^ n15656 ;
  assign n15659 = n15658 ^ x29 ;
  assign n15655 = n2429 & ~n9261 ;
  assign n15660 = n15659 ^ n15655 ;
  assign n15654 = x121 & n2435 ;
  assign n15661 = n15660 ^ n15654 ;
  assign n15647 = x117 & n2890 ;
  assign n15646 = x119 & n2893 ;
  assign n15648 = n15647 ^ n15646 ;
  assign n15649 = n15648 ^ x32 ;
  assign n15645 = n2894 & n8405 ;
  assign n15650 = n15649 ^ n15645 ;
  assign n15644 = x118 & n2899 ;
  assign n15651 = n15650 ^ n15644 ;
  assign n15637 = x114 & n3387 ;
  assign n15636 = x116 & n3390 ;
  assign n15638 = n15637 ^ n15636 ;
  assign n15639 = n15638 ^ x35 ;
  assign n15635 = n3391 & ~n7604 ;
  assign n15640 = n15639 ^ n15635 ;
  assign n15634 = x115 & n3395 ;
  assign n15641 = n15640 ^ n15634 ;
  assign n15627 = x111 & n3932 ;
  assign n15626 = x113 & n3935 ;
  assign n15628 = n15627 ^ n15626 ;
  assign n15629 = n15628 ^ x38 ;
  assign n15625 = n3936 & ~n6849 ;
  assign n15630 = n15629 ^ n15625 ;
  assign n15624 = x112 & n3940 ;
  assign n15631 = n15630 ^ n15624 ;
  assign n15616 = x108 & n4482 ;
  assign n15615 = x110 & n4478 ;
  assign n15617 = n15616 ^ n15615 ;
  assign n15618 = n15617 ^ x41 ;
  assign n15614 = n4479 & n6145 ;
  assign n15619 = n15618 ^ n15614 ;
  assign n15613 = x109 & n4475 ;
  assign n15620 = n15619 ^ n15613 ;
  assign n15607 = x105 & n5113 ;
  assign n15606 = x107 & n5116 ;
  assign n15608 = n15607 ^ n15606 ;
  assign n15609 = n15608 ^ x44 ;
  assign n15605 = n5117 & ~n5459 ;
  assign n15610 = n15609 ^ n15605 ;
  assign n15604 = x106 & n5121 ;
  assign n15611 = n15610 ^ n15604 ;
  assign n15594 = n15337 ^ n15281 ;
  assign n15595 = ~n15338 & ~n15594 ;
  assign n15596 = n15595 ^ n15337 ;
  assign n15588 = x99 & n6687 ;
  assign n15587 = x101 & n6444 ;
  assign n15589 = n15588 ^ n15587 ;
  assign n15590 = n15589 ^ x50 ;
  assign n15586 = n4223 & n6445 ;
  assign n15591 = n15590 ^ n15586 ;
  assign n15585 = x100 & n6449 ;
  assign n15592 = n15591 ^ n15585 ;
  assign n15578 = x96 & n7183 ;
  assign n15577 = x98 & n7186 ;
  assign n15579 = n15578 ^ n15577 ;
  assign n15580 = n15579 ^ x53 ;
  assign n15576 = n3673 & n7187 ;
  assign n15581 = n15580 ^ n15576 ;
  assign n15575 = x97 & n7191 ;
  assign n15582 = n15581 ^ n15575 ;
  assign n15571 = n15318 ^ n15292 ;
  assign n15572 = n15297 & ~n15571 ;
  assign n15573 = n15572 ^ n15292 ;
  assign n15569 = x94 & n7947 ;
  assign n15564 = x93 & n7954 ;
  assign n15563 = x95 & n7950 ;
  assign n15565 = n15564 ^ n15563 ;
  assign n15566 = n15565 ^ x56 ;
  assign n15562 = n3166 & n7951 ;
  assign n15567 = n15566 ^ n15562 ;
  assign n15555 = x90 & n8750 ;
  assign n15554 = x92 & n8746 ;
  assign n15556 = n15555 ^ n15554 ;
  assign n15557 = n15556 ^ x59 ;
  assign n15553 = n2696 & n8747 ;
  assign n15558 = n15557 ^ n15553 ;
  assign n15552 = x91 & n8743 ;
  assign n15559 = n15558 ^ n15552 ;
  assign n15549 = x86 & n9956 ;
  assign n15550 = n15549 ^ n15298 ;
  assign n15546 = n2255 & n9652 ;
  assign n15544 = x87 & n9655 ;
  assign n15537 = x84 ^ x20 ;
  assign n15540 = n15302 & ~n15537 ;
  assign n15541 = n15540 ^ x84 ;
  assign n15542 = n12206 & n15541 ;
  assign n15535 = x89 & n9651 ;
  assign n15536 = n15535 ^ x62 ;
  assign n15543 = n15542 ^ n15536 ;
  assign n15545 = n15544 ^ n15543 ;
  assign n15547 = n15546 ^ n15545 ;
  assign n15534 = x88 & n9648 ;
  assign n15548 = n15547 ^ n15534 ;
  assign n15551 = n15550 ^ n15548 ;
  assign n15560 = n15559 ^ n15551 ;
  assign n15531 = n15317 ^ n15311 ;
  assign n15532 = n15313 & n15531 ;
  assign n15533 = n15532 ^ n15317 ;
  assign n15561 = n15560 ^ n15533 ;
  assign n15568 = n15567 ^ n15561 ;
  assign n15570 = n15569 ^ n15568 ;
  assign n15574 = n15573 ^ n15570 ;
  assign n15583 = n15582 ^ n15574 ;
  assign n15528 = n15327 ^ n15284 ;
  assign n15529 = ~n15328 & n15528 ;
  assign n15530 = n15529 ^ n15327 ;
  assign n15584 = n15583 ^ n15530 ;
  assign n15593 = n15592 ^ n15584 ;
  assign n15597 = n15596 ^ n15593 ;
  assign n15525 = ~n4830 & n5749 ;
  assign n15523 = x102 & n5981 ;
  assign n15519 = n15339 ^ n15273 ;
  assign n15520 = ~n15278 & n15519 ;
  assign n15521 = n15520 ^ n15273 ;
  assign n15517 = x104 & n5748 ;
  assign n15518 = n15517 ^ x47 ;
  assign n15522 = n15521 ^ n15518 ;
  assign n15524 = n15523 ^ n15522 ;
  assign n15526 = n15525 ^ n15524 ;
  assign n15516 = x103 & n5755 ;
  assign n15527 = n15526 ^ n15516 ;
  assign n15598 = n15597 ^ n15527 ;
  assign n15600 = n15598 ^ n15340 ;
  assign n15599 = n15598 ^ n15353 ;
  assign n15601 = n15600 ^ n15599 ;
  assign n15602 = n15345 & ~n15601 ;
  assign n15603 = n15602 ^ n15600 ;
  assign n15612 = n15611 ^ n15603 ;
  assign n15621 = n15620 ^ n15612 ;
  assign n15513 = n15366 ^ n15362 ;
  assign n15514 = ~n15363 & ~n15513 ;
  assign n15515 = n15514 ^ n15366 ;
  assign n15622 = n15621 ^ n15515 ;
  assign n15510 = n15379 ^ n15367 ;
  assign n15511 = ~n15376 & ~n15510 ;
  assign n15512 = n15511 ^ n15367 ;
  assign n15623 = n15622 ^ n15512 ;
  assign n15632 = n15631 ^ n15623 ;
  assign n15507 = n15380 ^ n15265 ;
  assign n15508 = ~n15389 & n15507 ;
  assign n15509 = n15508 ^ n15388 ;
  assign n15633 = n15632 ^ n15509 ;
  assign n15642 = n15641 ^ n15633 ;
  assign n15504 = n15402 ^ n15398 ;
  assign n15505 = n15399 & ~n15504 ;
  assign n15506 = n15505 ^ n15402 ;
  assign n15643 = n15642 ^ n15506 ;
  assign n15652 = n15651 ^ n15643 ;
  assign n15501 = n15415 ^ n15411 ;
  assign n15502 = ~n15412 & ~n15501 ;
  assign n15503 = n15502 ^ n15415 ;
  assign n15653 = n15652 ^ n15503 ;
  assign n15662 = n15661 ^ n15653 ;
  assign n15663 = n15662 ^ n15428 ;
  assign n15664 = n15663 ^ n15419 ;
  assign n15665 = n15664 ^ n15662 ;
  assign n15666 = ~n15420 & ~n15665 ;
  assign n15667 = n15666 ^ n15663 ;
  assign n15676 = n15675 ^ n15667 ;
  assign n15498 = n15437 ^ n15262 ;
  assign n15499 = n15438 & n15498 ;
  assign n15500 = n15499 ^ n15437 ;
  assign n15677 = n15676 ^ n15500 ;
  assign n15684 = n15683 ^ n15677 ;
  assign n15495 = n15451 ^ n15447 ;
  assign n15496 = ~n15448 & ~n15495 ;
  assign n15497 = n15496 ^ n15451 ;
  assign n15685 = n15684 ^ n15497 ;
  assign n15457 = n15452 ^ n15059 ;
  assign n15458 = n15457 ^ n15452 ;
  assign n15459 = n15452 ^ n15056 ;
  assign n15460 = n15459 ^ n15452 ;
  assign n15461 = n15458 & ~n15460 ;
  assign n15462 = n15461 ^ n15452 ;
  assign n15470 = n15460 ^ n15458 ;
  assign n15471 = n15470 ^ n15452 ;
  assign n15464 = n15452 ^ n15063 ;
  assign n15463 = n15452 ^ n15253 ;
  assign n15465 = n15464 ^ n15463 ;
  assign n15466 = n15463 ^ n15459 ;
  assign n15467 = n15466 ^ n15457 ;
  assign n15468 = n15467 ^ n15452 ;
  assign n15469 = n15465 & ~n15468 ;
  assign n15472 = n15471 ^ n15469 ;
  assign n15473 = n15462 & ~n15472 ;
  assign n15474 = n15473 ^ n15452 ;
  assign n15477 = n15253 ^ n15059 ;
  assign n15478 = n15477 ^ n15056 ;
  assign n15479 = n15478 ^ n15063 ;
  assign n15480 = n15479 ^ n15060 ;
  assign n15481 = n15480 ^ n15452 ;
  assign n15482 = n15060 & ~n15481 ;
  assign n15483 = n15479 ^ n15056 ;
  assign n15484 = ~n15482 & ~n15483 ;
  assign n15485 = n15484 ^ n15056 ;
  assign n15486 = n15485 ^ n15482 ;
  assign n15489 = n15464 & n15480 ;
  assign n15490 = ~n15486 & n15489 ;
  assign n15491 = n15490 ^ n15485 ;
  assign n15492 = n15046 & ~n15491 ;
  assign n15493 = ~n15474 & n15492 ;
  assign n15494 = n15493 ^ n15474 ;
  assign n15686 = n15685 ^ n15494 ;
  assign n15873 = x127 & n1664 ;
  assign n15874 = n15873 ^ n1662 ;
  assign n15879 = n1442 & n11285 ;
  assign n15880 = n15879 ^ n15873 ;
  assign n15881 = n15874 & ~n15880 ;
  assign n15882 = n15881 ^ x22 ;
  assign n15862 = x124 & n2032 ;
  assign n15861 = x126 & n2028 ;
  assign n15863 = n15862 ^ n15861 ;
  assign n15864 = n15863 ^ x26 ;
  assign n15860 = n2029 & n10461 ;
  assign n15865 = n15864 ^ n15860 ;
  assign n15859 = x125 & n2025 ;
  assign n15866 = n15865 ^ n15859 ;
  assign n15848 = x121 & n2593 ;
  assign n15847 = x123 & n2428 ;
  assign n15849 = n15848 ^ n15847 ;
  assign n15850 = n15849 ^ x29 ;
  assign n15846 = n2429 & ~n9804 ;
  assign n15851 = n15850 ^ n15846 ;
  assign n15845 = x122 & n2435 ;
  assign n15852 = n15851 ^ n15845 ;
  assign n15838 = x118 & n2890 ;
  assign n15837 = x120 & n2893 ;
  assign n15839 = n15838 ^ n15837 ;
  assign n15840 = n15839 ^ x32 ;
  assign n15836 = n2894 & n8904 ;
  assign n15841 = n15840 ^ n15836 ;
  assign n15835 = x119 & n2899 ;
  assign n15842 = n15841 ^ n15835 ;
  assign n15831 = n15641 ^ n15509 ;
  assign n15832 = ~n15633 & n15831 ;
  assign n15833 = n15832 ^ n15641 ;
  assign n15825 = x115 & n3387 ;
  assign n15824 = x117 & n3390 ;
  assign n15826 = n15825 ^ n15824 ;
  assign n15827 = n15826 ^ x35 ;
  assign n15823 = n3391 & ~n7860 ;
  assign n15828 = n15827 ^ n15823 ;
  assign n15822 = x116 & n3395 ;
  assign n15829 = n15828 ^ n15822 ;
  assign n15811 = x112 & n3932 ;
  assign n15810 = x114 & n3935 ;
  assign n15812 = n15811 ^ n15810 ;
  assign n15813 = n15812 ^ x38 ;
  assign n15809 = n3936 & ~n7108 ;
  assign n15814 = n15813 ^ n15809 ;
  assign n15808 = x113 & n3940 ;
  assign n15815 = n15814 ^ n15808 ;
  assign n15804 = n15620 ^ n15515 ;
  assign n15805 = n15621 & ~n15804 ;
  assign n15806 = n15805 ^ n15620 ;
  assign n15798 = x109 & n4482 ;
  assign n15797 = x111 & n4478 ;
  assign n15799 = n15798 ^ n15797 ;
  assign n15800 = n15799 ^ x41 ;
  assign n15796 = n4479 & ~n6370 ;
  assign n15801 = n15800 ^ n15796 ;
  assign n15795 = x110 & n4475 ;
  assign n15802 = n15801 ^ n15795 ;
  assign n15791 = n15611 ^ n15598 ;
  assign n15792 = n15603 & ~n15791 ;
  assign n15793 = n15792 ^ n15598 ;
  assign n15785 = x106 & n5113 ;
  assign n15784 = x108 & n5116 ;
  assign n15786 = n15785 ^ n15784 ;
  assign n15787 = n15786 ^ x44 ;
  assign n15783 = n5117 & n5687 ;
  assign n15788 = n15787 ^ n15783 ;
  assign n15782 = x107 & n5121 ;
  assign n15789 = n15788 ^ n15782 ;
  assign n15770 = x88 & n9655 ;
  assign n15769 = x90 & n9651 ;
  assign n15771 = n15770 ^ n15769 ;
  assign n15772 = n15771 ^ x62 ;
  assign n15768 = n2398 & n9652 ;
  assign n15773 = n15772 ^ n15768 ;
  assign n15767 = x89 & n9648 ;
  assign n15774 = n15773 ^ n15767 ;
  assign n15763 = x63 & n1616 ;
  assign n15764 = n15763 ^ n1732 ;
  assign n15765 = ~n9956 & n15764 ;
  assign n15766 = n15765 ^ n1732 ;
  assign n15775 = n15774 ^ n15766 ;
  assign n15756 = n2842 & n8747 ;
  assign n15754 = x91 & n8750 ;
  assign n15750 = n15550 ^ n15542 ;
  assign n15751 = ~n15548 & ~n15750 ;
  assign n15752 = n15751 ^ n15550 ;
  assign n15748 = x93 & n8746 ;
  assign n15749 = n15748 ^ x59 ;
  assign n15753 = n15752 ^ n15749 ;
  assign n15755 = n15754 ^ n15753 ;
  assign n15757 = n15756 ^ n15755 ;
  assign n15747 = x92 & n8743 ;
  assign n15758 = n15757 ^ n15747 ;
  assign n15776 = n15775 ^ n15758 ;
  assign n15745 = x95 & n7947 ;
  assign n15743 = n3336 & n7951 ;
  assign n15741 = x94 & n7954 ;
  assign n15737 = n15551 ^ n15533 ;
  assign n15738 = ~n15560 & n15737 ;
  assign n15739 = n15738 ^ n15559 ;
  assign n15735 = x96 & n7950 ;
  assign n15736 = n15735 ^ x56 ;
  assign n15740 = n15739 ^ n15736 ;
  assign n15742 = n15741 ^ n15740 ;
  assign n15744 = n15743 ^ n15742 ;
  assign n15746 = n15745 ^ n15744 ;
  assign n15777 = n15776 ^ n15746 ;
  assign n15733 = x98 & n7191 ;
  assign n15731 = n3851 & n7187 ;
  assign n15729 = x97 & n7183 ;
  assign n15725 = n15573 ^ n15561 ;
  assign n15726 = ~n15570 & ~n15725 ;
  assign n15727 = n15726 ^ n15561 ;
  assign n15723 = x99 & n7186 ;
  assign n15724 = n15723 ^ x53 ;
  assign n15728 = n15727 ^ n15724 ;
  assign n15730 = n15729 ^ n15728 ;
  assign n15732 = n15731 ^ n15730 ;
  assign n15734 = n15733 ^ n15732 ;
  assign n15778 = n15777 ^ n15734 ;
  assign n15720 = n4425 & n6445 ;
  assign n15718 = x100 & n6687 ;
  assign n15716 = x102 & n6444 ;
  assign n15712 = n15582 ^ n15530 ;
  assign n15713 = ~n15583 & n15712 ;
  assign n15714 = n15713 ^ n15582 ;
  assign n15715 = n15714 ^ x50 ;
  assign n15717 = n15716 ^ n15715 ;
  assign n15719 = n15718 ^ n15717 ;
  assign n15721 = n15720 ^ n15719 ;
  assign n15711 = x101 & n6449 ;
  assign n15722 = n15721 ^ n15711 ;
  assign n15779 = n15778 ^ n15722 ;
  assign n15708 = ~n5034 & n5749 ;
  assign n15706 = x103 & n5981 ;
  assign n15702 = n15596 ^ n15592 ;
  assign n15703 = n15593 & n15702 ;
  assign n15704 = n15703 ^ n15596 ;
  assign n15700 = x105 & n5748 ;
  assign n15701 = n15700 ^ x47 ;
  assign n15705 = n15704 ^ n15701 ;
  assign n15707 = n15706 ^ n15705 ;
  assign n15709 = n15708 ^ n15707 ;
  assign n15699 = x104 & n5755 ;
  assign n15710 = n15709 ^ n15699 ;
  assign n15780 = n15779 ^ n15710 ;
  assign n15696 = n15597 ^ n15521 ;
  assign n15697 = ~n15527 & ~n15696 ;
  assign n15698 = n15697 ^ n15597 ;
  assign n15781 = n15780 ^ n15698 ;
  assign n15790 = n15789 ^ n15781 ;
  assign n15794 = n15793 ^ n15790 ;
  assign n15803 = n15802 ^ n15794 ;
  assign n15807 = n15806 ^ n15803 ;
  assign n15816 = n15815 ^ n15807 ;
  assign n15817 = n15816 ^ n15631 ;
  assign n15818 = n15817 ^ n15816 ;
  assign n15819 = n15818 ^ n15512 ;
  assign n15820 = ~n15623 & ~n15819 ;
  assign n15821 = n15820 ^ n15817 ;
  assign n15830 = n15829 ^ n15821 ;
  assign n15834 = n15833 ^ n15830 ;
  assign n15843 = n15842 ^ n15834 ;
  assign n15693 = n15651 ^ n15506 ;
  assign n15694 = n15643 & ~n15693 ;
  assign n15695 = n15694 ^ n15651 ;
  assign n15844 = n15843 ^ n15695 ;
  assign n15853 = n15852 ^ n15844 ;
  assign n15854 = n15853 ^ n15661 ;
  assign n15855 = n15854 ^ n15853 ;
  assign n15856 = n15855 ^ n15503 ;
  assign n15857 = ~n15653 & ~n15856 ;
  assign n15858 = n15857 ^ n15854 ;
  assign n15867 = n15866 ^ n15858 ;
  assign n15869 = n15867 ^ n15662 ;
  assign n15868 = n15867 ^ n15675 ;
  assign n15870 = n15869 ^ n15868 ;
  assign n15871 = n15667 & n15870 ;
  assign n15872 = n15871 ^ n15869 ;
  assign n15883 = n15882 ^ n15872 ;
  assign n15690 = n15683 ^ n15500 ;
  assign n15691 = ~n15677 & n15690 ;
  assign n15692 = n15691 ^ n15683 ;
  assign n15884 = n15883 ^ n15692 ;
  assign n15687 = n15497 ^ n15494 ;
  assign n15688 = n15685 & n15687 ;
  assign n15689 = n15688 ^ n15494 ;
  assign n15885 = n15884 ^ n15689 ;
  assign n16067 = n15882 ^ n15867 ;
  assign n16068 = ~n15872 & ~n16067 ;
  assign n16069 = n16068 ^ n15867 ;
  assign n16063 = n15866 ^ n15853 ;
  assign n16064 = ~n15858 & ~n16063 ;
  assign n16065 = n16064 ^ n15853 ;
  assign n16057 = x125 & n2032 ;
  assign n16056 = x127 & n2028 ;
  assign n16058 = n16057 ^ n16056 ;
  assign n16059 = n16058 ^ x26 ;
  assign n16055 = n2029 & n10986 ;
  assign n16060 = n16059 ^ n16055 ;
  assign n16054 = x126 & n2025 ;
  assign n16061 = n16060 ^ n16054 ;
  assign n16047 = x122 & n2593 ;
  assign n16046 = x124 & n2428 ;
  assign n16048 = n16047 ^ n16046 ;
  assign n16049 = n16048 ^ x29 ;
  assign n16045 = n2429 & n10117 ;
  assign n16050 = n16049 ^ n16045 ;
  assign n16044 = x123 & n2435 ;
  assign n16051 = n16050 ^ n16044 ;
  assign n16038 = x119 & n2890 ;
  assign n16037 = x121 & n2893 ;
  assign n16039 = n16038 ^ n16037 ;
  assign n16040 = n16039 ^ x32 ;
  assign n16036 = n2894 & n8979 ;
  assign n16041 = n16040 ^ n16036 ;
  assign n16035 = x120 & n2899 ;
  assign n16042 = n16041 ^ n16035 ;
  assign n16026 = n15829 ^ n15816 ;
  assign n16027 = ~n15821 & ~n16026 ;
  assign n16028 = n16027 ^ n15816 ;
  assign n16020 = x116 & n3387 ;
  assign n16019 = x118 & n3390 ;
  assign n16021 = n16020 ^ n16019 ;
  assign n16022 = n16021 ^ x35 ;
  assign n16018 = n3391 & ~n8140 ;
  assign n16023 = n16022 ^ n16018 ;
  assign n16017 = x117 & n3395 ;
  assign n16024 = n16023 ^ n16017 ;
  assign n16010 = x113 & n3932 ;
  assign n16009 = x115 & n3935 ;
  assign n16011 = n16010 ^ n16009 ;
  assign n16012 = n16011 ^ x38 ;
  assign n16008 = n3936 & ~n7353 ;
  assign n16013 = n16012 ^ n16008 ;
  assign n16007 = x114 & n3940 ;
  assign n16014 = n16013 ^ n16007 ;
  assign n16003 = n15802 ^ n15793 ;
  assign n16004 = n15794 & ~n16003 ;
  assign n16005 = n16004 ^ n15802 ;
  assign n16001 = x111 & n4475 ;
  assign n15996 = x110 & n4482 ;
  assign n15995 = x112 & n4478 ;
  assign n15997 = n15996 ^ n15995 ;
  assign n15998 = n15997 ^ x41 ;
  assign n15994 = n4479 & ~n6616 ;
  assign n15999 = n15998 ^ n15994 ;
  assign n15990 = n15789 ^ n15698 ;
  assign n15991 = ~n15781 & ~n15990 ;
  assign n15992 = n15991 ^ n15789 ;
  assign n15988 = x108 & n5121 ;
  assign n15983 = x107 & n5113 ;
  assign n15982 = x109 & n5116 ;
  assign n15984 = n15983 ^ n15982 ;
  assign n15985 = n15984 ^ x44 ;
  assign n15981 = n5117 & n5912 ;
  assign n15986 = n15985 ^ n15981 ;
  assign n15975 = x104 & n5981 ;
  assign n15974 = x106 & n5748 ;
  assign n15976 = n15975 ^ n15974 ;
  assign n15977 = n15976 ^ x47 ;
  assign n15973 = ~n5257 & n5749 ;
  assign n15978 = n15977 ^ n15973 ;
  assign n15972 = x105 & n5755 ;
  assign n15979 = n15978 ^ n15972 ;
  assign n15968 = n15779 ^ n15704 ;
  assign n15969 = ~n15710 & ~n15968 ;
  assign n15970 = n15969 ^ n15779 ;
  assign n15963 = x96 & n7947 ;
  assign n15950 = x89 & n9655 ;
  assign n15949 = x91 & n9651 ;
  assign n15951 = n15950 ^ n15949 ;
  assign n15952 = n15951 ^ x62 ;
  assign n15948 = n2548 & n9652 ;
  assign n15953 = n15952 ^ n15948 ;
  assign n15947 = x90 & n9648 ;
  assign n15954 = n15953 ^ n15947 ;
  assign n15955 = n15954 ^ x23 ;
  assign n15943 = x88 ^ x86 ;
  assign n15944 = ~n11895 & n15943 ;
  assign n15945 = n15944 ^ n1732 ;
  assign n15946 = n12206 & n15945 ;
  assign n15956 = n15955 ^ n15946 ;
  assign n15939 = n15774 ^ n9956 ;
  assign n15940 = n15939 ^ x86 ;
  assign n15941 = n15766 & ~n15940 ;
  assign n15942 = n15941 ^ n15774 ;
  assign n15957 = n15956 ^ n15942 ;
  assign n15929 = x92 & n8750 ;
  assign n15928 = x94 & n8746 ;
  assign n15930 = n15929 ^ n15928 ;
  assign n15931 = n15930 ^ x59 ;
  assign n15927 = n3010 & n8747 ;
  assign n15932 = n15931 ^ n15927 ;
  assign n15926 = x93 & n8743 ;
  assign n15933 = n15932 ^ n15926 ;
  assign n15934 = n15933 ^ n15775 ;
  assign n15935 = n15934 ^ n15752 ;
  assign n15936 = n15935 ^ n15933 ;
  assign n15937 = n15758 & n15936 ;
  assign n15938 = n15937 ^ n15934 ;
  assign n15958 = n15957 ^ n15938 ;
  assign n15959 = n15958 ^ x56 ;
  assign n15925 = x95 & n7954 ;
  assign n15960 = n15959 ^ n15925 ;
  assign n15924 = x97 & n7950 ;
  assign n15961 = n15960 ^ n15924 ;
  assign n15923 = n3501 & n7951 ;
  assign n15962 = n15961 ^ n15923 ;
  assign n15964 = n15963 ^ n15962 ;
  assign n15920 = n15776 ^ n15739 ;
  assign n15921 = ~n15746 & n15920 ;
  assign n15922 = n15921 ^ n15776 ;
  assign n15965 = n15964 ^ n15922 ;
  assign n15910 = x98 & n7183 ;
  assign n15909 = x100 & n7186 ;
  assign n15911 = n15910 ^ n15909 ;
  assign n15912 = n15911 ^ x53 ;
  assign n15908 = n4048 & n7187 ;
  assign n15913 = n15912 ^ n15908 ;
  assign n15907 = x99 & n7191 ;
  assign n15914 = n15913 ^ n15907 ;
  assign n15916 = n15914 ^ n15777 ;
  assign n15915 = n15914 ^ n15727 ;
  assign n15917 = n15916 ^ n15915 ;
  assign n15918 = n15734 & ~n15917 ;
  assign n15919 = n15918 ^ n15916 ;
  assign n15966 = n15965 ^ n15919 ;
  assign n15904 = ~n4624 & n6445 ;
  assign n15902 = x101 & n6687 ;
  assign n15898 = n15778 ^ n15714 ;
  assign n15899 = ~n15722 & ~n15898 ;
  assign n15900 = n15899 ^ n15778 ;
  assign n15896 = x103 & n6444 ;
  assign n15897 = n15896 ^ x50 ;
  assign n15901 = n15900 ^ n15897 ;
  assign n15903 = n15902 ^ n15901 ;
  assign n15905 = n15904 ^ n15903 ;
  assign n15895 = x102 & n6449 ;
  assign n15906 = n15905 ^ n15895 ;
  assign n15967 = n15966 ^ n15906 ;
  assign n15971 = n15970 ^ n15967 ;
  assign n15980 = n15979 ^ n15971 ;
  assign n15987 = n15986 ^ n15980 ;
  assign n15989 = n15988 ^ n15987 ;
  assign n15993 = n15992 ^ n15989 ;
  assign n16000 = n15999 ^ n15993 ;
  assign n16002 = n16001 ^ n16000 ;
  assign n16006 = n16005 ^ n16002 ;
  assign n16015 = n16014 ^ n16006 ;
  assign n15892 = n15815 ^ n15806 ;
  assign n15893 = n15807 & n15892 ;
  assign n15894 = n15893 ^ n15815 ;
  assign n16016 = n16015 ^ n15894 ;
  assign n16025 = n16024 ^ n16016 ;
  assign n16029 = n16028 ^ n16025 ;
  assign n16030 = n16029 ^ n15842 ;
  assign n16031 = n16030 ^ n15833 ;
  assign n16032 = n16031 ^ n16029 ;
  assign n16033 = n15834 & n16032 ;
  assign n16034 = n16033 ^ n16030 ;
  assign n16043 = n16042 ^ n16034 ;
  assign n16052 = n16051 ^ n16043 ;
  assign n15889 = n15852 ^ n15695 ;
  assign n15890 = n15844 & n15889 ;
  assign n15891 = n15890 ^ n15852 ;
  assign n16053 = n16052 ^ n15891 ;
  assign n16062 = n16061 ^ n16053 ;
  assign n16066 = n16065 ^ n16062 ;
  assign n16070 = n16069 ^ n16066 ;
  assign n15886 = n15692 ^ n15689 ;
  assign n15887 = ~n15884 & ~n15886 ;
  assign n15888 = n15887 ^ n15692 ;
  assign n16071 = n16070 ^ n15888 ;
  assign n16252 = n16061 & ~n16065 ;
  assign n16251 = n16065 ^ n16061 ;
  assign n16253 = n16252 ^ n16251 ;
  assign n16246 = n2029 & n10155 ;
  assign n16245 = x126 & n2032 ;
  assign n16247 = n16246 ^ n16245 ;
  assign n16248 = n16247 ^ x26 ;
  assign n16244 = x127 & n2025 ;
  assign n16249 = n16248 ^ n16244 ;
  assign n16237 = x123 & n2593 ;
  assign n16236 = x125 & n2428 ;
  assign n16238 = n16237 ^ n16236 ;
  assign n16239 = n16238 ^ x29 ;
  assign n16235 = n2429 & n10416 ;
  assign n16240 = n16239 ^ n16235 ;
  assign n16234 = x124 & n2435 ;
  assign n16241 = n16240 ^ n16234 ;
  assign n16223 = x120 & n2890 ;
  assign n16222 = x122 & n2893 ;
  assign n16224 = n16223 ^ n16222 ;
  assign n16225 = n16224 ^ x32 ;
  assign n16221 = n2894 & ~n9261 ;
  assign n16226 = n16225 ^ n16221 ;
  assign n16220 = x121 & n2899 ;
  assign n16227 = n16226 ^ n16220 ;
  assign n16212 = x114 & n3932 ;
  assign n16211 = x116 & n3935 ;
  assign n16213 = n16212 ^ n16211 ;
  assign n16214 = n16213 ^ x38 ;
  assign n16210 = n3936 & ~n7604 ;
  assign n16215 = n16214 ^ n16210 ;
  assign n16209 = x115 & n3940 ;
  assign n16216 = n16215 ^ n16209 ;
  assign n16202 = x111 & n4482 ;
  assign n16201 = x113 & n4478 ;
  assign n16203 = n16202 ^ n16201 ;
  assign n16204 = n16203 ^ x41 ;
  assign n16200 = n4479 & ~n6849 ;
  assign n16205 = n16204 ^ n16200 ;
  assign n16199 = x112 & n4475 ;
  assign n16206 = n16205 ^ n16199 ;
  assign n16191 = x108 & n5113 ;
  assign n16190 = x110 & n5116 ;
  assign n16192 = n16191 ^ n16190 ;
  assign n16193 = n16192 ^ x44 ;
  assign n16189 = n5117 & n6145 ;
  assign n16194 = n16193 ^ n16189 ;
  assign n16188 = x109 & n5121 ;
  assign n16195 = n16194 ^ n16188 ;
  assign n16182 = x105 & n5981 ;
  assign n16181 = x107 & n5748 ;
  assign n16183 = n16182 ^ n16181 ;
  assign n16184 = n16183 ^ x47 ;
  assign n16180 = ~n5459 & n5749 ;
  assign n16185 = n16184 ^ n16180 ;
  assign n16179 = x106 & n5755 ;
  assign n16186 = n16185 ^ n16179 ;
  assign n16169 = x97 & n7947 ;
  assign n16167 = n3673 & n7951 ;
  assign n16163 = x96 & n7954 ;
  assign n16162 = x98 & n7950 ;
  assign n16164 = n16163 ^ n16162 ;
  assign n16165 = n16164 ^ x56 ;
  assign n16159 = x94 & n8743 ;
  assign n16157 = n3166 & n8747 ;
  assign n16153 = x93 & n8750 ;
  assign n16152 = x95 & n8746 ;
  assign n16154 = n16153 ^ n16152 ;
  assign n16155 = n16154 ^ x59 ;
  assign n16146 = x90 & n9655 ;
  assign n16145 = x92 & n9651 ;
  assign n16147 = n16146 ^ n16145 ;
  assign n16148 = n16147 ^ x62 ;
  assign n16144 = n2696 & n9652 ;
  assign n16149 = n16148 ^ n16144 ;
  assign n16143 = x91 & n9648 ;
  assign n16150 = n16149 ^ n16143 ;
  assign n16140 = x88 & n11895 ;
  assign n16134 = x87 ^ x23 ;
  assign n16137 = n15945 & ~n16134 ;
  assign n16138 = n16137 ^ x87 ;
  assign n16139 = n12206 & n16138 ;
  assign n16141 = n16140 ^ n16139 ;
  assign n16133 = x89 & n9956 ;
  assign n16142 = n16141 ^ n16133 ;
  assign n16151 = n16150 ^ n16142 ;
  assign n16156 = n16155 ^ n16151 ;
  assign n16158 = n16157 ^ n16156 ;
  assign n16160 = n16159 ^ n16158 ;
  assign n16130 = n15954 ^ n15942 ;
  assign n16131 = ~n15956 & n16130 ;
  assign n16132 = n16131 ^ n15954 ;
  assign n16161 = n16160 ^ n16132 ;
  assign n16166 = n16165 ^ n16161 ;
  assign n16168 = n16167 ^ n16166 ;
  assign n16170 = n16169 ^ n16168 ;
  assign n16127 = n15957 ^ n15933 ;
  assign n16128 = ~n15938 & ~n16127 ;
  assign n16129 = n16128 ^ n15933 ;
  assign n16171 = n16170 ^ n16129 ;
  assign n16124 = n4223 & n7187 ;
  assign n16122 = x99 & n7183 ;
  assign n16118 = n15958 ^ n15922 ;
  assign n16119 = n15964 & n16118 ;
  assign n16120 = n16119 ^ n15958 ;
  assign n16116 = x101 & n7186 ;
  assign n16117 = n16116 ^ x53 ;
  assign n16121 = n16120 ^ n16117 ;
  assign n16123 = n16122 ^ n16121 ;
  assign n16125 = n16124 ^ n16123 ;
  assign n16115 = x100 & n7191 ;
  assign n16126 = n16125 ^ n16115 ;
  assign n16172 = n16171 ^ n16126 ;
  assign n16112 = ~n4830 & n6445 ;
  assign n16110 = x102 & n6687 ;
  assign n16106 = n15965 ^ n15914 ;
  assign n16107 = n15919 & n16106 ;
  assign n16108 = n16107 ^ n15914 ;
  assign n16104 = x104 & n6444 ;
  assign n16105 = n16104 ^ x50 ;
  assign n16109 = n16108 ^ n16105 ;
  assign n16111 = n16110 ^ n16109 ;
  assign n16113 = n16112 ^ n16111 ;
  assign n16103 = x103 & n6449 ;
  assign n16114 = n16113 ^ n16103 ;
  assign n16173 = n16172 ^ n16114 ;
  assign n16174 = n16173 ^ n15966 ;
  assign n16175 = n16174 ^ n15900 ;
  assign n16176 = n16175 ^ n16173 ;
  assign n16177 = n15906 & ~n16176 ;
  assign n16178 = n16177 ^ n16174 ;
  assign n16187 = n16186 ^ n16178 ;
  assign n16196 = n16195 ^ n16187 ;
  assign n16100 = n15979 ^ n15970 ;
  assign n16101 = ~n15971 & ~n16100 ;
  assign n16102 = n16101 ^ n15979 ;
  assign n16197 = n16196 ^ n16102 ;
  assign n16097 = n15992 ^ n15980 ;
  assign n16098 = n15989 & n16097 ;
  assign n16099 = n16098 ^ n15980 ;
  assign n16198 = n16197 ^ n16099 ;
  assign n16207 = n16206 ^ n16198 ;
  assign n16094 = n16005 ^ n15993 ;
  assign n16095 = n16002 & n16094 ;
  assign n16096 = n16095 ^ n15993 ;
  assign n16208 = n16207 ^ n16096 ;
  assign n16217 = n16216 ^ n16208 ;
  assign n16084 = x117 & n3387 ;
  assign n16083 = x119 & n3390 ;
  assign n16085 = n16084 ^ n16083 ;
  assign n16086 = n16085 ^ x35 ;
  assign n16082 = n3391 & n8405 ;
  assign n16087 = n16086 ^ n16082 ;
  assign n16081 = x118 & n3395 ;
  assign n16088 = n16087 ^ n16081 ;
  assign n16089 = n16088 ^ n16014 ;
  assign n16090 = n16089 ^ n15894 ;
  assign n16091 = n16090 ^ n16088 ;
  assign n16092 = n16015 & n16091 ;
  assign n16093 = n16092 ^ n16089 ;
  assign n16218 = n16217 ^ n16093 ;
  assign n16078 = n16028 ^ n16024 ;
  assign n16079 = ~n16025 & ~n16078 ;
  assign n16080 = n16079 ^ n16028 ;
  assign n16219 = n16218 ^ n16080 ;
  assign n16228 = n16227 ^ n16219 ;
  assign n16230 = n16228 ^ n16029 ;
  assign n16229 = n16228 ^ n16042 ;
  assign n16231 = n16230 ^ n16229 ;
  assign n16232 = ~n16034 & ~n16231 ;
  assign n16233 = n16232 ^ n16230 ;
  assign n16242 = n16241 ^ n16233 ;
  assign n16075 = n16051 ^ n15891 ;
  assign n16076 = ~n16052 & n16075 ;
  assign n16077 = n16076 ^ n16051 ;
  assign n16243 = n16242 ^ n16077 ;
  assign n16250 = n16249 ^ n16243 ;
  assign n16254 = n16253 ^ n16250 ;
  assign n16073 = n16066 ^ n15888 ;
  assign n16074 = ~n16070 & n16073 ;
  assign n16255 = n16254 ^ n16074 ;
  assign n16072 = ~n16053 & n16066 ;
  assign n16256 = n16255 ^ n16072 ;
  assign n16431 = n16053 & n16069 ;
  assign n16432 = n16431 ^ n16250 ;
  assign n16430 = n16069 ^ n16053 ;
  assign n16433 = n16432 ^ n16430 ;
  assign n16434 = ~n16253 & n16433 ;
  assign n16435 = n15888 & n16434 ;
  assign n16436 = n16431 ^ n16061 ;
  assign n16437 = ~n16251 & ~n16436 ;
  assign n16438 = n16437 ^ n16061 ;
  assign n16439 = ~n16250 & n16438 ;
  assign n16440 = ~n16435 & ~n16439 ;
  assign n16441 = n16252 ^ n16250 ;
  assign n16442 = n16053 ^ n15888 ;
  assign n16443 = n16430 & ~n16442 ;
  assign n16444 = n16443 ^ n16053 ;
  assign n16445 = ~n16441 & ~n16444 ;
  assign n16446 = n16440 & ~n16445 ;
  assign n16425 = n16241 ^ n16228 ;
  assign n16426 = ~n16233 & n16425 ;
  assign n16427 = n16426 ^ n16228 ;
  assign n16418 = x124 & n2593 ;
  assign n16417 = x126 & n2428 ;
  assign n16419 = n16418 ^ n16417 ;
  assign n16420 = n16419 ^ x29 ;
  assign n16416 = n2429 & n10461 ;
  assign n16421 = n16420 ^ n16416 ;
  assign n16415 = x125 & n2435 ;
  assign n16422 = n16421 ^ n16415 ;
  assign n16408 = x121 & n2890 ;
  assign n16407 = x123 & n2893 ;
  assign n16409 = n16408 ^ n16407 ;
  assign n16410 = n16409 ^ x32 ;
  assign n16406 = n2894 & ~n9804 ;
  assign n16411 = n16410 ^ n16406 ;
  assign n16405 = x122 & n2899 ;
  assign n16412 = n16411 ^ n16405 ;
  assign n16398 = x118 & n3387 ;
  assign n16397 = x120 & n3390 ;
  assign n16399 = n16398 ^ n16397 ;
  assign n16400 = n16399 ^ x35 ;
  assign n16396 = n3391 & n8904 ;
  assign n16401 = n16400 ^ n16396 ;
  assign n16395 = x119 & n3395 ;
  assign n16402 = n16401 ^ n16395 ;
  assign n16391 = n16216 ^ n16096 ;
  assign n16392 = n16208 & n16391 ;
  assign n16393 = n16392 ^ n16216 ;
  assign n16385 = x115 & n3932 ;
  assign n16384 = x117 & n3935 ;
  assign n16386 = n16385 ^ n16384 ;
  assign n16387 = n16386 ^ x38 ;
  assign n16383 = n3936 & ~n7860 ;
  assign n16388 = n16387 ^ n16383 ;
  assign n16382 = x116 & n3940 ;
  assign n16389 = n16388 ^ n16382 ;
  assign n16371 = x112 & n4482 ;
  assign n16370 = x114 & n4478 ;
  assign n16372 = n16371 ^ n16370 ;
  assign n16373 = n16372 ^ x41 ;
  assign n16369 = n4479 & ~n7108 ;
  assign n16374 = n16373 ^ n16369 ;
  assign n16368 = x113 & n4475 ;
  assign n16375 = n16374 ^ n16368 ;
  assign n16365 = n16195 ^ n16102 ;
  assign n16366 = ~n16196 & n16365 ;
  assign n16357 = x109 & n5113 ;
  assign n16356 = x111 & n5116 ;
  assign n16358 = n16357 ^ n16356 ;
  assign n16359 = n16358 ^ x44 ;
  assign n16355 = n5117 & ~n6370 ;
  assign n16360 = n16359 ^ n16355 ;
  assign n16354 = x110 & n5121 ;
  assign n16361 = n16360 ^ n16354 ;
  assign n16350 = n16186 ^ n16173 ;
  assign n16351 = ~n16178 & ~n16350 ;
  assign n16352 = n16351 ^ n16173 ;
  assign n16343 = x106 & n5981 ;
  assign n16342 = x108 & n5748 ;
  assign n16344 = n16343 ^ n16342 ;
  assign n16345 = n16344 ^ x47 ;
  assign n16341 = n5687 & n5749 ;
  assign n16346 = n16345 ^ n16341 ;
  assign n16340 = x107 & n5755 ;
  assign n16347 = n16346 ^ n16340 ;
  assign n16334 = x103 & n6687 ;
  assign n16333 = x105 & n6444 ;
  assign n16335 = n16334 ^ n16333 ;
  assign n16336 = n16335 ^ x50 ;
  assign n16332 = ~n5034 & n6445 ;
  assign n16337 = n16336 ^ n16332 ;
  assign n16331 = x104 & n6449 ;
  assign n16338 = n16337 ^ n16331 ;
  assign n16328 = n16171 ^ n16120 ;
  assign n16329 = ~n16126 & ~n16328 ;
  assign n16319 = x100 & n7183 ;
  assign n16318 = x102 & n7186 ;
  assign n16320 = n16319 ^ n16318 ;
  assign n16321 = n16320 ^ x53 ;
  assign n16317 = n4425 & n7187 ;
  assign n16322 = n16321 ^ n16317 ;
  assign n16316 = x101 & n7191 ;
  assign n16323 = n16322 ^ n16316 ;
  assign n16312 = n16151 ^ n16132 ;
  assign n16313 = ~n16160 & ~n16312 ;
  assign n16314 = n16313 ^ n16151 ;
  assign n16306 = x97 & n7954 ;
  assign n16305 = x99 & n7950 ;
  assign n16307 = n16306 ^ n16305 ;
  assign n16308 = n16307 ^ x56 ;
  assign n16304 = n3851 & n7951 ;
  assign n16309 = n16308 ^ n16304 ;
  assign n16303 = x98 & n7947 ;
  assign n16310 = n16309 ^ n16303 ;
  assign n16297 = x94 & n8750 ;
  assign n16296 = x96 & n8746 ;
  assign n16298 = n16297 ^ n16296 ;
  assign n16299 = n16298 ^ x59 ;
  assign n16295 = n3336 & n8747 ;
  assign n16300 = n16299 ^ n16295 ;
  assign n16294 = x95 & n8743 ;
  assign n16301 = n16300 ^ n16294 ;
  assign n16287 = x91 & n9655 ;
  assign n16286 = x93 & n9651 ;
  assign n16288 = n16287 ^ n16286 ;
  assign n16289 = n16288 ^ x62 ;
  assign n16285 = n2842 & n9652 ;
  assign n16290 = n16289 ^ n16285 ;
  assign n16284 = x92 & n9648 ;
  assign n16291 = n16290 ^ n16284 ;
  assign n16280 = ~x90 & n9956 ;
  assign n16281 = n16280 ^ n16140 ;
  assign n16282 = n16281 ^ n9956 ;
  assign n16279 = x89 & n12206 ;
  assign n16283 = n16282 ^ n16279 ;
  assign n16292 = n16291 ^ n16283 ;
  assign n16276 = n16150 ^ n16139 ;
  assign n16277 = n16142 & n16276 ;
  assign n16278 = n16277 ^ n16150 ;
  assign n16293 = n16292 ^ n16278 ;
  assign n16302 = n16301 ^ n16293 ;
  assign n16311 = n16310 ^ n16302 ;
  assign n16315 = n16314 ^ n16311 ;
  assign n16324 = n16323 ^ n16315 ;
  assign n16273 = n16161 ^ n16129 ;
  assign n16274 = ~n16170 & ~n16273 ;
  assign n16275 = n16274 ^ n16161 ;
  assign n16325 = n16324 ^ n16275 ;
  assign n16326 = n16325 ^ n16171 ;
  assign n16330 = n16329 ^ n16326 ;
  assign n16339 = n16338 ^ n16330 ;
  assign n16348 = n16347 ^ n16339 ;
  assign n16270 = n16172 ^ n16108 ;
  assign n16271 = ~n16114 & ~n16270 ;
  assign n16272 = n16271 ^ n16172 ;
  assign n16349 = n16348 ^ n16272 ;
  assign n16353 = n16352 ^ n16349 ;
  assign n16362 = n16361 ^ n16353 ;
  assign n16363 = n16362 ^ n16195 ;
  assign n16367 = n16366 ^ n16363 ;
  assign n16376 = n16375 ^ n16367 ;
  assign n16377 = n16376 ^ n16206 ;
  assign n16378 = n16377 ^ n16376 ;
  assign n16379 = n16378 ^ n16099 ;
  assign n16380 = n16198 & n16379 ;
  assign n16381 = n16380 ^ n16377 ;
  assign n16390 = n16389 ^ n16381 ;
  assign n16394 = n16393 ^ n16390 ;
  assign n16403 = n16402 ^ n16394 ;
  assign n16267 = n16217 ^ n16088 ;
  assign n16268 = n16093 & ~n16267 ;
  assign n16269 = n16268 ^ n16088 ;
  assign n16404 = n16403 ^ n16269 ;
  assign n16413 = n16412 ^ n16404 ;
  assign n16264 = n16227 ^ n16080 ;
  assign n16265 = ~n16219 & ~n16264 ;
  assign n16266 = n16265 ^ n16227 ;
  assign n16414 = n16413 ^ n16266 ;
  assign n16423 = n16422 ^ n16414 ;
  assign n2033 = n2032 ^ n2029 ;
  assign n16261 = x127 & n2033 ;
  assign n16260 = n2029 & n10154 ;
  assign n16262 = n16261 ^ n16260 ;
  assign n16263 = n16262 ^ x26 ;
  assign n16424 = n16423 ^ n16263 ;
  assign n16428 = n16427 ^ n16424 ;
  assign n16257 = n16249 ^ n16077 ;
  assign n16258 = n16243 & n16257 ;
  assign n16259 = n16258 ^ n16249 ;
  assign n16429 = n16428 ^ n16259 ;
  assign n16447 = n16446 ^ n16429 ;
  assign n16614 = x125 & n2593 ;
  assign n16613 = x127 & n2428 ;
  assign n16615 = n16614 ^ n16613 ;
  assign n16616 = n16615 ^ x29 ;
  assign n16612 = n2429 & n10986 ;
  assign n16617 = n16616 ^ n16612 ;
  assign n16611 = x126 & n2435 ;
  assign n16618 = n16617 ^ n16611 ;
  assign n16604 = x122 & n2890 ;
  assign n16603 = x124 & n2893 ;
  assign n16605 = n16604 ^ n16603 ;
  assign n16606 = n16605 ^ x32 ;
  assign n16602 = n2894 & n10117 ;
  assign n16607 = n16606 ^ n16602 ;
  assign n16601 = x123 & n2899 ;
  assign n16608 = n16607 ^ n16601 ;
  assign n16595 = x119 & n3387 ;
  assign n16594 = x121 & n3390 ;
  assign n16596 = n16595 ^ n16594 ;
  assign n16597 = n16596 ^ x35 ;
  assign n16593 = n3391 & n8979 ;
  assign n16598 = n16597 ^ n16593 ;
  assign n16592 = x120 & n3395 ;
  assign n16599 = n16598 ^ n16592 ;
  assign n16587 = n16389 ^ n16376 ;
  assign n16588 = n16381 & n16587 ;
  assign n16589 = n16588 ^ n16376 ;
  assign n16581 = x116 & n3932 ;
  assign n16580 = x118 & n3935 ;
  assign n16582 = n16581 ^ n16580 ;
  assign n16583 = n16582 ^ x38 ;
  assign n16579 = n3936 & ~n8140 ;
  assign n16584 = n16583 ^ n16579 ;
  assign n16578 = x117 & n3940 ;
  assign n16585 = n16584 ^ n16578 ;
  assign n16574 = n16375 ^ n16362 ;
  assign n16575 = n16367 & n16574 ;
  assign n16576 = n16575 ^ n16362 ;
  assign n16568 = x113 & n4482 ;
  assign n16567 = x115 & n4478 ;
  assign n16569 = n16568 ^ n16567 ;
  assign n16570 = n16569 ^ x41 ;
  assign n16566 = n4479 & ~n7353 ;
  assign n16571 = n16570 ^ n16566 ;
  assign n16565 = x114 & n4475 ;
  assign n16572 = n16571 ^ n16565 ;
  assign n16561 = n16361 ^ n16352 ;
  assign n16562 = ~n16353 & ~n16561 ;
  assign n16563 = n16562 ^ n16361 ;
  assign n16559 = x111 & n5121 ;
  assign n16554 = x110 & n5113 ;
  assign n16553 = x112 & n5116 ;
  assign n16555 = n16554 ^ n16553 ;
  assign n16556 = n16555 ^ x44 ;
  assign n16552 = n5117 & ~n6616 ;
  assign n16557 = n16556 ^ n16552 ;
  assign n16548 = n16347 ^ n16272 ;
  assign n16549 = n16348 & ~n16548 ;
  assign n16550 = n16549 ^ n16347 ;
  assign n16542 = x107 & n5981 ;
  assign n16541 = x109 & n5748 ;
  assign n16543 = n16542 ^ n16541 ;
  assign n16544 = n16543 ^ x47 ;
  assign n16540 = n5749 & n5912 ;
  assign n16545 = n16544 ^ n16540 ;
  assign n16539 = x108 & n5755 ;
  assign n16546 = n16545 ^ n16539 ;
  assign n16534 = ~n4624 & n7187 ;
  assign n16532 = x101 & n7183 ;
  assign n16530 = x103 & n7186 ;
  assign n16526 = n16323 ^ n16275 ;
  assign n16527 = n16324 & ~n16526 ;
  assign n16528 = n16527 ^ n16323 ;
  assign n16529 = n16528 ^ x53 ;
  assign n16531 = n16530 ^ n16529 ;
  assign n16533 = n16532 ^ n16531 ;
  assign n16535 = n16534 ^ n16533 ;
  assign n16525 = x102 & n7191 ;
  assign n16536 = n16535 ^ n16525 ;
  assign n16518 = x98 & n7954 ;
  assign n16517 = x100 & n7950 ;
  assign n16519 = n16518 ^ n16517 ;
  assign n16520 = n16519 ^ x56 ;
  assign n16516 = n4048 & n7951 ;
  assign n16521 = n16520 ^ n16516 ;
  assign n16515 = x99 & n7947 ;
  assign n16522 = n16521 ^ n16515 ;
  assign n16512 = x96 & n8743 ;
  assign n16510 = n3501 & n8747 ;
  assign n16506 = x95 & n8750 ;
  assign n16505 = x97 & n8746 ;
  assign n16507 = n16506 ^ n16505 ;
  assign n16508 = n16507 ^ x59 ;
  assign n16499 = ~n16283 & n16291 ;
  assign n16498 = x89 & n16281 ;
  assign n16500 = n16499 ^ n16498 ;
  assign n16501 = n16500 ^ n16140 ;
  assign n16502 = n16501 ^ x26 ;
  assign n16494 = x91 ^ x89 ;
  assign n16495 = ~n11895 & n16494 ;
  assign n16496 = n16495 ^ n2112 ;
  assign n16497 = n12206 & n16496 ;
  assign n16503 = n16502 ^ n16497 ;
  assign n16489 = x92 & n9655 ;
  assign n16488 = x94 & n9651 ;
  assign n16490 = n16489 ^ n16488 ;
  assign n16491 = n16490 ^ x62 ;
  assign n16487 = n3010 & n9652 ;
  assign n16492 = n16491 ^ n16487 ;
  assign n16486 = x93 & n9648 ;
  assign n16493 = n16492 ^ n16486 ;
  assign n16504 = n16503 ^ n16493 ;
  assign n16509 = n16508 ^ n16504 ;
  assign n16511 = n16510 ^ n16509 ;
  assign n16513 = n16512 ^ n16511 ;
  assign n16483 = n16301 ^ n16278 ;
  assign n16484 = n16293 & n16483 ;
  assign n16485 = n16484 ^ n16301 ;
  assign n16514 = n16513 ^ n16485 ;
  assign n16523 = n16522 ^ n16514 ;
  assign n16480 = n16314 ^ n16310 ;
  assign n16481 = n16311 & ~n16480 ;
  assign n16482 = n16481 ^ n16314 ;
  assign n16524 = n16523 ^ n16482 ;
  assign n16537 = n16536 ^ n16524 ;
  assign n16470 = x104 & n6687 ;
  assign n16469 = x106 & n6444 ;
  assign n16471 = n16470 ^ n16469 ;
  assign n16472 = n16471 ^ x50 ;
  assign n16468 = ~n5257 & n6445 ;
  assign n16473 = n16472 ^ n16468 ;
  assign n16467 = x105 & n6449 ;
  assign n16474 = n16473 ^ n16467 ;
  assign n16476 = n16474 ^ n16325 ;
  assign n16475 = n16474 ^ n16338 ;
  assign n16477 = n16476 ^ n16475 ;
  assign n16478 = n16330 & ~n16477 ;
  assign n16479 = n16478 ^ n16476 ;
  assign n16538 = n16537 ^ n16479 ;
  assign n16547 = n16546 ^ n16538 ;
  assign n16551 = n16550 ^ n16547 ;
  assign n16558 = n16557 ^ n16551 ;
  assign n16560 = n16559 ^ n16558 ;
  assign n16564 = n16563 ^ n16560 ;
  assign n16573 = n16572 ^ n16564 ;
  assign n16577 = n16576 ^ n16573 ;
  assign n16586 = n16585 ^ n16577 ;
  assign n16590 = n16589 ^ n16586 ;
  assign n16464 = n16402 ^ n16393 ;
  assign n16465 = ~n16394 & n16464 ;
  assign n16466 = n16465 ^ n16402 ;
  assign n16591 = n16590 ^ n16466 ;
  assign n16600 = n16599 ^ n16591 ;
  assign n16609 = n16608 ^ n16600 ;
  assign n16461 = n16412 ^ n16269 ;
  assign n16462 = ~n16404 & n16461 ;
  assign n16463 = n16462 ^ n16412 ;
  assign n16610 = n16609 ^ n16463 ;
  assign n16619 = n16618 ^ n16610 ;
  assign n16458 = n16422 ^ n16266 ;
  assign n16459 = ~n16414 & n16458 ;
  assign n16460 = n16459 ^ n16422 ;
  assign n16620 = n16619 ^ n16460 ;
  assign n16452 = ~n16259 & ~n16427 ;
  assign n16621 = n16620 ^ n16452 ;
  assign n16449 = n16427 ^ n16259 ;
  assign n16453 = n16452 ^ n16449 ;
  assign n16454 = n16453 ^ n16452 ;
  assign n16455 = n16454 ^ n16446 ;
  assign n16456 = n16455 ^ n16423 ;
  assign n16457 = n16263 & ~n16456 ;
  assign n16622 = n16621 ^ n16457 ;
  assign n16448 = n16446 ^ n16423 ;
  assign n16450 = n16449 ^ n16423 ;
  assign n16451 = n16448 & n16450 ;
  assign n16623 = n16622 ^ n16451 ;
  assign n16796 = ~n16263 & ~n16423 ;
  assign n16797 = n16796 ^ n16424 ;
  assign n16798 = n16797 ^ n16620 ;
  assign n16800 = n16452 ^ n16263 ;
  assign n16801 = n16424 & n16800 ;
  assign n16802 = n16801 ^ n16423 ;
  assign n16803 = n16802 ^ n16620 ;
  assign n16855 = n16803 ^ n16453 ;
  assign n16808 = n16796 ^ n16453 ;
  assign n16799 = n16453 ^ n16446 ;
  assign n16804 = n16803 ^ n16799 ;
  assign n16845 = n16808 ^ n16804 ;
  assign n16859 = n16855 ^ n16845 ;
  assign n16861 = n16859 ^ n16855 ;
  assign n16860 = n16859 ^ n16802 ;
  assign n16862 = n16861 ^ n16860 ;
  assign n16847 = n16845 ^ n16802 ;
  assign n16805 = n16804 ^ n16803 ;
  assign n16806 = n16805 ^ n16796 ;
  assign n16807 = n16806 ^ n16803 ;
  assign n16850 = n16847 ^ n16807 ;
  assign n16852 = n16850 ^ n16804 ;
  assign n16853 = n16852 ^ n16802 ;
  assign n16813 = n16807 ^ n16803 ;
  assign n16817 = n16813 ^ n16803 ;
  assign n16814 = n16813 ^ n16796 ;
  assign n16815 = n16814 ^ n16803 ;
  assign n16809 = n16808 ^ n16807 ;
  assign n16810 = n16809 ^ n16802 ;
  assign n16811 = n16810 ^ n16803 ;
  assign n16812 = n16811 ^ n16803 ;
  assign n16816 = n16815 ^ n16812 ;
  assign n16818 = n16817 ^ n16816 ;
  assign n16820 = n16818 ^ n16802 ;
  assign n16825 = n16820 ^ n16817 ;
  assign n16823 = n16815 ^ n16811 ;
  assign n16826 = n16825 ^ n16823 ;
  assign n16827 = ~n16803 & n16826 ;
  assign n16828 = n16827 ^ n16811 ;
  assign n16829 = n16828 ^ n16817 ;
  assign n16830 = n16829 ^ n16802 ;
  assign n16831 = n16823 ^ n16817 ;
  assign n16832 = n16831 ^ n16802 ;
  assign n16833 = n16830 & ~n16832 ;
  assign n16834 = n16818 ^ n16815 ;
  assign n16835 = n16834 ^ n16820 ;
  assign n16836 = n16818 ^ n16811 ;
  assign n16837 = n16836 ^ n16820 ;
  assign n16838 = n16835 & ~n16837 ;
  assign n16839 = n16833 & n16838 ;
  assign n16840 = n16839 ^ n16827 ;
  assign n16841 = n16840 ^ n16823 ;
  assign n16819 = n16818 ^ n16817 ;
  assign n16821 = n16820 ^ n16819 ;
  assign n16842 = n16841 ^ n16821 ;
  assign n16843 = n16842 ^ n16809 ;
  assign n16844 = n16843 ^ n16820 ;
  assign n16846 = n16845 ^ n16844 ;
  assign n16854 = n16853 ^ n16846 ;
  assign n16863 = n16862 ^ n16854 ;
  assign n16864 = n16863 ^ n16620 ;
  assign n16865 = n16864 ^ n16860 ;
  assign n16866 = n16446 ^ n16427 ;
  assign n16869 = n16449 & ~n16866 ;
  assign n16870 = n16869 ^ n16427 ;
  assign n16871 = ~n16865 & n16870 ;
  assign n16872 = n16798 & n16871 ;
  assign n16873 = n16872 ^ n16865 ;
  assign n16790 = n2429 & n10155 ;
  assign n16789 = x126 & n2593 ;
  assign n16791 = n16790 ^ n16789 ;
  assign n16792 = n16791 ^ x29 ;
  assign n16788 = x127 & n2435 ;
  assign n16793 = n16792 ^ n16788 ;
  assign n16784 = n16608 ^ n16463 ;
  assign n16785 = ~n16609 & n16784 ;
  assign n16786 = n16785 ^ n16608 ;
  assign n16778 = x123 & n2890 ;
  assign n16777 = x125 & n2893 ;
  assign n16779 = n16778 ^ n16777 ;
  assign n16780 = n16779 ^ x32 ;
  assign n16776 = n2894 & n10416 ;
  assign n16781 = n16780 ^ n16776 ;
  assign n16775 = x124 & n2899 ;
  assign n16782 = n16781 ^ n16775 ;
  assign n16764 = x120 & n3387 ;
  assign n16763 = x122 & n3390 ;
  assign n16765 = n16764 ^ n16763 ;
  assign n16766 = n16765 ^ x35 ;
  assign n16762 = n3391 & ~n9261 ;
  assign n16767 = n16766 ^ n16762 ;
  assign n16761 = x121 & n3395 ;
  assign n16768 = n16767 ^ n16761 ;
  assign n16754 = x117 & n3932 ;
  assign n16753 = x119 & n3935 ;
  assign n16755 = n16754 ^ n16753 ;
  assign n16756 = n16755 ^ x38 ;
  assign n16752 = n3936 & n8405 ;
  assign n16757 = n16756 ^ n16752 ;
  assign n16751 = x118 & n3940 ;
  assign n16758 = n16757 ^ n16751 ;
  assign n16744 = x114 & n4482 ;
  assign n16743 = x116 & n4478 ;
  assign n16745 = n16744 ^ n16743 ;
  assign n16746 = n16745 ^ x41 ;
  assign n16742 = n4479 & ~n7604 ;
  assign n16747 = n16746 ^ n16742 ;
  assign n16741 = x115 & n4475 ;
  assign n16748 = n16747 ^ n16741 ;
  assign n16734 = x111 & n5113 ;
  assign n16733 = x113 & n5116 ;
  assign n16735 = n16734 ^ n16733 ;
  assign n16736 = n16735 ^ x44 ;
  assign n16732 = n5117 & ~n6849 ;
  assign n16737 = n16736 ^ n16732 ;
  assign n16731 = x112 & n5121 ;
  assign n16738 = n16737 ^ n16731 ;
  assign n16720 = x108 & n5981 ;
  assign n16719 = x110 & n5748 ;
  assign n16721 = n16720 ^ n16719 ;
  assign n16722 = n16721 ^ x47 ;
  assign n16718 = n5749 & n6145 ;
  assign n16723 = n16722 ^ n16718 ;
  assign n16717 = x109 & n5755 ;
  assign n16724 = n16723 ^ n16717 ;
  assign n16706 = x105 & n6687 ;
  assign n16705 = x107 & n6444 ;
  assign n16707 = n16706 ^ n16705 ;
  assign n16708 = n16707 ^ x50 ;
  assign n16704 = ~n5459 & n6445 ;
  assign n16709 = n16708 ^ n16704 ;
  assign n16703 = x106 & n6449 ;
  assign n16710 = n16709 ^ n16703 ;
  assign n16698 = n16522 ^ n16482 ;
  assign n16699 = ~n16523 & ~n16698 ;
  assign n16700 = n16699 ^ n16522 ;
  assign n16692 = x102 & n7183 ;
  assign n16691 = x104 & n7186 ;
  assign n16693 = n16692 ^ n16691 ;
  assign n16694 = n16693 ^ x53 ;
  assign n16690 = ~n4830 & n7187 ;
  assign n16695 = n16694 ^ n16690 ;
  assign n16689 = x103 & n7191 ;
  assign n16696 = n16695 ^ n16689 ;
  assign n16685 = x97 & n8743 ;
  assign n16683 = n3673 & n8747 ;
  assign n16679 = x96 & n8750 ;
  assign n16678 = x98 & n8746 ;
  assign n16680 = n16679 ^ n16678 ;
  assign n16681 = n16680 ^ x59 ;
  assign n16672 = x93 & n9655 ;
  assign n16671 = x95 & n9651 ;
  assign n16673 = n16672 ^ n16671 ;
  assign n16674 = n16673 ^ x62 ;
  assign n16670 = n3166 & n9652 ;
  assign n16675 = n16674 ^ n16670 ;
  assign n16669 = x94 & n9648 ;
  assign n16676 = n16675 ^ n16669 ;
  assign n16665 = ~x63 & x91 ;
  assign n16666 = n16665 ^ n2379 ;
  assign n16667 = ~n9956 & n16666 ;
  assign n16654 = x90 ^ x26 ;
  assign n16657 = n16496 & ~n16654 ;
  assign n16658 = n16657 ^ x90 ;
  assign n16659 = n12206 & n16658 ;
  assign n16660 = n16659 ^ x92 ;
  assign n16668 = n16667 ^ n16660 ;
  assign n16677 = n16676 ^ n16668 ;
  assign n16682 = n16681 ^ n16677 ;
  assign n16684 = n16683 ^ n16682 ;
  assign n16686 = n16685 ^ n16684 ;
  assign n16651 = n16501 ^ n16493 ;
  assign n16652 = ~n16503 & n16651 ;
  assign n16653 = n16652 ^ n16501 ;
  assign n16687 = n16686 ^ n16653 ;
  assign n16648 = n4223 & n7951 ;
  assign n16646 = x99 & n7954 ;
  assign n16642 = n16504 ^ n16485 ;
  assign n16643 = ~n16513 & ~n16642 ;
  assign n16644 = n16643 ^ n16504 ;
  assign n16640 = x101 & n7950 ;
  assign n16641 = n16640 ^ x56 ;
  assign n16645 = n16644 ^ n16641 ;
  assign n16647 = n16646 ^ n16645 ;
  assign n16649 = n16648 ^ n16647 ;
  assign n16639 = x100 & n7947 ;
  assign n16650 = n16649 ^ n16639 ;
  assign n16688 = n16687 ^ n16650 ;
  assign n16697 = n16696 ^ n16688 ;
  assign n16701 = n16700 ^ n16697 ;
  assign n16636 = n16528 ^ n16524 ;
  assign n16637 = n16536 & n16636 ;
  assign n16638 = n16637 ^ n16528 ;
  assign n16702 = n16701 ^ n16638 ;
  assign n16711 = n16710 ^ n16702 ;
  assign n16713 = n16711 ^ n16474 ;
  assign n16712 = n16711 ^ n16537 ;
  assign n16714 = n16713 ^ n16712 ;
  assign n16715 = ~n16479 & n16714 ;
  assign n16716 = n16715 ^ n16713 ;
  assign n16725 = n16724 ^ n16716 ;
  assign n16726 = n16725 ^ n16550 ;
  assign n16727 = n16726 ^ n16538 ;
  assign n16728 = n16727 ^ n16725 ;
  assign n16729 = n16547 & ~n16728 ;
  assign n16730 = n16729 ^ n16726 ;
  assign n16739 = n16738 ^ n16730 ;
  assign n16633 = n16563 ^ n16551 ;
  assign n16634 = ~n16560 & ~n16633 ;
  assign n16635 = n16634 ^ n16551 ;
  assign n16740 = n16739 ^ n16635 ;
  assign n16749 = n16748 ^ n16740 ;
  assign n16630 = n16576 ^ n16572 ;
  assign n16631 = n16573 & n16630 ;
  assign n16632 = n16631 ^ n16576 ;
  assign n16750 = n16749 ^ n16632 ;
  assign n16759 = n16758 ^ n16750 ;
  assign n16627 = n16589 ^ n16585 ;
  assign n16628 = n16586 & n16627 ;
  assign n16629 = n16628 ^ n16589 ;
  assign n16760 = n16759 ^ n16629 ;
  assign n16769 = n16768 ^ n16760 ;
  assign n16770 = n16769 ^ n16599 ;
  assign n16771 = n16770 ^ n16769 ;
  assign n16772 = n16771 ^ n16466 ;
  assign n16773 = n16591 & n16772 ;
  assign n16774 = n16773 ^ n16770 ;
  assign n16783 = n16782 ^ n16774 ;
  assign n16787 = n16786 ^ n16783 ;
  assign n16794 = n16793 ^ n16787 ;
  assign n16624 = n16618 ^ n16460 ;
  assign n16625 = ~n16619 & n16624 ;
  assign n16626 = n16625 ^ n16618 ;
  assign n16795 = n16794 ^ n16626 ;
  assign n16874 = n16873 ^ n16795 ;
  assign n17046 = n16873 ^ n16626 ;
  assign n17047 = n16795 & n17046 ;
  assign n17048 = n17047 ^ n16873 ;
  assign n17034 = x127 & n2592 ;
  assign n17035 = n17034 ^ n2427 ;
  assign n17040 = n2170 & n11285 ;
  assign n17041 = n17040 ^ n17034 ;
  assign n17042 = n17035 & ~n17041 ;
  assign n17043 = n17042 ^ x28 ;
  assign n17023 = x124 & n2890 ;
  assign n17022 = x126 & n2893 ;
  assign n17024 = n17023 ^ n17022 ;
  assign n17025 = n17024 ^ x32 ;
  assign n17021 = n2894 & n10461 ;
  assign n17026 = n17025 ^ n17021 ;
  assign n17020 = x125 & n2899 ;
  assign n17027 = n17026 ^ n17020 ;
  assign n17009 = x121 & n3387 ;
  assign n17008 = x123 & n3390 ;
  assign n17010 = n17009 ^ n17008 ;
  assign n17011 = n17010 ^ x35 ;
  assign n17007 = n3391 & ~n9804 ;
  assign n17012 = n17011 ^ n17007 ;
  assign n17006 = x122 & n3395 ;
  assign n17013 = n17012 ^ n17006 ;
  assign n17002 = n16758 ^ n16632 ;
  assign n17003 = n16750 & n17002 ;
  assign n17004 = n17003 ^ n16758 ;
  assign n16996 = x118 & n3932 ;
  assign n16995 = x120 & n3935 ;
  assign n16997 = n16996 ^ n16995 ;
  assign n16998 = n16997 ^ x38 ;
  assign n16994 = n3936 & n8904 ;
  assign n16999 = n16998 ^ n16994 ;
  assign n16993 = x119 & n3940 ;
  assign n17000 = n16999 ^ n16993 ;
  assign n16982 = x115 & n4482 ;
  assign n16981 = x117 & n4478 ;
  assign n16983 = n16982 ^ n16981 ;
  assign n16984 = n16983 ^ x41 ;
  assign n16980 = n4479 & ~n7860 ;
  assign n16985 = n16984 ^ n16980 ;
  assign n16979 = x116 & n4475 ;
  assign n16986 = n16985 ^ n16979 ;
  assign n16968 = x112 & n5113 ;
  assign n16967 = x114 & n5116 ;
  assign n16969 = n16968 ^ n16967 ;
  assign n16970 = n16969 ^ x44 ;
  assign n16966 = n5117 & ~n7108 ;
  assign n16971 = n16970 ^ n16966 ;
  assign n16965 = x113 & n5121 ;
  assign n16972 = n16971 ^ n16965 ;
  assign n16954 = x109 & n5981 ;
  assign n16953 = x111 & n5748 ;
  assign n16955 = n16954 ^ n16953 ;
  assign n16956 = n16955 ^ x47 ;
  assign n16952 = n5749 & ~n6370 ;
  assign n16957 = n16956 ^ n16952 ;
  assign n16951 = x110 & n5755 ;
  assign n16958 = n16957 ^ n16951 ;
  assign n16941 = x97 & n8750 ;
  assign n16940 = x99 & n8746 ;
  assign n16942 = n16941 ^ n16940 ;
  assign n16943 = n16942 ^ x59 ;
  assign n16939 = n3851 & n8747 ;
  assign n16944 = n16943 ^ n16939 ;
  assign n16938 = x98 & n8743 ;
  assign n16945 = n16944 ^ n16938 ;
  assign n16936 = x95 & n9648 ;
  assign n16927 = x63 & n2379 ;
  assign n16928 = n16927 ^ n2529 ;
  assign n16929 = ~n9956 & n16928 ;
  assign n16930 = n16929 ^ n2529 ;
  assign n16920 = n16676 ^ n16659 ;
  assign n16921 = n16668 & n16920 ;
  assign n16922 = n16921 ^ n16676 ;
  assign n16931 = n16930 ^ n16922 ;
  assign n16932 = n16931 ^ x62 ;
  assign n16919 = x94 & n9655 ;
  assign n16933 = n16932 ^ n16919 ;
  assign n16918 = x96 & n9651 ;
  assign n16934 = n16933 ^ n16918 ;
  assign n16917 = n3336 & n9652 ;
  assign n16935 = n16934 ^ n16917 ;
  assign n16937 = n16936 ^ n16935 ;
  assign n16946 = n16945 ^ n16937 ;
  assign n16914 = n4425 & n7951 ;
  assign n16912 = x100 & n7954 ;
  assign n16908 = n16677 ^ n16653 ;
  assign n16909 = ~n16686 & ~n16908 ;
  assign n16910 = n16909 ^ n16677 ;
  assign n16906 = x102 & n7950 ;
  assign n16907 = n16906 ^ x56 ;
  assign n16911 = n16910 ^ n16907 ;
  assign n16913 = n16912 ^ n16911 ;
  assign n16915 = n16914 ^ n16913 ;
  assign n16905 = x101 & n7947 ;
  assign n16916 = n16915 ^ n16905 ;
  assign n16947 = n16946 ^ n16916 ;
  assign n16902 = ~n5034 & n7187 ;
  assign n16900 = x103 & n7183 ;
  assign n16896 = n16687 ^ n16644 ;
  assign n16897 = n16650 & n16896 ;
  assign n16898 = n16897 ^ n16687 ;
  assign n16894 = x105 & n7186 ;
  assign n16895 = n16894 ^ x53 ;
  assign n16899 = n16898 ^ n16895 ;
  assign n16901 = n16900 ^ n16899 ;
  assign n16903 = n16902 ^ n16901 ;
  assign n16893 = x104 & n7191 ;
  assign n16904 = n16903 ^ n16893 ;
  assign n16948 = n16947 ^ n16904 ;
  assign n16890 = n5687 & n6445 ;
  assign n16888 = x106 & n6687 ;
  assign n16884 = n16700 ^ n16696 ;
  assign n16885 = ~n16697 & n16884 ;
  assign n16886 = n16885 ^ n16700 ;
  assign n16882 = x108 & n6444 ;
  assign n16883 = n16882 ^ x50 ;
  assign n16887 = n16886 ^ n16883 ;
  assign n16889 = n16888 ^ n16887 ;
  assign n16891 = n16890 ^ n16889 ;
  assign n16881 = x107 & n6449 ;
  assign n16892 = n16891 ^ n16881 ;
  assign n16949 = n16948 ^ n16892 ;
  assign n16878 = n16710 ^ n16638 ;
  assign n16879 = ~n16702 & n16878 ;
  assign n16880 = n16879 ^ n16710 ;
  assign n16950 = n16949 ^ n16880 ;
  assign n16959 = n16958 ^ n16950 ;
  assign n16961 = n16959 ^ n16711 ;
  assign n16960 = n16959 ^ n16724 ;
  assign n16962 = n16961 ^ n16960 ;
  assign n16963 = n16716 & n16962 ;
  assign n16964 = n16963 ^ n16961 ;
  assign n16973 = n16972 ^ n16964 ;
  assign n16975 = n16973 ^ n16725 ;
  assign n16974 = n16973 ^ n16738 ;
  assign n16976 = n16975 ^ n16974 ;
  assign n16977 = n16730 & n16976 ;
  assign n16978 = n16977 ^ n16975 ;
  assign n16987 = n16986 ^ n16978 ;
  assign n16988 = n16987 ^ n16748 ;
  assign n16989 = n16988 ^ n16987 ;
  assign n16990 = n16989 ^ n16635 ;
  assign n16991 = n16740 & ~n16990 ;
  assign n16992 = n16991 ^ n16988 ;
  assign n17001 = n17000 ^ n16992 ;
  assign n17005 = n17004 ^ n17001 ;
  assign n17014 = n17013 ^ n17005 ;
  assign n17015 = n17014 ^ n16768 ;
  assign n17016 = n17015 ^ n17014 ;
  assign n17017 = n17016 ^ n16629 ;
  assign n17018 = n16760 & n17017 ;
  assign n17019 = n17018 ^ n17015 ;
  assign n17028 = n17027 ^ n17019 ;
  assign n17030 = n17028 ^ n16769 ;
  assign n17029 = n17028 ^ n16782 ;
  assign n17031 = n17030 ^ n17029 ;
  assign n17032 = ~n16774 & ~n17031 ;
  assign n17033 = n17032 ^ n17030 ;
  assign n17044 = n17043 ^ n17033 ;
  assign n16875 = n16793 ^ n16786 ;
  assign n16876 = n16787 & n16875 ;
  assign n16877 = n16876 ^ n16793 ;
  assign n17045 = n17044 ^ n16877 ;
  assign n17049 = n17048 ^ n17045 ;
  assign n17208 = n17027 ^ n17014 ;
  assign n17209 = ~n17019 & ~n17208 ;
  assign n17210 = n17209 ^ n17014 ;
  assign n17205 = n17043 ^ n17028 ;
  assign n17206 = n17033 & ~n17205 ;
  assign n17207 = n17206 ^ n17028 ;
  assign n17211 = n17210 ^ n17207 ;
  assign n17199 = x125 & n2890 ;
  assign n17198 = x127 & n2893 ;
  assign n17200 = n17199 ^ n17198 ;
  assign n17201 = n17200 ^ x32 ;
  assign n17197 = n2894 & n10986 ;
  assign n17202 = n17201 ^ n17197 ;
  assign n17196 = x126 & n2899 ;
  assign n17203 = n17202 ^ n17196 ;
  assign n17189 = x122 & n3387 ;
  assign n17188 = x124 & n3390 ;
  assign n17190 = n17189 ^ n17188 ;
  assign n17191 = n17190 ^ x35 ;
  assign n17187 = n3391 & n10117 ;
  assign n17192 = n17191 ^ n17187 ;
  assign n17186 = x123 & n3395 ;
  assign n17193 = n17192 ^ n17186 ;
  assign n17180 = x119 & n3932 ;
  assign n17179 = x121 & n3935 ;
  assign n17181 = n17180 ^ n17179 ;
  assign n17182 = n17181 ^ x38 ;
  assign n17178 = n3936 & n8979 ;
  assign n17183 = n17182 ^ n17178 ;
  assign n17177 = x120 & n3940 ;
  assign n17184 = n17183 ^ n17177 ;
  assign n17168 = n16986 ^ n16973 ;
  assign n17169 = ~n16978 & ~n17168 ;
  assign n17170 = n17169 ^ n16973 ;
  assign n17162 = x116 & n4482 ;
  assign n17161 = x118 & n4478 ;
  assign n17163 = n17162 ^ n17161 ;
  assign n17164 = n17163 ^ x41 ;
  assign n17160 = n4479 & ~n8140 ;
  assign n17165 = n17164 ^ n17160 ;
  assign n17159 = x117 & n4475 ;
  assign n17166 = n17165 ^ n17159 ;
  assign n17155 = n16972 ^ n16959 ;
  assign n17156 = ~n16964 & ~n17155 ;
  assign n17157 = n17156 ^ n16959 ;
  assign n17149 = x113 & n5113 ;
  assign n17148 = x115 & n5116 ;
  assign n17150 = n17149 ^ n17148 ;
  assign n17151 = n17150 ^ x44 ;
  assign n17147 = n5117 & ~n7353 ;
  assign n17152 = n17151 ^ n17147 ;
  assign n17146 = x114 & n5121 ;
  assign n17153 = n17152 ^ n17146 ;
  assign n17139 = x110 & n5981 ;
  assign n17138 = x112 & n5748 ;
  assign n17140 = n17139 ^ n17138 ;
  assign n17141 = n17140 ^ x47 ;
  assign n17137 = n5749 & ~n6616 ;
  assign n17142 = n17141 ^ n17137 ;
  assign n17136 = x111 & n5755 ;
  assign n17143 = n17142 ^ n17136 ;
  assign n17124 = x95 & n9655 ;
  assign n17123 = x97 & n9651 ;
  assign n17125 = n17124 ^ n17123 ;
  assign n17126 = n17125 ^ x62 ;
  assign n17122 = n3501 & n9652 ;
  assign n17127 = n17126 ^ n17122 ;
  assign n17121 = x96 & n9648 ;
  assign n17128 = n17127 ^ n17121 ;
  assign n17129 = n17128 ^ x29 ;
  assign n17117 = x94 ^ x92 ;
  assign n17118 = ~n11895 & n17117 ;
  assign n17119 = n17118 ^ n2529 ;
  assign n17120 = n12206 & n17119 ;
  assign n17130 = n17129 ^ n17120 ;
  assign n17115 = ~n16922 & ~n16930 ;
  assign n17109 = n9956 ^ x92 ;
  assign n17110 = x63 & ~x91 ;
  assign n17111 = n17110 ^ x93 ;
  assign n17112 = x92 & n17111 ;
  assign n17113 = n17112 ^ x93 ;
  assign n17114 = n17109 & n17113 ;
  assign n17116 = n17115 ^ n17114 ;
  assign n17131 = n17130 ^ n17116 ;
  assign n17099 = x98 & n8750 ;
  assign n17098 = x100 & n8746 ;
  assign n17100 = n17099 ^ n17098 ;
  assign n17101 = n17100 ^ x59 ;
  assign n17097 = n4048 & n8747 ;
  assign n17102 = n17101 ^ n17097 ;
  assign n17096 = x99 & n8743 ;
  assign n17103 = n17102 ^ n17096 ;
  assign n17104 = n17103 ^ n16945 ;
  assign n17105 = n17104 ^ n16931 ;
  assign n17106 = n17105 ^ n17103 ;
  assign n17107 = n16937 & ~n17106 ;
  assign n17108 = n17107 ^ n17104 ;
  assign n17132 = n17131 ^ n17108 ;
  assign n17093 = ~n4624 & n7951 ;
  assign n17091 = x101 & n7954 ;
  assign n17087 = n16946 ^ n16910 ;
  assign n17088 = n16916 & n17087 ;
  assign n17089 = n17088 ^ n16946 ;
  assign n17085 = x103 & n7950 ;
  assign n17086 = n17085 ^ x56 ;
  assign n17090 = n17089 ^ n17086 ;
  assign n17092 = n17091 ^ n17090 ;
  assign n17094 = n17093 ^ n17092 ;
  assign n17084 = x102 & n7947 ;
  assign n17095 = n17094 ^ n17084 ;
  assign n17133 = n17132 ^ n17095 ;
  assign n17074 = x104 & n7183 ;
  assign n17073 = x106 & n7186 ;
  assign n17075 = n17074 ^ n17073 ;
  assign n17076 = n17075 ^ x53 ;
  assign n17072 = ~n5257 & n7187 ;
  assign n17077 = n17076 ^ n17072 ;
  assign n17071 = x105 & n7191 ;
  assign n17078 = n17077 ^ n17071 ;
  assign n17079 = n17078 ^ n16947 ;
  assign n17080 = n17079 ^ n17078 ;
  assign n17081 = n17080 ^ n16898 ;
  assign n17082 = n16904 & ~n17081 ;
  assign n17083 = n17082 ^ n17079 ;
  assign n17134 = n17133 ^ n17083 ;
  assign n17068 = n5912 & n6445 ;
  assign n17066 = x107 & n6687 ;
  assign n17064 = x109 & n6444 ;
  assign n17060 = n16948 ^ n16886 ;
  assign n17061 = ~n16892 & ~n17060 ;
  assign n17062 = n17061 ^ n16948 ;
  assign n17063 = n17062 ^ x50 ;
  assign n17065 = n17064 ^ n17063 ;
  assign n17067 = n17066 ^ n17065 ;
  assign n17069 = n17068 ^ n17067 ;
  assign n17059 = x108 & n6449 ;
  assign n17070 = n17069 ^ n17059 ;
  assign n17135 = n17134 ^ n17070 ;
  assign n17144 = n17143 ^ n17135 ;
  assign n17056 = n16958 ^ n16880 ;
  assign n17057 = n16950 & n17056 ;
  assign n17058 = n17057 ^ n16958 ;
  assign n17145 = n17144 ^ n17058 ;
  assign n17154 = n17153 ^ n17145 ;
  assign n17158 = n17157 ^ n17154 ;
  assign n17167 = n17166 ^ n17158 ;
  assign n17171 = n17170 ^ n17167 ;
  assign n17173 = n17171 ^ n16987 ;
  assign n17172 = n17171 ^ n17000 ;
  assign n17174 = n17173 ^ n17172 ;
  assign n17175 = ~n16992 & ~n17174 ;
  assign n17176 = n17175 ^ n17173 ;
  assign n17185 = n17184 ^ n17176 ;
  assign n17194 = n17193 ^ n17185 ;
  assign n17053 = n17013 ^ n17004 ;
  assign n17054 = n17005 & n17053 ;
  assign n17055 = n17054 ^ n17013 ;
  assign n17195 = n17194 ^ n17055 ;
  assign n17204 = n17203 ^ n17195 ;
  assign n17212 = n17211 ^ n17204 ;
  assign n17050 = n17048 ^ n16877 ;
  assign n17051 = ~n17045 & n17050 ;
  assign n17052 = n17051 ^ n17048 ;
  assign n17213 = n17212 ^ n17052 ;
  assign n17365 = ~n17195 & n17203 ;
  assign n17364 = n17207 & n17210 ;
  assign n17366 = n17365 ^ n17364 ;
  assign n17359 = n2894 & n10155 ;
  assign n17358 = x126 & n2890 ;
  assign n17360 = n17359 ^ n17358 ;
  assign n17361 = n17360 ^ x32 ;
  assign n17357 = x127 & n2899 ;
  assign n17362 = n17361 ^ n17357 ;
  assign n17353 = n17193 ^ n17055 ;
  assign n17354 = ~n17194 & n17353 ;
  assign n17355 = n17354 ^ n17193 ;
  assign n17347 = x123 & n3387 ;
  assign n17346 = x125 & n3390 ;
  assign n17348 = n17347 ^ n17346 ;
  assign n17349 = n17348 ^ x35 ;
  assign n17345 = n3391 & n10416 ;
  assign n17350 = n17349 ^ n17345 ;
  assign n17344 = x124 & n3395 ;
  assign n17351 = n17350 ^ n17344 ;
  assign n17340 = n17184 ^ n17171 ;
  assign n17341 = ~n17176 & n17340 ;
  assign n17342 = n17341 ^ n17171 ;
  assign n17334 = x120 & n3932 ;
  assign n17333 = x122 & n3935 ;
  assign n17335 = n17334 ^ n17333 ;
  assign n17336 = n17335 ^ x38 ;
  assign n17332 = n3936 & ~n9261 ;
  assign n17337 = n17336 ^ n17332 ;
  assign n17331 = x121 & n3940 ;
  assign n17338 = n17337 ^ n17331 ;
  assign n17324 = x117 & n4482 ;
  assign n17323 = x119 & n4478 ;
  assign n17325 = n17324 ^ n17323 ;
  assign n17326 = n17325 ^ x41 ;
  assign n17322 = n4479 & n8405 ;
  assign n17327 = n17326 ^ n17322 ;
  assign n17321 = x118 & n4475 ;
  assign n17328 = n17327 ^ n17321 ;
  assign n17314 = x114 & n5113 ;
  assign n17313 = x116 & n5116 ;
  assign n17315 = n17314 ^ n17313 ;
  assign n17316 = n17315 ^ x44 ;
  assign n17312 = n5117 & ~n7604 ;
  assign n17317 = n17316 ^ n17312 ;
  assign n17311 = x115 & n5121 ;
  assign n17318 = n17317 ^ n17311 ;
  assign n17304 = x111 & n5981 ;
  assign n17303 = x113 & n5748 ;
  assign n17305 = n17304 ^ n17303 ;
  assign n17306 = n17305 ^ x47 ;
  assign n17302 = n5749 & ~n6849 ;
  assign n17307 = n17306 ^ n17302 ;
  assign n17301 = x112 & n5755 ;
  assign n17308 = n17307 ^ n17301 ;
  assign n17291 = ~n5459 & n7187 ;
  assign n17289 = x105 & n7183 ;
  assign n17285 = n17132 ^ n17089 ;
  assign n17286 = n17095 & ~n17285 ;
  assign n17287 = n17286 ^ n17132 ;
  assign n17283 = x107 & n7186 ;
  assign n17284 = n17283 ^ x53 ;
  assign n17288 = n17287 ^ n17284 ;
  assign n17290 = n17289 ^ n17288 ;
  assign n17292 = n17291 ^ n17290 ;
  assign n17282 = x106 & n7191 ;
  assign n17293 = n17292 ^ n17282 ;
  assign n17279 = x103 & n7947 ;
  assign n17277 = ~n4830 & n7951 ;
  assign n17273 = x102 & n7954 ;
  assign n17272 = x104 & n7950 ;
  assign n17274 = n17273 ^ n17272 ;
  assign n17275 = n17274 ^ x56 ;
  assign n17268 = n4223 & n8747 ;
  assign n17266 = x99 & n8750 ;
  assign n17262 = x94 & n11895 ;
  assign n17261 = x95 & n9956 ;
  assign n17263 = n17262 ^ n17261 ;
  assign n17258 = n3673 & n9652 ;
  assign n17256 = x96 & n9655 ;
  assign n17249 = x93 ^ x29 ;
  assign n17252 = n17119 & ~n17249 ;
  assign n17253 = n17252 ^ x93 ;
  assign n17254 = n12206 & n17253 ;
  assign n17247 = x98 & n9651 ;
  assign n17248 = n17247 ^ x62 ;
  assign n17255 = n17254 ^ n17248 ;
  assign n17257 = n17256 ^ n17255 ;
  assign n17259 = n17258 ^ n17257 ;
  assign n17246 = x97 & n9648 ;
  assign n17260 = n17259 ^ n17246 ;
  assign n17264 = n17263 ^ n17260 ;
  assign n17244 = x101 & n8746 ;
  assign n17245 = n17244 ^ x59 ;
  assign n17265 = n17264 ^ n17245 ;
  assign n17267 = n17266 ^ n17265 ;
  assign n17269 = n17268 ^ n17267 ;
  assign n17243 = x100 & n8743 ;
  assign n17270 = n17269 ^ n17243 ;
  assign n17240 = n17128 ^ n17116 ;
  assign n17241 = ~n17130 & ~n17240 ;
  assign n17242 = n17241 ^ n17128 ;
  assign n17271 = n17270 ^ n17242 ;
  assign n17276 = n17275 ^ n17271 ;
  assign n17278 = n17277 ^ n17276 ;
  assign n17280 = n17279 ^ n17278 ;
  assign n17237 = n17131 ^ n17103 ;
  assign n17238 = n17108 & n17237 ;
  assign n17239 = n17238 ^ n17103 ;
  assign n17281 = n17280 ^ n17239 ;
  assign n17294 = n17293 ^ n17281 ;
  assign n17234 = n6145 & n6445 ;
  assign n17232 = x108 & n6687 ;
  assign n17228 = n17133 ^ n17078 ;
  assign n17229 = n17083 & ~n17228 ;
  assign n17230 = n17229 ^ n17078 ;
  assign n17226 = x110 & n6444 ;
  assign n17227 = n17226 ^ x50 ;
  assign n17231 = n17230 ^ n17227 ;
  assign n17233 = n17232 ^ n17231 ;
  assign n17235 = n17234 ^ n17233 ;
  assign n17225 = x109 & n6449 ;
  assign n17236 = n17235 ^ n17225 ;
  assign n17295 = n17294 ^ n17236 ;
  assign n17296 = n17295 ^ n17134 ;
  assign n17297 = n17296 ^ n17062 ;
  assign n17298 = n17297 ^ n17295 ;
  assign n17299 = n17070 & n17298 ;
  assign n17300 = n17299 ^ n17296 ;
  assign n17309 = n17308 ^ n17300 ;
  assign n17222 = n17143 ^ n17058 ;
  assign n17223 = n17144 & n17222 ;
  assign n17224 = n17223 ^ n17143 ;
  assign n17310 = n17309 ^ n17224 ;
  assign n17319 = n17318 ^ n17310 ;
  assign n17219 = n17157 ^ n17153 ;
  assign n17220 = ~n17154 & ~n17219 ;
  assign n17221 = n17220 ^ n17157 ;
  assign n17320 = n17319 ^ n17221 ;
  assign n17329 = n17328 ^ n17320 ;
  assign n17216 = n17170 ^ n17166 ;
  assign n17217 = n17167 & ~n17216 ;
  assign n17218 = n17217 ^ n17170 ;
  assign n17330 = n17329 ^ n17218 ;
  assign n17339 = n17338 ^ n17330 ;
  assign n17343 = n17342 ^ n17339 ;
  assign n17352 = n17351 ^ n17343 ;
  assign n17356 = n17355 ^ n17352 ;
  assign n17363 = n17362 ^ n17356 ;
  assign n17367 = n17366 ^ n17363 ;
  assign n17214 = n17204 ^ n17052 ;
  assign n17215 = ~n17212 & n17214 ;
  assign n17368 = n17367 ^ n17215 ;
  assign n17552 = n17211 ^ n17203 ;
  assign n17553 = n17552 ^ n17195 ;
  assign n17534 = n17363 ^ n17195 ;
  assign n17532 = n17363 ^ n17207 ;
  assign n17554 = n17534 ^ n17532 ;
  assign n17538 = n17363 ^ n17203 ;
  assign n17555 = n17538 ^ n17532 ;
  assign n17556 = n17554 & ~n17555 ;
  assign n17557 = n17556 ^ n17532 ;
  assign n17558 = ~n17553 & ~n17557 ;
  assign n17559 = n17052 & n17558 ;
  assign n17533 = n17532 ^ n17363 ;
  assign n17535 = n17534 ^ n17363 ;
  assign n17536 = ~n17533 & ~n17535 ;
  assign n17537 = n17536 ^ n17363 ;
  assign n17545 = n17535 ^ n17533 ;
  assign n17546 = n17545 ^ n17363 ;
  assign n17539 = n17363 ^ n17210 ;
  assign n17540 = n17539 ^ n17538 ;
  assign n17541 = n17539 ^ n17534 ;
  assign n17542 = n17541 ^ n17532 ;
  assign n17543 = n17542 ^ n17363 ;
  assign n17544 = n17540 & ~n17543 ;
  assign n17547 = n17546 ^ n17544 ;
  assign n17548 = n17537 & n17547 ;
  assign n17549 = n17548 ^ n17363 ;
  assign n17560 = n17559 ^ n17549 ;
  assign n17527 = n17351 ^ n17342 ;
  assign n17528 = ~n17343 & n17527 ;
  assign n17529 = n17528 ^ n17351 ;
  assign n17511 = n2746 ^ x31 ;
  assign n17512 = x127 & n2887 ;
  assign n17513 = n17511 & n17512 ;
  assign n17514 = n17513 ^ x32 ;
  assign n17520 = ~x31 & ~x127 ;
  assign n17521 = n17520 ^ n2887 ;
  assign n17522 = ~n10154 & n17521 ;
  assign n17523 = n17522 ^ x32 ;
  assign n17524 = n2747 & ~n17523 ;
  assign n17525 = n17514 & n17524 ;
  assign n17505 = x124 & n3387 ;
  assign n17504 = x126 & n3390 ;
  assign n17506 = n17505 ^ n17504 ;
  assign n17507 = n17506 ^ x35 ;
  assign n17503 = n3391 & n10461 ;
  assign n17508 = n17507 ^ n17503 ;
  assign n17502 = x125 & n3395 ;
  assign n17509 = n17508 ^ n17502 ;
  assign n17491 = x121 & n3932 ;
  assign n17490 = x123 & n3935 ;
  assign n17492 = n17491 ^ n17490 ;
  assign n17493 = n17492 ^ x38 ;
  assign n17489 = n3936 & ~n9804 ;
  assign n17494 = n17493 ^ n17489 ;
  assign n17488 = x122 & n3940 ;
  assign n17495 = n17494 ^ n17488 ;
  assign n17481 = x118 & n4482 ;
  assign n17480 = x120 & n4478 ;
  assign n17482 = n17481 ^ n17480 ;
  assign n17483 = n17482 ^ x41 ;
  assign n17479 = n4479 & n8904 ;
  assign n17484 = n17483 ^ n17479 ;
  assign n17478 = x119 & n4475 ;
  assign n17485 = n17484 ^ n17478 ;
  assign n17467 = x115 & n5113 ;
  assign n17466 = x117 & n5116 ;
  assign n17468 = n17467 ^ n17466 ;
  assign n17469 = n17468 ^ x44 ;
  assign n17465 = n5117 & ~n7860 ;
  assign n17470 = n17469 ^ n17465 ;
  assign n17464 = x116 & n5121 ;
  assign n17471 = n17470 ^ n17464 ;
  assign n17453 = x112 & n5981 ;
  assign n17452 = x114 & n5748 ;
  assign n17454 = n17453 ^ n17452 ;
  assign n17455 = n17454 ^ x47 ;
  assign n17451 = n5749 & ~n7108 ;
  assign n17456 = n17455 ^ n17451 ;
  assign n17450 = x113 & n5755 ;
  assign n17457 = n17456 ^ n17450 ;
  assign n17443 = x109 & n6687 ;
  assign n17442 = x111 & n6444 ;
  assign n17444 = n17443 ^ n17442 ;
  assign n17445 = n17444 ^ x50 ;
  assign n17441 = ~n6370 & n6445 ;
  assign n17446 = n17445 ^ n17441 ;
  assign n17440 = x110 & n6449 ;
  assign n17447 = n17446 ^ n17440 ;
  assign n17436 = n17287 ^ n17281 ;
  assign n17437 = ~n17293 & ~n17436 ;
  assign n17438 = n17437 ^ n17281 ;
  assign n17432 = n5687 & n7187 ;
  assign n17430 = x106 & n7183 ;
  assign n17426 = n17271 ^ n17239 ;
  assign n17427 = ~n17280 & ~n17426 ;
  assign n17428 = n17427 ^ n17271 ;
  assign n17424 = x108 & n7186 ;
  assign n17425 = n17424 ^ x53 ;
  assign n17429 = n17428 ^ n17425 ;
  assign n17431 = n17430 ^ n17429 ;
  assign n17433 = n17432 ^ n17431 ;
  assign n17423 = x107 & n7191 ;
  assign n17434 = n17433 ^ n17423 ;
  assign n17416 = x100 & n8750 ;
  assign n17415 = x102 & n8746 ;
  assign n17417 = n17416 ^ n17415 ;
  assign n17418 = n17417 ^ x59 ;
  assign n17414 = n4425 & n8747 ;
  assign n17419 = n17418 ^ n17414 ;
  assign n17413 = x101 & n8743 ;
  assign n17420 = n17419 ^ n17413 ;
  assign n17407 = x97 & n9655 ;
  assign n17406 = x99 & n9651 ;
  assign n17408 = n17407 ^ n17406 ;
  assign n17409 = n17408 ^ x62 ;
  assign n17405 = n3851 & n9652 ;
  assign n17410 = n17409 ^ n17405 ;
  assign n17404 = x98 & n9648 ;
  assign n17411 = n17410 ^ n17404 ;
  assign n17400 = n17263 ^ n17254 ;
  assign n17401 = ~n17260 & ~n17400 ;
  assign n17402 = n17401 ^ n17263 ;
  assign n17394 = n9956 ^ x95 ;
  assign n17390 = ~x96 & n9956 ;
  assign n17391 = n17390 ^ n17262 ;
  assign n17395 = n17391 ^ n12206 ;
  assign n17396 = n17394 & n17395 ;
  assign n17397 = n17396 ^ n2988 ;
  assign n17392 = x95 & n17391 ;
  assign n17393 = n17392 ^ n17262 ;
  assign n17398 = n17397 ^ n17393 ;
  assign n17399 = n17398 ^ n2988 ;
  assign n17403 = n17402 ^ n17399 ;
  assign n17412 = n17411 ^ n17403 ;
  assign n17421 = n17420 ^ n17412 ;
  assign n17387 = ~n5034 & n7951 ;
  assign n17385 = x103 & n7954 ;
  assign n17381 = n17264 ^ n17242 ;
  assign n17382 = ~n17270 & ~n17381 ;
  assign n17383 = n17382 ^ n17264 ;
  assign n17379 = x105 & n7950 ;
  assign n17380 = n17379 ^ x56 ;
  assign n17384 = n17383 ^ n17380 ;
  assign n17386 = n17385 ^ n17384 ;
  assign n17388 = n17387 ^ n17386 ;
  assign n17378 = x104 & n7947 ;
  assign n17389 = n17388 ^ n17378 ;
  assign n17422 = n17421 ^ n17389 ;
  assign n17435 = n17434 ^ n17422 ;
  assign n17439 = n17438 ^ n17435 ;
  assign n17448 = n17447 ^ n17439 ;
  assign n17375 = n17294 ^ n17230 ;
  assign n17376 = ~n17236 & ~n17375 ;
  assign n17377 = n17376 ^ n17294 ;
  assign n17449 = n17448 ^ n17377 ;
  assign n17458 = n17457 ^ n17449 ;
  assign n17460 = n17458 ^ n17295 ;
  assign n17459 = n17458 ^ n17308 ;
  assign n17461 = n17460 ^ n17459 ;
  assign n17462 = n17300 & ~n17461 ;
  assign n17463 = n17462 ^ n17460 ;
  assign n17472 = n17471 ^ n17463 ;
  assign n17473 = n17472 ^ n17318 ;
  assign n17474 = n17473 ^ n17472 ;
  assign n17475 = n17474 ^ n17224 ;
  assign n17476 = ~n17310 & n17475 ;
  assign n17477 = n17476 ^ n17473 ;
  assign n17486 = n17485 ^ n17477 ;
  assign n17372 = n17328 ^ n17221 ;
  assign n17373 = n17320 & ~n17372 ;
  assign n17374 = n17373 ^ n17328 ;
  assign n17487 = n17486 ^ n17374 ;
  assign n17496 = n17495 ^ n17487 ;
  assign n17497 = n17496 ^ n17338 ;
  assign n17498 = n17497 ^ n17496 ;
  assign n17499 = n17498 ^ n17218 ;
  assign n17500 = ~n17330 & ~n17499 ;
  assign n17501 = n17500 ^ n17497 ;
  assign n17510 = n17509 ^ n17501 ;
  assign n17515 = n17514 ^ n17510 ;
  assign n17526 = n17525 ^ n17515 ;
  assign n17530 = n17529 ^ n17526 ;
  assign n17369 = n17362 ^ n17355 ;
  assign n17370 = ~n17356 & n17369 ;
  assign n17371 = n17370 ^ n17362 ;
  assign n17531 = n17530 ^ n17371 ;
  assign n17561 = n17560 ^ n17531 ;
  assign n17703 = n17509 ^ n17496 ;
  assign n17704 = ~n17501 & ~n17703 ;
  assign n17705 = n17704 ^ n17496 ;
  assign n17697 = x125 & n3387 ;
  assign n17696 = x127 & n3390 ;
  assign n17698 = n17697 ^ n17696 ;
  assign n17699 = n17698 ^ x35 ;
  assign n17695 = n3391 & n10986 ;
  assign n17700 = n17699 ^ n17695 ;
  assign n17694 = x126 & n3395 ;
  assign n17701 = n17700 ^ n17694 ;
  assign n17687 = x122 & n3932 ;
  assign n17686 = x124 & n3935 ;
  assign n17688 = n17687 ^ n17686 ;
  assign n17689 = n17688 ^ x38 ;
  assign n17685 = n3936 & n10117 ;
  assign n17690 = n17689 ^ n17685 ;
  assign n17684 = x123 & n3940 ;
  assign n17691 = n17690 ^ n17684 ;
  assign n17678 = x119 & n4482 ;
  assign n17677 = x121 & n4478 ;
  assign n17679 = n17678 ^ n17677 ;
  assign n17680 = n17679 ^ x41 ;
  assign n17676 = n4479 & n8979 ;
  assign n17681 = n17680 ^ n17676 ;
  assign n17675 = x120 & n4475 ;
  assign n17682 = n17681 ^ n17675 ;
  assign n17671 = n17485 ^ n17472 ;
  assign n17672 = ~n17477 & ~n17671 ;
  assign n17673 = n17672 ^ n17472 ;
  assign n17665 = x116 & n5113 ;
  assign n17664 = x118 & n5116 ;
  assign n17666 = n17665 ^ n17664 ;
  assign n17667 = n17666 ^ x44 ;
  assign n17663 = n5117 & ~n8140 ;
  assign n17668 = n17667 ^ n17663 ;
  assign n17662 = x117 & n5121 ;
  assign n17669 = n17668 ^ n17662 ;
  assign n17653 = n17457 ^ n17377 ;
  assign n17654 = ~n17449 & ~n17653 ;
  assign n17655 = n17654 ^ n17457 ;
  assign n17651 = x114 & n5755 ;
  assign n17646 = x113 & n5981 ;
  assign n17645 = x115 & n5748 ;
  assign n17647 = n17646 ^ n17645 ;
  assign n17648 = n17647 ^ x47 ;
  assign n17644 = n5749 & ~n7353 ;
  assign n17649 = n17648 ^ n17644 ;
  assign n17632 = x98 & n9655 ;
  assign n17631 = x100 & n9651 ;
  assign n17633 = n17632 ^ n17631 ;
  assign n17634 = n17633 ^ x62 ;
  assign n17630 = n4048 & n9652 ;
  assign n17635 = n17634 ^ n17630 ;
  assign n17629 = x99 & n9648 ;
  assign n17636 = n17635 ^ n17629 ;
  assign n17637 = n17636 ^ x32 ;
  assign n17625 = x97 ^ x95 ;
  assign n17626 = ~n11895 & n17625 ;
  assign n17627 = n17626 ^ n2988 ;
  assign n17628 = n12206 & n17627 ;
  assign n17638 = n17637 ^ n17628 ;
  assign n17622 = ~n17396 & n17402 ;
  assign n17623 = ~n17393 & n17622 ;
  assign n17624 = n17623 ^ n17396 ;
  assign n17639 = n17638 ^ n17624 ;
  assign n17619 = ~n4624 & n8747 ;
  assign n17617 = x101 & n8750 ;
  assign n17613 = n17420 ^ n17411 ;
  assign n17614 = ~n17412 & n17613 ;
  assign n17615 = n17614 ^ n17420 ;
  assign n17611 = x103 & n8746 ;
  assign n17612 = n17611 ^ x59 ;
  assign n17616 = n17615 ^ n17612 ;
  assign n17618 = n17617 ^ n17616 ;
  assign n17620 = n17619 ^ n17618 ;
  assign n17610 = x102 & n8743 ;
  assign n17621 = n17620 ^ n17610 ;
  assign n17640 = n17639 ^ n17621 ;
  assign n17600 = x104 & n7954 ;
  assign n17599 = x106 & n7950 ;
  assign n17601 = n17600 ^ n17599 ;
  assign n17602 = n17601 ^ x56 ;
  assign n17598 = ~n5257 & n7951 ;
  assign n17603 = n17602 ^ n17598 ;
  assign n17597 = x105 & n7947 ;
  assign n17604 = n17603 ^ n17597 ;
  assign n17605 = n17604 ^ n17421 ;
  assign n17606 = n17605 ^ n17383 ;
  assign n17607 = n17606 ^ n17604 ;
  assign n17608 = n17389 & ~n17607 ;
  assign n17609 = n17608 ^ n17605 ;
  assign n17641 = n17640 ^ n17609 ;
  assign n17594 = n17428 ^ n17422 ;
  assign n17595 = n17434 & n17594 ;
  assign n17587 = x107 & n7183 ;
  assign n17586 = x109 & n7186 ;
  assign n17588 = n17587 ^ n17586 ;
  assign n17589 = n17588 ^ x53 ;
  assign n17585 = n5912 & n7187 ;
  assign n17590 = n17589 ^ n17585 ;
  assign n17584 = x108 & n7191 ;
  assign n17591 = n17590 ^ n17584 ;
  assign n17592 = n17591 ^ n17422 ;
  assign n17596 = n17595 ^ n17592 ;
  assign n17642 = n17641 ^ n17596 ;
  assign n17574 = x110 & n6687 ;
  assign n17573 = x112 & n6444 ;
  assign n17575 = n17574 ^ n17573 ;
  assign n17576 = n17575 ^ x50 ;
  assign n17572 = n6445 & ~n6616 ;
  assign n17577 = n17576 ^ n17572 ;
  assign n17571 = x111 & n6449 ;
  assign n17578 = n17577 ^ n17571 ;
  assign n17579 = n17578 ^ n17447 ;
  assign n17580 = n17579 ^ n17438 ;
  assign n17581 = n17580 ^ n17578 ;
  assign n17582 = n17439 & ~n17581 ;
  assign n17583 = n17582 ^ n17579 ;
  assign n17643 = n17642 ^ n17583 ;
  assign n17650 = n17649 ^ n17643 ;
  assign n17652 = n17651 ^ n17650 ;
  assign n17656 = n17655 ^ n17652 ;
  assign n17658 = n17656 ^ n17458 ;
  assign n17657 = n17656 ^ n17471 ;
  assign n17659 = n17658 ^ n17657 ;
  assign n17660 = ~n17463 & n17659 ;
  assign n17661 = n17660 ^ n17658 ;
  assign n17670 = n17669 ^ n17661 ;
  assign n17674 = n17673 ^ n17670 ;
  assign n17683 = n17682 ^ n17674 ;
  assign n17692 = n17691 ^ n17683 ;
  assign n17568 = n17495 ^ n17374 ;
  assign n17569 = n17487 & n17568 ;
  assign n17570 = n17569 ^ n17495 ;
  assign n17693 = n17692 ^ n17570 ;
  assign n17702 = n17701 ^ n17693 ;
  assign n17706 = n17705 ^ n17702 ;
  assign n17565 = n17529 ^ n17510 ;
  assign n17566 = ~n17526 & ~n17565 ;
  assign n17567 = n17566 ^ n17510 ;
  assign n17707 = n17706 ^ n17567 ;
  assign n17562 = n17560 ^ n17371 ;
  assign n17563 = n17531 & n17562 ;
  assign n17564 = n17563 ^ n17560 ;
  assign n17708 = n17707 ^ n17564 ;
  assign n17847 = n17691 ^ n17570 ;
  assign n17848 = n17692 & n17847 ;
  assign n17849 = n17848 ^ n17691 ;
  assign n17844 = n17705 ^ n17701 ;
  assign n17845 = ~n17702 & ~n17844 ;
  assign n17846 = n17845 ^ n17705 ;
  assign n17854 = n17849 ^ n17846 ;
  assign n17850 = n17846 & ~n17849 ;
  assign n17855 = n17854 ^ n17850 ;
  assign n17839 = n3391 & n10155 ;
  assign n17838 = x126 & n3387 ;
  assign n17840 = n17839 ^ n17838 ;
  assign n17841 = n17840 ^ x35 ;
  assign n17837 = x127 & n3395 ;
  assign n17842 = n17841 ^ n17837 ;
  assign n17831 = x123 & n3932 ;
  assign n17830 = x125 & n3935 ;
  assign n17832 = n17831 ^ n17830 ;
  assign n17833 = n17832 ^ x38 ;
  assign n17829 = n3936 & n10416 ;
  assign n17834 = n17833 ^ n17829 ;
  assign n17828 = x124 & n3940 ;
  assign n17835 = n17834 ^ n17828 ;
  assign n17817 = x120 & n4482 ;
  assign n17816 = x122 & n4478 ;
  assign n17818 = n17817 ^ n17816 ;
  assign n17819 = n17818 ^ x41 ;
  assign n17815 = n4479 & ~n9261 ;
  assign n17820 = n17819 ^ n17815 ;
  assign n17814 = x121 & n4475 ;
  assign n17821 = n17820 ^ n17814 ;
  assign n17810 = n17669 ^ n17656 ;
  assign n17811 = ~n17661 & ~n17810 ;
  assign n17812 = n17811 ^ n17656 ;
  assign n17804 = x117 & n5113 ;
  assign n17803 = x119 & n5116 ;
  assign n17805 = n17804 ^ n17803 ;
  assign n17806 = n17805 ^ x44 ;
  assign n17802 = n5117 & n8405 ;
  assign n17807 = n17806 ^ n17802 ;
  assign n17801 = x118 & n5121 ;
  assign n17808 = n17807 ^ n17801 ;
  assign n17789 = x114 & n5981 ;
  assign n17788 = x116 & n5748 ;
  assign n17790 = n17789 ^ n17788 ;
  assign n17791 = n17790 ^ x47 ;
  assign n17787 = n5749 & ~n7604 ;
  assign n17792 = n17791 ^ n17787 ;
  assign n17786 = x115 & n5755 ;
  assign n17793 = n17792 ^ n17786 ;
  assign n17779 = n17636 ^ n17624 ;
  assign n17780 = ~n17638 & ~n17779 ;
  assign n17781 = n17780 ^ n17636 ;
  assign n17773 = x102 & n8750 ;
  assign n17772 = x104 & n8746 ;
  assign n17774 = n17773 ^ n17772 ;
  assign n17775 = n17774 ^ x59 ;
  assign n17771 = ~n4830 & n8747 ;
  assign n17776 = n17775 ^ n17771 ;
  assign n17770 = x103 & n8743 ;
  assign n17777 = n17776 ^ n17770 ;
  assign n17767 = x97 & n11895 ;
  assign n17766 = x98 & n9956 ;
  assign n17768 = n17767 ^ n17766 ;
  assign n17763 = n4223 & n9652 ;
  assign n17761 = x99 & n9655 ;
  assign n17754 = x96 ^ x32 ;
  assign n17757 = n17627 & ~n17754 ;
  assign n17758 = n17757 ^ x96 ;
  assign n17759 = n12206 & n17758 ;
  assign n17752 = x101 & n9651 ;
  assign n17753 = n17752 ^ x62 ;
  assign n17760 = n17759 ^ n17753 ;
  assign n17762 = n17761 ^ n17760 ;
  assign n17764 = n17763 ^ n17762 ;
  assign n17751 = x100 & n9648 ;
  assign n17765 = n17764 ^ n17751 ;
  assign n17769 = n17768 ^ n17765 ;
  assign n17778 = n17777 ^ n17769 ;
  assign n17782 = n17781 ^ n17778 ;
  assign n17748 = ~n5459 & n7951 ;
  assign n17746 = x105 & n7954 ;
  assign n17742 = n17639 ^ n17615 ;
  assign n17743 = ~n17621 & n17742 ;
  assign n17744 = n17743 ^ n17639 ;
  assign n17740 = x107 & n7950 ;
  assign n17741 = n17740 ^ x56 ;
  assign n17745 = n17744 ^ n17741 ;
  assign n17747 = n17746 ^ n17745 ;
  assign n17749 = n17748 ^ n17747 ;
  assign n17739 = x106 & n7947 ;
  assign n17750 = n17749 ^ n17739 ;
  assign n17783 = n17782 ^ n17750 ;
  assign n17736 = n6145 & n7187 ;
  assign n17734 = x108 & n7183 ;
  assign n17730 = n17640 ^ n17604 ;
  assign n17731 = n17609 & n17730 ;
  assign n17732 = n17731 ^ n17604 ;
  assign n17728 = x110 & n7186 ;
  assign n17729 = n17728 ^ x53 ;
  assign n17733 = n17732 ^ n17729 ;
  assign n17735 = n17734 ^ n17733 ;
  assign n17737 = n17736 ^ n17735 ;
  assign n17727 = x109 & n7191 ;
  assign n17738 = n17737 ^ n17727 ;
  assign n17784 = n17783 ^ n17738 ;
  assign n17724 = n6445 & ~n6849 ;
  assign n17722 = x111 & n6687 ;
  assign n17718 = n17641 ^ n17591 ;
  assign n17719 = ~n17596 & n17718 ;
  assign n17720 = n17719 ^ n17591 ;
  assign n17716 = x113 & n6444 ;
  assign n17717 = n17716 ^ x50 ;
  assign n17721 = n17720 ^ n17717 ;
  assign n17723 = n17722 ^ n17721 ;
  assign n17725 = n17724 ^ n17723 ;
  assign n17715 = x112 & n6449 ;
  assign n17726 = n17725 ^ n17715 ;
  assign n17785 = n17784 ^ n17726 ;
  assign n17794 = n17793 ^ n17785 ;
  assign n17712 = n17642 ^ n17578 ;
  assign n17713 = n17583 & ~n17712 ;
  assign n17714 = n17713 ^ n17578 ;
  assign n17795 = n17794 ^ n17714 ;
  assign n17797 = n17795 ^ n17655 ;
  assign n17796 = n17795 ^ n17643 ;
  assign n17798 = n17797 ^ n17796 ;
  assign n17799 = ~n17652 & ~n17798 ;
  assign n17800 = n17799 ^ n17796 ;
  assign n17809 = n17808 ^ n17800 ;
  assign n17813 = n17812 ^ n17809 ;
  assign n17822 = n17821 ^ n17813 ;
  assign n17823 = n17822 ^ n17682 ;
  assign n17824 = n17823 ^ n17673 ;
  assign n17825 = n17824 ^ n17822 ;
  assign n17826 = ~n17674 & ~n17825 ;
  assign n17827 = n17826 ^ n17823 ;
  assign n17836 = n17835 ^ n17827 ;
  assign n17852 = n17842 ^ n17836 ;
  assign n17843 = ~n17836 & n17842 ;
  assign n17853 = n17852 ^ n17843 ;
  assign n17856 = n17855 ^ n17853 ;
  assign n17851 = n17850 ^ n17843 ;
  assign n17857 = n17856 ^ n17851 ;
  assign n17709 = n17567 ^ n17564 ;
  assign n17710 = ~n17707 & ~n17709 ;
  assign n17711 = n17710 ^ n17564 ;
  assign n17858 = n17857 ^ n17711 ;
  assign n17992 = x127 & n3386 ;
  assign n17993 = n17992 ^ n3384 ;
  assign n17998 = n3051 & n11285 ;
  assign n17999 = n17998 ^ n17992 ;
  assign n18000 = n17993 & ~n17999 ;
  assign n18001 = n18000 ^ x34 ;
  assign n17981 = x124 & n3932 ;
  assign n17980 = x126 & n3935 ;
  assign n17982 = n17981 ^ n17980 ;
  assign n17983 = n17982 ^ x38 ;
  assign n17979 = n3936 & n10461 ;
  assign n17984 = n17983 ^ n17979 ;
  assign n17978 = x125 & n3940 ;
  assign n17985 = n17984 ^ n17978 ;
  assign n17967 = x121 & n4482 ;
  assign n17966 = x123 & n4478 ;
  assign n17968 = n17967 ^ n17966 ;
  assign n17969 = n17968 ^ x41 ;
  assign n17965 = n4479 & ~n9804 ;
  assign n17970 = n17969 ^ n17965 ;
  assign n17964 = x122 & n4475 ;
  assign n17971 = n17970 ^ n17964 ;
  assign n17960 = n17808 ^ n17795 ;
  assign n17961 = n17800 & ~n17960 ;
  assign n17962 = n17961 ^ n17795 ;
  assign n17954 = x118 & n5113 ;
  assign n17953 = x120 & n5116 ;
  assign n17955 = n17954 ^ n17953 ;
  assign n17956 = n17955 ^ x44 ;
  assign n17952 = n5117 & n8904 ;
  assign n17957 = n17956 ^ n17952 ;
  assign n17951 = x119 & n5121 ;
  assign n17958 = n17957 ^ n17951 ;
  assign n17944 = x115 & n5981 ;
  assign n17943 = x117 & n5748 ;
  assign n17945 = n17944 ^ n17943 ;
  assign n17946 = n17945 ^ x47 ;
  assign n17942 = n5749 & ~n7860 ;
  assign n17947 = n17946 ^ n17942 ;
  assign n17941 = x116 & n5755 ;
  assign n17948 = n17947 ^ n17941 ;
  assign n17927 = x103 & n8750 ;
  assign n17926 = x105 & n8746 ;
  assign n17928 = n17927 ^ n17926 ;
  assign n17929 = n17928 ^ x59 ;
  assign n17925 = ~n5034 & n8747 ;
  assign n17930 = n17929 ^ n17925 ;
  assign n17924 = x104 & n8743 ;
  assign n17931 = n17930 ^ n17924 ;
  assign n17922 = x101 & n9648 ;
  assign n17914 = n17768 ^ n17759 ;
  assign n17915 = ~n17765 & ~n17914 ;
  assign n17916 = n17915 ^ n17768 ;
  assign n17908 = n9956 ^ x98 ;
  assign n17904 = ~x99 & n9956 ;
  assign n17905 = n17904 ^ n17767 ;
  assign n17909 = n17905 ^ n12206 ;
  assign n17910 = n17908 & n17909 ;
  assign n17911 = n17910 ^ n3485 ;
  assign n17906 = x98 & n17905 ;
  assign n17907 = n17906 ^ n17767 ;
  assign n17912 = n17911 ^ n17907 ;
  assign n17913 = n17912 ^ n3485 ;
  assign n17917 = n17916 ^ n17913 ;
  assign n17918 = n17917 ^ x62 ;
  assign n17903 = x100 & n9655 ;
  assign n17919 = n17918 ^ n17903 ;
  assign n17902 = x102 & n9651 ;
  assign n17920 = n17919 ^ n17902 ;
  assign n17901 = n4425 & n9652 ;
  assign n17921 = n17920 ^ n17901 ;
  assign n17923 = n17922 ^ n17921 ;
  assign n17932 = n17931 ^ n17923 ;
  assign n17898 = n5687 & n7951 ;
  assign n17896 = x106 & n7954 ;
  assign n17892 = n17781 ^ n17777 ;
  assign n17893 = n17778 & n17892 ;
  assign n17894 = n17893 ^ n17781 ;
  assign n17890 = x108 & n7950 ;
  assign n17891 = n17890 ^ x56 ;
  assign n17895 = n17894 ^ n17891 ;
  assign n17897 = n17896 ^ n17895 ;
  assign n17899 = n17898 ^ n17897 ;
  assign n17889 = x107 & n7947 ;
  assign n17900 = n17899 ^ n17889 ;
  assign n17933 = n17932 ^ n17900 ;
  assign n17887 = x110 & n7191 ;
  assign n17885 = ~n6370 & n7187 ;
  assign n17883 = x109 & n7183 ;
  assign n17879 = n17782 ^ n17744 ;
  assign n17880 = ~n17750 & ~n17879 ;
  assign n17881 = n17880 ^ n17782 ;
  assign n17877 = x111 & n7186 ;
  assign n17878 = n17877 ^ x53 ;
  assign n17882 = n17881 ^ n17878 ;
  assign n17884 = n17883 ^ n17882 ;
  assign n17886 = n17885 ^ n17884 ;
  assign n17888 = n17887 ^ n17886 ;
  assign n17934 = n17933 ^ n17888 ;
  assign n17875 = x113 & n6449 ;
  assign n17873 = n6445 & ~n7108 ;
  assign n17871 = x112 & n6687 ;
  assign n17867 = n17783 ^ n17732 ;
  assign n17868 = ~n17738 & ~n17867 ;
  assign n17869 = n17868 ^ n17783 ;
  assign n17865 = x114 & n6444 ;
  assign n17866 = n17865 ^ x50 ;
  assign n17870 = n17869 ^ n17866 ;
  assign n17872 = n17871 ^ n17870 ;
  assign n17874 = n17873 ^ n17872 ;
  assign n17876 = n17875 ^ n17874 ;
  assign n17935 = n17934 ^ n17876 ;
  assign n17936 = n17935 ^ n17784 ;
  assign n17937 = n17936 ^ n17720 ;
  assign n17938 = n17937 ^ n17935 ;
  assign n17939 = ~n17726 & ~n17938 ;
  assign n17940 = n17939 ^ n17936 ;
  assign n17949 = n17948 ^ n17940 ;
  assign n17862 = n17793 ^ n17714 ;
  assign n17863 = ~n17794 & n17862 ;
  assign n17864 = n17863 ^ n17793 ;
  assign n17950 = n17949 ^ n17864 ;
  assign n17959 = n17958 ^ n17950 ;
  assign n17963 = n17962 ^ n17959 ;
  assign n17972 = n17971 ^ n17963 ;
  assign n17973 = n17972 ^ n17821 ;
  assign n17974 = n17973 ^ n17812 ;
  assign n17975 = n17974 ^ n17972 ;
  assign n17976 = n17813 & ~n17975 ;
  assign n17977 = n17976 ^ n17973 ;
  assign n17986 = n17985 ^ n17977 ;
  assign n17988 = n17986 ^ n17822 ;
  assign n17987 = n17986 ^ n17835 ;
  assign n17989 = n17988 ^ n17987 ;
  assign n17990 = ~n17827 & ~n17989 ;
  assign n17991 = n17990 ^ n17988 ;
  assign n18002 = n18001 ^ n17991 ;
  assign n18003 = n18002 ^ n17851 ;
  assign n17859 = n17854 ^ n17852 ;
  assign n17860 = n17852 ^ n17711 ;
  assign n17861 = n17859 & n17860 ;
  assign n18004 = n18003 ^ n17861 ;
  assign n18178 = n18001 ^ n17986 ;
  assign n18179 = ~n17991 & n18178 ;
  assign n18180 = n18179 ^ n17986 ;
  assign n18174 = n17985 ^ n17972 ;
  assign n18175 = n17977 & n18174 ;
  assign n18176 = n18175 ^ n17972 ;
  assign n18168 = x125 & n3932 ;
  assign n18167 = x127 & n3935 ;
  assign n18169 = n18168 ^ n18167 ;
  assign n18170 = n18169 ^ x38 ;
  assign n18166 = n3936 & n10986 ;
  assign n18171 = n18170 ^ n18166 ;
  assign n18165 = x126 & n3940 ;
  assign n18172 = n18171 ^ n18165 ;
  assign n18158 = x122 & n4482 ;
  assign n18157 = x124 & n4478 ;
  assign n18159 = n18158 ^ n18157 ;
  assign n18160 = n18159 ^ x41 ;
  assign n18156 = n4479 & n10117 ;
  assign n18161 = n18160 ^ n18156 ;
  assign n18155 = x123 & n4475 ;
  assign n18162 = n18161 ^ n18155 ;
  assign n18148 = x119 & n5113 ;
  assign n18147 = x121 & n5116 ;
  assign n18149 = n18148 ^ n18147 ;
  assign n18150 = n18149 ^ x44 ;
  assign n18146 = n5117 & n8979 ;
  assign n18151 = n18150 ^ n18146 ;
  assign n18145 = x120 & n5121 ;
  assign n18152 = n18151 ^ n18145 ;
  assign n18141 = n17948 ^ n17935 ;
  assign n18142 = ~n17940 & n18141 ;
  assign n18143 = n18142 ^ n17935 ;
  assign n18135 = x116 & n5981 ;
  assign n18134 = x118 & n5748 ;
  assign n18136 = n18135 ^ n18134 ;
  assign n18137 = n18136 ^ x47 ;
  assign n18133 = n5749 & ~n8140 ;
  assign n18138 = n18137 ^ n18133 ;
  assign n18132 = x117 & n5755 ;
  assign n18139 = n18138 ^ n18132 ;
  assign n18126 = x113 & n6687 ;
  assign n18125 = x115 & n6444 ;
  assign n18127 = n18126 ^ n18125 ;
  assign n18128 = n18127 ^ x50 ;
  assign n18124 = n6445 & ~n7353 ;
  assign n18129 = n18128 ^ n18124 ;
  assign n18123 = x114 & n6449 ;
  assign n18130 = n18129 ^ n18123 ;
  assign n18111 = x110 & n7183 ;
  assign n18110 = x112 & n7186 ;
  assign n18112 = n18111 ^ n18110 ;
  assign n18113 = n18112 ^ x53 ;
  assign n18109 = ~n6616 & n7187 ;
  assign n18114 = n18113 ^ n18109 ;
  assign n18108 = x111 & n7191 ;
  assign n18115 = n18114 ^ n18108 ;
  assign n18098 = x101 & n9655 ;
  assign n18097 = x103 & n9651 ;
  assign n18099 = n18098 ^ n18097 ;
  assign n18100 = n18099 ^ x62 ;
  assign n18096 = ~n4624 & n9652 ;
  assign n18101 = n18100 ^ n18096 ;
  assign n18095 = x102 & n9648 ;
  assign n18102 = n18101 ^ n18095 ;
  assign n18103 = n18102 ^ x35 ;
  assign n18091 = x100 ^ x98 ;
  assign n18092 = ~n11895 & n18091 ;
  assign n18093 = n18092 ^ n3485 ;
  assign n18094 = n12206 & n18093 ;
  assign n18104 = n18103 ^ n18094 ;
  assign n18088 = ~n17910 & n17916 ;
  assign n18089 = ~n17907 & n18088 ;
  assign n18090 = n18089 ^ n17910 ;
  assign n18105 = n18104 ^ n18090 ;
  assign n18078 = x104 & n8750 ;
  assign n18077 = x106 & n8746 ;
  assign n18079 = n18078 ^ n18077 ;
  assign n18080 = n18079 ^ x59 ;
  assign n18076 = ~n5257 & n8747 ;
  assign n18081 = n18080 ^ n18076 ;
  assign n18075 = x105 & n8743 ;
  assign n18082 = n18081 ^ n18075 ;
  assign n18083 = n18082 ^ n17931 ;
  assign n18084 = n18083 ^ n17917 ;
  assign n18085 = n18084 ^ n18082 ;
  assign n18086 = ~n17923 & n18085 ;
  assign n18087 = n18086 ^ n18083 ;
  assign n18106 = n18105 ^ n18087 ;
  assign n18072 = n17932 ^ n17894 ;
  assign n18073 = ~n17900 & n18072 ;
  assign n18065 = x107 & n7954 ;
  assign n18064 = x109 & n7950 ;
  assign n18066 = n18065 ^ n18064 ;
  assign n18067 = n18066 ^ x56 ;
  assign n18063 = n5912 & n7951 ;
  assign n18068 = n18067 ^ n18063 ;
  assign n18062 = x108 & n7947 ;
  assign n18069 = n18068 ^ n18062 ;
  assign n18070 = n18069 ^ n17932 ;
  assign n18074 = n18073 ^ n18070 ;
  assign n18107 = n18106 ^ n18074 ;
  assign n18116 = n18115 ^ n18107 ;
  assign n18059 = n17933 ^ n17881 ;
  assign n18060 = n17888 & ~n18059 ;
  assign n18061 = n18060 ^ n17933 ;
  assign n18117 = n18116 ^ n18061 ;
  assign n18119 = n18117 ^ n17934 ;
  assign n18118 = n18117 ^ n17869 ;
  assign n18120 = n18119 ^ n18118 ;
  assign n18121 = n17876 & n18120 ;
  assign n18122 = n18121 ^ n18119 ;
  assign n18131 = n18130 ^ n18122 ;
  assign n18140 = n18139 ^ n18131 ;
  assign n18144 = n18143 ^ n18140 ;
  assign n18153 = n18152 ^ n18144 ;
  assign n18056 = n17958 ^ n17864 ;
  assign n18057 = n17950 & n18056 ;
  assign n18058 = n18057 ^ n17958 ;
  assign n18154 = n18153 ^ n18058 ;
  assign n18163 = n18162 ^ n18154 ;
  assign n18053 = n17971 ^ n17962 ;
  assign n18054 = ~n17963 & ~n18053 ;
  assign n18055 = n18054 ^ n17971 ;
  assign n18164 = n18163 ^ n18055 ;
  assign n18173 = n18172 ^ n18164 ;
  assign n18177 = n18176 ^ n18173 ;
  assign n18181 = n18180 ^ n18177 ;
  assign n18005 = n18002 ^ n17842 ;
  assign n18006 = n18005 ^ n18002 ;
  assign n18007 = n18002 ^ n17836 ;
  assign n18008 = n18007 ^ n18002 ;
  assign n18009 = ~n18006 & n18008 ;
  assign n18010 = n18009 ^ n18002 ;
  assign n18018 = n18008 ^ n18006 ;
  assign n18019 = n18018 ^ n18002 ;
  assign n18012 = n18002 ^ n17846 ;
  assign n18011 = n18002 ^ n17849 ;
  assign n18013 = n18012 ^ n18011 ;
  assign n18014 = n18012 ^ n18005 ;
  assign n18015 = n18014 ^ n18007 ;
  assign n18016 = n18015 ^ n18002 ;
  assign n18017 = n18013 & ~n18016 ;
  assign n18020 = n18019 ^ n18017 ;
  assign n18021 = n18010 & ~n18020 ;
  assign n18022 = n18021 ^ n18002 ;
  assign n18025 = n18002 ^ n17854 ;
  assign n18026 = n18025 ^ n17850 ;
  assign n18034 = n18002 & ~n18026 ;
  assign n18027 = n18026 ^ n18005 ;
  assign n18028 = n18027 ^ n17836 ;
  assign n18029 = n18028 ^ n18025 ;
  assign n18030 = n18029 ^ n18026 ;
  assign n18036 = n18034 ^ n18030 ;
  assign n18037 = ~n17842 & n18036 ;
  assign n18044 = n18037 ^ n18034 ;
  assign n18038 = n18037 ^ n18029 ;
  assign n18039 = n18026 ^ n18007 ;
  assign n18040 = n18039 ^ n17842 ;
  assign n18041 = n18040 ^ n18026 ;
  assign n18042 = n18041 ^ n18002 ;
  assign n18043 = ~n18038 & ~n18042 ;
  assign n18045 = n18044 ^ n18043 ;
  assign n18048 = n18045 ^ n18025 ;
  assign n18049 = n18048 ^ n18030 ;
  assign n18050 = ~n17711 & ~n18049 ;
  assign n18051 = ~n18022 & n18050 ;
  assign n18052 = n18051 ^ n18022 ;
  assign n18182 = n18181 ^ n18052 ;
  assign n18307 = n3936 & n10155 ;
  assign n18306 = x126 & n3932 ;
  assign n18308 = n18307 ^ n18306 ;
  assign n18309 = n18308 ^ x38 ;
  assign n18305 = x127 & n3940 ;
  assign n18310 = n18309 ^ n18305 ;
  assign n18298 = x123 & n4482 ;
  assign n18297 = x125 & n4478 ;
  assign n18299 = n18298 ^ n18297 ;
  assign n18300 = n18299 ^ x41 ;
  assign n18296 = n4479 & n10416 ;
  assign n18301 = n18300 ^ n18296 ;
  assign n18295 = x124 & n4475 ;
  assign n18302 = n18301 ^ n18295 ;
  assign n18288 = x120 & n5113 ;
  assign n18287 = x122 & n5116 ;
  assign n18289 = n18288 ^ n18287 ;
  assign n18290 = n18289 ^ x44 ;
  assign n18286 = n5117 & ~n9261 ;
  assign n18291 = n18290 ^ n18286 ;
  assign n18285 = x121 & n5121 ;
  assign n18292 = n18291 ^ n18285 ;
  assign n18278 = x117 & n5981 ;
  assign n18277 = x119 & n5748 ;
  assign n18279 = n18278 ^ n18277 ;
  assign n18280 = n18279 ^ x47 ;
  assign n18276 = n5749 & n8405 ;
  assign n18281 = n18280 ^ n18276 ;
  assign n18275 = x118 & n5755 ;
  assign n18282 = n18281 ^ n18275 ;
  assign n18260 = x102 & n9655 ;
  assign n18259 = x104 & n9651 ;
  assign n18261 = n18260 ^ n18259 ;
  assign n18262 = n18261 ^ x62 ;
  assign n18258 = ~n4830 & n9652 ;
  assign n18263 = n18262 ^ n18258 ;
  assign n18257 = x103 & n9648 ;
  assign n18264 = n18263 ^ n18257 ;
  assign n18254 = x100 & n11895 ;
  assign n18253 = x101 & n9956 ;
  assign n18255 = n18254 ^ n18253 ;
  assign n18247 = x99 ^ x35 ;
  assign n18250 = n18093 & ~n18247 ;
  assign n18251 = n18250 ^ x99 ;
  assign n18252 = n12206 & n18251 ;
  assign n18256 = n18255 ^ n18252 ;
  assign n18265 = n18264 ^ n18256 ;
  assign n18244 = ~n5459 & n8747 ;
  assign n18242 = x105 & n8750 ;
  assign n18238 = n18102 ^ n18090 ;
  assign n18239 = ~n18104 & ~n18238 ;
  assign n18240 = n18239 ^ n18102 ;
  assign n18236 = x107 & n8746 ;
  assign n18237 = n18236 ^ x59 ;
  assign n18241 = n18240 ^ n18237 ;
  assign n18243 = n18242 ^ n18241 ;
  assign n18245 = n18244 ^ n18243 ;
  assign n18235 = x106 & n8743 ;
  assign n18246 = n18245 ^ n18235 ;
  assign n18266 = n18265 ^ n18246 ;
  assign n18232 = n6145 & n7951 ;
  assign n18230 = x108 & n7954 ;
  assign n18226 = n18105 ^ n18082 ;
  assign n18227 = n18087 & n18226 ;
  assign n18228 = n18227 ^ n18082 ;
  assign n18224 = x110 & n7950 ;
  assign n18225 = n18224 ^ x56 ;
  assign n18229 = n18228 ^ n18225 ;
  assign n18231 = n18230 ^ n18229 ;
  assign n18233 = n18232 ^ n18231 ;
  assign n18223 = x109 & n7947 ;
  assign n18234 = n18233 ^ n18223 ;
  assign n18267 = n18266 ^ n18234 ;
  assign n18220 = ~n6849 & n7187 ;
  assign n18218 = x111 & n7183 ;
  assign n18214 = n18106 ^ n18069 ;
  assign n18215 = n18074 & n18214 ;
  assign n18216 = n18215 ^ n18069 ;
  assign n18212 = x113 & n7186 ;
  assign n18213 = n18212 ^ x53 ;
  assign n18217 = n18216 ^ n18213 ;
  assign n18219 = n18218 ^ n18217 ;
  assign n18221 = n18220 ^ n18219 ;
  assign n18211 = x112 & n7191 ;
  assign n18222 = n18221 ^ n18211 ;
  assign n18268 = n18267 ^ n18222 ;
  assign n18208 = n18115 ^ n18061 ;
  assign n18209 = n18116 & n18208 ;
  assign n18201 = x114 & n6687 ;
  assign n18200 = x116 & n6444 ;
  assign n18202 = n18201 ^ n18200 ;
  assign n18203 = n18202 ^ x50 ;
  assign n18199 = n6445 & ~n7604 ;
  assign n18204 = n18203 ^ n18199 ;
  assign n18198 = x115 & n6449 ;
  assign n18205 = n18204 ^ n18198 ;
  assign n18206 = n18205 ^ n18115 ;
  assign n18210 = n18209 ^ n18206 ;
  assign n18269 = n18268 ^ n18210 ;
  assign n18271 = n18269 ^ n18117 ;
  assign n18270 = n18269 ^ n18130 ;
  assign n18272 = n18271 ^ n18270 ;
  assign n18273 = ~n18122 & n18272 ;
  assign n18274 = n18273 ^ n18271 ;
  assign n18283 = n18282 ^ n18274 ;
  assign n18195 = n18143 ^ n18139 ;
  assign n18196 = n18140 & n18195 ;
  assign n18197 = n18196 ^ n18143 ;
  assign n18284 = n18283 ^ n18197 ;
  assign n18293 = n18292 ^ n18284 ;
  assign n18192 = n18152 ^ n18058 ;
  assign n18193 = ~n18153 & n18192 ;
  assign n18194 = n18193 ^ n18152 ;
  assign n18294 = n18293 ^ n18194 ;
  assign n18303 = n18302 ^ n18294 ;
  assign n18189 = n18162 ^ n18055 ;
  assign n18190 = ~n18163 & n18189 ;
  assign n18191 = n18190 ^ n18162 ;
  assign n18304 = n18303 ^ n18191 ;
  assign n18311 = n18310 ^ n18304 ;
  assign n18186 = n18176 ^ n18172 ;
  assign n18187 = n18173 & n18186 ;
  assign n18188 = n18187 ^ n18176 ;
  assign n18312 = n18311 ^ n18188 ;
  assign n18183 = n18180 ^ n18052 ;
  assign n18184 = ~n18181 & ~n18183 ;
  assign n18185 = n18184 ^ n18180 ;
  assign n18313 = n18312 ^ n18185 ;
  assign n18434 = x127 & n3931 ;
  assign n18435 = n18434 ^ n3929 ;
  assign n18440 = n3542 & n11285 ;
  assign n18441 = n18440 ^ n18434 ;
  assign n18442 = n18435 & ~n18441 ;
  assign n18443 = n18442 ^ x37 ;
  assign n18423 = x124 & n4482 ;
  assign n18422 = x126 & n4478 ;
  assign n18424 = n18423 ^ n18422 ;
  assign n18425 = n18424 ^ x41 ;
  assign n18421 = n4479 & n10461 ;
  assign n18426 = n18425 ^ n18421 ;
  assign n18420 = x125 & n4475 ;
  assign n18427 = n18426 ^ n18420 ;
  assign n18413 = x121 & n5113 ;
  assign n18412 = x123 & n5116 ;
  assign n18414 = n18413 ^ n18412 ;
  assign n18415 = n18414 ^ x44 ;
  assign n18411 = n5117 & ~n9804 ;
  assign n18416 = n18415 ^ n18411 ;
  assign n18410 = x122 & n5121 ;
  assign n18417 = n18416 ^ n18410 ;
  assign n18406 = n18282 ^ n18269 ;
  assign n18407 = ~n18274 & ~n18406 ;
  assign n18408 = n18407 ^ n18269 ;
  assign n18400 = x118 & n5981 ;
  assign n18399 = x120 & n5748 ;
  assign n18401 = n18400 ^ n18399 ;
  assign n18402 = n18401 ^ x47 ;
  assign n18398 = n5749 & n8904 ;
  assign n18403 = n18402 ^ n18398 ;
  assign n18397 = x119 & n5755 ;
  assign n18404 = n18403 ^ n18397 ;
  assign n18385 = x115 & n6687 ;
  assign n18384 = x117 & n6444 ;
  assign n18386 = n18385 ^ n18384 ;
  assign n18387 = n18386 ^ x50 ;
  assign n18383 = n6445 & ~n7860 ;
  assign n18388 = n18387 ^ n18383 ;
  assign n18382 = x116 & n6449 ;
  assign n18389 = n18388 ^ n18382 ;
  assign n18376 = x112 & n7183 ;
  assign n18375 = x114 & n7186 ;
  assign n18377 = n18376 ^ n18375 ;
  assign n18378 = n18377 ^ x53 ;
  assign n18374 = ~n7108 & n7187 ;
  assign n18379 = n18378 ^ n18374 ;
  assign n18373 = x113 & n7191 ;
  assign n18380 = n18379 ^ n18373 ;
  assign n18365 = x103 & n9655 ;
  assign n18364 = x105 & n9651 ;
  assign n18366 = n18365 ^ n18364 ;
  assign n18367 = n18366 ^ x62 ;
  assign n18363 = ~n5034 & n9652 ;
  assign n18368 = n18367 ^ n18363 ;
  assign n18362 = x104 & n9648 ;
  assign n18369 = n18368 ^ n18362 ;
  assign n18356 = x106 & n8750 ;
  assign n18355 = x108 & n8746 ;
  assign n18357 = n18356 ^ n18355 ;
  assign n18358 = n18357 ^ x59 ;
  assign n18354 = n5687 & n8747 ;
  assign n18359 = n18358 ^ n18354 ;
  assign n18353 = x107 & n8743 ;
  assign n18360 = n18359 ^ n18353 ;
  assign n18348 = x63 & n3829 ;
  assign n4025 = x102 ^ x101 ;
  assign n18349 = n18348 ^ n4025 ;
  assign n18350 = ~n9956 & n18349 ;
  assign n18351 = n18350 ^ n4025 ;
  assign n18341 = n18264 ^ n18255 ;
  assign n18342 = n18256 & ~n18341 ;
  assign n18343 = n18342 ^ n18264 ;
  assign n18352 = n18351 ^ n18343 ;
  assign n18361 = n18360 ^ n18352 ;
  assign n18370 = n18369 ^ n18361 ;
  assign n18339 = x110 & n7947 ;
  assign n18337 = ~n6370 & n7951 ;
  assign n18335 = x109 & n7954 ;
  assign n18331 = n18265 ^ n18240 ;
  assign n18332 = ~n18246 & ~n18331 ;
  assign n18333 = n18332 ^ n18265 ;
  assign n18329 = x111 & n7950 ;
  assign n18330 = n18329 ^ x56 ;
  assign n18334 = n18333 ^ n18330 ;
  assign n18336 = n18335 ^ n18334 ;
  assign n18338 = n18337 ^ n18336 ;
  assign n18340 = n18339 ^ n18338 ;
  assign n18371 = n18370 ^ n18340 ;
  assign n18326 = n18266 ^ n18228 ;
  assign n18327 = ~n18234 & ~n18326 ;
  assign n18328 = n18327 ^ n18266 ;
  assign n18372 = n18371 ^ n18328 ;
  assign n18381 = n18380 ^ n18372 ;
  assign n18390 = n18389 ^ n18381 ;
  assign n18323 = n18267 ^ n18216 ;
  assign n18324 = ~n18222 & ~n18323 ;
  assign n18325 = n18324 ^ n18267 ;
  assign n18391 = n18390 ^ n18325 ;
  assign n18393 = n18391 ^ n18205 ;
  assign n18392 = n18391 ^ n18268 ;
  assign n18394 = n18393 ^ n18392 ;
  assign n18395 = n18210 & ~n18394 ;
  assign n18396 = n18395 ^ n18393 ;
  assign n18405 = n18404 ^ n18396 ;
  assign n18409 = n18408 ^ n18405 ;
  assign n18418 = n18417 ^ n18409 ;
  assign n18320 = n18292 ^ n18197 ;
  assign n18321 = n18284 & n18320 ;
  assign n18322 = n18321 ^ n18292 ;
  assign n18419 = n18418 ^ n18322 ;
  assign n18428 = n18427 ^ n18419 ;
  assign n18429 = n18428 ^ n18302 ;
  assign n18430 = n18429 ^ n18428 ;
  assign n18431 = n18430 ^ n18194 ;
  assign n18432 = n18294 & n18431 ;
  assign n18433 = n18432 ^ n18429 ;
  assign n18444 = n18443 ^ n18433 ;
  assign n18317 = n18310 ^ n18191 ;
  assign n18318 = n18304 & n18317 ;
  assign n18319 = n18318 ^ n18310 ;
  assign n18445 = n18444 ^ n18319 ;
  assign n18314 = n18188 ^ n18185 ;
  assign n18315 = n18312 & n18314 ;
  assign n18316 = n18315 ^ n18185 ;
  assign n18446 = n18445 ^ n18316 ;
  assign n18578 = n18319 ^ n18316 ;
  assign n18579 = ~n18445 & n18578 ;
  assign n18580 = n18579 ^ n18319 ;
  assign n18573 = n18443 ^ n18428 ;
  assign n18574 = ~n18433 & ~n18573 ;
  assign n18575 = n18574 ^ n18428 ;
  assign n18567 = x122 & n5113 ;
  assign n18566 = x124 & n5116 ;
  assign n18568 = n18567 ^ n18566 ;
  assign n18569 = n18568 ^ x44 ;
  assign n18565 = n5117 & n10117 ;
  assign n18570 = n18569 ^ n18565 ;
  assign n18564 = x123 & n5121 ;
  assign n18571 = n18570 ^ n18564 ;
  assign n18555 = n18404 ^ n18391 ;
  assign n18556 = n18396 & n18555 ;
  assign n18557 = n18556 ^ n18391 ;
  assign n18549 = x119 & n5981 ;
  assign n18548 = x121 & n5748 ;
  assign n18550 = n18549 ^ n18548 ;
  assign n18551 = n18550 ^ x47 ;
  assign n18547 = n5749 & n8979 ;
  assign n18552 = n18551 ^ n18547 ;
  assign n18546 = x120 & n5755 ;
  assign n18553 = n18552 ^ n18546 ;
  assign n18539 = ~n18343 & ~n18351 ;
  assign n18535 = ~x102 & n9956 ;
  assign n18536 = n18535 ^ n18254 ;
  assign n18537 = x101 & n18536 ;
  assign n18538 = n18537 ^ n18254 ;
  assign n18540 = n18539 ^ n18538 ;
  assign n18525 = x104 & n9655 ;
  assign n18524 = x106 & n9651 ;
  assign n18526 = n18525 ^ n18524 ;
  assign n18527 = n18526 ^ x62 ;
  assign n18523 = ~n5257 & n9652 ;
  assign n18528 = n18527 ^ n18523 ;
  assign n18522 = x105 & n9648 ;
  assign n18529 = n18528 ^ n18522 ;
  assign n18517 = x63 & x102 ;
  assign n18518 = n18517 ^ x103 ;
  assign n18519 = ~n9956 & n18518 ;
  assign n18511 = n18255 ^ x103 ;
  assign n18520 = n18519 ^ n18511 ;
  assign n18521 = n18520 ^ x38 ;
  assign n18530 = n18529 ^ n18521 ;
  assign n18541 = n18540 ^ n18530 ;
  assign n18501 = x107 & n8750 ;
  assign n18500 = x109 & n8746 ;
  assign n18502 = n18501 ^ n18500 ;
  assign n18503 = n18502 ^ x59 ;
  assign n18499 = n5912 & n8747 ;
  assign n18504 = n18503 ^ n18499 ;
  assign n18498 = x108 & n8743 ;
  assign n18505 = n18504 ^ n18498 ;
  assign n18506 = n18505 ^ n18369 ;
  assign n18507 = n18506 ^ n18360 ;
  assign n18508 = n18507 ^ n18505 ;
  assign n18509 = n18361 & n18508 ;
  assign n18510 = n18509 ^ n18506 ;
  assign n18542 = n18541 ^ n18510 ;
  assign n18488 = x110 & n7954 ;
  assign n18487 = x112 & n7950 ;
  assign n18489 = n18488 ^ n18487 ;
  assign n18490 = n18489 ^ x56 ;
  assign n18486 = ~n6616 & n7951 ;
  assign n18491 = n18490 ^ n18486 ;
  assign n18485 = x111 & n7947 ;
  assign n18492 = n18491 ^ n18485 ;
  assign n18494 = n18492 ^ n18370 ;
  assign n18493 = n18492 ^ n18333 ;
  assign n18495 = n18494 ^ n18493 ;
  assign n18496 = n18340 & n18495 ;
  assign n18497 = n18496 ^ n18494 ;
  assign n18543 = n18542 ^ n18497 ;
  assign n18482 = n18380 ^ n18328 ;
  assign n18483 = n18372 & ~n18482 ;
  assign n18475 = x113 & n7183 ;
  assign n18474 = x115 & n7186 ;
  assign n18476 = n18475 ^ n18474 ;
  assign n18477 = n18476 ^ x53 ;
  assign n18473 = n7187 & ~n7353 ;
  assign n18478 = n18477 ^ n18473 ;
  assign n18472 = x114 & n7191 ;
  assign n18479 = n18478 ^ n18472 ;
  assign n18480 = n18479 ^ n18380 ;
  assign n18484 = n18483 ^ n18480 ;
  assign n18544 = n18543 ^ n18484 ;
  assign n18469 = n18389 ^ n18325 ;
  assign n18470 = ~n18390 & ~n18469 ;
  assign n18462 = x116 & n6687 ;
  assign n18461 = x118 & n6444 ;
  assign n18463 = n18462 ^ n18461 ;
  assign n18464 = n18463 ^ x50 ;
  assign n18460 = n6445 & ~n8140 ;
  assign n18465 = n18464 ^ n18460 ;
  assign n18459 = x117 & n6449 ;
  assign n18466 = n18465 ^ n18459 ;
  assign n18467 = n18466 ^ n18389 ;
  assign n18471 = n18470 ^ n18467 ;
  assign n18545 = n18544 ^ n18471 ;
  assign n18554 = n18553 ^ n18545 ;
  assign n18558 = n18557 ^ n18554 ;
  assign n18559 = n18558 ^ n18417 ;
  assign n18560 = n18559 ^ n18408 ;
  assign n18561 = n18560 ^ n18558 ;
  assign n18562 = n18409 & ~n18561 ;
  assign n18563 = n18562 ^ n18559 ;
  assign n18572 = n18571 ^ n18563 ;
  assign n18576 = n18575 ^ n18572 ;
  assign n18453 = x125 & n4482 ;
  assign n18452 = x127 & n4478 ;
  assign n18454 = n18453 ^ n18452 ;
  assign n18455 = n18454 ^ x41 ;
  assign n18451 = n4479 & n10986 ;
  assign n18456 = n18455 ^ n18451 ;
  assign n18450 = x126 & n4475 ;
  assign n18457 = n18456 ^ n18450 ;
  assign n18447 = n18427 ^ n18322 ;
  assign n18448 = n18419 & n18447 ;
  assign n18449 = n18448 ^ n18427 ;
  assign n18458 = n18457 ^ n18449 ;
  assign n18577 = n18576 ^ n18458 ;
  assign n18581 = n18580 ^ n18577 ;
  assign n18698 = n18580 ^ n18576 ;
  assign n18699 = n18577 & ~n18698 ;
  assign n18694 = n18572 & n18575 ;
  assign n18695 = n18694 ^ n18576 ;
  assign n18692 = n18449 & n18457 ;
  assign n18693 = n18692 ^ n18458 ;
  assign n18696 = n18695 ^ n18693 ;
  assign n18687 = n4479 & n10155 ;
  assign n18686 = x126 & n4482 ;
  assign n18688 = n18687 ^ n18686 ;
  assign n18689 = n18688 ^ x41 ;
  assign n18685 = x127 & n4475 ;
  assign n18690 = n18689 ^ n18685 ;
  assign n18676 = n5117 & n10416 ;
  assign n18674 = x123 & n5113 ;
  assign n18670 = x121 & n5755 ;
  assign n18668 = n5749 & ~n9261 ;
  assign n18664 = x120 & n5981 ;
  assign n18663 = x122 & n5748 ;
  assign n18665 = n18664 ^ n18663 ;
  assign n18666 = n18665 ^ x47 ;
  assign n18659 = n18543 ^ n18479 ;
  assign n18660 = n18484 & ~n18659 ;
  assign n18661 = n18660 ^ n18479 ;
  assign n18657 = x118 & n6449 ;
  assign n18652 = x117 & n6687 ;
  assign n18651 = x119 & n6444 ;
  assign n18653 = n18652 ^ n18651 ;
  assign n18654 = n18653 ^ x50 ;
  assign n18650 = n6445 & n8405 ;
  assign n18655 = n18654 ^ n18650 ;
  assign n18641 = x108 & n8750 ;
  assign n18640 = x110 & n8746 ;
  assign n18642 = n18641 ^ n18640 ;
  assign n18643 = n18642 ^ x59 ;
  assign n18639 = n6145 & n8747 ;
  assign n18644 = n18643 ^ n18639 ;
  assign n18638 = x109 & n8743 ;
  assign n18645 = n18644 ^ n18638 ;
  assign n18632 = x105 & n9655 ;
  assign n18631 = x107 & n9651 ;
  assign n18633 = n18632 ^ n18631 ;
  assign n18634 = n18633 ^ x62 ;
  assign n18630 = ~n5459 & n9652 ;
  assign n18635 = n18634 ^ n18630 ;
  assign n18629 = x106 & n9648 ;
  assign n18636 = n18635 ^ n18629 ;
  assign n18625 = n18255 ^ x38 ;
  assign n18626 = ~n18520 & ~n18625 ;
  assign n18627 = n18626 ^ x38 ;
  assign n18621 = x63 & x103 ;
  assign n18622 = n18621 ^ x104 ;
  assign n18623 = ~n9956 & n18622 ;
  assign n18624 = n18623 ^ x104 ;
  assign n18628 = n18627 ^ n18624 ;
  assign n18637 = n18636 ^ n18628 ;
  assign n18646 = n18645 ^ n18637 ;
  assign n18616 = n18540 ^ n18529 ;
  assign n18617 = n18530 & ~n18616 ;
  assign n18618 = n18617 ^ n18540 ;
  assign n18647 = n18646 ^ n18618 ;
  assign n18613 = ~n6849 & n7951 ;
  assign n18611 = x111 & n7954 ;
  assign n18607 = n18541 ^ n18505 ;
  assign n18608 = n18510 & n18607 ;
  assign n18609 = n18608 ^ n18505 ;
  assign n18605 = x113 & n7950 ;
  assign n18606 = n18605 ^ x56 ;
  assign n18610 = n18609 ^ n18606 ;
  assign n18612 = n18611 ^ n18610 ;
  assign n18614 = n18613 ^ n18612 ;
  assign n18604 = x112 & n7947 ;
  assign n18615 = n18614 ^ n18604 ;
  assign n18648 = n18647 ^ n18615 ;
  assign n18594 = x114 & n7183 ;
  assign n18593 = x116 & n7186 ;
  assign n18595 = n18594 ^ n18593 ;
  assign n18596 = n18595 ^ x53 ;
  assign n18592 = n7187 & ~n7604 ;
  assign n18597 = n18596 ^ n18592 ;
  assign n18591 = x115 & n7191 ;
  assign n18598 = n18597 ^ n18591 ;
  assign n18600 = n18598 ^ n18492 ;
  assign n18599 = n18598 ^ n18542 ;
  assign n18601 = n18600 ^ n18599 ;
  assign n18602 = ~n18497 & n18601 ;
  assign n18603 = n18602 ^ n18600 ;
  assign n18649 = n18648 ^ n18603 ;
  assign n18656 = n18655 ^ n18649 ;
  assign n18658 = n18657 ^ n18656 ;
  assign n18662 = n18661 ^ n18658 ;
  assign n18667 = n18666 ^ n18662 ;
  assign n18669 = n18668 ^ n18667 ;
  assign n18671 = n18670 ^ n18669 ;
  assign n18588 = n18544 ^ n18466 ;
  assign n18589 = n18471 & ~n18588 ;
  assign n18590 = n18589 ^ n18466 ;
  assign n18672 = n18671 ^ n18590 ;
  assign n18586 = x125 & n5116 ;
  assign n18587 = n18586 ^ x44 ;
  assign n18673 = n18672 ^ n18587 ;
  assign n18675 = n18674 ^ n18673 ;
  assign n18677 = n18676 ^ n18675 ;
  assign n18585 = x124 & n5121 ;
  assign n18678 = n18677 ^ n18585 ;
  assign n18582 = n18557 ^ n18553 ;
  assign n18583 = n18554 & n18582 ;
  assign n18584 = n18583 ^ n18557 ;
  assign n18679 = n18678 ^ n18584 ;
  assign n18681 = n18679 ^ n18558 ;
  assign n18680 = n18679 ^ n18571 ;
  assign n18682 = n18681 ^ n18680 ;
  assign n18683 = ~n18563 & ~n18682 ;
  assign n18684 = n18683 ^ n18681 ;
  assign n18691 = n18690 ^ n18684 ;
  assign n18697 = n18696 ^ n18691 ;
  assign n18700 = n18699 ^ n18697 ;
  assign n18807 = n18695 ^ n18691 ;
  assign n18882 = n18692 ^ n18580 ;
  assign n18808 = n18693 ^ n18572 ;
  assign n18809 = n18576 & n18808 ;
  assign n18810 = n18809 ^ n18575 ;
  assign n18812 = n18810 ^ n18691 ;
  assign n18811 = n18694 ^ n18692 ;
  assign n18813 = n18812 ^ n18811 ;
  assign n18885 = n18882 ^ n18813 ;
  assign n18881 = n18812 ^ n18692 ;
  assign n18886 = n18885 ^ n18881 ;
  assign n18887 = n18886 ^ n18810 ;
  assign n18889 = n18887 ^ n18885 ;
  assign n18828 = n18810 ^ n18692 ;
  assign n18834 = n18828 ^ n18694 ;
  assign n18829 = n18828 ^ n18580 ;
  assign n18830 = n18829 ^ n18810 ;
  assign n18870 = n18834 ^ n18830 ;
  assign n18868 = n18828 ^ n18810 ;
  assign n18871 = n18870 ^ n18868 ;
  assign n18872 = n18871 ^ n18691 ;
  assign n18874 = n18872 ^ n18870 ;
  assign n18835 = n18834 ^ n18810 ;
  assign n18838 = n18835 ^ n18812 ;
  assign n18831 = n18830 ^ n18694 ;
  assign n18832 = n18831 ^ n18812 ;
  assign n18846 = n18838 ^ n18832 ;
  assign n18840 = n18830 ^ n18812 ;
  assign n18833 = n18832 ^ n18812 ;
  assign n18839 = n18838 ^ n18833 ;
  assign n18841 = n18840 ^ n18839 ;
  assign n18842 = n18841 ^ n18840 ;
  assign n18847 = n18846 ^ n18842 ;
  assign n18848 = n18840 ^ n18828 ;
  assign n18849 = n18848 ^ n18846 ;
  assign n18850 = ~n18847 & ~n18849 ;
  assign n18851 = n18850 ^ n18832 ;
  assign n18852 = n18851 ^ n18840 ;
  assign n18853 = n18852 ^ n18810 ;
  assign n18854 = n18846 ^ n18840 ;
  assign n18855 = n18854 ^ n18810 ;
  assign n18856 = n18853 & n18855 ;
  assign n18857 = n18841 ^ n18838 ;
  assign n18858 = n18857 ^ n18828 ;
  assign n18859 = n18841 ^ n18832 ;
  assign n18860 = n18859 ^ n18828 ;
  assign n18861 = n18858 & ~n18860 ;
  assign n18862 = n18856 & n18861 ;
  assign n18863 = n18862 ^ n18850 ;
  assign n18864 = n18863 ^ n18846 ;
  assign n18844 = n18842 ^ n18828 ;
  assign n18865 = n18864 ^ n18844 ;
  assign n18836 = n18835 ^ n18830 ;
  assign n18866 = n18865 ^ n18836 ;
  assign n18867 = n18866 ^ n18828 ;
  assign n18875 = n18874 ^ n18867 ;
  assign n18876 = n18875 ^ n18692 ;
  assign n18877 = n18876 ^ n18872 ;
  assign n18819 = n18813 ^ n18812 ;
  assign n18823 = n18819 ^ n18812 ;
  assign n18820 = n18819 ^ n18580 ;
  assign n18821 = n18820 ^ n18812 ;
  assign n18814 = n18813 ^ n18692 ;
  assign n18815 = n18814 ^ n18580 ;
  assign n18816 = n18815 ^ n18810 ;
  assign n18817 = n18816 ^ n18812 ;
  assign n18818 = n18817 ^ n18812 ;
  assign n18822 = n18821 ^ n18818 ;
  assign n18824 = n18823 ^ n18822 ;
  assign n18826 = n18824 ^ n18810 ;
  assign n18825 = n18824 ^ n18823 ;
  assign n18827 = n18826 ^ n18825 ;
  assign n18878 = n18877 ^ n18827 ;
  assign n18879 = n18878 ^ n18815 ;
  assign n18880 = n18879 ^ n18826 ;
  assign n18890 = n18889 ^ n18880 ;
  assign n18891 = n18890 ^ n18691 ;
  assign n18892 = n18891 ^ n18887 ;
  assign n18893 = n18580 ^ n18457 ;
  assign n18896 = n18458 & n18893 ;
  assign n18897 = n18896 ^ n18457 ;
  assign n18898 = n18892 & n18897 ;
  assign n18899 = ~n18807 & n18898 ;
  assign n18900 = n18899 ^ n18892 ;
  assign n18803 = n18690 ^ n18679 ;
  assign n18804 = n18684 & ~n18803 ;
  assign n18805 = n18804 ^ n18679 ;
  assign n4483 = n4482 ^ n4479 ;
  assign n18798 = x127 & n4483 ;
  assign n18797 = n4479 & n10154 ;
  assign n18799 = n18798 ^ n18797 ;
  assign n18800 = n18799 ^ x41 ;
  assign n18794 = n18672 ^ n18584 ;
  assign n18795 = ~n18678 & ~n18794 ;
  assign n18796 = n18795 ^ n18672 ;
  assign n18801 = n18800 ^ n18796 ;
  assign n18788 = x124 & n5113 ;
  assign n18787 = x126 & n5116 ;
  assign n18789 = n18788 ^ n18787 ;
  assign n18790 = n18789 ^ x44 ;
  assign n18786 = n5117 & n10461 ;
  assign n18791 = n18790 ^ n18786 ;
  assign n18785 = x125 & n5121 ;
  assign n18792 = n18791 ^ n18785 ;
  assign n18778 = x121 & n5981 ;
  assign n18777 = x123 & n5748 ;
  assign n18779 = n18778 ^ n18777 ;
  assign n18780 = n18779 ^ x47 ;
  assign n18776 = n5749 & ~n9804 ;
  assign n18781 = n18780 ^ n18776 ;
  assign n18775 = x122 & n5755 ;
  assign n18782 = n18781 ^ n18775 ;
  assign n18765 = n7187 & ~n7860 ;
  assign n18763 = x115 & n7183 ;
  assign n18759 = n18647 ^ n18609 ;
  assign n18760 = ~n18615 & ~n18759 ;
  assign n18761 = n18760 ^ n18647 ;
  assign n18757 = x117 & n7186 ;
  assign n18758 = n18757 ^ x53 ;
  assign n18762 = n18761 ^ n18758 ;
  assign n18764 = n18763 ^ n18762 ;
  assign n18766 = n18765 ^ n18764 ;
  assign n18756 = x116 & n7191 ;
  assign n18767 = n18766 ^ n18756 ;
  assign n18749 = x109 & n8750 ;
  assign n18748 = x111 & n8746 ;
  assign n18750 = n18749 ^ n18748 ;
  assign n18751 = n18750 ^ x59 ;
  assign n18747 = ~n6370 & n8747 ;
  assign n18752 = n18751 ^ n18747 ;
  assign n18746 = x110 & n8743 ;
  assign n18753 = n18752 ^ n18746 ;
  assign n18744 = x107 & n9648 ;
  assign n18737 = n18636 ^ n18627 ;
  assign n18738 = n18628 & n18737 ;
  assign n18733 = x63 & x104 ;
  assign n18734 = n18733 ^ x105 ;
  assign n18735 = ~n9956 & n18734 ;
  assign n18736 = n18735 ^ x105 ;
  assign n18739 = n18738 ^ n18736 ;
  assign n18740 = n18739 ^ x62 ;
  assign n18730 = x106 & n9655 ;
  assign n18741 = n18740 ^ n18730 ;
  assign n18729 = x108 & n9651 ;
  assign n18742 = n18741 ^ n18729 ;
  assign n18728 = n5687 & n9652 ;
  assign n18743 = n18742 ^ n18728 ;
  assign n18745 = n18744 ^ n18743 ;
  assign n18754 = n18753 ^ n18745 ;
  assign n18726 = x113 & n7947 ;
  assign n18721 = x112 & n7954 ;
  assign n18720 = x114 & n7950 ;
  assign n18722 = n18721 ^ n18720 ;
  assign n18723 = n18722 ^ x56 ;
  assign n18719 = ~n7108 & n7951 ;
  assign n18724 = n18723 ^ n18719 ;
  assign n18716 = n18645 ^ n18618 ;
  assign n18717 = n18646 & ~n18716 ;
  assign n18718 = n18717 ^ n18645 ;
  assign n18725 = n18724 ^ n18718 ;
  assign n18727 = n18726 ^ n18725 ;
  assign n18755 = n18754 ^ n18727 ;
  assign n18768 = n18767 ^ n18755 ;
  assign n18713 = n6445 & n8904 ;
  assign n18711 = x118 & n6687 ;
  assign n18707 = n18648 ^ n18598 ;
  assign n18708 = n18603 & ~n18707 ;
  assign n18709 = n18708 ^ n18598 ;
  assign n18705 = x120 & n6444 ;
  assign n18706 = n18705 ^ x50 ;
  assign n18710 = n18709 ^ n18706 ;
  assign n18712 = n18711 ^ n18710 ;
  assign n18714 = n18713 ^ n18712 ;
  assign n18704 = x119 & n6449 ;
  assign n18715 = n18714 ^ n18704 ;
  assign n18769 = n18768 ^ n18715 ;
  assign n18771 = n18769 ^ n18661 ;
  assign n18770 = n18769 ^ n18649 ;
  assign n18772 = n18771 ^ n18770 ;
  assign n18773 = ~n18658 & ~n18772 ;
  assign n18774 = n18773 ^ n18770 ;
  assign n18783 = n18782 ^ n18774 ;
  assign n18701 = n18662 ^ n18590 ;
  assign n18702 = ~n18671 & ~n18701 ;
  assign n18703 = n18702 ^ n18662 ;
  assign n18784 = n18783 ^ n18703 ;
  assign n18793 = n18792 ^ n18784 ;
  assign n18802 = n18801 ^ n18793 ;
  assign n18806 = n18805 ^ n18802 ;
  assign n18901 = n18900 ^ n18806 ;
  assign n19019 = x125 & n5113 ;
  assign n19018 = x127 & n5116 ;
  assign n19020 = n19019 ^ n19018 ;
  assign n19021 = n19020 ^ x44 ;
  assign n19017 = n5117 & n10986 ;
  assign n19022 = n19021 ^ n19017 ;
  assign n19016 = x126 & n5121 ;
  assign n19023 = n19022 ^ n19016 ;
  assign n19012 = n18782 ^ n18769 ;
  assign n19013 = n18774 & ~n19012 ;
  assign n19014 = n19013 ^ n18769 ;
  assign n19006 = x122 & n5981 ;
  assign n19005 = x124 & n5748 ;
  assign n19007 = n19006 ^ n19005 ;
  assign n19008 = n19007 ^ x47 ;
  assign n19004 = n5749 & n10117 ;
  assign n19009 = n19008 ^ n19004 ;
  assign n19003 = x123 & n5755 ;
  assign n19010 = n19009 ^ n19003 ;
  assign n18994 = x113 & n7954 ;
  assign n18993 = x115 & n7950 ;
  assign n18995 = n18994 ^ n18993 ;
  assign n18996 = n18995 ^ x56 ;
  assign n18992 = ~n7353 & n7951 ;
  assign n18997 = n18996 ^ n18992 ;
  assign n18991 = x114 & n7947 ;
  assign n18998 = n18997 ^ n18991 ;
  assign n18984 = x110 & n8750 ;
  assign n18983 = x112 & n8746 ;
  assign n18985 = n18984 ^ n18983 ;
  assign n18986 = n18985 ^ x59 ;
  assign n18982 = ~n6616 & n8747 ;
  assign n18987 = n18986 ^ n18982 ;
  assign n18981 = x111 & n8743 ;
  assign n18988 = n18987 ^ n18981 ;
  assign n18975 = x63 & x105 ;
  assign n18976 = n18975 ^ x106 ;
  assign n18977 = ~n9956 & n18976 ;
  assign n18969 = n18624 ^ x106 ;
  assign n18978 = n18977 ^ n18969 ;
  assign n18979 = n18978 ^ x41 ;
  assign n18966 = n5912 & n9652 ;
  assign n18964 = x107 & n9655 ;
  assign n18960 = n18736 ^ n18624 ;
  assign n18961 = n18738 & ~n18960 ;
  assign n18962 = n18961 ^ n18624 ;
  assign n18958 = x109 & n9651 ;
  assign n18959 = n18958 ^ x62 ;
  assign n18963 = n18962 ^ n18959 ;
  assign n18965 = n18964 ^ n18963 ;
  assign n18967 = n18966 ^ n18965 ;
  assign n18957 = x108 & n9648 ;
  assign n18968 = n18967 ^ n18957 ;
  assign n18980 = n18979 ^ n18968 ;
  assign n18989 = n18988 ^ n18980 ;
  assign n18954 = n18753 ^ n18739 ;
  assign n18955 = ~n18745 & n18954 ;
  assign n18956 = n18955 ^ n18753 ;
  assign n18990 = n18989 ^ n18956 ;
  assign n18999 = n18998 ^ n18990 ;
  assign n18951 = n18754 ^ n18718 ;
  assign n18952 = n18727 & n18951 ;
  assign n18953 = n18952 ^ n18718 ;
  assign n19000 = n18999 ^ n18953 ;
  assign n18948 = n18761 ^ n18755 ;
  assign n18949 = n18767 & ~n18948 ;
  assign n18941 = x116 & n7183 ;
  assign n18940 = x118 & n7186 ;
  assign n18942 = n18941 ^ n18940 ;
  assign n18943 = n18942 ^ x53 ;
  assign n18939 = n7187 & ~n8140 ;
  assign n18944 = n18943 ^ n18939 ;
  assign n18938 = x117 & n7191 ;
  assign n18945 = n18944 ^ n18938 ;
  assign n18946 = n18945 ^ n18755 ;
  assign n18950 = n18949 ^ n18946 ;
  assign n19001 = n19000 ^ n18950 ;
  assign n18928 = x119 & n6687 ;
  assign n18927 = x121 & n6444 ;
  assign n18929 = n18928 ^ n18927 ;
  assign n18930 = n18929 ^ x50 ;
  assign n18926 = n6445 & n8979 ;
  assign n18931 = n18930 ^ n18926 ;
  assign n18925 = x120 & n6449 ;
  assign n18932 = n18931 ^ n18925 ;
  assign n18933 = n18932 ^ n18768 ;
  assign n18934 = n18933 ^ n18709 ;
  assign n18935 = n18934 ^ n18932 ;
  assign n18936 = ~n18715 & ~n18935 ;
  assign n18937 = n18936 ^ n18933 ;
  assign n19002 = n19001 ^ n18937 ;
  assign n19011 = n19010 ^ n19002 ;
  assign n19015 = n19014 ^ n19011 ;
  assign n19024 = n19023 ^ n19015 ;
  assign n18922 = n18792 ^ n18703 ;
  assign n18923 = n18784 & ~n18922 ;
  assign n18924 = n18923 ^ n18792 ;
  assign n19025 = n19024 ^ n18924 ;
  assign n18905 = n18800 ^ n18793 ;
  assign n18906 = ~n18801 & n18905 ;
  assign n18907 = n18906 ^ n18905 ;
  assign n18902 = ~n18793 & n18800 ;
  assign n18903 = ~n18796 & n18902 ;
  assign n18908 = n18907 ^ n18903 ;
  assign n18909 = n18805 & n18908 ;
  assign n18904 = ~n18805 & n18903 ;
  assign n18910 = n18909 ^ n18904 ;
  assign n18911 = n18906 ^ n18796 ;
  assign n18912 = n18903 ^ n18805 ;
  assign n18913 = n18912 ^ n18904 ;
  assign n18914 = ~n18911 & ~n18913 ;
  assign n18915 = n18914 ^ n18806 ;
  assign n18916 = n18915 ^ n18914 ;
  assign n18917 = n18914 ^ n18900 ;
  assign n18918 = n18917 ^ n18914 ;
  assign n18919 = ~n18916 & n18918 ;
  assign n18920 = n18919 ^ n18914 ;
  assign n18921 = ~n18910 & ~n18920 ;
  assign n19026 = n19025 ^ n18921 ;
  assign n19131 = n5117 & n10155 ;
  assign n19130 = x126 & n5113 ;
  assign n19132 = n19131 ^ n19130 ;
  assign n19133 = n19132 ^ x44 ;
  assign n19129 = x127 & n5121 ;
  assign n19134 = n19133 ^ n19129 ;
  assign n19121 = x120 & n6687 ;
  assign n19120 = x122 & n6444 ;
  assign n19122 = n19121 ^ n19120 ;
  assign n19123 = n19122 ^ x50 ;
  assign n19119 = n6445 & ~n9261 ;
  assign n19124 = n19123 ^ n19119 ;
  assign n19118 = x121 & n6449 ;
  assign n19125 = n19124 ^ n19118 ;
  assign n19109 = n18998 ^ n18953 ;
  assign n19110 = n18999 & n19109 ;
  assign n19111 = n19110 ^ n18998 ;
  assign n19103 = x117 & n7183 ;
  assign n19102 = x119 & n7186 ;
  assign n19104 = n19103 ^ n19102 ;
  assign n19105 = n19104 ^ x53 ;
  assign n19101 = n7187 & n8405 ;
  assign n19106 = n19105 ^ n19101 ;
  assign n19100 = x118 & n7191 ;
  assign n19107 = n19106 ^ n19100 ;
  assign n19092 = x108 & n9655 ;
  assign n19091 = x110 & n9651 ;
  assign n19093 = n19092 ^ n19091 ;
  assign n19094 = n19093 ^ x62 ;
  assign n19090 = n6145 & n9652 ;
  assign n19095 = n19094 ^ n19090 ;
  assign n19089 = x109 & n9648 ;
  assign n19096 = n19095 ^ n19089 ;
  assign n19085 = n18624 ^ x41 ;
  assign n19086 = ~n18978 & ~n19085 ;
  assign n19087 = n19086 ^ x41 ;
  assign n19081 = x63 & x106 ;
  assign n19082 = n19081 ^ x107 ;
  assign n19083 = ~n9956 & n19082 ;
  assign n19084 = n19083 ^ x107 ;
  assign n19088 = n19087 ^ n19084 ;
  assign n19097 = n19096 ^ n19088 ;
  assign n19076 = ~n6849 & n8747 ;
  assign n19074 = x111 & n8750 ;
  assign n19070 = n18979 ^ n18962 ;
  assign n19071 = n18968 & n19070 ;
  assign n19072 = n19071 ^ n18979 ;
  assign n19068 = x113 & n8746 ;
  assign n19069 = n19068 ^ x59 ;
  assign n19073 = n19072 ^ n19069 ;
  assign n19075 = n19074 ^ n19073 ;
  assign n19077 = n19076 ^ n19075 ;
  assign n19067 = x112 & n8743 ;
  assign n19078 = n19077 ^ n19067 ;
  assign n19098 = n19097 ^ n19078 ;
  assign n19064 = n18988 ^ n18956 ;
  assign n19065 = n18989 & n19064 ;
  assign n19057 = x114 & n7954 ;
  assign n19056 = x116 & n7950 ;
  assign n19058 = n19057 ^ n19056 ;
  assign n19059 = n19058 ^ x56 ;
  assign n19055 = ~n7604 & n7951 ;
  assign n19060 = n19059 ^ n19055 ;
  assign n19054 = x115 & n7947 ;
  assign n19061 = n19060 ^ n19054 ;
  assign n19062 = n19061 ^ n18988 ;
  assign n19066 = n19065 ^ n19062 ;
  assign n19099 = n19098 ^ n19066 ;
  assign n19108 = n19107 ^ n19099 ;
  assign n19112 = n19111 ^ n19108 ;
  assign n19114 = n19112 ^ n18945 ;
  assign n19113 = n19112 ^ n19000 ;
  assign n19115 = n19114 ^ n19113 ;
  assign n19116 = n18950 & n19115 ;
  assign n19117 = n19116 ^ n19114 ;
  assign n19126 = n19125 ^ n19117 ;
  assign n19051 = n5749 & n10416 ;
  assign n19049 = x123 & n5981 ;
  assign n19045 = n19001 ^ n18932 ;
  assign n19046 = ~n18937 & n19045 ;
  assign n19047 = n19046 ^ n18932 ;
  assign n19043 = x125 & n5748 ;
  assign n19044 = n19043 ^ x47 ;
  assign n19048 = n19047 ^ n19044 ;
  assign n19050 = n19049 ^ n19048 ;
  assign n19052 = n19051 ^ n19050 ;
  assign n19042 = x124 & n5755 ;
  assign n19053 = n19052 ^ n19042 ;
  assign n19127 = n19126 ^ n19053 ;
  assign n19039 = n19014 ^ n19010 ;
  assign n19040 = n19011 & ~n19039 ;
  assign n19041 = n19040 ^ n19014 ;
  assign n19128 = n19127 ^ n19041 ;
  assign n19135 = n19134 ^ n19128 ;
  assign n19036 = n19023 ^ n18924 ;
  assign n19037 = n19024 & n19036 ;
  assign n19038 = n19037 ^ n19023 ;
  assign n19136 = n19135 ^ n19038 ;
  assign n19027 = ~n18900 & ~n18909 ;
  assign n19028 = n18915 ^ n18910 ;
  assign n19029 = ~n18904 & n19025 ;
  assign n19030 = n19028 & n19029 ;
  assign n19031 = n19030 ^ n18904 ;
  assign n19032 = n19025 ^ n18914 ;
  assign n19033 = ~n19031 & n19032 ;
  assign n19034 = n19027 & n19033 ;
  assign n19035 = n19034 ^ n19031 ;
  assign n19137 = n19136 ^ n19035 ;
  assign n19239 = n19135 ^ n19035 ;
  assign n19240 = n19038 ^ n19035 ;
  assign n19241 = n19239 & ~n19240 ;
  assign n19242 = n19241 ^ n19135 ;
  assign n19226 = x127 & n5112 ;
  assign n19227 = n19226 ^ n5110 ;
  assign n19232 = n4685 & n11285 ;
  assign n19233 = n19232 ^ n19226 ;
  assign n19234 = n19227 & ~n19233 ;
  assign n19235 = n19234 ^ x43 ;
  assign n19223 = n19126 ^ n19047 ;
  assign n19224 = ~n19053 & ~n19223 ;
  assign n19225 = n19224 ^ n19126 ;
  assign n19236 = n19235 ^ n19225 ;
  assign n19220 = x125 & n5755 ;
  assign n19218 = n5749 & n10461 ;
  assign n19214 = x124 & n5981 ;
  assign n19213 = x126 & n5748 ;
  assign n19215 = n19214 ^ n19213 ;
  assign n19216 = n19215 ^ x47 ;
  assign n19210 = x122 & n6449 ;
  assign n19208 = n6445 & ~n9804 ;
  assign n19204 = x121 & n6687 ;
  assign n19203 = x123 & n6444 ;
  assign n19205 = n19204 ^ n19203 ;
  assign n19206 = n19205 ^ x50 ;
  assign n19200 = x119 & n7191 ;
  assign n19198 = n7187 & n8904 ;
  assign n19194 = x118 & n7183 ;
  assign n19193 = x120 & n7186 ;
  assign n19195 = n19194 ^ n19193 ;
  assign n19196 = n19195 ^ x53 ;
  assign n19186 = x115 & n7954 ;
  assign n19185 = x117 & n7950 ;
  assign n19187 = n19186 ^ n19185 ;
  assign n19188 = n19187 ^ x56 ;
  assign n19184 = ~n7860 & n7951 ;
  assign n19189 = n19188 ^ n19184 ;
  assign n19183 = x116 & n7947 ;
  assign n19190 = n19189 ^ n19183 ;
  assign n19177 = x112 & n8750 ;
  assign n19176 = x114 & n8746 ;
  assign n19178 = n19177 ^ n19176 ;
  assign n19179 = n19178 ^ x59 ;
  assign n19175 = ~n7108 & n8747 ;
  assign n19180 = n19179 ^ n19175 ;
  assign n19174 = x113 & n8743 ;
  assign n19181 = n19180 ^ n19174 ;
  assign n19168 = ~n6370 & n9652 ;
  assign n19167 = x110 & n9648 ;
  assign n19169 = n19168 ^ n19167 ;
  assign n19165 = x109 & n9655 ;
  assign n19164 = x111 & n9651 ;
  assign n19166 = n19165 ^ n19164 ;
  assign n19170 = n19169 ^ n19166 ;
  assign n19163 = n5232 ^ x62 ;
  assign n19171 = n19170 ^ n19163 ;
  assign n19160 = n19096 ^ n19087 ;
  assign n19161 = ~n19088 & ~n19160 ;
  assign n19162 = n19161 ^ n19096 ;
  assign n19172 = n19171 ^ n19162 ;
  assign n19157 = x63 & n5012 ;
  assign n19158 = n19157 ^ n5232 ;
  assign n19159 = ~n9956 & n19158 ;
  assign n19173 = n19172 ^ n19159 ;
  assign n19182 = n19181 ^ n19173 ;
  assign n19191 = n19190 ^ n19182 ;
  assign n19150 = n19097 ^ n19072 ;
  assign n19151 = n19078 & ~n19150 ;
  assign n19152 = n19151 ^ n19097 ;
  assign n19192 = n19191 ^ n19152 ;
  assign n19197 = n19196 ^ n19192 ;
  assign n19199 = n19198 ^ n19197 ;
  assign n19201 = n19200 ^ n19199 ;
  assign n19147 = n19098 ^ n19061 ;
  assign n19148 = n19066 & ~n19147 ;
  assign n19149 = n19148 ^ n19061 ;
  assign n19202 = n19201 ^ n19149 ;
  assign n19207 = n19206 ^ n19202 ;
  assign n19209 = n19208 ^ n19207 ;
  assign n19211 = n19210 ^ n19209 ;
  assign n19144 = n19111 ^ n19107 ;
  assign n19145 = n19108 & n19144 ;
  assign n19146 = n19145 ^ n19111 ;
  assign n19212 = n19211 ^ n19146 ;
  assign n19217 = n19216 ^ n19212 ;
  assign n19219 = n19218 ^ n19217 ;
  assign n19221 = n19220 ^ n19219 ;
  assign n19141 = n19125 ^ n19112 ;
  assign n19142 = ~n19117 & ~n19141 ;
  assign n19143 = n19142 ^ n19112 ;
  assign n19222 = n19221 ^ n19143 ;
  assign n19237 = n19236 ^ n19222 ;
  assign n19138 = n19134 ^ n19041 ;
  assign n19139 = ~n19128 & ~n19138 ;
  assign n19140 = n19139 ^ n19134 ;
  assign n19238 = n19237 ^ n19140 ;
  assign n19243 = n19242 ^ n19238 ;
  assign n19244 = n19242 ^ n19222 ;
  assign n19377 = n19235 ^ n19222 ;
  assign n19378 = ~n19244 & ~n19377 ;
  assign n19372 = n19212 ^ n19143 ;
  assign n19373 = ~n19221 & n19372 ;
  assign n19374 = n19373 ^ n19212 ;
  assign n19366 = x125 & n5981 ;
  assign n19365 = x127 & n5748 ;
  assign n19367 = n19366 ^ n19365 ;
  assign n19368 = n19367 ^ x47 ;
  assign n19364 = n5749 & n10986 ;
  assign n19369 = n19368 ^ n19364 ;
  assign n19363 = x126 & n5755 ;
  assign n19370 = n19369 ^ n19363 ;
  assign n19359 = n19202 ^ n19146 ;
  assign n19360 = ~n19211 & ~n19359 ;
  assign n19361 = n19360 ^ n19202 ;
  assign n19353 = x122 & n6687 ;
  assign n19352 = x124 & n6444 ;
  assign n19354 = n19353 ^ n19352 ;
  assign n19355 = n19354 ^ x50 ;
  assign n19351 = n6445 & n10117 ;
  assign n19356 = n19355 ^ n19351 ;
  assign n19350 = x123 & n6449 ;
  assign n19357 = n19356 ^ n19350 ;
  assign n19345 = n19190 ^ n19152 ;
  assign n19346 = ~n19191 & n19345 ;
  assign n19347 = n19346 ^ n19190 ;
  assign n19343 = x117 & n7947 ;
  assign n19331 = x110 & n9655 ;
  assign n19330 = x112 & n9651 ;
  assign n19332 = n19331 ^ n19330 ;
  assign n19333 = n19332 ^ x62 ;
  assign n19329 = ~n6616 & n9652 ;
  assign n19334 = n19333 ^ n19329 ;
  assign n19328 = x111 & n9648 ;
  assign n19335 = n19334 ^ n19328 ;
  assign n19323 = ~x63 & x108 ;
  assign n19324 = n19323 ^ n5441 ;
  assign n19325 = ~n9956 & n19324 ;
  assign n19318 = n19084 ^ x109 ;
  assign n19326 = n19325 ^ n19318 ;
  assign n19327 = n19326 ^ x44 ;
  assign n19336 = n19335 ^ n19327 ;
  assign n19278 = x108 ^ x63 ;
  assign n19279 = n19278 ^ n19170 ;
  assign n19282 = n5232 & ~n19279 ;
  assign n19283 = n19282 ^ n19170 ;
  assign n19284 = n9956 & n19283 ;
  assign n19310 = n19284 ^ x62 ;
  assign n19293 = x107 & ~x108 ;
  assign n19295 = n19293 ^ x106 ;
  assign n19294 = n19293 ^ n19170 ;
  assign n19296 = n19295 ^ n19294 ;
  assign n19299 = ~n5012 & n19296 ;
  assign n19300 = n19299 ^ n19295 ;
  assign n19301 = x62 & n19300 ;
  assign n19302 = n19301 ^ n19293 ;
  assign n19311 = n19310 ^ n19302 ;
  assign n19303 = n19302 ^ x63 ;
  assign n19312 = n19311 ^ n19303 ;
  assign n19290 = n19170 & ~n19284 ;
  assign n19291 = n19290 ^ x63 ;
  assign n19292 = n19291 & ~n19310 ;
  assign n19313 = n19312 ^ n19292 ;
  assign n19314 = n19313 ^ n19302 ;
  assign n19315 = ~n19292 & n19311 ;
  assign n19316 = ~n19314 & n19315 ;
  assign n19317 = n19316 ^ n19313 ;
  assign n19337 = n19336 ^ n19317 ;
  assign n19275 = n19181 ^ n19162 ;
  assign n19276 = n19173 & n19275 ;
  assign n19268 = x113 & n8750 ;
  assign n19267 = x115 & n8746 ;
  assign n19269 = n19268 ^ n19267 ;
  assign n19270 = n19269 ^ x59 ;
  assign n19266 = ~n7353 & n8747 ;
  assign n19271 = n19270 ^ n19266 ;
  assign n19265 = x114 & n8743 ;
  assign n19272 = n19271 ^ n19265 ;
  assign n19273 = n19272 ^ n19181 ;
  assign n19277 = n19276 ^ n19273 ;
  assign n19338 = n19337 ^ n19277 ;
  assign n19339 = n19338 ^ x56 ;
  assign n19264 = x116 & n7954 ;
  assign n19340 = n19339 ^ n19264 ;
  assign n19263 = x118 & n7950 ;
  assign n19341 = n19340 ^ n19263 ;
  assign n19262 = n7951 & ~n8140 ;
  assign n19342 = n19341 ^ n19262 ;
  assign n19344 = n19343 ^ n19342 ;
  assign n19348 = n19347 ^ n19344 ;
  assign n19252 = x119 & n7183 ;
  assign n19251 = x121 & n7186 ;
  assign n19253 = n19252 ^ n19251 ;
  assign n19254 = n19253 ^ x53 ;
  assign n19250 = n7187 & n8979 ;
  assign n19255 = n19254 ^ n19250 ;
  assign n19249 = x120 & n7191 ;
  assign n19256 = n19255 ^ n19249 ;
  assign n19257 = n19256 ^ n19192 ;
  assign n19258 = n19257 ^ n19149 ;
  assign n19259 = n19258 ^ n19256 ;
  assign n19260 = ~n19201 & ~n19259 ;
  assign n19261 = n19260 ^ n19257 ;
  assign n19349 = n19348 ^ n19261 ;
  assign n19358 = n19357 ^ n19349 ;
  assign n19362 = n19361 ^ n19358 ;
  assign n19371 = n19370 ^ n19362 ;
  assign n19375 = n19374 ^ n19371 ;
  assign n19245 = n19244 ^ n19235 ;
  assign n19246 = n19245 ^ n19225 ;
  assign n19247 = n19225 ^ n19140 ;
  assign n19248 = ~n19246 & n19247 ;
  assign n19376 = n19375 ^ n19248 ;
  assign n19379 = n19378 ^ n19376 ;
  assign n19554 = n5749 & n10155 ;
  assign n19553 = x126 & n5981 ;
  assign n19555 = n19554 ^ n19553 ;
  assign n19556 = n19555 ^ x47 ;
  assign n19552 = x127 & n5755 ;
  assign n19557 = n19556 ^ n19552 ;
  assign n19549 = x124 & n6449 ;
  assign n19547 = n6445 & n10416 ;
  assign n19543 = x123 & n6687 ;
  assign n19542 = x125 & n6444 ;
  assign n19544 = n19543 ^ n19542 ;
  assign n19545 = n19544 ^ x50 ;
  assign n19535 = x120 & n7183 ;
  assign n19534 = x122 & n7186 ;
  assign n19536 = n19535 ^ n19534 ;
  assign n19537 = n19536 ^ x53 ;
  assign n19533 = n7187 & ~n9261 ;
  assign n19538 = n19537 ^ n19533 ;
  assign n19532 = x121 & n7191 ;
  assign n19539 = n19538 ^ n19532 ;
  assign n19528 = n19337 ^ n19272 ;
  assign n19529 = n19277 & ~n19528 ;
  assign n19530 = n19529 ^ n19272 ;
  assign n19522 = x117 & n7954 ;
  assign n19521 = x119 & n7950 ;
  assign n19523 = n19522 ^ n19521 ;
  assign n19524 = n19523 ^ x56 ;
  assign n19520 = n7951 & n8405 ;
  assign n19525 = n19524 ^ n19520 ;
  assign n19519 = x118 & n7947 ;
  assign n19526 = n19525 ^ n19519 ;
  assign n19512 = x114 & n8750 ;
  assign n19511 = x116 & n8746 ;
  assign n19513 = n19512 ^ n19511 ;
  assign n19514 = n19513 ^ x59 ;
  assign n19510 = ~n7604 & n8747 ;
  assign n19515 = n19514 ^ n19510 ;
  assign n19509 = x115 & n8743 ;
  assign n19516 = n19515 ^ n19509 ;
  assign n19506 = x109 & n11895 ;
  assign n19505 = x110 & n9956 ;
  assign n19507 = n19506 ^ n19505 ;
  assign n19502 = ~n6849 & n9652 ;
  assign n19500 = x111 & n9655 ;
  assign n19496 = n19084 ^ x44 ;
  assign n19497 = ~n19326 & ~n19496 ;
  assign n19498 = n19497 ^ x44 ;
  assign n19494 = x113 & n9651 ;
  assign n19495 = n19494 ^ x62 ;
  assign n19499 = n19498 ^ n19495 ;
  assign n19501 = n19500 ^ n19499 ;
  assign n19503 = n19502 ^ n19501 ;
  assign n19493 = x112 & n9648 ;
  assign n19504 = n19503 ^ n19493 ;
  assign n19508 = n19507 ^ n19504 ;
  assign n19517 = n19516 ^ n19508 ;
  assign n19490 = n19335 ^ n19317 ;
  assign n19491 = ~n19336 & n19490 ;
  assign n19492 = n19491 ^ n19335 ;
  assign n19518 = n19517 ^ n19492 ;
  assign n19527 = n19526 ^ n19518 ;
  assign n19531 = n19530 ^ n19527 ;
  assign n19540 = n19539 ^ n19531 ;
  assign n19487 = n19347 ^ n19338 ;
  assign n19488 = n19344 & ~n19487 ;
  assign n19489 = n19488 ^ n19347 ;
  assign n19541 = n19540 ^ n19489 ;
  assign n19546 = n19545 ^ n19541 ;
  assign n19548 = n19547 ^ n19546 ;
  assign n19550 = n19549 ^ n19548 ;
  assign n19484 = n19348 ^ n19256 ;
  assign n19485 = ~n19261 & ~n19484 ;
  assign n19486 = n19485 ^ n19256 ;
  assign n19551 = n19550 ^ n19486 ;
  assign n19558 = n19557 ^ n19551 ;
  assign n19481 = n19361 ^ n19357 ;
  assign n19482 = ~n19358 & ~n19481 ;
  assign n19483 = n19482 ^ n19361 ;
  assign n19559 = n19558 ^ n19483 ;
  assign n19478 = n19374 ^ n19370 ;
  assign n19479 = n19371 & ~n19478 ;
  assign n19480 = n19479 ^ n19374 ;
  assign n19560 = n19559 ^ n19480 ;
  assign n19380 = n19140 & ~n19225 ;
  assign n19385 = n19380 ^ n19247 ;
  assign n19457 = n19385 ^ n19242 ;
  assign n19381 = n19380 ^ n19222 ;
  assign n19382 = n19377 & ~n19381 ;
  assign n19383 = n19382 ^ n19235 ;
  assign n19387 = n19383 ^ n19375 ;
  assign n19384 = n19222 & n19235 ;
  assign n19386 = n19385 ^ n19384 ;
  assign n19388 = n19387 ^ n19386 ;
  assign n19460 = n19457 ^ n19388 ;
  assign n19456 = n19387 ^ n19385 ;
  assign n19461 = n19460 ^ n19456 ;
  assign n19462 = n19461 ^ n19383 ;
  assign n19464 = n19462 ^ n19460 ;
  assign n19403 = n19385 ^ n19383 ;
  assign n19409 = n19403 ^ n19384 ;
  assign n19404 = n19403 ^ n19242 ;
  assign n19405 = n19404 ^ n19383 ;
  assign n19445 = n19409 ^ n19405 ;
  assign n19446 = n19445 ^ n19385 ;
  assign n19447 = n19446 ^ n19375 ;
  assign n19449 = n19447 ^ n19445 ;
  assign n19410 = n19409 ^ n19383 ;
  assign n19413 = n19410 ^ n19387 ;
  assign n19406 = n19405 ^ n19384 ;
  assign n19407 = n19406 ^ n19387 ;
  assign n19421 = n19413 ^ n19407 ;
  assign n19415 = n19405 ^ n19387 ;
  assign n19417 = n19415 ^ n19385 ;
  assign n19422 = n19421 ^ n19417 ;
  assign n19423 = n19415 ^ n19403 ;
  assign n19424 = n19423 ^ n19421 ;
  assign n19425 = n19422 & n19424 ;
  assign n19426 = n19425 ^ n19407 ;
  assign n19427 = n19426 ^ n19415 ;
  assign n19428 = n19427 ^ n19383 ;
  assign n19429 = n19421 ^ n19415 ;
  assign n19430 = n19429 ^ n19383 ;
  assign n19431 = n19428 & ~n19430 ;
  assign n19432 = n19413 ^ n19385 ;
  assign n19433 = n19432 ^ n19403 ;
  assign n19434 = n19407 ^ n19385 ;
  assign n19435 = n19434 ^ n19403 ;
  assign n19436 = ~n19433 & ~n19435 ;
  assign n19437 = n19431 & n19436 ;
  assign n19438 = n19437 ^ n19425 ;
  assign n19439 = n19438 ^ n19421 ;
  assign n19419 = n19417 ^ n19403 ;
  assign n19440 = n19439 ^ n19419 ;
  assign n19411 = n19410 ^ n19405 ;
  assign n19441 = n19440 ^ n19411 ;
  assign n19442 = n19441 ^ n19403 ;
  assign n19450 = n19449 ^ n19442 ;
  assign n19451 = n19450 ^ n19385 ;
  assign n19452 = n19451 ^ n19447 ;
  assign n19394 = n19388 ^ n19387 ;
  assign n19398 = n19394 ^ n19387 ;
  assign n19395 = n19394 ^ n19242 ;
  assign n19396 = n19395 ^ n19387 ;
  assign n19389 = n19388 ^ n19385 ;
  assign n19390 = n19389 ^ n19242 ;
  assign n19391 = n19390 ^ n19383 ;
  assign n19392 = n19391 ^ n19387 ;
  assign n19393 = n19392 ^ n19387 ;
  assign n19397 = n19396 ^ n19393 ;
  assign n19399 = n19398 ^ n19397 ;
  assign n19401 = n19399 ^ n19383 ;
  assign n19400 = n19399 ^ n19398 ;
  assign n19402 = n19401 ^ n19400 ;
  assign n19453 = n19452 ^ n19402 ;
  assign n19454 = n19453 ^ n19390 ;
  assign n19455 = n19454 ^ n19401 ;
  assign n19465 = n19464 ^ n19455 ;
  assign n19466 = n19465 ^ n19375 ;
  assign n19467 = n19466 ^ n19462 ;
  assign n19468 = n19242 ^ n19140 ;
  assign n19471 = n19247 & n19468 ;
  assign n19472 = n19471 ^ n19242 ;
  assign n19473 = n19467 & ~n19472 ;
  assign n19474 = n19384 ^ n19375 ;
  assign n19475 = n19474 ^ n19377 ;
  assign n19476 = n19473 & n19475 ;
  assign n19477 = n19476 ^ n19467 ;
  assign n19561 = n19560 ^ n19477 ;
  assign n19562 = n19483 ^ n19480 ;
  assign n19656 = n19480 ^ n19477 ;
  assign n19657 = ~n19562 & n19656 ;
  assign n19651 = n19541 ^ n19486 ;
  assign n19652 = n19550 & n19651 ;
  assign n19653 = n19652 ^ n19541 ;
  assign n19566 = x127 & n5980 ;
  assign n19567 = n19566 ^ n5323 ;
  assign n19568 = n19567 ^ n19566 ;
  assign n19571 = n11285 & n19568 ;
  assign n19572 = n19571 ^ n19566 ;
  assign n19642 = x125 & n6449 ;
  assign n19640 = n6445 & n10461 ;
  assign n19636 = x124 & n6687 ;
  assign n19635 = x126 & n6444 ;
  assign n19637 = n19636 ^ n19635 ;
  assign n19638 = n19637 ^ x50 ;
  assign n19628 = x121 & n7183 ;
  assign n19627 = x123 & n7186 ;
  assign n19629 = n19628 ^ n19627 ;
  assign n19630 = n19629 ^ x53 ;
  assign n19626 = n7187 & ~n9804 ;
  assign n19631 = n19630 ^ n19626 ;
  assign n19625 = x122 & n7191 ;
  assign n19632 = n19631 ^ n19625 ;
  assign n19612 = ~x111 & n9956 ;
  assign n19613 = n19612 ^ n19506 ;
  assign n19614 = x110 & n19613 ;
  assign n19615 = n19614 ^ n19506 ;
  assign n19616 = n9956 ^ x110 ;
  assign n19617 = n19613 ^ n12206 ;
  assign n19618 = n19616 & n19617 ;
  assign n19675 = ~n19615 & ~n19618 ;
  assign n19609 = n19507 ^ n19498 ;
  assign n19610 = n19504 & n19609 ;
  assign n19611 = n19610 ^ n19507 ;
  assign n19622 = ~n19675 ^ n19611 ;
  assign n19606 = ~n7860 & n8747 ;
  assign n19604 = x115 & n8750 ;
  assign n19598 = x112 & n9655 ;
  assign n19597 = x114 & n9651 ;
  assign n19599 = n19598 ^ n19597 ;
  assign n19600 = n19599 ^ x62 ;
  assign n19596 = ~n7108 & n9652 ;
  assign n19601 = n19600 ^ n19596 ;
  assign n19595 = x113 & n9648 ;
  assign n19602 = n19601 ^ n19595 ;
  assign n19593 = x117 & n8746 ;
  assign n19594 = n19593 ^ x59 ;
  assign n19603 = n19602 ^ n19594 ;
  assign n19605 = n19604 ^ n19603 ;
  assign n19607 = n19606 ^ n19605 ;
  assign n19592 = x116 & n8743 ;
  assign n19608 = n19607 ^ n19592 ;
  assign n19623 = n19622 ^ n19608 ;
  assign n19582 = x118 & n7954 ;
  assign n19581 = x120 & n7950 ;
  assign n19583 = n19582 ^ n19581 ;
  assign n19584 = n19583 ^ x56 ;
  assign n19580 = n7951 & n8904 ;
  assign n19585 = n19584 ^ n19580 ;
  assign n19579 = x119 & n7947 ;
  assign n19586 = n19585 ^ n19579 ;
  assign n19587 = n19586 ^ n19516 ;
  assign n19588 = n19587 ^ n19586 ;
  assign n19589 = n19588 ^ n19492 ;
  assign n19590 = n19517 & n19589 ;
  assign n19591 = n19590 ^ n19587 ;
  assign n19624 = n19623 ^ n19591 ;
  assign n19633 = n19632 ^ n19624 ;
  assign n19576 = n19530 ^ n19526 ;
  assign n19577 = ~n19527 & n19576 ;
  assign n19578 = n19577 ^ n19530 ;
  assign n19634 = n19633 ^ n19578 ;
  assign n19639 = n19638 ^ n19634 ;
  assign n19641 = n19640 ^ n19639 ;
  assign n19643 = n19642 ^ n19641 ;
  assign n19573 = n19539 ^ n19489 ;
  assign n19574 = n19540 & n19573 ;
  assign n19575 = n19574 ^ n19539 ;
  assign n19644 = n19643 ^ n19575 ;
  assign n19647 = n19644 ^ x46 ;
  assign n19645 = n19644 ^ x47 ;
  assign n19646 = n19645 ^ n19566 ;
  assign n19648 = n19647 ^ n19646 ;
  assign n19649 = ~n19572 & n19648 ;
  assign n19650 = n19649 ^ n19647 ;
  assign n19654 = n19653 ^ n19650 ;
  assign n19563 = n19562 ^ n19551 ;
  assign n19564 = n19563 ^ n19477 ;
  assign n19565 = ~n19558 & n19564 ;
  assign n19655 = n19654 ^ n19565 ;
  assign n19658 = n19657 ^ n19655 ;
  assign n19734 = ~n19551 & ~n19557 ;
  assign n19735 = n19734 ^ n19558 ;
  assign n19736 = n19480 & n19483 ;
  assign n19737 = n19736 ^ n19654 ;
  assign n19738 = n19735 & ~n19737 ;
  assign n19739 = n19735 ^ n19477 ;
  assign n19740 = n19736 ^ n19562 ;
  assign n19741 = ~n19734 & ~n19740 ;
  assign n19742 = n19741 ^ n19654 ;
  assign n19743 = ~n19739 & n19742 ;
  assign n19744 = n19738 & ~n19743 ;
  assign n19745 = ~n19562 & ~n19656 ;
  assign n19746 = n19745 ^ n19477 ;
  assign n19747 = n19654 & ~n19734 ;
  assign n19748 = ~n19746 & n19747 ;
  assign n19749 = n19748 ^ n19746 ;
  assign n19750 = ~n19744 & n19749 ;
  assign n19729 = n19653 ^ n19644 ;
  assign n19730 = n19650 & n19729 ;
  assign n19731 = n19730 ^ n19644 ;
  assign n19726 = n19634 ^ n19575 ;
  assign n19727 = n19643 & n19726 ;
  assign n19728 = n19727 ^ n19634 ;
  assign n19732 = n19731 ^ n19728 ;
  assign n19720 = x125 & n6687 ;
  assign n19719 = x127 & n6444 ;
  assign n19721 = n19720 ^ n19719 ;
  assign n19722 = n19721 ^ x50 ;
  assign n19718 = n6445 & n10986 ;
  assign n19723 = n19722 ^ n19718 ;
  assign n19717 = x126 & n6449 ;
  assign n19724 = n19723 ^ n19717 ;
  assign n19710 = x122 & n7183 ;
  assign n19709 = x124 & n7186 ;
  assign n19711 = n19710 ^ n19709 ;
  assign n19712 = n19711 ^ x53 ;
  assign n19708 = n7187 & n10117 ;
  assign n19713 = n19712 ^ n19708 ;
  assign n19707 = x123 & n7191 ;
  assign n19714 = n19713 ^ n19707 ;
  assign n19703 = n19623 ^ n19586 ;
  assign n19704 = n19591 & n19703 ;
  assign n19705 = n19704 ^ n19586 ;
  assign n19701 = x120 & n7947 ;
  assign n19696 = x119 & n7954 ;
  assign n19695 = x121 & n7950 ;
  assign n19697 = n19696 ^ n19695 ;
  assign n19698 = n19697 ^ x56 ;
  assign n19694 = n7951 & n8979 ;
  assign n19699 = n19698 ^ n19694 ;
  assign n19685 = x113 & n9655 ;
  assign n19684 = x115 & n9651 ;
  assign n19686 = n19685 ^ n19684 ;
  assign n19687 = n19686 ^ x62 ;
  assign n19683 = ~n7353 & n9652 ;
  assign n19688 = n19687 ^ n19683 ;
  assign n19682 = x114 & n9648 ;
  assign n19689 = n19688 ^ n19682 ;
  assign n19690 = n19689 ^ x47 ;
  assign n19678 = x112 ^ x110 ;
  assign n19679 = ~n11895 & n19678 ;
  assign n5894 = x111 ^ x110 ;
  assign n19680 = n19679 ^ n5894 ;
  assign n19681 = n12206 & n19680 ;
  assign n19691 = n19690 ^ n19681 ;
  assign n19676 = n19611 & n19675 ;
  assign n19677 = n19676 ^ n19618 ;
  assign n19692 = n19691 ^ n19677 ;
  assign n19665 = x116 & n8750 ;
  assign n19664 = x118 & n8746 ;
  assign n19666 = n19665 ^ n19664 ;
  assign n19667 = n19666 ^ x59 ;
  assign n19663 = ~n8140 & n8747 ;
  assign n19668 = n19667 ^ n19663 ;
  assign n19662 = x117 & n8743 ;
  assign n19669 = n19668 ^ n19662 ;
  assign n19670 = n19669 ^ n19622 ;
  assign n19671 = n19670 ^ n19602 ;
  assign n19672 = n19671 ^ n19669 ;
  assign n19673 = ~n19608 & n19672 ;
  assign n19674 = n19673 ^ n19670 ;
  assign n19693 = n19692 ^ n19674 ;
  assign n19700 = n19699 ^ n19693 ;
  assign n19702 = n19701 ^ n19700 ;
  assign n19706 = n19705 ^ n19702 ;
  assign n19715 = n19714 ^ n19706 ;
  assign n19659 = n19624 ^ n19578 ;
  assign n19660 = n19633 & ~n19659 ;
  assign n19661 = n19660 ^ n19632 ;
  assign n19716 = n19715 ^ n19661 ;
  assign n19725 = n19724 ^ n19716 ;
  assign n19733 = n19732 ^ n19725 ;
  assign n19751 = n19750 ^ n19733 ;
  assign n19827 = ~n19728 & ~n19731 ;
  assign n19826 = n19716 & n19724 ;
  assign n19828 = n19827 ^ n19826 ;
  assign n19821 = n6445 & n10155 ;
  assign n19820 = x126 & n6687 ;
  assign n19822 = n19821 ^ n19820 ;
  assign n19823 = n19822 ^ x50 ;
  assign n19819 = x127 & n6449 ;
  assign n19824 = n19823 ^ n19819 ;
  assign n19815 = n19714 ^ n19661 ;
  assign n19816 = n19715 & n19815 ;
  assign n19817 = n19816 ^ n19714 ;
  assign n19809 = n19689 ^ n19677 ;
  assign n19810 = ~n19691 & ~n19809 ;
  assign n19811 = n19810 ^ n19689 ;
  assign n19803 = x117 & n8750 ;
  assign n19802 = x119 & n8746 ;
  assign n19804 = n19803 ^ n19802 ;
  assign n19805 = n19804 ^ x59 ;
  assign n19801 = n8405 & n8747 ;
  assign n19806 = n19805 ^ n19801 ;
  assign n19800 = x118 & n8743 ;
  assign n19807 = n19806 ^ n19800 ;
  assign n19794 = x114 & n9655 ;
  assign n19793 = x116 & n9651 ;
  assign n19795 = n19794 ^ n19793 ;
  assign n19796 = n19795 ^ x62 ;
  assign n19792 = ~n7604 & n9652 ;
  assign n19797 = n19796 ^ n19792 ;
  assign n19791 = x115 & n9648 ;
  assign n19798 = n19797 ^ n19791 ;
  assign n19784 = x111 ^ x47 ;
  assign n19787 = n19680 & ~n19784 ;
  assign n19788 = n19787 ^ x111 ;
  assign n19789 = n12206 & n19788 ;
  assign n19780 = x63 & x112 ;
  assign n19781 = n19780 ^ x113 ;
  assign n19782 = ~n9956 & n19781 ;
  assign n19783 = n19782 ^ x113 ;
  assign n19790 = n19789 ^ n19783 ;
  assign n19799 = n19798 ^ n19790 ;
  assign n19808 = n19807 ^ n19799 ;
  assign n19812 = n19811 ^ n19808 ;
  assign n19775 = n7951 & ~n9261 ;
  assign n19773 = x120 & n7954 ;
  assign n19769 = n19692 ^ n19669 ;
  assign n19770 = n19674 & n19769 ;
  assign n19771 = n19770 ^ n19669 ;
  assign n19767 = x122 & n7950 ;
  assign n19768 = n19767 ^ x56 ;
  assign n19772 = n19771 ^ n19768 ;
  assign n19774 = n19773 ^ n19772 ;
  assign n19776 = n19775 ^ n19774 ;
  assign n19766 = x121 & n7947 ;
  assign n19777 = n19776 ^ n19766 ;
  assign n19813 = n19812 ^ n19777 ;
  assign n19763 = n7187 & n10416 ;
  assign n19761 = x123 & n7183 ;
  assign n19757 = n19705 ^ n19693 ;
  assign n19758 = n19702 & n19757 ;
  assign n19759 = n19758 ^ n19693 ;
  assign n19755 = x125 & n7186 ;
  assign n19756 = n19755 ^ x53 ;
  assign n19760 = n19759 ^ n19756 ;
  assign n19762 = n19761 ^ n19760 ;
  assign n19764 = n19763 ^ n19762 ;
  assign n19754 = x124 & n7191 ;
  assign n19765 = n19764 ^ n19754 ;
  assign n19814 = n19813 ^ n19765 ;
  assign n19818 = n19817 ^ n19814 ;
  assign n19825 = n19824 ^ n19818 ;
  assign n19829 = n19828 ^ n19825 ;
  assign n19752 = n19750 ^ n19732 ;
  assign n19753 = n19733 & n19752 ;
  assign n19830 = n19829 ^ n19753 ;
  assign n19963 = x121 & n7954 ;
  assign n19962 = x123 & n7950 ;
  assign n19964 = n19963 ^ n19962 ;
  assign n19965 = n19964 ^ x56 ;
  assign n19961 = n7951 & ~n9804 ;
  assign n19966 = n19965 ^ n19961 ;
  assign n19960 = x122 & n7947 ;
  assign n19967 = n19966 ^ n19960 ;
  assign n19954 = x118 & n8750 ;
  assign n19953 = x120 & n8746 ;
  assign n19955 = n19954 ^ n19953 ;
  assign n19956 = n19955 ^ x59 ;
  assign n19952 = n8747 & n8904 ;
  assign n19957 = n19956 ^ n19952 ;
  assign n19951 = x119 & n8743 ;
  assign n19958 = n19957 ^ n19951 ;
  assign n19946 = n19798 ^ n19783 ;
  assign n19947 = n19790 & ~n19946 ;
  assign n19948 = n19947 ^ n19798 ;
  assign n19942 = ~n7860 & n9652 ;
  assign n19941 = x116 & n9648 ;
  assign n19943 = n19942 ^ n19941 ;
  assign n19939 = x115 & n9655 ;
  assign n19938 = x117 & n9651 ;
  assign n19940 = n19939 ^ n19938 ;
  assign n19944 = n19943 ^ n19940 ;
  assign n6595 = x114 ^ x113 ;
  assign n19937 = n6595 ^ x62 ;
  assign n19945 = n19944 ^ n19937 ;
  assign n19949 = n19948 ^ n19945 ;
  assign n6352 = x113 ^ x112 ;
  assign n19934 = x63 & n6352 ;
  assign n19935 = n19934 ^ n6595 ;
  assign n19936 = ~n9956 & n19935 ;
  assign n19950 = n19949 ^ n19936 ;
  assign n19959 = n19958 ^ n19950 ;
  assign n19968 = n19967 ^ n19959 ;
  assign n19927 = n19811 ^ n19807 ;
  assign n19928 = n19808 & n19927 ;
  assign n19929 = n19928 ^ n19811 ;
  assign n19969 = n19968 ^ n19929 ;
  assign n19925 = x125 & n7191 ;
  assign n19923 = n7187 & n10461 ;
  assign n19921 = x124 & n7183 ;
  assign n19917 = n19812 ^ n19771 ;
  assign n19918 = ~n19777 & ~n19917 ;
  assign n19919 = n19918 ^ n19812 ;
  assign n19915 = x126 & n7186 ;
  assign n19916 = n19915 ^ x53 ;
  assign n19920 = n19919 ^ n19916 ;
  assign n19922 = n19921 ^ n19920 ;
  assign n19924 = n19923 ^ n19922 ;
  assign n19926 = n19925 ^ n19924 ;
  assign n19970 = n19969 ^ n19926 ;
  assign n19912 = n19824 ^ n19817 ;
  assign n19913 = n19818 & n19912 ;
  assign n19914 = n19913 ^ n19824 ;
  assign n19971 = n19970 ^ n19914 ;
  assign n19908 = n19813 ^ n19759 ;
  assign n19909 = ~n19765 & ~n19908 ;
  assign n19910 = n19909 ^ n19813 ;
  assign n19898 = x127 & n6686 ;
  assign n19899 = n19898 ^ n6443 ;
  assign n19904 = n5986 & n11285 ;
  assign n19905 = n19904 ^ n19898 ;
  assign n19906 = n19899 & ~n19905 ;
  assign n19907 = n19906 ^ x49 ;
  assign n19911 = n19910 ^ n19907 ;
  assign n19972 = n19971 ^ n19911 ;
  assign n19837 = n19826 ^ n19750 ;
  assign n19831 = n19728 ^ n19725 ;
  assign n19832 = n19831 ^ n19826 ;
  assign n19833 = n19732 & ~n19832 ;
  assign n19834 = n19833 ^ n19731 ;
  assign n19835 = n19834 ^ n19825 ;
  assign n19838 = n19837 ^ n19835 ;
  assign n19884 = n19838 ^ n19828 ;
  assign n19881 = n19835 ^ n19826 ;
  assign n19885 = n19884 ^ n19881 ;
  assign n19886 = n19885 ^ n19834 ;
  assign n19836 = n19835 ^ n19827 ;
  assign n19839 = n19838 ^ n19836 ;
  assign n19868 = n19839 ^ n19835 ;
  assign n19869 = n19868 ^ n19837 ;
  assign n19840 = n19839 ^ n19834 ;
  assign n19841 = n19840 ^ n19750 ;
  assign n19843 = n19841 ^ n19825 ;
  assign n19862 = n19843 ^ n19835 ;
  assign n19870 = n19869 ^ n19862 ;
  assign n19871 = n19870 ^ n19825 ;
  assign n19873 = n19871 ^ n19869 ;
  assign n19853 = n19826 ^ n19825 ;
  assign n19854 = ~n19825 & ~n19834 ;
  assign n19855 = n19854 ^ n19825 ;
  assign n19856 = ~n19853 & n19855 ;
  assign n19857 = n19854 ^ n19827 ;
  assign n19858 = n19857 ^ n19826 ;
  assign n19859 = n19750 & n19858 ;
  assign n19860 = n19856 & n19859 ;
  assign n19861 = n19860 ^ n19857 ;
  assign n19874 = n19873 ^ n19861 ;
  assign n19863 = n19843 ^ n19838 ;
  assign n19875 = n19874 ^ n19863 ;
  assign n19876 = n19875 ^ n19871 ;
  assign n19848 = n19840 ^ n19825 ;
  assign n19847 = n19841 ^ n19838 ;
  assign n19849 = n19848 ^ n19847 ;
  assign n19850 = n19849 ^ n19848 ;
  assign n19852 = n19850 ^ n19826 ;
  assign n19877 = n19876 ^ n19852 ;
  assign n19878 = n19877 ^ n19839 ;
  assign n19879 = n19878 ^ n19826 ;
  assign n19880 = n19879 ^ n19825 ;
  assign n19887 = n19886 ^ n19880 ;
  assign n19888 = n19750 ^ n19724 ;
  assign n19891 = n19725 & n19888 ;
  assign n19892 = n19891 ^ n19724 ;
  assign n19893 = n19887 & n19892 ;
  assign n19894 = n19825 ^ n19732 ;
  assign n19895 = n19894 ^ n19827 ;
  assign n19896 = n19893 & n19895 ;
  assign n19897 = n19896 ^ n19887 ;
  assign n19973 = n19972 ^ n19897 ;
  assign n20072 = n19914 & n19970 ;
  assign n20071 = ~n19907 & n19910 ;
  assign n20073 = n20072 ^ n20071 ;
  assign n20067 = n19969 ^ n19919 ;
  assign n20068 = n19926 & n20067 ;
  assign n20069 = n20068 ^ n19969 ;
  assign n20061 = x125 & n7183 ;
  assign n20060 = x127 & n7186 ;
  assign n20062 = n20061 ^ n20060 ;
  assign n20063 = n20062 ^ x53 ;
  assign n20059 = n7187 & n10986 ;
  assign n20064 = n20063 ^ n20059 ;
  assign n20058 = x126 & n7191 ;
  assign n20065 = n20064 ^ n20058 ;
  assign n20054 = n19967 ^ n19929 ;
  assign n20055 = ~n19968 & n20054 ;
  assign n20056 = n20055 ^ n19967 ;
  assign n20048 = x122 & n7954 ;
  assign n20047 = x124 & n7950 ;
  assign n20049 = n20048 ^ n20047 ;
  assign n20050 = n20049 ^ x56 ;
  assign n20046 = n7951 & n10117 ;
  assign n20051 = n20050 ^ n20046 ;
  assign n20045 = x123 & n7947 ;
  assign n20052 = n20051 ^ n20045 ;
  assign n20037 = x116 & n9655 ;
  assign n20036 = x118 & n9651 ;
  assign n20038 = n20037 ^ n20036 ;
  assign n20039 = n20038 ^ x62 ;
  assign n20035 = ~n8140 & n9652 ;
  assign n20040 = n20039 ^ n20035 ;
  assign n20034 = x117 & n9648 ;
  assign n20041 = n20040 ^ n20034 ;
  assign n20028 = x63 & x114 ;
  assign n20029 = n20028 ^ x115 ;
  assign n20030 = ~n9956 & n20029 ;
  assign n20031 = n20030 ^ x115 ;
  assign n20032 = n20031 ^ x50 ;
  assign n20033 = n20032 ^ n19783 ;
  assign n20042 = n20041 ^ n20033 ;
  assign n19989 = x114 ^ x63 ;
  assign n19990 = n19989 ^ n19944 ;
  assign n19993 = n6595 & ~n19990 ;
  assign n19994 = n19993 ^ n19944 ;
  assign n19995 = n9956 & n19994 ;
  assign n20014 = n19995 ^ x62 ;
  assign n20020 = n19944 & ~n19995 ;
  assign n20002 = x113 & ~x114 ;
  assign n20001 = n19995 ^ n9956 ;
  assign n20011 = n20002 ^ n20001 ;
  assign n20004 = n20002 ^ x112 ;
  assign n20003 = n20002 ^ n19944 ;
  assign n20005 = n20004 ^ n20003 ;
  assign n20008 = ~n6352 & n20005 ;
  assign n20009 = n20008 ^ n20004 ;
  assign n20010 = x62 & n20009 ;
  assign n20012 = n20011 ^ n20010 ;
  assign n20015 = n20012 ^ x63 ;
  assign n20021 = n20020 ^ n20015 ;
  assign n20022 = ~n20014 & n20021 ;
  assign n20024 = n20022 ^ n20015 ;
  assign n20013 = n20001 & ~n20012 ;
  assign n20023 = n20013 & ~n20022 ;
  assign n20025 = n20024 ^ n20023 ;
  assign n20043 = n20042 ^ n20025 ;
  assign n19979 = x119 & n8750 ;
  assign n19978 = x121 & n8746 ;
  assign n19980 = n19979 ^ n19978 ;
  assign n19981 = n19980 ^ x59 ;
  assign n19977 = n8747 & n8979 ;
  assign n19982 = n19981 ^ n19977 ;
  assign n19976 = x120 & n8743 ;
  assign n19983 = n19982 ^ n19976 ;
  assign n19984 = n19983 ^ n19958 ;
  assign n19985 = n19984 ^ n19948 ;
  assign n19986 = n19985 ^ n19983 ;
  assign n19987 = n19950 & n19986 ;
  assign n19988 = n19987 ^ n19984 ;
  assign n20044 = n20043 ^ n19988 ;
  assign n20053 = n20052 ^ n20044 ;
  assign n20057 = n20056 ^ n20053 ;
  assign n20066 = n20065 ^ n20057 ;
  assign n20070 = n20069 ^ n20066 ;
  assign n20074 = n20073 ^ n20070 ;
  assign n19974 = n19911 ^ n19897 ;
  assign n19975 = ~n19972 & n19974 ;
  assign n20075 = n20074 ^ n19975 ;
  assign n20189 = n7187 & n10155 ;
  assign n20188 = x126 & n7183 ;
  assign n20190 = n20189 ^ n20188 ;
  assign n20191 = n20190 ^ x53 ;
  assign n20187 = x127 & n7191 ;
  assign n20192 = n20191 ^ n20187 ;
  assign n20178 = x120 & n8750 ;
  assign n20177 = x122 & n8746 ;
  assign n20179 = n20178 ^ n20177 ;
  assign n20180 = n20179 ^ x59 ;
  assign n20176 = n8747 & ~n9261 ;
  assign n20181 = n20180 ^ n20176 ;
  assign n20175 = x121 & n8743 ;
  assign n20182 = n20181 ^ n20175 ;
  assign n20172 = x115 & n11895 ;
  assign n20171 = x116 & n9956 ;
  assign n20173 = n20172 ^ n20171 ;
  assign n20168 = n8405 & n9652 ;
  assign n20166 = x117 & n9655 ;
  assign n20162 = n20031 ^ n19783 ;
  assign n20163 = ~n20032 & ~n20162 ;
  assign n20164 = n20163 ^ x50 ;
  assign n20160 = x119 & n9651 ;
  assign n20161 = n20160 ^ x62 ;
  assign n20165 = n20164 ^ n20161 ;
  assign n20167 = n20166 ^ n20165 ;
  assign n20169 = n20168 ^ n20167 ;
  assign n20159 = x118 & n9648 ;
  assign n20170 = n20169 ^ n20159 ;
  assign n20174 = n20173 ^ n20170 ;
  assign n20183 = n20182 ^ n20174 ;
  assign n20156 = n20041 ^ n20025 ;
  assign n20157 = ~n20042 & n20156 ;
  assign n20158 = n20157 ^ n20041 ;
  assign n20184 = n20183 ^ n20158 ;
  assign n20146 = x123 & n7954 ;
  assign n20145 = x125 & n7950 ;
  assign n20147 = n20146 ^ n20145 ;
  assign n20148 = n20147 ^ x56 ;
  assign n20144 = n7951 & n10416 ;
  assign n20149 = n20148 ^ n20144 ;
  assign n20143 = x124 & n7947 ;
  assign n20150 = n20149 ^ n20143 ;
  assign n20152 = n20150 ^ n19983 ;
  assign n20151 = n20150 ^ n20043 ;
  assign n20153 = n20152 ^ n20151 ;
  assign n20154 = n19988 & ~n20153 ;
  assign n20155 = n20154 ^ n20152 ;
  assign n20185 = n20184 ^ n20155 ;
  assign n20140 = n20056 ^ n20052 ;
  assign n20141 = n20053 & n20140 ;
  assign n20142 = n20141 ^ n20056 ;
  assign n20186 = n20185 ^ n20142 ;
  assign n20193 = n20192 ^ n20186 ;
  assign n20137 = n20069 ^ n20065 ;
  assign n20138 = n20066 & ~n20137 ;
  assign n20139 = n20138 ^ n20069 ;
  assign n20194 = n20193 ^ n20139 ;
  assign n20097 = n20071 ^ n19897 ;
  assign n20076 = n20071 ^ n19911 ;
  assign n20077 = n20076 ^ n19914 ;
  assign n20078 = n19971 & ~n20077 ;
  assign n20079 = n20078 ^ n19970 ;
  assign n20080 = n20079 ^ n20070 ;
  assign n20081 = n20080 ^ n20073 ;
  assign n20121 = n20097 ^ n20081 ;
  assign n20084 = n20080 ^ n20071 ;
  assign n20122 = n20121 ^ n20084 ;
  assign n20123 = n20122 ^ n20079 ;
  assign n20125 = n20123 ^ n20121 ;
  assign n20098 = n20097 ^ n20080 ;
  assign n20119 = n20098 ^ n20081 ;
  assign n20094 = n20072 ^ n19897 ;
  assign n20095 = n20094 ^ n20071 ;
  assign n20096 = n20095 ^ n20080 ;
  assign n20100 = n20097 ^ n20096 ;
  assign n20101 = n20100 ^ n20084 ;
  assign n20102 = n20101 ^ n20079 ;
  assign n20113 = n20102 ^ n20100 ;
  assign n20110 = n20098 ^ n20096 ;
  assign n20103 = n20102 ^ n20080 ;
  assign n20093 = n20070 & ~n20079 ;
  assign n20104 = n20096 ^ n20093 ;
  assign n20105 = ~n20103 & ~n20104 ;
  assign n20106 = n20098 ^ n20079 ;
  assign n20107 = ~n20072 & n20106 ;
  assign n20108 = n20105 & n20107 ;
  assign n20109 = n20108 ^ n20093 ;
  assign n20111 = n20110 ^ n20109 ;
  assign n20114 = n20113 ^ n20111 ;
  assign n20115 = n20114 ^ n20094 ;
  assign n20116 = n20115 ^ n20102 ;
  assign n20085 = n20084 ^ n19897 ;
  assign n20086 = n20085 ^ n20080 ;
  assign n20087 = n20086 ^ n20081 ;
  assign n20089 = n20087 ^ n20071 ;
  assign n20091 = n20089 ^ n20070 ;
  assign n20092 = n20091 ^ n20087 ;
  assign n20117 = n20116 ^ n20092 ;
  assign n20118 = n20117 ^ n20091 ;
  assign n20120 = n20119 ^ n20118 ;
  assign n20126 = n20125 ^ n20120 ;
  assign n20127 = n20126 ^ n20070 ;
  assign n20128 = n20127 ^ n20123 ;
  assign n20129 = n19907 ^ n19897 ;
  assign n20130 = ~n19911 & ~n20129 ;
  assign n20131 = n20130 ^ n19907 ;
  assign n20132 = n20128 & ~n20131 ;
  assign n20133 = n20070 ^ n19971 ;
  assign n20134 = n20133 ^ n20072 ;
  assign n20135 = n20132 & n20134 ;
  assign n20136 = n20135 ^ n20128 ;
  assign n20195 = n20194 ^ n20136 ;
  assign n20253 = x124 & n7954 ;
  assign n20252 = x126 & n7950 ;
  assign n20254 = n20253 ^ n20252 ;
  assign n20255 = n20254 ^ x56 ;
  assign n20251 = n7951 & n10461 ;
  assign n20256 = n20255 ^ n20251 ;
  assign n20250 = x125 & n7947 ;
  assign n20257 = n20256 ^ n20250 ;
  assign n20246 = n20182 ^ n20158 ;
  assign n20247 = n20183 & n20246 ;
  assign n20248 = n20247 ^ n20182 ;
  assign n20239 = n9956 ^ x116 ;
  assign n20236 = ~x117 & n9956 ;
  assign n20237 = n20236 ^ n20172 ;
  assign n20240 = n20237 ^ n12206 ;
  assign n20241 = n20239 & n20240 ;
  assign n20242 = n20241 ^ n20172 ;
  assign n20238 = x116 & n20237 ;
  assign n20243 = n20242 ^ n20238 ;
  assign n20233 = n20173 ^ n20164 ;
  assign n20234 = n20170 & n20233 ;
  assign n20235 = n20234 ^ n20173 ;
  assign n20244 = n20243 ^ n20235 ;
  assign n20230 = n8747 & ~n9804 ;
  assign n20228 = x121 & n8750 ;
  assign n20222 = x118 & n9655 ;
  assign n20221 = x120 & n9651 ;
  assign n20223 = n20222 ^ n20221 ;
  assign n20224 = n20223 ^ x62 ;
  assign n20220 = n8904 & n9652 ;
  assign n20225 = n20224 ^ n20220 ;
  assign n20219 = x119 & n9648 ;
  assign n20226 = n20225 ^ n20219 ;
  assign n20217 = x123 & n8746 ;
  assign n20218 = n20217 ^ x59 ;
  assign n20227 = n20226 ^ n20218 ;
  assign n20229 = n20228 ^ n20227 ;
  assign n20231 = n20230 ^ n20229 ;
  assign n20216 = x122 & n8743 ;
  assign n20232 = n20231 ^ n20216 ;
  assign n20245 = n20244 ^ n20232 ;
  assign n20249 = n20248 ^ n20245 ;
  assign n20258 = n20257 ^ n20249 ;
  assign n20206 = x127 & n7182 ;
  assign n20207 = n20206 ^ n7180 ;
  assign n20208 = n20206 ^ n6680 ;
  assign n20209 = n20208 ^ n20206 ;
  assign n20212 = n11285 & n20209 ;
  assign n20213 = n20212 ^ n20206 ;
  assign n20214 = n20207 & ~n20213 ;
  assign n20215 = n20214 ^ x52 ;
  assign n20259 = n20258 ^ n20215 ;
  assign n20203 = n20184 ^ n20150 ;
  assign n20204 = n20155 & n20203 ;
  assign n20205 = n20204 ^ n20150 ;
  assign n20260 = n20259 ^ n20205 ;
  assign n20200 = n20192 ^ n20142 ;
  assign n20201 = ~n20186 & n20200 ;
  assign n20202 = n20201 ^ n20192 ;
  assign n20261 = n20260 ^ n20202 ;
  assign n20196 = n20139 ^ n20136 ;
  assign n20197 = n20193 ^ n20136 ;
  assign n20198 = n20196 & n20197 ;
  assign n20199 = n20198 ^ n20193 ;
  assign n20262 = n20261 ^ n20199 ;
  assign n20310 = n20257 ^ n20248 ;
  assign n20311 = ~n20249 & n20310 ;
  assign n20312 = n20311 ^ n20257 ;
  assign n20307 = n20215 ^ n20205 ;
  assign n20308 = n20259 & n20307 ;
  assign n20309 = n20308 ^ n20215 ;
  assign n20313 = n20312 ^ n20309 ;
  assign n20301 = x125 & n7954 ;
  assign n20300 = x127 & n7950 ;
  assign n20302 = n20301 ^ n20300 ;
  assign n20303 = n20302 ^ x56 ;
  assign n20299 = n7951 & n10986 ;
  assign n20304 = n20303 ^ n20299 ;
  assign n20298 = x126 & n7947 ;
  assign n20305 = n20304 ^ n20298 ;
  assign n20289 = x119 & n9655 ;
  assign n20288 = x121 & n9651 ;
  assign n20290 = n20289 ^ n20288 ;
  assign n20291 = n20290 ^ x62 ;
  assign n20287 = n8979 & n9652 ;
  assign n20292 = n20291 ^ n20287 ;
  assign n20286 = x120 & n9648 ;
  assign n20293 = n20292 ^ n20286 ;
  assign n20294 = n20293 ^ x53 ;
  assign n20282 = x118 ^ x116 ;
  assign n20283 = ~n11895 & n20282 ;
  assign n7335 = x117 ^ x116 ;
  assign n20284 = n20283 ^ n7335 ;
  assign n20285 = n12206 & n20284 ;
  assign n20295 = n20294 ^ n20285 ;
  assign n20280 = n20235 & ~n20243 ;
  assign n20281 = n20280 ^ n20241 ;
  assign n20296 = n20295 ^ n20281 ;
  assign n20270 = x122 & n8750 ;
  assign n20269 = x124 & n8746 ;
  assign n20271 = n20270 ^ n20269 ;
  assign n20272 = n20271 ^ x59 ;
  assign n20268 = n8747 & n10117 ;
  assign n20273 = n20272 ^ n20268 ;
  assign n20267 = x123 & n8743 ;
  assign n20274 = n20273 ^ n20267 ;
  assign n20275 = n20274 ^ n20244 ;
  assign n20276 = n20275 ^ n20226 ;
  assign n20277 = n20276 ^ n20274 ;
  assign n20278 = ~n20232 & n20277 ;
  assign n20279 = n20278 ^ n20275 ;
  assign n20297 = n20296 ^ n20279 ;
  assign n20306 = n20305 ^ n20297 ;
  assign n20314 = n20313 ^ n20306 ;
  assign n20263 = n20202 ^ n20199 ;
  assign n20264 = n20260 ^ n20199 ;
  assign n20265 = ~n20263 & n20264 ;
  assign n20266 = n20265 ^ n20260 ;
  assign n20315 = n20314 ^ n20266 ;
  assign n20316 = n20312 ^ n20305 ;
  assign n20319 = ~n20306 & n20316 ;
  assign n20317 = n20309 ^ n20306 ;
  assign n20321 = n20319 ^ n20317 ;
  assign n20322 = ~n20266 & ~n20321 ;
  assign n20329 = n20322 ^ n20319 ;
  assign n20323 = n20322 ^ n20309 ;
  assign n20325 = n20309 ^ n20305 ;
  assign n20326 = n20325 ^ n20306 ;
  assign n20327 = n20326 ^ n20316 ;
  assign n20328 = n20323 & ~n20327 ;
  assign n20330 = n20329 ^ n20328 ;
  assign n20331 = n20330 ^ n20317 ;
  assign n20381 = ~n20297 & ~n20305 ;
  assign n20382 = n20381 ^ n20306 ;
  assign n20383 = ~n20266 & n20382 ;
  assign n20384 = n20381 ^ n20309 ;
  assign n20385 = n20381 ^ n20312 ;
  assign n20386 = n20384 & ~n20385 ;
  assign n20387 = n20386 ^ n20312 ;
  assign n20388 = n20383 & ~n20387 ;
  assign n20389 = n20331 & n20388 ;
  assign n20374 = n7951 & n10155 ;
  assign n20373 = x126 & n7954 ;
  assign n20375 = n20374 ^ n20373 ;
  assign n20376 = n20375 ^ x56 ;
  assign n20372 = x127 & n7947 ;
  assign n20377 = n20376 ^ n20372 ;
  assign n20360 = x120 & n9655 ;
  assign n20359 = x122 & n9651 ;
  assign n20361 = n20360 ^ n20359 ;
  assign n20362 = n20361 ^ x62 ;
  assign n20358 = ~n9261 & n9652 ;
  assign n20363 = n20362 ^ n20358 ;
  assign n20357 = x121 & n9648 ;
  assign n20364 = n20363 ^ n20357 ;
  assign n20352 = x63 & x118 ;
  assign n20353 = n20352 ^ x119 ;
  assign n20354 = ~n9956 & n20353 ;
  assign n20355 = n20354 ^ x119 ;
  assign n20344 = x117 ^ x53 ;
  assign n20347 = n20284 & ~n20344 ;
  assign n20348 = n20347 ^ x117 ;
  assign n20349 = n12206 & n20348 ;
  assign n20356 = n20355 ^ n20349 ;
  assign n20365 = n20364 ^ n20356 ;
  assign n20342 = x124 & n8743 ;
  assign n20340 = n8747 & n10416 ;
  assign n20338 = x123 & n8750 ;
  assign n20334 = n20293 ^ n20281 ;
  assign n20335 = ~n20295 & ~n20334 ;
  assign n20336 = n20335 ^ n20293 ;
  assign n20332 = x125 & n8746 ;
  assign n20333 = n20332 ^ x59 ;
  assign n20337 = n20336 ^ n20333 ;
  assign n20339 = n20338 ^ n20337 ;
  assign n20341 = n20340 ^ n20339 ;
  assign n20343 = n20342 ^ n20341 ;
  assign n20366 = n20365 ^ n20343 ;
  assign n20368 = n20366 ^ n20274 ;
  assign n20367 = n20366 ^ n20296 ;
  assign n20369 = n20368 ^ n20367 ;
  assign n20370 = n20279 & n20369 ;
  assign n20371 = n20370 ^ n20368 ;
  assign n20378 = n20377 ^ n20371 ;
  assign n20379 = n20378 ^ n20331 ;
  assign n20390 = n20389 ^ n20379 ;
  assign n20519 = n20377 ^ n20366 ;
  assign n20520 = ~n20371 & ~n20519 ;
  assign n20521 = n20520 ^ n20366 ;
  assign n20513 = x124 & n8750 ;
  assign n20512 = x126 & n8746 ;
  assign n20514 = n20513 ^ n20512 ;
  assign n20515 = n20514 ^ x59 ;
  assign n20511 = n8747 & n10461 ;
  assign n20516 = n20515 ^ n20511 ;
  assign n20510 = x125 & n8743 ;
  assign n20517 = n20516 ^ n20510 ;
  assign n20503 = x121 & n9655 ;
  assign n20502 = x123 & n9651 ;
  assign n20504 = n20503 ^ n20502 ;
  assign n20505 = n20504 ^ x62 ;
  assign n20501 = n9652 & ~n9804 ;
  assign n20506 = n20505 ^ n20501 ;
  assign n20500 = x122 & n9648 ;
  assign n20507 = n20506 ^ n20500 ;
  assign n20496 = x63 & n7838 ;
  assign n20497 = n20496 ^ n8114 ;
  assign n20498 = ~n9956 & n20497 ;
  assign n20499 = n20498 ^ n8114 ;
  assign n20508 = n20507 ^ n20499 ;
  assign n20489 = n20364 ^ n20355 ;
  assign n20490 = n20356 & ~n20489 ;
  assign n20491 = n20490 ^ n20364 ;
  assign n20509 = n20508 ^ n20491 ;
  assign n20518 = n20517 ^ n20509 ;
  assign n20522 = n20521 ^ n20518 ;
  assign n20485 = n20365 ^ n20336 ;
  assign n20486 = ~n20343 & ~n20485 ;
  assign n20487 = n20486 ^ n20365 ;
  assign n7955 = n7954 ^ n7951 ;
  assign n20482 = x127 & n7955 ;
  assign n20481 = n7951 & n10154 ;
  assign n20483 = n20482 ^ n20481 ;
  assign n20484 = n20483 ^ x56 ;
  assign n20488 = n20487 ^ n20484 ;
  assign n20523 = n20522 ^ n20488 ;
  assign n20392 = ~n20309 & ~n20312 ;
  assign n20477 = n20392 ^ n20313 ;
  assign n20391 = ~n20381 & ~n20383 ;
  assign n20464 = n20382 ^ n20266 ;
  assign n20394 = n20387 ^ n20378 ;
  assign n20393 = n20392 ^ n20382 ;
  assign n20395 = n20394 ^ n20393 ;
  assign n20467 = n20464 ^ n20395 ;
  assign n20463 = n20394 ^ n20382 ;
  assign n20468 = n20467 ^ n20463 ;
  assign n20469 = n20468 ^ n20387 ;
  assign n20471 = n20469 ^ n20467 ;
  assign n20410 = n20387 ^ n20382 ;
  assign n20416 = n20410 ^ n20392 ;
  assign n20411 = n20410 ^ n20266 ;
  assign n20412 = n20411 ^ n20387 ;
  assign n20452 = n20416 ^ n20412 ;
  assign n20453 = n20452 ^ n20382 ;
  assign n20454 = n20453 ^ n20378 ;
  assign n20456 = n20454 ^ n20452 ;
  assign n20422 = n20412 ^ n20394 ;
  assign n20424 = n20422 ^ n20382 ;
  assign n20429 = n20424 ^ n20266 ;
  assign n20430 = n20422 ^ n20410 ;
  assign n20431 = n20430 ^ n20266 ;
  assign n20432 = ~n20429 & n20431 ;
  assign n20413 = n20412 ^ n20392 ;
  assign n20414 = n20413 ^ n20394 ;
  assign n20433 = n20432 ^ n20414 ;
  assign n20434 = n20433 ^ n20422 ;
  assign n20435 = n20434 ^ n20387 ;
  assign n20436 = n20422 ^ n20266 ;
  assign n20437 = n20436 ^ n20387 ;
  assign n20438 = ~n20435 & n20437 ;
  assign n20417 = n20416 ^ n20387 ;
  assign n20420 = n20417 ^ n20394 ;
  assign n20439 = n20420 ^ n20382 ;
  assign n20440 = n20439 ^ n20410 ;
  assign n20441 = n20414 ^ n20382 ;
  assign n20442 = n20441 ^ n20410 ;
  assign n20443 = n20440 & ~n20442 ;
  assign n20444 = n20438 & n20443 ;
  assign n20445 = n20444 ^ n20432 ;
  assign n20446 = n20445 ^ n20266 ;
  assign n20426 = n20424 ^ n20410 ;
  assign n20447 = n20446 ^ n20426 ;
  assign n20418 = n20417 ^ n20412 ;
  assign n20448 = n20447 ^ n20418 ;
  assign n20449 = n20448 ^ n20410 ;
  assign n20457 = n20456 ^ n20449 ;
  assign n20458 = n20457 ^ n20382 ;
  assign n20459 = n20458 ^ n20454 ;
  assign n20402 = n20393 ^ n20266 ;
  assign n20403 = n20402 ^ n20394 ;
  assign n20396 = n20395 ^ n20382 ;
  assign n20397 = n20396 ^ n20266 ;
  assign n20398 = n20397 ^ n20387 ;
  assign n20404 = n20403 ^ n20398 ;
  assign n20406 = n20404 ^ n20395 ;
  assign n20408 = n20406 ^ n20387 ;
  assign n20409 = n20408 ^ n20404 ;
  assign n20460 = n20459 ^ n20409 ;
  assign n20461 = n20460 ^ n20397 ;
  assign n20462 = n20461 ^ n20408 ;
  assign n20472 = n20471 ^ n20462 ;
  assign n20473 = n20472 ^ n20378 ;
  assign n20474 = n20473 ^ n20469 ;
  assign n20475 = n20391 & ~n20474 ;
  assign n20478 = n20378 & n20475 ;
  assign n20479 = n20477 & n20478 ;
  assign n20476 = n20475 ^ n20474 ;
  assign n20480 = n20479 ^ n20476 ;
  assign n20524 = n20523 ^ n20480 ;
  assign n20573 = ~n20499 & n20507 ;
  assign n20567 = n9956 ^ x119 ;
  assign n20568 = x63 & ~x118 ;
  assign n20569 = n20568 ^ x120 ;
  assign n20570 = x119 & n20569 ;
  assign n20571 = n20570 ^ x120 ;
  assign n20572 = n20567 & n20571 ;
  assign n20574 = n20573 ^ n20572 ;
  assign n20561 = x122 & n9655 ;
  assign n20560 = x124 & n9651 ;
  assign n20562 = n20561 ^ n20560 ;
  assign n20563 = n20562 ^ x62 ;
  assign n20559 = n9652 & n10117 ;
  assign n20564 = n20563 ^ n20559 ;
  assign n20558 = x123 & n9648 ;
  assign n20565 = n20564 ^ n20558 ;
  assign n20552 = x63 & x120 ;
  assign n20553 = n20552 ^ x121 ;
  assign n20554 = ~n9956 & n20553 ;
  assign n20555 = n20554 ^ x121 ;
  assign n20556 = n20555 ^ x56 ;
  assign n20557 = n20556 ^ n20355 ;
  assign n20566 = n20565 ^ n20557 ;
  assign n20575 = n20574 ^ n20566 ;
  assign n20540 = x125 & n8750 ;
  assign n20539 = x127 & n8746 ;
  assign n20541 = n20540 ^ n20539 ;
  assign n20542 = n20541 ^ x59 ;
  assign n20538 = n8747 & n10986 ;
  assign n20543 = n20542 ^ n20538 ;
  assign n20537 = x126 & n8743 ;
  assign n20544 = n20543 ^ n20537 ;
  assign n20545 = n20544 ^ n20517 ;
  assign n20546 = n20545 ^ n20491 ;
  assign n20547 = n20546 ^ n20544 ;
  assign n20548 = n20509 & n20547 ;
  assign n20549 = n20548 ^ n20545 ;
  assign n20576 = n20575 ^ n20549 ;
  assign n20532 = ~n20484 & n20487 ;
  assign n20533 = n20532 ^ n20518 ;
  assign n20534 = n20522 & ~n20533 ;
  assign n20535 = n20534 ^ n20521 ;
  assign n20536 = n20535 ^ n20522 ;
  assign n20577 = n20576 ^ n20536 ;
  assign n20578 = n20577 ^ n20532 ;
  assign n20529 = ~n20487 & n20488 ;
  assign n20530 = n20529 ^ n20480 ;
  assign n20531 = ~n20523 & ~n20530 ;
  assign n20579 = n20578 ^ n20531 ;
  assign n20693 = n8747 & n10155 ;
  assign n20692 = x126 & n8750 ;
  assign n20694 = n20693 ^ n20692 ;
  assign n20695 = n20694 ^ x59 ;
  assign n20691 = x127 & n8743 ;
  assign n20696 = n20695 ^ n20691 ;
  assign n20687 = x121 & n11895 ;
  assign n20686 = x122 & n9956 ;
  assign n20688 = n20687 ^ n20686 ;
  assign n20683 = n9652 & n10416 ;
  assign n20681 = x123 & n9655 ;
  assign n20677 = n20555 ^ n20355 ;
  assign n20678 = ~n20556 & ~n20677 ;
  assign n20679 = n20678 ^ x56 ;
  assign n20675 = x125 & n9651 ;
  assign n20676 = n20675 ^ x62 ;
  assign n20680 = n20679 ^ n20676 ;
  assign n20682 = n20681 ^ n20680 ;
  assign n20684 = n20683 ^ n20682 ;
  assign n20674 = x124 & n9648 ;
  assign n20685 = n20684 ^ n20674 ;
  assign n20689 = n20688 ^ n20685 ;
  assign n20671 = n20574 ^ n20565 ;
  assign n20672 = n20566 & n20671 ;
  assign n20673 = n20672 ^ n20574 ;
  assign n20690 = n20689 ^ n20673 ;
  assign n20697 = n20696 ^ n20690 ;
  assign n20668 = n20575 ^ n20544 ;
  assign n20669 = n20549 & ~n20668 ;
  assign n20670 = n20669 ^ n20544 ;
  assign n20698 = n20697 ^ n20670 ;
  assign n20581 = n20518 & n20521 ;
  assign n20664 = n20581 ^ n20522 ;
  assign n20580 = n20532 ^ n20488 ;
  assign n20648 = n20580 ^ n20480 ;
  assign n20583 = n20576 ^ n20535 ;
  assign n20582 = n20581 ^ n20580 ;
  assign n20584 = n20583 ^ n20582 ;
  assign n20651 = n20648 ^ n20584 ;
  assign n20603 = n20583 ^ n20580 ;
  assign n20652 = n20651 ^ n20603 ;
  assign n20653 = n20652 ^ n20535 ;
  assign n20655 = n20653 ^ n20651 ;
  assign n20641 = n20582 ^ n20535 ;
  assign n20631 = n20581 ^ n20480 ;
  assign n20632 = n20631 ^ n20580 ;
  assign n20642 = n20641 ^ n20632 ;
  assign n20643 = n20642 ^ n20580 ;
  assign n20644 = n20643 ^ n20576 ;
  assign n20597 = n20576 ^ n20480 ;
  assign n20600 = n20597 ^ n20583 ;
  assign n20609 = n20600 ^ n20584 ;
  assign n20602 = n20597 ^ n20584 ;
  assign n20610 = n20609 ^ n20602 ;
  assign n20613 = n20576 & n20610 ;
  assign n20614 = n20613 ^ n20600 ;
  assign n20615 = n20614 ^ n20603 ;
  assign n20616 = n20615 ^ n20535 ;
  assign n20617 = n20609 ^ n20603 ;
  assign n20618 = n20617 ^ n20535 ;
  assign n20619 = ~n20616 & n20618 ;
  assign n20604 = n20603 ^ n20602 ;
  assign n20620 = n20604 ^ n20584 ;
  assign n20606 = n20604 ^ n20535 ;
  assign n20621 = n20620 ^ n20606 ;
  assign n20624 = n20480 & ~n20621 ;
  assign n20625 = n20619 & n20624 ;
  assign n20626 = n20625 ^ n20613 ;
  assign n20627 = n20626 ^ n20609 ;
  assign n20607 = n20606 ^ n20602 ;
  assign n20628 = n20627 ^ n20607 ;
  assign n20598 = n20597 ^ n20580 ;
  assign n20629 = n20628 ^ n20598 ;
  assign n20630 = n20629 ^ n20606 ;
  assign n20633 = n20632 ^ n20630 ;
  assign n20645 = n20644 ^ n20633 ;
  assign n20585 = n20584 ^ n20580 ;
  assign n20586 = n20585 ^ n20480 ;
  assign n20646 = n20645 ^ n20586 ;
  assign n20587 = n20586 ^ n20535 ;
  assign n20594 = n20587 ^ n20583 ;
  assign n20588 = n20587 ^ n20480 ;
  assign n20593 = n20588 ^ n20584 ;
  assign n20595 = n20594 ^ n20593 ;
  assign n20596 = n20595 ^ n20535 ;
  assign n20647 = n20646 ^ n20596 ;
  assign n20656 = n20655 ^ n20647 ;
  assign n20657 = n20656 ^ n20576 ;
  assign n20658 = n20657 ^ n20653 ;
  assign n20659 = n20484 ^ n20480 ;
  assign n20660 = ~n20488 & n20659 ;
  assign n20661 = n20660 ^ n20484 ;
  assign n20662 = n20658 & n20661 ;
  assign n20665 = n20576 & n20662 ;
  assign n20666 = n20664 & n20665 ;
  assign n20663 = n20662 ^ n20658 ;
  assign n20667 = n20666 ^ n20663 ;
  assign n20699 = n20698 ^ n20667 ;
  assign n8751 = n8750 ^ n8747 ;
  assign n20728 = x127 & n8751 ;
  assign n20727 = n8747 & n10154 ;
  assign n20729 = n20728 ^ n20727 ;
  assign n20730 = n20729 ^ x59 ;
  assign n20724 = n20696 ^ n20673 ;
  assign n20725 = ~n20690 & n20724 ;
  assign n20726 = n20725 ^ n20696 ;
  assign n20731 = n20730 ^ n20726 ;
  assign n20718 = x124 & n9655 ;
  assign n20717 = x126 & n9651 ;
  assign n20719 = n20718 ^ n20717 ;
  assign n20720 = n20719 ^ x62 ;
  assign n20716 = n9652 & n10461 ;
  assign n20721 = n20720 ^ n20716 ;
  assign n20715 = x125 & n9648 ;
  assign n20722 = n20721 ^ n20715 ;
  assign n20709 = n9956 ^ x122 ;
  assign n20706 = ~x123 & n9956 ;
  assign n20707 = n20706 ^ n20687 ;
  assign n20710 = n20707 ^ n12206 ;
  assign n20711 = n20709 & n20710 ;
  assign n20712 = n20711 ^ n20687 ;
  assign n20708 = x122 & n20707 ;
  assign n20713 = n20712 ^ n20708 ;
  assign n20703 = n20688 ^ n20679 ;
  assign n20704 = n20685 & n20703 ;
  assign n20705 = n20704 ^ n20688 ;
  assign n20714 = n20713 ^ n20705 ;
  assign n20723 = n20722 ^ n20714 ;
  assign n20732 = n20731 ^ n20723 ;
  assign n20700 = n20670 ^ n20667 ;
  assign n20701 = n20698 & ~n20700 ;
  assign n20702 = n20701 ^ n20670 ;
  assign n20733 = n20732 ^ n20702 ;
  assign n20748 = x125 & n9655 ;
  assign n20747 = x127 & n9651 ;
  assign n20749 = n20748 ^ n20747 ;
  assign n20750 = n20749 ^ x62 ;
  assign n20746 = n9652 & n10986 ;
  assign n20751 = n20750 ^ n20746 ;
  assign n20745 = x126 & n9648 ;
  assign n20752 = n20751 ^ n20745 ;
  assign n20753 = n20752 ^ x59 ;
  assign n20741 = x124 ^ x122 ;
  assign n20742 = ~n11895 & n20741 ;
  assign n20743 = n20742 ^ n8961 ;
  assign n20744 = n12206 & n20743 ;
  assign n20754 = n20753 ^ n20744 ;
  assign n20739 = n20705 & ~n20713 ;
  assign n20740 = n20739 ^ n20711 ;
  assign n20755 = n20754 ^ n20740 ;
  assign n20736 = n20731 ^ n20714 ;
  assign n20737 = n20736 ^ n20702 ;
  assign n20738 = ~n20723 & n20737 ;
  assign n20756 = n20755 ^ n20738 ;
  assign n20734 = n20726 ^ n20702 ;
  assign n20735 = ~n20731 & ~n20734 ;
  assign n20757 = n20756 ^ n20735 ;
  assign n20798 = n20723 & n20726 ;
  assign n20780 = n20714 & n20722 ;
  assign n20781 = n20780 ^ n20755 ;
  assign n20799 = n20798 ^ n20781 ;
  assign n20800 = n20702 & n20799 ;
  assign n20801 = n20732 & n20800 ;
  assign n20802 = n20801 ^ n20755 ;
  assign n20782 = n20755 ^ n20730 ;
  assign n20783 = n20782 ^ n20731 ;
  assign n20784 = n20783 ^ n20782 ;
  assign n20785 = n20782 ^ n20726 ;
  assign n20786 = n20726 ^ n20723 ;
  assign n20787 = n20786 ^ n20782 ;
  assign n20788 = ~n20785 & ~n20787 ;
  assign n20789 = n20788 ^ n20782 ;
  assign n20790 = n20784 & n20789 ;
  assign n20791 = n20790 ^ n20782 ;
  assign n20792 = n20781 & n20791 ;
  assign n20803 = n20802 ^ n20792 ;
  assign n20772 = n9537 & n11895 ;
  assign n20771 = x125 & n12206 ;
  assign n20773 = n20772 ^ n20771 ;
  assign n20768 = x126 & n9655 ;
  assign n20766 = n9652 & n10155 ;
  assign n20759 = x123 ^ x59 ;
  assign n20762 = n20743 & ~n20759 ;
  assign n20763 = n20762 ^ x123 ;
  assign n20764 = n12206 & n20763 ;
  assign n20765 = n20764 ^ x62 ;
  assign n20767 = n20766 ^ n20765 ;
  assign n20769 = n20768 ^ n20767 ;
  assign n20758 = x127 & n9648 ;
  assign n20770 = n20769 ^ n20758 ;
  assign n20774 = n20773 ^ n20770 ;
  assign n20775 = n20774 ^ n20752 ;
  assign n20776 = n20775 ^ n20740 ;
  assign n20777 = n20776 ^ n20774 ;
  assign n20778 = ~n20754 & ~n20777 ;
  assign n20779 = n20778 ^ n20775 ;
  assign n20804 = n20803 ^ n20779 ;
  assign n20817 = n9848 & n9956 ;
  assign n20813 = n20773 ^ n20764 ;
  assign n20814 = ~n20770 & ~n20813 ;
  assign n20815 = n20814 ^ n20773 ;
  assign n9656 = n9655 ^ n9652 ;
  assign n20810 = x127 & n9656 ;
  assign n20809 = n9652 & n10154 ;
  assign n20811 = n20810 ^ n20809 ;
  assign n20808 = n20772 ^ x62 ;
  assign n20812 = n20811 ^ n20808 ;
  assign n20816 = n20815 ^ n20812 ;
  assign n20818 = n20817 ^ n20816 ;
  assign n20805 = n20803 ^ n20774 ;
  assign n20806 = ~n20779 & ~n20805 ;
  assign n20807 = n20806 ^ n20774 ;
  assign n20819 = n20818 ^ n20807 ;
  assign n20853 = n20815 ^ n20807 ;
  assign n20854 = n20818 & n20853 ;
  assign n20855 = n20854 ^ n20815 ;
  assign n20820 = x126 ^ x124 ;
  assign n20826 = x63 & n20820 ;
  assign n20821 = x127 ^ x125 ;
  assign n20827 = n20826 ^ n20821 ;
  assign n20851 = ~n9956 & n20827 ;
  assign n20843 = n20811 ^ x126 ;
  assign n20844 = x63 & n9848 ;
  assign n20845 = n20843 & n20844 ;
  assign n20830 = n20811 ^ x62 ;
  assign n20829 = x125 ^ x63 ;
  assign n20831 = n20830 ^ n20829 ;
  assign n20833 = n20820 ^ x125 ;
  assign n20834 = n20833 ^ n20830 ;
  assign n20835 = n20834 ^ n20820 ;
  assign n20838 = n9537 & ~n20835 ;
  assign n20839 = n20838 ^ n20820 ;
  assign n20840 = x62 & n20839 ;
  assign n20841 = ~n20831 & n20840 ;
  assign n20842 = n20841 ^ n20830 ;
  assign n20846 = n20845 ^ n20842 ;
  assign n20828 = n20821 ^ x62 ;
  assign n20847 = n20846 ^ n20828 ;
  assign n20852 = n20851 ^ n20847 ;
  assign n20856 = n20855 ^ n20852 ;
  assign n20870 = n20855 ^ n20846 ;
  assign n20871 = ~n20852 & ~n20870 ;
  assign n20867 = x124 & x126 ;
  assign n20868 = n11895 & n20867 ;
  assign n20857 = x127 ^ x62 ;
  assign n20860 = ~x125 & ~n20857 ;
  assign n20861 = n20860 ^ x62 ;
  assign n20862 = n20846 ^ x63 ;
  assign n20863 = n20862 ^ x127 ;
  assign n20864 = n20863 ^ n20846 ;
  assign n20865 = n20861 & n20864 ;
  assign n20866 = n20865 ^ n20862 ;
  assign n20869 = n20868 ^ n20866 ;
  assign n20872 = n20871 ^ n20869 ;
  assign y0 = n129 ;
  assign y1 = n132 ;
  assign y2 = n149 ;
  assign y3 = n184 ;
  assign y4 = n218 ;
  assign y5 = n272 ;
  assign y6 = n310 ;
  assign y7 = n359 ;
  assign y8 = ~n416 ;
  assign y9 = n473 ;
  assign y10 = n539 ;
  assign y11 = n617 ;
  assign y12 = n683 ;
  assign y13 = n759 ;
  assign y14 = n840 ;
  assign y15 = n920 ;
  assign y16 = n1013 ;
  assign y17 = n1106 ;
  assign y18 = n1194 ;
  assign y19 = n1293 ;
  assign y20 = n1399 ;
  assign y21 = n1500 ;
  assign y22 = n1612 ;
  assign y23 = n1731 ;
  assign y24 = n1845 ;
  assign y25 = n1970 ;
  assign y26 = n2108 ;
  assign y27 = n2238 ;
  assign y28 = n2375 ;
  assign y29 = ~n2528 ;
  assign y30 = n2673 ;
  assign y31 = n2825 ;
  assign y32 = n2984 ;
  assign y33 = n3140 ;
  assign y34 = ~n3313 ;
  assign y35 = ~n3484 ;
  assign y36 = ~n3650 ;
  assign y37 = ~n3828 ;
  assign y38 = ~n4021 ;
  assign y39 = ~n4204 ;
  assign y40 = n4400 ;
  assign y41 = n4605 ;
  assign y42 = n4805 ;
  assign y43 = n5011 ;
  assign y44 = n5228 ;
  assign y45 = n5440 ;
  assign y46 = n5660 ;
  assign y47 = ~n5893 ;
  assign y48 = ~n6120 ;
  assign y49 = n6351 ;
  assign y50 = n6591 ;
  assign y51 = n6830 ;
  assign y52 = n7083 ;
  assign y53 = n7334 ;
  assign y54 = n7581 ;
  assign y55 = ~n7837 ;
  assign y56 = n8110 ;
  assign y57 = ~n8382 ;
  assign y58 = ~n8652 ;
  assign y59 = ~n8937 ;
  assign y60 = n9232 ;
  assign y61 = n9530 ;
  assign y62 = n9841 ;
  assign y63 = n10140 ;
  assign y64 = ~n10443 ;
  assign y65 = n10728 ;
  assign y66 = n11003 ;
  assign y67 = n11273 ;
  assign y68 = ~n11547 ;
  assign y69 = ~n11824 ;
  assign y70 = ~n12099 ;
  assign y71 = n12368 ;
  assign y72 = n12618 ;
  assign y73 = ~n12878 ;
  assign y74 = ~n13134 ;
  assign y75 = n13380 ;
  assign y76 = ~n13613 ;
  assign y77 = n13853 ;
  assign y78 = ~n14087 ;
  assign y79 = n14326 ;
  assign y80 = ~n14556 ;
  assign y81 = ~n14809 ;
  assign y82 = n15024 ;
  assign y83 = ~n15256 ;
  assign y84 = n15456 ;
  assign y85 = n15686 ;
  assign y86 = n15885 ;
  assign y87 = ~n16071 ;
  assign y88 = n16256 ;
  assign y89 = ~n16447 ;
  assign y90 = n16623 ;
  assign y91 = ~n16874 ;
  assign y92 = n17049 ;
  assign y93 = ~n17213 ;
  assign y94 = ~n17368 ;
  assign y95 = ~n17561 ;
  assign y96 = n17708 ;
  assign y97 = n17858 ;
  assign y98 = n18004 ;
  assign y99 = n18182 ;
  assign y100 = ~n18313 ;
  assign y101 = ~n18446 ;
  assign y102 = n18581 ;
  assign y103 = ~n18700 ;
  assign y104 = n18901 ;
  assign y105 = n19026 ;
  assign y106 = n19137 ;
  assign y107 = ~n19243 ;
  assign y108 = ~n19379 ;
  assign y109 = n19561 ;
  assign y110 = ~n19658 ;
  assign y111 = n19751 ;
  assign y112 = n19830 ;
  assign y113 = n19973 ;
  assign y114 = ~n20075 ;
  assign y115 = ~n20195 ;
  assign y116 = n20262 ;
  assign y117 = n20315 ;
  assign y118 = ~n20390 ;
  assign y119 = ~n20524 ;
  assign y120 = ~n20579 ;
  assign y121 = ~n20699 ;
  assign y122 = n20733 ;
  assign y123 = ~n20757 ;
  assign y124 = ~n20804 ;
  assign y125 = ~n20819 ;
  assign y126 = n20856 ;
  assign y127 = ~n20872 ;
endmodule
