module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n545 , n546 , n547 , n550 , n551 , n553 , n555 , n556 , n558 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n573 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n583 , n585 , n586 , n588 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n608 , n610 , n611 , n613 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n623 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n638 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n648 , n650 , n651 , n653 , n655 , n656 , n658 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n678 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n693 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n713 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n728 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n781 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n791 , n793 , n794 , n796 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n806 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n816 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n826 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n892 , n894 , n895 , n897 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n907 , n909 , n910 , n912 , n914 , n915 , n917 , n919 , n920 , n922 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n942 , n944 , n945 , n947 , n949 , n950 , n952 , n954 , n955 , n957 , n959 , n960 , n962 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n982 , n984 , n985 , n987 , n989 , n990 , n992 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1042 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1057 , n1059 , n1060 , n1062 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1092 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1107 , n1109 , n1110 , n1112 , n1114 , n1115 , n1117 , n1119 , n1120 , n1122 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1152 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1223 , n1224 , n1225 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1241 , n1243 , n1244 , n1246 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1256 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1271 , n1273 , n1274 , n1276 , n1278 , n1279 , n1281 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1296 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1306 , n1308 , n1309 , n1311 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1321 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1341 , n1343 , n1344 , n1346 , n1348 , n1349 , n1351 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1361 , n1363 , n1364 , n1366 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1376 , n1378 , n1379 , n1381 , n1383 , n1384 , n1386 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1396 , n1398 , n1399 , n1401 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1436 , n1438 , n1439 , n1441 , n1443 , n1444 , n1446 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1456 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1471 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1481 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1491 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1552 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1567 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1592 , n1594 , n1595 , n1597 , n1599 , n1600 , n1602 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1632 , n1634 , n1635 , n1637 , n1639 , n1640 , n1642 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1662 , n1664 , n1665 , n1667 , n1669 , n1670 , n1672 , n1674 , n1675 , n1677 , n1679 , n1680 , n1682 , n1684 , n1685 , n1687 , n1689 , n1690 , n1692 , n1694 , n1695 , n1697 , n1699 , n1700 , n1702 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1712 , n1714 , n1715 , n1717 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1732 , n1734 , n1735 , n1737 , n1739 , n1740 , n1742 , n1744 , n1745 , n1747 , n1749 , n1750 , n1752 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1762 , n1764 , n1765 , n1767 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1792 , n1794 , n1795 , n1797 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1815 , n1816 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2355 , n2356 , n2357 , n2358 , n2359 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 ;
  assign n1164 = x384 ^ x256 ;
  assign n1165 = x511 ^ x383 ;
  assign n1822 = x511 ^ x382 ;
  assign n1166 = ~x380 & x508 ;
  assign n1167 = x509 ^ x381 ;
  assign n1168 = x507 ^ x379 ;
  assign n1169 = x455 ^ x327 ;
  assign n1172 = x454 ^ x326 ;
  assign n1173 = x453 ^ x325 ;
  assign n1174 = ~n1172 & ~n1173 ;
  assign n1176 = x451 ^ x323 ;
  assign n1175 = x323 & ~x451 ;
  assign n1177 = n1176 ^ n1175 ;
  assign n1179 = x324 & ~x452 ;
  assign n1178 = x452 ^ x324 ;
  assign n1180 = n1179 ^ n1178 ;
  assign n1181 = ~n1177 & ~n1180 ;
  assign n1182 = n1174 & n1181 ;
  assign n1183 = x450 ^ x322 ;
  assign n1187 = x448 ^ x320 ;
  assign n1186 = x320 & ~x448 ;
  assign n1188 = n1187 ^ n1186 ;
  assign n1190 = x444 ^ x316 ;
  assign n1189 = x316 & ~x444 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1192 = ~x319 & x447 ;
  assign n1194 = x445 ^ x317 ;
  assign n1193 = x317 & ~x445 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1197 = x446 ^ x318 ;
  assign n1196 = x318 & ~x446 ;
  assign n1198 = n1197 ^ n1196 ;
  assign n1199 = ~n1195 & ~n1198 ;
  assign n1200 = n1192 & n1199 ;
  assign n1201 = n1200 ^ n1199 ;
  assign n1202 = x443 ^ x315 ;
  assign n1204 = x300 & ~x428 ;
  assign n1203 = x428 ^ x300 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1206 = x427 ^ x299 ;
  assign n1207 = x425 ^ x297 ;
  assign n1208 = x426 ^ x298 ;
  assign n1209 = ~n1207 & ~n1208 ;
  assign n1211 = x423 ^ x295 ;
  assign n1210 = x295 & ~x423 ;
  assign n1212 = n1211 ^ n1210 ;
  assign n1214 = x424 ^ x296 ;
  assign n1213 = x296 & ~x424 ;
  assign n1215 = n1214 ^ n1213 ;
  assign n1216 = ~n1212 & ~n1215 ;
  assign n1217 = n1209 & n1216 ;
  assign n1218 = x422 ^ x294 ;
  assign n1223 = x256 & ~x384 ;
  assign n1224 = n1223 ^ x385 ;
  assign n1994 = x385 ^ x257 ;
  assign n1228 = n1224 & ~n1994 ;
  assign n1225 = x386 ^ x257 ;
  assign n1229 = n1228 ^ n1225 ;
  assign n1231 = x387 ^ x258 ;
  assign n1230 = x387 ^ x386 ;
  assign n1232 = n1231 ^ n1230 ;
  assign n1233 = n1229 & ~n1232 ;
  assign n1234 = n1233 ^ n1231 ;
  assign n1236 = x388 ^ x259 ;
  assign n1235 = x388 ^ x387 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1238 = n1234 & ~n1237 ;
  assign n1239 = n1238 ^ n1236 ;
  assign n1987 = x388 ^ x260 ;
  assign n1243 = n1239 & ~n1987 ;
  assign n1241 = x389 ^ x260 ;
  assign n1244 = n1243 ^ n1241 ;
  assign n1990 = x389 ^ x261 ;
  assign n1248 = n1244 & ~n1990 ;
  assign n1246 = x390 ^ x261 ;
  assign n1249 = n1248 ^ n1246 ;
  assign n1251 = x391 ^ x262 ;
  assign n1250 = x391 ^ x390 ;
  assign n1252 = n1251 ^ n1250 ;
  assign n1253 = n1249 & ~n1252 ;
  assign n1254 = n1253 ^ n1251 ;
  assign n2056 = x391 ^ x263 ;
  assign n1258 = n1254 & ~n2056 ;
  assign n1256 = x392 ^ x263 ;
  assign n1259 = n1258 ^ n1256 ;
  assign n1261 = x393 ^ x264 ;
  assign n1260 = x393 ^ x392 ;
  assign n1262 = n1261 ^ n1260 ;
  assign n1263 = n1259 & ~n1262 ;
  assign n1264 = n1263 ^ n1261 ;
  assign n1266 = x394 ^ x265 ;
  assign n1265 = x394 ^ x393 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1268 = n1264 & ~n1267 ;
  assign n1269 = n1268 ^ n1266 ;
  assign n1983 = x394 ^ x266 ;
  assign n1273 = n1269 & ~n1983 ;
  assign n1271 = x395 ^ x266 ;
  assign n1274 = n1273 ^ n1271 ;
  assign n1976 = x395 ^ x267 ;
  assign n1278 = n1274 & ~n1976 ;
  assign n1276 = x396 ^ x267 ;
  assign n1279 = n1278 ^ n1276 ;
  assign n1979 = x396 ^ x268 ;
  assign n1283 = n1279 & ~n1979 ;
  assign n1281 = x397 ^ x268 ;
  assign n1284 = n1283 ^ n1281 ;
  assign n1286 = x398 ^ x269 ;
  assign n1285 = x398 ^ x397 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1288 = n1284 & ~n1287 ;
  assign n1289 = n1288 ^ n1286 ;
  assign n1291 = x399 ^ x270 ;
  assign n1290 = x399 ^ x398 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1293 = n1289 & ~n1292 ;
  assign n1294 = n1293 ^ n1291 ;
  assign n2133 = x399 ^ x271 ;
  assign n1298 = n1294 & ~n2133 ;
  assign n1296 = x400 ^ x271 ;
  assign n1299 = n1298 ^ n1296 ;
  assign n1301 = x401 ^ x272 ;
  assign n1300 = x401 ^ x400 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1303 = n1299 & ~n1302 ;
  assign n1304 = n1303 ^ n1301 ;
  assign n1969 = x401 ^ x273 ;
  assign n1308 = n1304 & ~n1969 ;
  assign n1306 = x402 ^ x273 ;
  assign n1309 = n1308 ^ n1306 ;
  assign n1972 = x402 ^ x274 ;
  assign n1313 = n1309 & ~n1972 ;
  assign n1311 = x403 ^ x274 ;
  assign n1314 = n1313 ^ n1311 ;
  assign n1316 = x404 ^ x275 ;
  assign n1315 = x404 ^ x403 ;
  assign n1317 = n1316 ^ n1315 ;
  assign n1318 = n1314 & ~n1317 ;
  assign n1319 = n1318 ^ n1316 ;
  assign n2181 = x404 ^ x276 ;
  assign n1323 = n1319 & ~n2181 ;
  assign n1321 = x405 ^ x276 ;
  assign n1324 = n1323 ^ n1321 ;
  assign n1326 = x406 ^ x277 ;
  assign n1325 = x406 ^ x405 ;
  assign n1327 = n1326 ^ n1325 ;
  assign n1328 = n1324 & ~n1327 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1331 = x407 ^ x278 ;
  assign n1330 = x407 ^ x406 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1333 = n1329 & ~n1332 ;
  assign n1334 = n1333 ^ n1331 ;
  assign n1336 = x408 ^ x279 ;
  assign n1335 = x408 ^ x407 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1338 = n1334 & ~n1337 ;
  assign n1339 = n1338 ^ n1336 ;
  assign n1965 = x408 ^ x280 ;
  assign n1343 = n1339 & ~n1965 ;
  assign n1341 = x409 ^ x280 ;
  assign n1344 = n1343 ^ n1341 ;
  assign n1958 = x409 ^ x281 ;
  assign n1348 = n1344 & ~n1958 ;
  assign n1346 = x410 ^ x281 ;
  assign n1349 = n1348 ^ n1346 ;
  assign n1961 = x410 ^ x282 ;
  assign n1353 = n1349 & ~n1961 ;
  assign n1351 = x411 ^ x282 ;
  assign n1354 = n1353 ^ n1351 ;
  assign n1356 = x412 ^ x283 ;
  assign n1355 = x412 ^ x411 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1358 = n1354 & ~n1357 ;
  assign n1359 = n1358 ^ n1356 ;
  assign n1951 = x412 ^ x284 ;
  assign n1363 = n1359 & ~n1951 ;
  assign n1361 = x413 ^ x284 ;
  assign n1364 = n1363 ^ n1361 ;
  assign n1954 = x413 ^ x285 ;
  assign n1368 = n1364 & ~n1954 ;
  assign n1366 = x414 ^ x285 ;
  assign n1369 = n1368 ^ n1366 ;
  assign n1371 = x415 ^ x286 ;
  assign n1370 = x415 ^ x414 ;
  assign n1372 = n1371 ^ n1370 ;
  assign n1373 = n1369 & ~n1372 ;
  assign n1374 = n1373 ^ n1371 ;
  assign n1947 = x415 ^ x287 ;
  assign n1378 = n1374 & ~n1947 ;
  assign n1376 = x416 ^ x287 ;
  assign n1379 = n1378 ^ n1376 ;
  assign n1940 = x416 ^ x288 ;
  assign n1383 = n1379 & ~n1940 ;
  assign n1381 = x417 ^ x288 ;
  assign n1384 = n1383 ^ n1381 ;
  assign n1943 = x417 ^ x289 ;
  assign n1388 = n1384 & ~n1943 ;
  assign n1386 = x418 ^ x289 ;
  assign n1389 = n1388 ^ n1386 ;
  assign n1391 = x419 ^ x290 ;
  assign n1390 = x419 ^ x418 ;
  assign n1392 = n1391 ^ n1390 ;
  assign n1393 = n1389 & ~n1392 ;
  assign n1394 = n1393 ^ n1391 ;
  assign n1933 = x419 ^ x291 ;
  assign n1398 = n1394 & ~n1933 ;
  assign n1396 = x420 ^ x291 ;
  assign n1399 = n1398 ^ n1396 ;
  assign n1936 = x420 ^ x292 ;
  assign n1403 = n1399 & ~n1936 ;
  assign n1401 = x421 ^ x292 ;
  assign n1404 = n1403 ^ n1401 ;
  assign n1406 = x422 ^ x293 ;
  assign n1405 = x422 ^ x421 ;
  assign n1407 = n1406 ^ n1405 ;
  assign n1408 = n1404 & ~n1407 ;
  assign n1409 = n1408 ^ n1406 ;
  assign n1410 = ~n1218 & n1409 ;
  assign n1411 = n1410 ^ x294 ;
  assign n1412 = ~n1210 & ~n1411 ;
  assign n1413 = n1217 & ~n1412 ;
  assign n1414 = x426 ^ x425 ;
  assign n1415 = n1414 ^ n1213 ;
  assign n1416 = n1415 ^ x297 ;
  assign n1417 = n1416 ^ n1414 ;
  assign n1418 = n1213 ^ x426 ;
  assign n1419 = n1418 ^ n1414 ;
  assign n1420 = ~n1417 & ~n1419 ;
  assign n1421 = n1420 ^ n1414 ;
  assign n1422 = ~n1208 & ~n1421 ;
  assign n1423 = n1422 ^ x298 ;
  assign n1424 = ~n1413 & ~n1423 ;
  assign n1425 = n1424 ^ x427 ;
  assign n1426 = ~n1206 & ~n1425 ;
  assign n1427 = n1426 ^ x299 ;
  assign n1428 = ~n1205 & n1427 ;
  assign n1429 = x302 ^ x301 ;
  assign n1430 = n1429 ^ x430 ;
  assign n1431 = n1430 ^ n1204 ;
  assign n1432 = n1431 ^ x429 ;
  assign n1433 = ~n1428 & ~n1432 ;
  assign n1434 = n1433 ^ n1430 ;
  assign n1915 = x429 ^ x301 ;
  assign n1438 = ~n1434 & ~n1915 ;
  assign n1436 = x430 ^ x301 ;
  assign n1439 = n1438 ^ n1436 ;
  assign n1908 = x430 ^ x302 ;
  assign n1443 = n1439 & ~n1908 ;
  assign n1441 = x431 ^ x302 ;
  assign n1444 = n1443 ^ n1441 ;
  assign n1911 = x431 ^ x303 ;
  assign n1448 = n1444 & ~n1911 ;
  assign n1446 = x432 ^ x303 ;
  assign n1449 = n1448 ^ n1446 ;
  assign n1451 = x433 ^ x304 ;
  assign n1450 = x433 ^ x432 ;
  assign n1452 = n1451 ^ n1450 ;
  assign n1453 = n1449 & ~n1452 ;
  assign n1454 = n1453 ^ n1451 ;
  assign n2432 = x433 ^ x305 ;
  assign n1458 = n1454 & ~n2432 ;
  assign n1456 = x434 ^ x305 ;
  assign n1459 = n1458 ^ n1456 ;
  assign n1461 = x435 ^ x306 ;
  assign n1460 = x435 ^ x434 ;
  assign n1462 = n1461 ^ n1460 ;
  assign n1463 = n1459 & ~n1462 ;
  assign n1464 = n1463 ^ n1461 ;
  assign n1466 = x436 ^ x307 ;
  assign n1465 = x436 ^ x435 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1468 = n1464 & ~n1467 ;
  assign n1469 = n1468 ^ n1466 ;
  assign n2465 = x436 ^ x308 ;
  assign n1473 = n1469 & ~n2465 ;
  assign n1471 = x437 ^ x308 ;
  assign n1474 = n1473 ^ n1471 ;
  assign n1476 = x438 ^ x309 ;
  assign n1475 = x438 ^ x437 ;
  assign n1477 = n1476 ^ n1475 ;
  assign n1478 = n1474 & ~n1477 ;
  assign n1479 = n1478 ^ n1476 ;
  assign n2487 = x438 ^ x310 ;
  assign n1483 = n1479 & ~n2487 ;
  assign n1481 = x439 ^ x310 ;
  assign n1484 = n1483 ^ n1481 ;
  assign n1486 = x440 ^ x311 ;
  assign n1485 = x440 ^ x439 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1488 = n1484 & ~n1487 ;
  assign n1489 = n1488 ^ n1486 ;
  assign n2509 = x440 ^ x312 ;
  assign n1493 = n1489 & ~n2509 ;
  assign n1491 = x441 ^ x312 ;
  assign n1494 = n1493 ^ n1491 ;
  assign n1496 = x442 ^ x313 ;
  assign n1495 = x442 ^ x441 ;
  assign n1497 = n1496 ^ n1495 ;
  assign n1498 = n1494 & ~n1497 ;
  assign n1499 = n1498 ^ n1496 ;
  assign n1501 = x443 ^ x314 ;
  assign n1500 = x443 ^ x442 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1503 = n1499 & ~n1502 ;
  assign n1504 = n1503 ^ n1501 ;
  assign n1505 = ~n1202 & n1504 ;
  assign n1506 = n1505 ^ x315 ;
  assign n1507 = n1201 & n1506 ;
  assign n1508 = ~n1191 & n1507 ;
  assign n1509 = x447 ^ x319 ;
  assign n1510 = n1196 ^ x447 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = n1511 ^ x447 ;
  assign n1513 = ~n1186 & n1512 ;
  assign n1514 = n1201 & n1513 ;
  assign n1521 = ~n1189 & ~n1193 ;
  assign n1522 = n1514 & n1521 ;
  assign n1523 = n1522 ^ n1514 ;
  assign n1524 = n1523 ^ n1513 ;
  assign n1525 = ~n1508 & n1524 ;
  assign n1526 = ~n1188 & ~n1525 ;
  assign n1184 = x450 ^ x449 ;
  assign n1185 = n1184 ^ x321 ;
  assign n1527 = n1526 ^ n1185 ;
  assign n1528 = n1527 ^ n1184 ;
  assign n1895 = x449 ^ x321 ;
  assign n1531 = ~n1528 & ~n1895 ;
  assign n1532 = n1531 ^ n1184 ;
  assign n1533 = ~n1183 & ~n1532 ;
  assign n1534 = n1533 ^ x322 ;
  assign n1535 = ~n1175 & ~n1534 ;
  assign n1536 = n1182 & ~n1535 ;
  assign n1537 = x454 ^ x453 ;
  assign n1538 = n1537 ^ n1179 ;
  assign n1539 = n1538 ^ x325 ;
  assign n1540 = n1539 ^ n1537 ;
  assign n1541 = n1179 ^ x454 ;
  assign n1542 = n1541 ^ n1537 ;
  assign n1543 = ~n1540 & ~n1542 ;
  assign n1544 = n1543 ^ n1537 ;
  assign n1545 = ~n1172 & ~n1544 ;
  assign n1546 = n1545 ^ x326 ;
  assign n1547 = ~n1536 & ~n1546 ;
  assign n1548 = n1547 ^ x327 ;
  assign n1549 = ~n1169 & ~n1548 ;
  assign n1170 = x456 ^ x327 ;
  assign n1550 = n1549 ^ n1170 ;
  assign n1880 = x456 ^ x328 ;
  assign n1554 = n1550 & ~n1880 ;
  assign n1552 = x457 ^ x328 ;
  assign n1555 = n1554 ^ n1552 ;
  assign n1557 = x458 ^ x329 ;
  assign n1556 = x458 ^ x457 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1559 = n1555 & ~n1558 ;
  assign n1560 = n1559 ^ n1557 ;
  assign n1562 = x459 ^ x330 ;
  assign n1561 = x459 ^ x458 ;
  assign n1563 = n1562 ^ n1561 ;
  assign n1564 = n1560 & ~n1563 ;
  assign n1565 = n1564 ^ n1562 ;
  assign n2673 = x459 ^ x331 ;
  assign n1569 = n1565 & ~n2673 ;
  assign n1567 = x460 ^ x331 ;
  assign n1570 = n1569 ^ n1567 ;
  assign n1572 = x461 ^ x332 ;
  assign n1571 = x461 ^ x460 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1574 = n1570 & ~n1573 ;
  assign n1575 = n1574 ^ n1572 ;
  assign n1577 = x462 ^ x333 ;
  assign n1576 = x462 ^ x461 ;
  assign n1578 = n1577 ^ n1576 ;
  assign n1579 = n1575 & ~n1578 ;
  assign n1580 = n1579 ^ n1577 ;
  assign n1582 = x463 ^ x334 ;
  assign n1581 = x463 ^ x462 ;
  assign n1583 = n1582 ^ n1581 ;
  assign n1584 = n1580 & ~n1583 ;
  assign n1585 = n1584 ^ n1582 ;
  assign n1587 = x464 ^ x335 ;
  assign n1586 = x464 ^ x463 ;
  assign n1588 = n1587 ^ n1586 ;
  assign n1589 = n1585 & ~n1588 ;
  assign n1590 = n1589 ^ n1587 ;
  assign n1871 = x464 ^ x336 ;
  assign n1594 = n1590 & ~n1871 ;
  assign n1592 = x465 ^ x336 ;
  assign n1595 = n1594 ^ n1592 ;
  assign n1874 = x465 ^ x337 ;
  assign n1599 = n1595 & ~n1874 ;
  assign n1597 = x466 ^ x337 ;
  assign n1600 = n1599 ^ n1597 ;
  assign n2743 = x466 ^ x338 ;
  assign n1604 = n1600 & ~n2743 ;
  assign n1602 = x467 ^ x338 ;
  assign n1605 = n1604 ^ n1602 ;
  assign n1607 = x468 ^ x339 ;
  assign n1606 = x468 ^ x467 ;
  assign n1608 = n1607 ^ n1606 ;
  assign n1609 = n1605 & ~n1608 ;
  assign n1610 = n1609 ^ n1607 ;
  assign n1612 = x469 ^ x340 ;
  assign n1611 = x469 ^ x468 ;
  assign n1613 = n1612 ^ n1611 ;
  assign n1614 = n1610 & ~n1613 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1617 = x470 ^ x341 ;
  assign n1616 = x470 ^ x469 ;
  assign n1618 = n1617 ^ n1616 ;
  assign n1619 = n1615 & ~n1618 ;
  assign n1620 = n1619 ^ n1617 ;
  assign n1622 = x471 ^ x342 ;
  assign n1621 = x471 ^ x470 ;
  assign n1623 = n1622 ^ n1621 ;
  assign n1624 = n1620 & ~n1623 ;
  assign n1625 = n1624 ^ n1622 ;
  assign n1627 = x472 ^ x343 ;
  assign n1626 = x472 ^ x471 ;
  assign n1628 = n1627 ^ n1626 ;
  assign n1629 = n1625 & ~n1628 ;
  assign n1630 = n1629 ^ n1627 ;
  assign n2809 = x472 ^ x344 ;
  assign n1634 = n1630 & ~n2809 ;
  assign n1632 = x473 ^ x344 ;
  assign n1635 = n1634 ^ n1632 ;
  assign n2820 = x473 ^ x345 ;
  assign n1639 = n1635 & ~n2820 ;
  assign n1637 = x474 ^ x345 ;
  assign n1640 = n1639 ^ n1637 ;
  assign n2831 = x474 ^ x346 ;
  assign n1644 = n1640 & ~n2831 ;
  assign n1642 = x475 ^ x346 ;
  assign n1645 = n1644 ^ n1642 ;
  assign n1647 = x476 ^ x347 ;
  assign n1646 = x476 ^ x475 ;
  assign n1648 = n1647 ^ n1646 ;
  assign n1649 = n1645 & ~n1648 ;
  assign n1650 = n1649 ^ n1647 ;
  assign n1652 = x477 ^ x348 ;
  assign n1651 = x477 ^ x476 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n1654 = n1650 & ~n1653 ;
  assign n1655 = n1654 ^ n1652 ;
  assign n1657 = x478 ^ x349 ;
  assign n1656 = x478 ^ x477 ;
  assign n1658 = n1657 ^ n1656 ;
  assign n1659 = n1655 & ~n1658 ;
  assign n1660 = n1659 ^ n1657 ;
  assign n2875 = x478 ^ x350 ;
  assign n1664 = n1660 & ~n2875 ;
  assign n1662 = x479 ^ x350 ;
  assign n1665 = n1664 ^ n1662 ;
  assign n2886 = x479 ^ x351 ;
  assign n1669 = n1665 & ~n2886 ;
  assign n1667 = x480 ^ x351 ;
  assign n1670 = n1669 ^ n1667 ;
  assign n1864 = x480 ^ x352 ;
  assign n1674 = n1670 & ~n1864 ;
  assign n1672 = x481 ^ x352 ;
  assign n1675 = n1674 ^ n1672 ;
  assign n1867 = x481 ^ x353 ;
  assign n1679 = n1675 & ~n1867 ;
  assign n1677 = x482 ^ x353 ;
  assign n1680 = n1679 ^ n1677 ;
  assign n2912 = x482 ^ x354 ;
  assign n1684 = n1680 & ~n2912 ;
  assign n1682 = x483 ^ x354 ;
  assign n1685 = n1684 ^ n1682 ;
  assign n2923 = x483 ^ x355 ;
  assign n1689 = n1685 & ~n2923 ;
  assign n1687 = x484 ^ x355 ;
  assign n1690 = n1689 ^ n1687 ;
  assign n1857 = x484 ^ x356 ;
  assign n1694 = n1690 & ~n1857 ;
  assign n1692 = x485 ^ x356 ;
  assign n1695 = n1694 ^ n1692 ;
  assign n1860 = x485 ^ x357 ;
  assign n1699 = n1695 & ~n1860 ;
  assign n1697 = x486 ^ x357 ;
  assign n1700 = n1699 ^ n1697 ;
  assign n2949 = x486 ^ x358 ;
  assign n1704 = n1700 & ~n2949 ;
  assign n1702 = x487 ^ x358 ;
  assign n1705 = n1704 ^ n1702 ;
  assign n1707 = x488 ^ x359 ;
  assign n1706 = x488 ^ x487 ;
  assign n1708 = n1707 ^ n1706 ;
  assign n1709 = n1705 & ~n1708 ;
  assign n1710 = n1709 ^ n1707 ;
  assign n2971 = x488 ^ x360 ;
  assign n1714 = n1710 & ~n2971 ;
  assign n1712 = x489 ^ x360 ;
  assign n1715 = n1714 ^ n1712 ;
  assign n2982 = x489 ^ x361 ;
  assign n1719 = n1715 & ~n2982 ;
  assign n1717 = x490 ^ x361 ;
  assign n1720 = n1719 ^ n1717 ;
  assign n1722 = x491 ^ x362 ;
  assign n1721 = x491 ^ x490 ;
  assign n1723 = n1722 ^ n1721 ;
  assign n1724 = n1720 & ~n1723 ;
  assign n1725 = n1724 ^ n1722 ;
  assign n1727 = x492 ^ x363 ;
  assign n1726 = x492 ^ x491 ;
  assign n1728 = n1727 ^ n1726 ;
  assign n1729 = n1725 & ~n1728 ;
  assign n1730 = n1729 ^ n1727 ;
  assign n1853 = x492 ^ x364 ;
  assign n1734 = n1730 & ~n1853 ;
  assign n1732 = x493 ^ x364 ;
  assign n1735 = n1734 ^ n1732 ;
  assign n1846 = x493 ^ x365 ;
  assign n1739 = n1735 & ~n1846 ;
  assign n1737 = x494 ^ x365 ;
  assign n1740 = n1739 ^ n1737 ;
  assign n1849 = x494 ^ x366 ;
  assign n1744 = n1740 & ~n1849 ;
  assign n1742 = x495 ^ x366 ;
  assign n1745 = n1744 ^ n1742 ;
  assign n3037 = x495 ^ x367 ;
  assign n1749 = n1745 & ~n3037 ;
  assign n1747 = x496 ^ x367 ;
  assign n1750 = n1749 ^ n1747 ;
  assign n3048 = x496 ^ x368 ;
  assign n1754 = n1750 & ~n3048 ;
  assign n1752 = x497 ^ x368 ;
  assign n1755 = n1754 ^ n1752 ;
  assign n1757 = x498 ^ x369 ;
  assign n1756 = x498 ^ x497 ;
  assign n1758 = n1757 ^ n1756 ;
  assign n1759 = n1755 & ~n1758 ;
  assign n1760 = n1759 ^ n1757 ;
  assign n3070 = x498 ^ x370 ;
  assign n1764 = n1760 & ~n3070 ;
  assign n1762 = x499 ^ x370 ;
  assign n1765 = n1764 ^ n1762 ;
  assign n3081 = x499 ^ x371 ;
  assign n1769 = n1765 & ~n3081 ;
  assign n1767 = x500 ^ x371 ;
  assign n1770 = n1769 ^ n1767 ;
  assign n1772 = x501 ^ x372 ;
  assign n1771 = x501 ^ x500 ;
  assign n1773 = n1772 ^ n1771 ;
  assign n1774 = n1770 & ~n1773 ;
  assign n1775 = n1774 ^ n1772 ;
  assign n1777 = x502 ^ x373 ;
  assign n1776 = x502 ^ x501 ;
  assign n1778 = n1777 ^ n1776 ;
  assign n1779 = n1775 & ~n1778 ;
  assign n1780 = n1779 ^ n1777 ;
  assign n1782 = x503 ^ x374 ;
  assign n1781 = x503 ^ x502 ;
  assign n1783 = n1782 ^ n1781 ;
  assign n1784 = n1780 & ~n1783 ;
  assign n1785 = n1784 ^ n1782 ;
  assign n1787 = x504 ^ x375 ;
  assign n1786 = x504 ^ x503 ;
  assign n1788 = n1787 ^ n1786 ;
  assign n1789 = n1785 & ~n1788 ;
  assign n1790 = n1789 ^ n1787 ;
  assign n1839 = x504 ^ x376 ;
  assign n1794 = n1790 & ~n1839 ;
  assign n1792 = x505 ^ x376 ;
  assign n1795 = n1794 ^ n1792 ;
  assign n1842 = x505 ^ x377 ;
  assign n1799 = n1795 & ~n1842 ;
  assign n1797 = x506 ^ x377 ;
  assign n1800 = n1799 ^ n1797 ;
  assign n1802 = x507 ^ x378 ;
  assign n1801 = x507 ^ x506 ;
  assign n1803 = n1802 ^ n1801 ;
  assign n1804 = n1800 & ~n1803 ;
  assign n1805 = n1804 ^ n1802 ;
  assign n1806 = ~n1168 & n1805 ;
  assign n1807 = n1806 ^ x379 ;
  assign n1808 = ~n1167 & n1807 ;
  assign n1809 = ~n1166 & n1808 ;
  assign n1810 = x508 ^ x380 ;
  assign n1811 = n1810 ^ x509 ;
  assign n1812 = n1811 ^ n1166 ;
  assign n1818 = ~n1167 & n1812 ;
  assign n1815 = x382 ^ x381 ;
  assign n1816 = n1815 ^ x510 ;
  assign n1819 = n1818 ^ n1816 ;
  assign n1820 = ~n1809 & ~n1819 ;
  assign n1821 = n1820 ^ x511 ;
  assign n1823 = n1822 ^ n1821 ;
  assign n1824 = x511 ^ x510 ;
  assign n1825 = n1824 ^ n1822 ;
  assign n1826 = ~n1823 & ~n1825 ;
  assign n1827 = n1826 ^ n1822 ;
  assign n1828 = ~n1165 & ~n1827 ;
  assign n1829 = n1828 ^ x383 ;
  assign n1830 = n1164 & n1829 ;
  assign n1831 = n1830 ^ x256 ;
  assign n513 = x128 ^ x0 ;
  assign n514 = x255 ^ x127 ;
  assign n515 = x123 & ~x251 ;
  assign n516 = x250 ^ x122 ;
  assign n869 = x197 ^ x68 ;
  assign n517 = x196 ^ x68 ;
  assign n518 = x191 ^ x63 ;
  assign n521 = x190 ^ x62 ;
  assign n522 = x189 ^ x61 ;
  assign n523 = ~n521 & ~n522 ;
  assign n525 = x187 ^ x59 ;
  assign n524 = x59 & ~x187 ;
  assign n526 = n525 ^ n524 ;
  assign n528 = x60 & ~x188 ;
  assign n527 = x188 ^ x60 ;
  assign n529 = n528 ^ n527 ;
  assign n530 = ~n526 & ~n529 ;
  assign n531 = n523 & n530 ;
  assign n532 = x186 ^ x58 ;
  assign n534 = x44 & ~x172 ;
  assign n533 = x172 ^ x44 ;
  assign n535 = n534 ^ n533 ;
  assign n536 = x171 ^ x43 ;
  assign n538 = x168 ^ x40 ;
  assign n537 = x40 & ~x168 ;
  assign n539 = n538 ^ n537 ;
  assign n540 = x167 ^ x39 ;
  assign n545 = x0 & ~x128 ;
  assign n546 = n545 ^ x129 ;
  assign n1997 = x129 ^ x1 ;
  assign n550 = n546 & ~n1997 ;
  assign n547 = x130 ^ x1 ;
  assign n551 = n550 ^ n547 ;
  assign n2008 = x130 ^ x2 ;
  assign n555 = n551 & ~n2008 ;
  assign n553 = x131 ^ x2 ;
  assign n556 = n555 ^ n553 ;
  assign n2019 = x131 ^ x3 ;
  assign n560 = n556 & ~n2019 ;
  assign n558 = x132 ^ x3 ;
  assign n561 = n560 ^ n558 ;
  assign n563 = x133 ^ x4 ;
  assign n562 = x133 ^ x132 ;
  assign n564 = n563 ^ n562 ;
  assign n565 = n561 & ~n564 ;
  assign n566 = n565 ^ n563 ;
  assign n568 = x134 ^ x5 ;
  assign n567 = x134 ^ x133 ;
  assign n569 = n568 ^ n567 ;
  assign n570 = n566 & ~n569 ;
  assign n571 = n570 ^ n568 ;
  assign n2045 = x134 ^ x6 ;
  assign n575 = n571 & ~n2045 ;
  assign n573 = x135 ^ x6 ;
  assign n576 = n575 ^ n573 ;
  assign n578 = x136 ^ x7 ;
  assign n577 = x136 ^ x135 ;
  assign n579 = n578 ^ n577 ;
  assign n580 = n576 & ~n579 ;
  assign n581 = n580 ^ n578 ;
  assign n2067 = x136 ^ x8 ;
  assign n585 = n581 & ~n2067 ;
  assign n583 = x137 ^ x8 ;
  assign n586 = n585 ^ n583 ;
  assign n2078 = x137 ^ x9 ;
  assign n590 = n586 & ~n2078 ;
  assign n588 = x138 ^ x9 ;
  assign n591 = n590 ^ n588 ;
  assign n593 = x139 ^ x10 ;
  assign n592 = x139 ^ x138 ;
  assign n594 = n593 ^ n592 ;
  assign n595 = n591 & ~n594 ;
  assign n596 = n595 ^ n593 ;
  assign n598 = x140 ^ x11 ;
  assign n597 = x140 ^ x139 ;
  assign n599 = n598 ^ n597 ;
  assign n600 = n596 & ~n599 ;
  assign n601 = n600 ^ n598 ;
  assign n603 = x141 ^ x12 ;
  assign n602 = x141 ^ x140 ;
  assign n604 = n603 ^ n602 ;
  assign n605 = n601 & ~n604 ;
  assign n606 = n605 ^ n603 ;
  assign n2111 = x141 ^ x13 ;
  assign n610 = n606 & ~n2111 ;
  assign n608 = x142 ^ x13 ;
  assign n611 = n610 ^ n608 ;
  assign n2122 = x142 ^ x14 ;
  assign n615 = n611 & ~n2122 ;
  assign n613 = x143 ^ x14 ;
  assign n616 = n615 ^ n613 ;
  assign n618 = x144 ^ x15 ;
  assign n617 = x144 ^ x143 ;
  assign n619 = n618 ^ n617 ;
  assign n620 = n616 & ~n619 ;
  assign n621 = n620 ^ n618 ;
  assign n2144 = x144 ^ x16 ;
  assign n625 = n621 & ~n2144 ;
  assign n623 = x145 ^ x16 ;
  assign n626 = n625 ^ n623 ;
  assign n628 = x146 ^ x17 ;
  assign n627 = x146 ^ x145 ;
  assign n629 = n628 ^ n627 ;
  assign n630 = n626 & ~n629 ;
  assign n631 = n630 ^ n628 ;
  assign n633 = x147 ^ x18 ;
  assign n632 = x147 ^ x146 ;
  assign n634 = n633 ^ n632 ;
  assign n635 = n631 & ~n634 ;
  assign n636 = n635 ^ n633 ;
  assign n2170 = x147 ^ x19 ;
  assign n640 = n636 & ~n2170 ;
  assign n638 = x148 ^ x19 ;
  assign n641 = n640 ^ n638 ;
  assign n643 = x149 ^ x20 ;
  assign n642 = x149 ^ x148 ;
  assign n644 = n643 ^ n642 ;
  assign n645 = n641 & ~n644 ;
  assign n646 = n645 ^ n643 ;
  assign n2192 = x149 ^ x21 ;
  assign n650 = n646 & ~n2192 ;
  assign n648 = x150 ^ x21 ;
  assign n651 = n650 ^ n648 ;
  assign n2203 = x150 ^ x22 ;
  assign n655 = n651 & ~n2203 ;
  assign n653 = x151 ^ x22 ;
  assign n656 = n655 ^ n653 ;
  assign n2214 = x151 ^ x23 ;
  assign n660 = n656 & ~n2214 ;
  assign n658 = x152 ^ x23 ;
  assign n661 = n660 ^ n658 ;
  assign n663 = x153 ^ x24 ;
  assign n662 = x153 ^ x152 ;
  assign n664 = n663 ^ n662 ;
  assign n665 = n661 & ~n664 ;
  assign n666 = n665 ^ n663 ;
  assign n668 = x154 ^ x25 ;
  assign n667 = x154 ^ x153 ;
  assign n669 = n668 ^ n667 ;
  assign n670 = n666 & ~n669 ;
  assign n671 = n670 ^ n668 ;
  assign n673 = x155 ^ x26 ;
  assign n672 = x155 ^ x154 ;
  assign n674 = n673 ^ n672 ;
  assign n675 = n671 & ~n674 ;
  assign n676 = n675 ^ n673 ;
  assign n2247 = x155 ^ x27 ;
  assign n680 = n676 & ~n2247 ;
  assign n678 = x156 ^ x27 ;
  assign n681 = n680 ^ n678 ;
  assign n683 = x157 ^ x28 ;
  assign n682 = x157 ^ x156 ;
  assign n684 = n683 ^ n682 ;
  assign n685 = n681 & ~n684 ;
  assign n686 = n685 ^ n683 ;
  assign n688 = x158 ^ x29 ;
  assign n687 = x158 ^ x157 ;
  assign n689 = n688 ^ n687 ;
  assign n690 = n686 & ~n689 ;
  assign n691 = n690 ^ n688 ;
  assign n2273 = x158 ^ x30 ;
  assign n695 = n691 & ~n2273 ;
  assign n693 = x159 ^ x30 ;
  assign n696 = n695 ^ n693 ;
  assign n698 = x160 ^ x31 ;
  assign n697 = x160 ^ x159 ;
  assign n699 = n698 ^ n697 ;
  assign n700 = n696 & ~n699 ;
  assign n701 = n700 ^ n698 ;
  assign n703 = x161 ^ x32 ;
  assign n702 = x161 ^ x160 ;
  assign n704 = n703 ^ n702 ;
  assign n705 = n701 & ~n704 ;
  assign n706 = n705 ^ n703 ;
  assign n708 = x162 ^ x33 ;
  assign n707 = x162 ^ x161 ;
  assign n709 = n708 ^ n707 ;
  assign n710 = n706 & ~n709 ;
  assign n711 = n710 ^ n708 ;
  assign n2306 = x162 ^ x34 ;
  assign n715 = n711 & ~n2306 ;
  assign n713 = x163 ^ x34 ;
  assign n716 = n715 ^ n713 ;
  assign n718 = x164 ^ x35 ;
  assign n717 = x164 ^ x163 ;
  assign n719 = n718 ^ n717 ;
  assign n720 = n716 & ~n719 ;
  assign n721 = n720 ^ n718 ;
  assign n723 = x165 ^ x36 ;
  assign n722 = x165 ^ x164 ;
  assign n724 = n723 ^ n722 ;
  assign n725 = n721 & ~n724 ;
  assign n726 = n725 ^ n723 ;
  assign n2332 = x165 ^ x37 ;
  assign n730 = n726 & ~n2332 ;
  assign n728 = x166 ^ x37 ;
  assign n731 = n730 ^ n728 ;
  assign n733 = x167 ^ x38 ;
  assign n732 = x167 ^ x166 ;
  assign n734 = n733 ^ n732 ;
  assign n735 = n731 & ~n734 ;
  assign n736 = n735 ^ n733 ;
  assign n737 = ~n540 & n736 ;
  assign n738 = n737 ^ x39 ;
  assign n739 = ~n539 & n738 ;
  assign n741 = x42 ^ x41 ;
  assign n742 = n741 ^ x170 ;
  assign n740 = n537 ^ x169 ;
  assign n743 = n742 ^ n740 ;
  assign n744 = ~n739 & ~n743 ;
  assign n745 = n744 ^ n742 ;
  assign n747 = x170 ^ x41 ;
  assign n746 = x170 ^ x169 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = ~n745 & ~n748 ;
  assign n750 = n749 ^ n747 ;
  assign n752 = x171 ^ x42 ;
  assign n751 = x171 ^ x170 ;
  assign n753 = n752 ^ n751 ;
  assign n754 = n750 & ~n753 ;
  assign n755 = n754 ^ n752 ;
  assign n756 = ~n536 & n755 ;
  assign n757 = n756 ^ x43 ;
  assign n758 = ~n535 & n757 ;
  assign n759 = x46 ^ x45 ;
  assign n760 = n759 ^ x174 ;
  assign n761 = n760 ^ n534 ;
  assign n762 = n761 ^ x173 ;
  assign n763 = ~n758 & ~n762 ;
  assign n764 = n763 ^ n760 ;
  assign n766 = x174 ^ x45 ;
  assign n765 = x174 ^ x173 ;
  assign n767 = n766 ^ n765 ;
  assign n768 = ~n764 & ~n767 ;
  assign n769 = n768 ^ n766 ;
  assign n771 = x175 ^ x46 ;
  assign n770 = x175 ^ x174 ;
  assign n772 = n771 ^ n770 ;
  assign n773 = n769 & ~n772 ;
  assign n774 = n773 ^ n771 ;
  assign n776 = x176 ^ x47 ;
  assign n775 = x176 ^ x175 ;
  assign n777 = n776 ^ n775 ;
  assign n778 = n774 & ~n777 ;
  assign n779 = n778 ^ n776 ;
  assign n2421 = x176 ^ x48 ;
  assign n783 = n779 & ~n2421 ;
  assign n781 = x177 ^ x48 ;
  assign n784 = n783 ^ n781 ;
  assign n786 = x178 ^ x49 ;
  assign n785 = x178 ^ x177 ;
  assign n787 = n786 ^ n785 ;
  assign n788 = n784 & ~n787 ;
  assign n789 = n788 ^ n786 ;
  assign n2443 = x178 ^ x50 ;
  assign n793 = n789 & ~n2443 ;
  assign n791 = x179 ^ x50 ;
  assign n794 = n793 ^ n791 ;
  assign n2454 = x179 ^ x51 ;
  assign n798 = n794 & ~n2454 ;
  assign n796 = x180 ^ x51 ;
  assign n799 = n798 ^ n796 ;
  assign n801 = x181 ^ x52 ;
  assign n800 = x181 ^ x180 ;
  assign n802 = n801 ^ n800 ;
  assign n803 = n799 & ~n802 ;
  assign n804 = n803 ^ n801 ;
  assign n2476 = x181 ^ x53 ;
  assign n808 = n804 & ~n2476 ;
  assign n806 = x182 ^ x53 ;
  assign n809 = n808 ^ n806 ;
  assign n811 = x183 ^ x54 ;
  assign n810 = x183 ^ x182 ;
  assign n812 = n811 ^ n810 ;
  assign n813 = n809 & ~n812 ;
  assign n814 = n813 ^ n811 ;
  assign n2498 = x183 ^ x55 ;
  assign n818 = n814 & ~n2498 ;
  assign n816 = x184 ^ x55 ;
  assign n819 = n818 ^ n816 ;
  assign n821 = x185 ^ x56 ;
  assign n820 = x185 ^ x184 ;
  assign n822 = n821 ^ n820 ;
  assign n823 = n819 & ~n822 ;
  assign n824 = n823 ^ n821 ;
  assign n2520 = x185 ^ x57 ;
  assign n828 = n824 & ~n2520 ;
  assign n826 = x186 ^ x57 ;
  assign n829 = n828 ^ n826 ;
  assign n830 = ~n532 & n829 ;
  assign n831 = n830 ^ x58 ;
  assign n832 = ~n524 & ~n831 ;
  assign n833 = n531 & ~n832 ;
  assign n834 = x190 ^ x189 ;
  assign n835 = n834 ^ n528 ;
  assign n836 = n835 ^ x61 ;
  assign n837 = n836 ^ n834 ;
  assign n838 = n528 ^ x190 ;
  assign n839 = n838 ^ n834 ;
  assign n840 = ~n837 & ~n839 ;
  assign n841 = n840 ^ n834 ;
  assign n842 = ~n521 & ~n841 ;
  assign n843 = n842 ^ x62 ;
  assign n844 = ~n833 & ~n843 ;
  assign n845 = n844 ^ x63 ;
  assign n846 = ~n518 & ~n845 ;
  assign n519 = x192 ^ x63 ;
  assign n847 = n846 ^ n519 ;
  assign n849 = x193 ^ x64 ;
  assign n848 = x193 ^ x192 ;
  assign n850 = n849 ^ n848 ;
  assign n851 = n847 & ~n850 ;
  assign n852 = n851 ^ n849 ;
  assign n854 = x194 ^ x65 ;
  assign n853 = x194 ^ x193 ;
  assign n855 = n854 ^ n853 ;
  assign n856 = n852 & ~n855 ;
  assign n857 = n856 ^ n854 ;
  assign n859 = x195 ^ x66 ;
  assign n858 = x195 ^ x194 ;
  assign n860 = n859 ^ n858 ;
  assign n861 = n857 & ~n860 ;
  assign n862 = n861 ^ n859 ;
  assign n864 = x68 ^ x67 ;
  assign n863 = x195 ^ x68 ;
  assign n865 = n864 ^ n863 ;
  assign n866 = n862 & ~n865 ;
  assign n867 = n866 ^ n864 ;
  assign n868 = ~n517 & n867 ;
  assign n870 = n869 ^ n868 ;
  assign n872 = x198 ^ x69 ;
  assign n871 = x198 ^ x197 ;
  assign n873 = n872 ^ n871 ;
  assign n874 = n870 & ~n873 ;
  assign n875 = n874 ^ n872 ;
  assign n877 = x199 ^ x70 ;
  assign n876 = x199 ^ x198 ;
  assign n878 = n877 ^ n876 ;
  assign n879 = n875 & ~n878 ;
  assign n880 = n879 ^ n877 ;
  assign n882 = x200 ^ x71 ;
  assign n881 = x200 ^ x199 ;
  assign n883 = n882 ^ n881 ;
  assign n884 = n880 & ~n883 ;
  assign n885 = n884 ^ n882 ;
  assign n887 = x201 ^ x72 ;
  assign n886 = x201 ^ x200 ;
  assign n888 = n887 ^ n886 ;
  assign n889 = n885 & ~n888 ;
  assign n890 = n889 ^ n887 ;
  assign n2651 = x201 ^ x73 ;
  assign n894 = n890 & ~n2651 ;
  assign n892 = x202 ^ x73 ;
  assign n895 = n894 ^ n892 ;
  assign n2662 = x202 ^ x74 ;
  assign n899 = n895 & ~n2662 ;
  assign n897 = x203 ^ x74 ;
  assign n900 = n899 ^ n897 ;
  assign n902 = x204 ^ x75 ;
  assign n901 = x204 ^ x203 ;
  assign n903 = n902 ^ n901 ;
  assign n904 = n900 & ~n903 ;
  assign n905 = n904 ^ n902 ;
  assign n2684 = x204 ^ x76 ;
  assign n909 = n905 & ~n2684 ;
  assign n907 = x205 ^ x76 ;
  assign n910 = n909 ^ n907 ;
  assign n2695 = x205 ^ x77 ;
  assign n914 = n910 & ~n2695 ;
  assign n912 = x206 ^ x77 ;
  assign n915 = n914 ^ n912 ;
  assign n2706 = x206 ^ x78 ;
  assign n919 = n915 & ~n2706 ;
  assign n917 = x207 ^ x78 ;
  assign n920 = n919 ^ n917 ;
  assign n2717 = x207 ^ x79 ;
  assign n924 = n920 & ~n2717 ;
  assign n922 = x208 ^ x79 ;
  assign n925 = n924 ^ n922 ;
  assign n927 = x209 ^ x80 ;
  assign n926 = x209 ^ x208 ;
  assign n928 = n927 ^ n926 ;
  assign n929 = n925 & ~n928 ;
  assign n930 = n929 ^ n927 ;
  assign n932 = x210 ^ x81 ;
  assign n931 = x210 ^ x209 ;
  assign n933 = n932 ^ n931 ;
  assign n934 = n930 & ~n933 ;
  assign n935 = n934 ^ n932 ;
  assign n937 = x211 ^ x82 ;
  assign n936 = x211 ^ x210 ;
  assign n938 = n937 ^ n936 ;
  assign n939 = n935 & ~n938 ;
  assign n940 = n939 ^ n937 ;
  assign n2754 = x211 ^ x83 ;
  assign n944 = n940 & ~n2754 ;
  assign n942 = x212 ^ x83 ;
  assign n945 = n944 ^ n942 ;
  assign n2765 = x212 ^ x84 ;
  assign n949 = n945 & ~n2765 ;
  assign n947 = x213 ^ x84 ;
  assign n950 = n949 ^ n947 ;
  assign n2776 = x213 ^ x85 ;
  assign n954 = n950 & ~n2776 ;
  assign n952 = x214 ^ x85 ;
  assign n955 = n954 ^ n952 ;
  assign n2787 = x214 ^ x86 ;
  assign n959 = n955 & ~n2787 ;
  assign n957 = x215 ^ x86 ;
  assign n960 = n959 ^ n957 ;
  assign n2798 = x215 ^ x87 ;
  assign n964 = n960 & ~n2798 ;
  assign n962 = x216 ^ x87 ;
  assign n965 = n964 ^ n962 ;
  assign n967 = x217 ^ x88 ;
  assign n966 = x217 ^ x216 ;
  assign n968 = n967 ^ n966 ;
  assign n969 = n965 & ~n968 ;
  assign n970 = n969 ^ n967 ;
  assign n972 = x218 ^ x89 ;
  assign n971 = x218 ^ x217 ;
  assign n973 = n972 ^ n971 ;
  assign n974 = n970 & ~n973 ;
  assign n975 = n974 ^ n972 ;
  assign n977 = x219 ^ x90 ;
  assign n976 = x219 ^ x218 ;
  assign n978 = n977 ^ n976 ;
  assign n979 = n975 & ~n978 ;
  assign n980 = n979 ^ n977 ;
  assign n2842 = x219 ^ x91 ;
  assign n984 = n980 & ~n2842 ;
  assign n982 = x220 ^ x91 ;
  assign n985 = n984 ^ n982 ;
  assign n2853 = x220 ^ x92 ;
  assign n989 = n985 & ~n2853 ;
  assign n987 = x221 ^ x92 ;
  assign n990 = n989 ^ n987 ;
  assign n2864 = x221 ^ x93 ;
  assign n994 = n990 & ~n2864 ;
  assign n992 = x222 ^ x93 ;
  assign n995 = n994 ^ n992 ;
  assign n997 = x223 ^ x94 ;
  assign n996 = x223 ^ x222 ;
  assign n998 = n997 ^ n996 ;
  assign n999 = n995 & ~n998 ;
  assign n1000 = n999 ^ n997 ;
  assign n1002 = x224 ^ x95 ;
  assign n1001 = x224 ^ x223 ;
  assign n1003 = n1002 ^ n1001 ;
  assign n1004 = n1000 & ~n1003 ;
  assign n1005 = n1004 ^ n1002 ;
  assign n1007 = x225 ^ x96 ;
  assign n1006 = x225 ^ x224 ;
  assign n1008 = n1007 ^ n1006 ;
  assign n1009 = n1005 & ~n1008 ;
  assign n1010 = n1009 ^ n1007 ;
  assign n1012 = x226 ^ x97 ;
  assign n1011 = x226 ^ x225 ;
  assign n1013 = n1012 ^ n1011 ;
  assign n1014 = n1010 & ~n1013 ;
  assign n1015 = n1014 ^ n1012 ;
  assign n1017 = x227 ^ x98 ;
  assign n1016 = x227 ^ x226 ;
  assign n1018 = n1017 ^ n1016 ;
  assign n1019 = n1015 & ~n1018 ;
  assign n1020 = n1019 ^ n1017 ;
  assign n1022 = x228 ^ x99 ;
  assign n1021 = x228 ^ x227 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = n1024 ^ n1022 ;
  assign n1027 = x229 ^ x100 ;
  assign n1026 = x229 ^ x228 ;
  assign n1028 = n1027 ^ n1026 ;
  assign n1029 = n1025 & ~n1028 ;
  assign n1030 = n1029 ^ n1027 ;
  assign n1032 = x230 ^ x101 ;
  assign n1031 = x230 ^ x229 ;
  assign n1033 = n1032 ^ n1031 ;
  assign n1034 = n1030 & ~n1033 ;
  assign n1035 = n1034 ^ n1032 ;
  assign n1037 = x231 ^ x102 ;
  assign n1036 = x231 ^ x230 ;
  assign n1038 = n1037 ^ n1036 ;
  assign n1039 = n1035 & ~n1038 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n2960 = x231 ^ x103 ;
  assign n1044 = n1040 & ~n2960 ;
  assign n1042 = x232 ^ x103 ;
  assign n1045 = n1044 ^ n1042 ;
  assign n1047 = x233 ^ x104 ;
  assign n1046 = x233 ^ x232 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1049 = n1045 & ~n1048 ;
  assign n1050 = n1049 ^ n1047 ;
  assign n1052 = x234 ^ x105 ;
  assign n1051 = x234 ^ x233 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1054 = n1050 & ~n1053 ;
  assign n1055 = n1054 ^ n1052 ;
  assign n2993 = x234 ^ x106 ;
  assign n1059 = n1055 & ~n2993 ;
  assign n1057 = x235 ^ x106 ;
  assign n1060 = n1059 ^ n1057 ;
  assign n3004 = x235 ^ x107 ;
  assign n1064 = n1060 & ~n3004 ;
  assign n1062 = x236 ^ x107 ;
  assign n1065 = n1064 ^ n1062 ;
  assign n1067 = x237 ^ x108 ;
  assign n1066 = x237 ^ x236 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n1069 = n1065 & ~n1068 ;
  assign n1070 = n1069 ^ n1067 ;
  assign n1072 = x238 ^ x109 ;
  assign n1071 = x238 ^ x237 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1074 = n1070 & ~n1073 ;
  assign n1075 = n1074 ^ n1072 ;
  assign n1077 = x239 ^ x110 ;
  assign n1076 = x239 ^ x238 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1079 = n1075 & ~n1078 ;
  assign n1080 = n1079 ^ n1077 ;
  assign n1082 = x240 ^ x111 ;
  assign n1081 = x240 ^ x239 ;
  assign n1083 = n1082 ^ n1081 ;
  assign n1084 = n1080 & ~n1083 ;
  assign n1085 = n1084 ^ n1082 ;
  assign n1087 = x241 ^ x112 ;
  assign n1086 = x241 ^ x240 ;
  assign n1088 = n1087 ^ n1086 ;
  assign n1089 = n1085 & ~n1088 ;
  assign n1090 = n1089 ^ n1087 ;
  assign n3059 = x241 ^ x113 ;
  assign n1094 = n1090 & ~n3059 ;
  assign n1092 = x242 ^ x113 ;
  assign n1095 = n1094 ^ n1092 ;
  assign n1097 = x243 ^ x114 ;
  assign n1096 = x243 ^ x242 ;
  assign n1098 = n1097 ^ n1096 ;
  assign n1099 = n1095 & ~n1098 ;
  assign n1100 = n1099 ^ n1097 ;
  assign n1102 = x244 ^ x115 ;
  assign n1101 = x244 ^ x243 ;
  assign n1103 = n1102 ^ n1101 ;
  assign n1104 = n1100 & ~n1103 ;
  assign n1105 = n1104 ^ n1102 ;
  assign n3092 = x244 ^ x116 ;
  assign n1109 = n1105 & ~n3092 ;
  assign n1107 = x245 ^ x116 ;
  assign n1110 = n1109 ^ n1107 ;
  assign n3103 = x245 ^ x117 ;
  assign n1114 = n1110 & ~n3103 ;
  assign n1112 = x246 ^ x117 ;
  assign n1115 = n1114 ^ n1112 ;
  assign n3114 = x246 ^ x118 ;
  assign n1119 = n1115 & ~n3114 ;
  assign n1117 = x247 ^ x118 ;
  assign n1120 = n1119 ^ n1117 ;
  assign n3125 = x247 ^ x119 ;
  assign n1124 = n1120 & ~n3125 ;
  assign n1122 = x248 ^ x119 ;
  assign n1125 = n1124 ^ n1122 ;
  assign n1127 = x249 ^ x120 ;
  assign n1126 = x249 ^ x248 ;
  assign n1128 = n1127 ^ n1126 ;
  assign n1129 = n1125 & ~n1128 ;
  assign n1130 = n1129 ^ n1127 ;
  assign n1132 = x250 ^ x121 ;
  assign n1131 = x250 ^ x249 ;
  assign n1133 = n1132 ^ n1131 ;
  assign n1134 = n1130 & ~n1133 ;
  assign n1135 = n1134 ^ n1132 ;
  assign n1136 = ~n516 & n1135 ;
  assign n1137 = n1136 ^ x122 ;
  assign n1138 = ~n515 & ~n1137 ;
  assign n1139 = ~x124 & x252 ;
  assign n1140 = x253 ^ x125 ;
  assign n1141 = ~n1139 & ~n1140 ;
  assign n1142 = x254 ^ x126 ;
  assign n1143 = x251 ^ x123 ;
  assign n1144 = n1143 ^ n515 ;
  assign n1145 = ~n1142 & ~n1144 ;
  assign n1146 = n1141 & n1145 ;
  assign n1147 = ~n1138 & n1146 ;
  assign n1149 = n1139 ^ x253 ;
  assign n1148 = x252 ^ x124 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1154 = ~n1140 & n1150 ;
  assign n1152 = x254 ^ x125 ;
  assign n1155 = n1154 ^ n1152 ;
  assign n1156 = ~n1142 & n1155 ;
  assign n1157 = n1156 ^ x126 ;
  assign n1158 = ~n1147 & ~n1157 ;
  assign n1159 = n1158 ^ x255 ;
  assign n1160 = ~n514 & n1159 ;
  assign n1161 = n1160 ^ x127 ;
  assign n1162 = n513 & n1161 ;
  assign n1163 = n1162 ^ x0 ;
  assign n1832 = n1831 ^ n1163 ;
  assign n1834 = x383 & x511 ;
  assign n1833 = x127 & x255 ;
  assign n1835 = n1834 ^ n1833 ;
  assign n3181 = n1140 & n1161 ;
  assign n3182 = n3181 ^ x125 ;
  assign n1836 = n1142 & n1161 ;
  assign n1837 = n1836 ^ x126 ;
  assign n3191 = n3182 ^ n1837 ;
  assign n3171 = n1810 & n1829 ;
  assign n3172 = n3171 ^ x380 ;
  assign n3183 = n3182 ^ n3172 ;
  assign n3161 = n1168 & n1829 ;
  assign n3162 = n3161 ^ x379 ;
  assign n3173 = n3172 ^ n3162 ;
  assign n3151 = n516 & n1161 ;
  assign n3152 = n3151 ^ x122 ;
  assign n3163 = n3162 ^ n3152 ;
  assign n1843 = n1829 & n1842 ;
  assign n1844 = n1843 ^ x377 ;
  assign n3153 = n3152 ^ n1844 ;
  assign n3126 = n1161 & n3125 ;
  assign n3127 = n3126 ^ x119 ;
  assign n1840 = n1829 & n1839 ;
  assign n1841 = n1840 ^ x376 ;
  assign n3136 = n3127 ^ n1841 ;
  assign n3115 = n1161 & n3114 ;
  assign n3116 = n3115 ^ x118 ;
  assign n3128 = n3127 ^ n3116 ;
  assign n3104 = n1161 & n3103 ;
  assign n3105 = n3104 ^ x117 ;
  assign n3117 = n3116 ^ n3105 ;
  assign n3093 = n1161 & n3092 ;
  assign n3094 = n3093 ^ x116 ;
  assign n3106 = n3105 ^ n3094 ;
  assign n3082 = n1829 & n3081 ;
  assign n3083 = n3082 ^ x371 ;
  assign n3095 = n3094 ^ n3083 ;
  assign n3071 = n1829 & n3070 ;
  assign n3072 = n3071 ^ x370 ;
  assign n3084 = n3083 ^ n3072 ;
  assign n3060 = n1161 & n3059 ;
  assign n3061 = n3060 ^ x113 ;
  assign n3073 = n3072 ^ n3061 ;
  assign n3049 = n1829 & n3048 ;
  assign n3050 = n3049 ^ x368 ;
  assign n3062 = n3061 ^ n3050 ;
  assign n3038 = n1829 & n3037 ;
  assign n3039 = n3038 ^ x367 ;
  assign n3051 = n3050 ^ n3039 ;
  assign n1850 = n1829 & n1849 ;
  assign n1851 = n1850 ^ x366 ;
  assign n3040 = n3039 ^ n1851 ;
  assign n3005 = n1161 & n3004 ;
  assign n3006 = n3005 ^ x107 ;
  assign n1854 = n1829 & n1853 ;
  assign n1855 = n1854 ^ x364 ;
  assign n3015 = n3006 ^ n1855 ;
  assign n2994 = n1161 & n2993 ;
  assign n2995 = n2994 ^ x106 ;
  assign n3007 = n3006 ^ n2995 ;
  assign n2983 = n1829 & n2982 ;
  assign n2984 = n2983 ^ x361 ;
  assign n2996 = n2995 ^ n2984 ;
  assign n2972 = n1829 & n2971 ;
  assign n2973 = n2972 ^ x360 ;
  assign n2985 = n2984 ^ n2973 ;
  assign n2961 = n1161 & n2960 ;
  assign n2962 = n2961 ^ x103 ;
  assign n2974 = n2973 ^ n2962 ;
  assign n2950 = n1829 & n2949 ;
  assign n2951 = n2950 ^ x358 ;
  assign n2963 = n2962 ^ n2951 ;
  assign n1861 = n1829 & n1860 ;
  assign n1862 = n1861 ^ x357 ;
  assign n2952 = n2951 ^ n1862 ;
  assign n2924 = n1829 & n2923 ;
  assign n2925 = n2924 ^ x355 ;
  assign n1858 = n1829 & n1857 ;
  assign n1859 = n1858 ^ x356 ;
  assign n2934 = n2925 ^ n1859 ;
  assign n2913 = n1829 & n2912 ;
  assign n2914 = n2913 ^ x354 ;
  assign n2926 = n2925 ^ n2914 ;
  assign n1868 = n1829 & n1867 ;
  assign n1869 = n1868 ^ x353 ;
  assign n2915 = n2914 ^ n1869 ;
  assign n2887 = n1829 & n2886 ;
  assign n2888 = n2887 ^ x351 ;
  assign n1865 = n1829 & n1864 ;
  assign n1866 = n1865 ^ x352 ;
  assign n2897 = n2888 ^ n1866 ;
  assign n2876 = n1829 & n2875 ;
  assign n2877 = n2876 ^ x350 ;
  assign n2889 = n2888 ^ n2877 ;
  assign n2865 = n1161 & n2864 ;
  assign n2866 = n2865 ^ x93 ;
  assign n2878 = n2877 ^ n2866 ;
  assign n2854 = n1161 & n2853 ;
  assign n2855 = n2854 ^ x92 ;
  assign n2867 = n2866 ^ n2855 ;
  assign n2843 = n1161 & n2842 ;
  assign n2844 = n2843 ^ x91 ;
  assign n2856 = n2855 ^ n2844 ;
  assign n2832 = n1829 & n2831 ;
  assign n2833 = n2832 ^ x346 ;
  assign n2845 = n2844 ^ n2833 ;
  assign n2821 = n1829 & n2820 ;
  assign n2822 = n2821 ^ x345 ;
  assign n2834 = n2833 ^ n2822 ;
  assign n2810 = n1829 & n2809 ;
  assign n2811 = n2810 ^ x344 ;
  assign n2823 = n2822 ^ n2811 ;
  assign n2799 = n1161 & n2798 ;
  assign n2800 = n2799 ^ x87 ;
  assign n2812 = n2811 ^ n2800 ;
  assign n2788 = n1161 & n2787 ;
  assign n2789 = n2788 ^ x86 ;
  assign n2801 = n2800 ^ n2789 ;
  assign n2777 = n1161 & n2776 ;
  assign n2778 = n2777 ^ x85 ;
  assign n2790 = n2789 ^ n2778 ;
  assign n2766 = n1161 & n2765 ;
  assign n2767 = n2766 ^ x84 ;
  assign n2779 = n2778 ^ n2767 ;
  assign n2755 = n1161 & n2754 ;
  assign n2756 = n2755 ^ x83 ;
  assign n2768 = n2767 ^ n2756 ;
  assign n2744 = n1829 & n2743 ;
  assign n2745 = n2744 ^ x338 ;
  assign n2757 = n2756 ^ n2745 ;
  assign n1875 = n1829 & n1874 ;
  assign n1876 = n1875 ^ x337 ;
  assign n2746 = n2745 ^ n1876 ;
  assign n2718 = n1161 & n2717 ;
  assign n2719 = n2718 ^ x79 ;
  assign n1872 = n1829 & n1871 ;
  assign n1873 = n1872 ^ x336 ;
  assign n2728 = n2719 ^ n1873 ;
  assign n2707 = n1161 & n2706 ;
  assign n2708 = n2707 ^ x78 ;
  assign n2720 = n2719 ^ n2708 ;
  assign n2696 = n1161 & n2695 ;
  assign n2697 = n2696 ^ x77 ;
  assign n2709 = n2708 ^ n2697 ;
  assign n2685 = n1161 & n2684 ;
  assign n2686 = n2685 ^ x76 ;
  assign n2698 = n2697 ^ n2686 ;
  assign n2674 = n1829 & n2673 ;
  assign n2675 = n2674 ^ x331 ;
  assign n2687 = n2686 ^ n2675 ;
  assign n2663 = n1161 & n2662 ;
  assign n2664 = n2663 ^ x74 ;
  assign n2676 = n2675 ^ n2664 ;
  assign n2652 = n1161 & n2651 ;
  assign n2653 = n2652 ^ x73 ;
  assign n2665 = n2664 ^ n2653 ;
  assign n1881 = n1829 & n1880 ;
  assign n1882 = n1881 ^ x328 ;
  assign n2654 = n2653 ^ n1882 ;
  assign n2612 = n517 & n1161 ;
  assign n2613 = n2612 ^ x68 ;
  assign n1887 = n1173 & n1829 ;
  assign n1888 = n1887 ^ x325 ;
  assign n2622 = n2613 ^ n1888 ;
  assign n1892 = n1176 & n1829 ;
  assign n1893 = n1892 ^ x323 ;
  assign n2614 = n2613 ^ n1893 ;
  assign n2561 = n522 & n1161 ;
  assign n2562 = n2561 ^ x61 ;
  assign n1905 = n1197 & n1829 ;
  assign n1906 = n1905 ^ x318 ;
  assign n2571 = n2562 ^ n1906 ;
  assign n2551 = n1190 & n1829 ;
  assign n2552 = n2551 ^ x316 ;
  assign n2563 = n2562 ^ n2552 ;
  assign n2541 = n525 & n1161 ;
  assign n2542 = n2541 ^ x59 ;
  assign n2553 = n2552 ^ n2542 ;
  assign n2531 = n532 & n1161 ;
  assign n2532 = n2531 ^ x58 ;
  assign n2543 = n2542 ^ n2532 ;
  assign n2521 = n1161 & n2520 ;
  assign n2522 = n2521 ^ x57 ;
  assign n2533 = n2532 ^ n2522 ;
  assign n2510 = n1829 & n2509 ;
  assign n2511 = n2510 ^ x312 ;
  assign n2523 = n2522 ^ n2511 ;
  assign n2499 = n1161 & n2498 ;
  assign n2500 = n2499 ^ x55 ;
  assign n2512 = n2511 ^ n2500 ;
  assign n2488 = n1829 & n2487 ;
  assign n2489 = n2488 ^ x310 ;
  assign n2501 = n2500 ^ n2489 ;
  assign n2477 = n1161 & n2476 ;
  assign n2478 = n2477 ^ x53 ;
  assign n2490 = n2489 ^ n2478 ;
  assign n2466 = n1829 & n2465 ;
  assign n2467 = n2466 ^ x308 ;
  assign n2479 = n2478 ^ n2467 ;
  assign n2455 = n1161 & n2454 ;
  assign n2456 = n2455 ^ x51 ;
  assign n2468 = n2467 ^ n2456 ;
  assign n2444 = n1161 & n2443 ;
  assign n2445 = n2444 ^ x50 ;
  assign n2457 = n2456 ^ n2445 ;
  assign n2433 = n1829 & n2432 ;
  assign n2434 = n2433 ^ x305 ;
  assign n2446 = n2445 ^ n2434 ;
  assign n2422 = n1161 & n2421 ;
  assign n2423 = n2422 ^ x48 ;
  assign n2435 = n2434 ^ n2423 ;
  assign n1912 = n1829 & n1911 ;
  assign n1913 = n1912 ^ x303 ;
  assign n2424 = n2423 ^ n1913 ;
  assign n2389 = n533 & n1161 ;
  assign n2390 = n2389 ^ x44 ;
  assign n1916 = n1829 & n1915 ;
  assign n1917 = n1916 ^ x301 ;
  assign n2399 = n2390 ^ n1917 ;
  assign n2379 = n536 & n1161 ;
  assign n2380 = n2379 ^ x43 ;
  assign n2391 = n2390 ^ n2380 ;
  assign n1921 = n1208 & n1829 ;
  assign n1922 = n1921 ^ x298 ;
  assign n2381 = n2380 ^ n1922 ;
  assign n2333 = n1161 & n2332 ;
  assign n2334 = n2333 ^ x37 ;
  assign n1930 = n1218 & n1829 ;
  assign n1931 = n1930 ^ x294 ;
  assign n2343 = n2334 ^ n1931 ;
  assign n1937 = n1829 & n1936 ;
  assign n1938 = n1937 ^ x292 ;
  assign n2335 = n2334 ^ n1938 ;
  assign n2307 = n1161 & n2306 ;
  assign n2308 = n2307 ^ x34 ;
  assign n1934 = n1829 & n1933 ;
  assign n1935 = n1934 ^ x291 ;
  assign n2317 = n2308 ^ n1935 ;
  assign n1944 = n1829 & n1943 ;
  assign n1945 = n1944 ^ x289 ;
  assign n2309 = n2308 ^ n1945 ;
  assign n2274 = n1161 & n2273 ;
  assign n2275 = n2274 ^ x30 ;
  assign n1948 = n1829 & n1947 ;
  assign n1949 = n1948 ^ x287 ;
  assign n2284 = n2275 ^ n1949 ;
  assign n1955 = n1829 & n1954 ;
  assign n1956 = n1955 ^ x285 ;
  assign n2276 = n2275 ^ n1956 ;
  assign n2248 = n1161 & n2247 ;
  assign n2249 = n2248 ^ x27 ;
  assign n1952 = n1829 & n1951 ;
  assign n1953 = n1952 ^ x284 ;
  assign n2258 = n2249 ^ n1953 ;
  assign n1962 = n1829 & n1961 ;
  assign n1963 = n1962 ^ x282 ;
  assign n2250 = n2249 ^ n1963 ;
  assign n2215 = n1161 & n2214 ;
  assign n2216 = n2215 ^ x23 ;
  assign n1966 = n1829 & n1965 ;
  assign n1967 = n1966 ^ x280 ;
  assign n2225 = n2216 ^ n1967 ;
  assign n2204 = n1161 & n2203 ;
  assign n2205 = n2204 ^ x22 ;
  assign n2217 = n2216 ^ n2205 ;
  assign n2193 = n1161 & n2192 ;
  assign n2194 = n2193 ^ x21 ;
  assign n2206 = n2205 ^ n2194 ;
  assign n2182 = n1829 & n2181 ;
  assign n2183 = n2182 ^ x276 ;
  assign n2195 = n2194 ^ n2183 ;
  assign n2171 = n1161 & n2170 ;
  assign n2172 = n2171 ^ x19 ;
  assign n2184 = n2183 ^ n2172 ;
  assign n1973 = n1829 & n1972 ;
  assign n1974 = n1973 ^ x274 ;
  assign n2173 = n2172 ^ n1974 ;
  assign n2145 = n1161 & n2144 ;
  assign n2146 = n2145 ^ x16 ;
  assign n1970 = n1829 & n1969 ;
  assign n1971 = n1970 ^ x273 ;
  assign n2155 = n2146 ^ n1971 ;
  assign n2134 = n1829 & n2133 ;
  assign n2135 = n2134 ^ x271 ;
  assign n2147 = n2146 ^ n2135 ;
  assign n2123 = n1161 & n2122 ;
  assign n2124 = n2123 ^ x14 ;
  assign n2136 = n2135 ^ n2124 ;
  assign n2112 = n1161 & n2111 ;
  assign n2113 = n2112 ^ x13 ;
  assign n2125 = n2124 ^ n2113 ;
  assign n1980 = n1829 & n1979 ;
  assign n1981 = n1980 ^ x268 ;
  assign n2114 = n2113 ^ n1981 ;
  assign n2079 = n1161 & n2078 ;
  assign n2080 = n2079 ^ x9 ;
  assign n1984 = n1829 & n1983 ;
  assign n1985 = n1984 ^ x266 ;
  assign n2089 = n2080 ^ n1985 ;
  assign n2068 = n1161 & n2067 ;
  assign n2069 = n2068 ^ x8 ;
  assign n2081 = n2080 ^ n2069 ;
  assign n2057 = n1829 & n2056 ;
  assign n2058 = n2057 ^ x263 ;
  assign n2070 = n2069 ^ n2058 ;
  assign n2046 = n1161 & n2045 ;
  assign n2047 = n2046 ^ x6 ;
  assign n2059 = n2058 ^ n2047 ;
  assign n1991 = n1829 & n1990 ;
  assign n1992 = n1991 ^ x261 ;
  assign n2048 = n2047 ^ n1992 ;
  assign n2020 = n1161 & n2019 ;
  assign n2021 = n2020 ^ x3 ;
  assign n1988 = n1829 & n1987 ;
  assign n1989 = n1988 ^ x260 ;
  assign n2030 = n2021 ^ n1989 ;
  assign n2009 = n1161 & n2008 ;
  assign n2010 = n2009 ^ x2 ;
  assign n2022 = n2021 ^ n2010 ;
  assign n1998 = n1161 & n1997 ;
  assign n1999 = n1998 ^ x1 ;
  assign n2011 = n2010 ^ n1999 ;
  assign n1995 = n1829 & n1994 ;
  assign n1996 = n1995 ^ x257 ;
  assign n2000 = n1999 ^ n1996 ;
  assign n2005 = n1163 & ~n1831 ;
  assign n2006 = n2005 ^ n1996 ;
  assign n2007 = ~n2000 & n2006 ;
  assign n2012 = n2011 ^ n2007 ;
  assign n2013 = n2010 ^ x258 ;
  assign n2014 = n2013 ^ x386 ;
  assign n2015 = n2014 ^ n2010 ;
  assign n2016 = n1829 & n2015 ;
  assign n2017 = n2016 ^ n2013 ;
  assign n2018 = n2012 & ~n2017 ;
  assign n2023 = n2022 ^ n2018 ;
  assign n2024 = n2021 ^ x259 ;
  assign n2025 = n2024 ^ x387 ;
  assign n2026 = n2025 ^ n2021 ;
  assign n2027 = n1829 & n2026 ;
  assign n2028 = n2027 ^ n2024 ;
  assign n2029 = n2023 & ~n2028 ;
  assign n2031 = n2030 ^ n2029 ;
  assign n2032 = n1989 ^ x4 ;
  assign n2033 = n2032 ^ x132 ;
  assign n2034 = n2033 ^ n1989 ;
  assign n2035 = n1161 & n2034 ;
  assign n2036 = n2035 ^ n2032 ;
  assign n2037 = ~n2031 & ~n2036 ;
  assign n1993 = n1992 ^ n1989 ;
  assign n2038 = n2037 ^ n1993 ;
  assign n2039 = n1992 ^ x5 ;
  assign n2040 = n2039 ^ x133 ;
  assign n2041 = n2040 ^ n1992 ;
  assign n2042 = n1161 & n2041 ;
  assign n2043 = n2042 ^ n2039 ;
  assign n2044 = n2038 & ~n2043 ;
  assign n2049 = n2048 ^ n2044 ;
  assign n2050 = n2047 ^ x262 ;
  assign n2051 = n2050 ^ x390 ;
  assign n2052 = n2051 ^ n2047 ;
  assign n2053 = n1829 & n2052 ;
  assign n2054 = n2053 ^ n2050 ;
  assign n2055 = ~n2049 & ~n2054 ;
  assign n2060 = n2059 ^ n2055 ;
  assign n2061 = n2058 ^ x7 ;
  assign n2062 = n2061 ^ x135 ;
  assign n2063 = n2062 ^ n2058 ;
  assign n2064 = n1161 & n2063 ;
  assign n2065 = n2064 ^ n2061 ;
  assign n2066 = ~n2060 & ~n2065 ;
  assign n2071 = n2070 ^ n2066 ;
  assign n2072 = n2069 ^ x264 ;
  assign n2073 = n2072 ^ x392 ;
  assign n2074 = n2073 ^ n2069 ;
  assign n2075 = n1829 & n2074 ;
  assign n2076 = n2075 ^ n2072 ;
  assign n2077 = ~n2071 & ~n2076 ;
  assign n2082 = n2081 ^ n2077 ;
  assign n2083 = n2080 ^ x265 ;
  assign n2084 = n2083 ^ x393 ;
  assign n2085 = n2084 ^ n2080 ;
  assign n2086 = n1829 & n2085 ;
  assign n2087 = n2086 ^ n2083 ;
  assign n2088 = n2082 & ~n2087 ;
  assign n2090 = n2089 ^ n2088 ;
  assign n2091 = n1985 ^ x10 ;
  assign n2092 = n2091 ^ x138 ;
  assign n2093 = n2092 ^ n1985 ;
  assign n2094 = n1161 & n2093 ;
  assign n2095 = n2094 ^ n2091 ;
  assign n2096 = ~n2090 & ~n2095 ;
  assign n1977 = n1829 & n1976 ;
  assign n1978 = n1977 ^ x267 ;
  assign n1986 = n1985 ^ n1978 ;
  assign n2097 = n2096 ^ n1986 ;
  assign n2098 = n1978 ^ x11 ;
  assign n2099 = n2098 ^ x139 ;
  assign n2100 = n2099 ^ n1978 ;
  assign n2101 = n1161 & n2100 ;
  assign n2102 = n2101 ^ n2098 ;
  assign n2103 = n2097 & ~n2102 ;
  assign n1982 = n1981 ^ n1978 ;
  assign n2104 = n2103 ^ n1982 ;
  assign n2105 = n1981 ^ x12 ;
  assign n2106 = n2105 ^ x140 ;
  assign n2107 = n2106 ^ n1981 ;
  assign n2108 = n1161 & n2107 ;
  assign n2109 = n2108 ^ n2105 ;
  assign n2110 = n2104 & ~n2109 ;
  assign n2115 = n2114 ^ n2110 ;
  assign n2116 = n2113 ^ x269 ;
  assign n2117 = n2116 ^ x397 ;
  assign n2118 = n2117 ^ n2113 ;
  assign n2119 = n1829 & n2118 ;
  assign n2120 = n2119 ^ n2116 ;
  assign n2121 = ~n2115 & ~n2120 ;
  assign n2126 = n2125 ^ n2121 ;
  assign n2127 = n2124 ^ x270 ;
  assign n2128 = n2127 ^ x398 ;
  assign n2129 = n2128 ^ n2124 ;
  assign n2130 = n1829 & n2129 ;
  assign n2131 = n2130 ^ n2127 ;
  assign n2132 = n2126 & ~n2131 ;
  assign n2137 = n2136 ^ n2132 ;
  assign n2138 = n2135 ^ x15 ;
  assign n2139 = n2138 ^ x143 ;
  assign n2140 = n2139 ^ n2135 ;
  assign n2141 = n1161 & n2140 ;
  assign n2142 = n2141 ^ n2138 ;
  assign n2143 = ~n2137 & ~n2142 ;
  assign n2148 = n2147 ^ n2143 ;
  assign n2149 = n2146 ^ x272 ;
  assign n2150 = n2149 ^ x400 ;
  assign n2151 = n2150 ^ n2146 ;
  assign n2152 = n1829 & n2151 ;
  assign n2153 = n2152 ^ n2149 ;
  assign n2154 = ~n2148 & ~n2153 ;
  assign n2156 = n2155 ^ n2154 ;
  assign n2157 = n1971 ^ x17 ;
  assign n2158 = n2157 ^ x145 ;
  assign n2159 = n2158 ^ n1971 ;
  assign n2160 = n1161 & n2159 ;
  assign n2161 = n2160 ^ n2157 ;
  assign n2162 = ~n2156 & ~n2161 ;
  assign n1975 = n1974 ^ n1971 ;
  assign n2163 = n2162 ^ n1975 ;
  assign n2164 = n1974 ^ x18 ;
  assign n2165 = n2164 ^ x146 ;
  assign n2166 = n2165 ^ n1974 ;
  assign n2167 = n1161 & n2166 ;
  assign n2168 = n2167 ^ n2164 ;
  assign n2169 = n2163 & ~n2168 ;
  assign n2174 = n2173 ^ n2169 ;
  assign n2175 = n2172 ^ x275 ;
  assign n2176 = n2175 ^ x403 ;
  assign n2177 = n2176 ^ n2172 ;
  assign n2178 = n1829 & n2177 ;
  assign n2179 = n2178 ^ n2175 ;
  assign n2180 = ~n2174 & ~n2179 ;
  assign n2185 = n2184 ^ n2180 ;
  assign n2186 = n2183 ^ x20 ;
  assign n2187 = n2186 ^ x148 ;
  assign n2188 = n2187 ^ n2183 ;
  assign n2189 = n1161 & n2188 ;
  assign n2190 = n2189 ^ n2186 ;
  assign n2191 = ~n2185 & ~n2190 ;
  assign n2196 = n2195 ^ n2191 ;
  assign n2197 = n2194 ^ x277 ;
  assign n2198 = n2197 ^ x405 ;
  assign n2199 = n2198 ^ n2194 ;
  assign n2200 = n1829 & n2199 ;
  assign n2201 = n2200 ^ n2197 ;
  assign n2202 = ~n2196 & ~n2201 ;
  assign n2207 = n2206 ^ n2202 ;
  assign n2208 = n2205 ^ x278 ;
  assign n2209 = n2208 ^ x406 ;
  assign n2210 = n2209 ^ n2205 ;
  assign n2211 = n1829 & n2210 ;
  assign n2212 = n2211 ^ n2208 ;
  assign n2213 = n2207 & ~n2212 ;
  assign n2218 = n2217 ^ n2213 ;
  assign n2219 = n2216 ^ x279 ;
  assign n2220 = n2219 ^ x407 ;
  assign n2221 = n2220 ^ n2216 ;
  assign n2222 = n1829 & n2221 ;
  assign n2223 = n2222 ^ n2219 ;
  assign n2224 = n2218 & ~n2223 ;
  assign n2226 = n2225 ^ n2224 ;
  assign n2227 = n1967 ^ x24 ;
  assign n2228 = n2227 ^ x152 ;
  assign n2229 = n2228 ^ n1967 ;
  assign n2230 = n1161 & n2229 ;
  assign n2231 = n2230 ^ n2227 ;
  assign n2232 = ~n2226 & ~n2231 ;
  assign n1959 = n1829 & n1958 ;
  assign n1960 = n1959 ^ x281 ;
  assign n1968 = n1967 ^ n1960 ;
  assign n2233 = n2232 ^ n1968 ;
  assign n2234 = n1960 ^ x25 ;
  assign n2235 = n2234 ^ x153 ;
  assign n2236 = n2235 ^ n1960 ;
  assign n2237 = n1161 & n2236 ;
  assign n2238 = n2237 ^ n2234 ;
  assign n2239 = n2233 & ~n2238 ;
  assign n1964 = n1963 ^ n1960 ;
  assign n2240 = n2239 ^ n1964 ;
  assign n2241 = n1963 ^ x26 ;
  assign n2242 = n2241 ^ x154 ;
  assign n2243 = n2242 ^ n1963 ;
  assign n2244 = n1161 & n2243 ;
  assign n2245 = n2244 ^ n2241 ;
  assign n2246 = n2240 & ~n2245 ;
  assign n2251 = n2250 ^ n2246 ;
  assign n2252 = n2249 ^ x283 ;
  assign n2253 = n2252 ^ x411 ;
  assign n2254 = n2253 ^ n2249 ;
  assign n2255 = n1829 & n2254 ;
  assign n2256 = n2255 ^ n2252 ;
  assign n2257 = ~n2251 & ~n2256 ;
  assign n2259 = n2258 ^ n2257 ;
  assign n2260 = n1953 ^ x28 ;
  assign n2261 = n2260 ^ x156 ;
  assign n2262 = n2261 ^ n1953 ;
  assign n2263 = n1161 & n2262 ;
  assign n2264 = n2263 ^ n2260 ;
  assign n2265 = ~n2259 & ~n2264 ;
  assign n1957 = n1956 ^ n1953 ;
  assign n2266 = n2265 ^ n1957 ;
  assign n2267 = n1956 ^ x29 ;
  assign n2268 = n2267 ^ x157 ;
  assign n2269 = n2268 ^ n1956 ;
  assign n2270 = n1161 & n2269 ;
  assign n2271 = n2270 ^ n2267 ;
  assign n2272 = n2266 & ~n2271 ;
  assign n2277 = n2276 ^ n2272 ;
  assign n2278 = n2275 ^ x286 ;
  assign n2279 = n2278 ^ x414 ;
  assign n2280 = n2279 ^ n2275 ;
  assign n2281 = n1829 & n2280 ;
  assign n2282 = n2281 ^ n2278 ;
  assign n2283 = ~n2277 & ~n2282 ;
  assign n2285 = n2284 ^ n2283 ;
  assign n2286 = n1949 ^ x31 ;
  assign n2287 = n2286 ^ x159 ;
  assign n2288 = n2287 ^ n1949 ;
  assign n2289 = n1161 & n2288 ;
  assign n2290 = n2289 ^ n2286 ;
  assign n2291 = ~n2285 & ~n2290 ;
  assign n1941 = n1829 & n1940 ;
  assign n1942 = n1941 ^ x288 ;
  assign n1950 = n1949 ^ n1942 ;
  assign n2292 = n2291 ^ n1950 ;
  assign n2293 = n1942 ^ x32 ;
  assign n2294 = n2293 ^ x160 ;
  assign n2295 = n2294 ^ n1942 ;
  assign n2296 = n1161 & n2295 ;
  assign n2297 = n2296 ^ n2293 ;
  assign n2298 = n2292 & ~n2297 ;
  assign n1946 = n1945 ^ n1942 ;
  assign n2299 = n2298 ^ n1946 ;
  assign n2300 = n1945 ^ x33 ;
  assign n2301 = n2300 ^ x161 ;
  assign n2302 = n2301 ^ n1945 ;
  assign n2303 = n1161 & n2302 ;
  assign n2304 = n2303 ^ n2300 ;
  assign n2305 = n2299 & ~n2304 ;
  assign n2310 = n2309 ^ n2305 ;
  assign n2311 = n2308 ^ x290 ;
  assign n2312 = n2311 ^ x418 ;
  assign n2313 = n2312 ^ n2308 ;
  assign n2314 = n1829 & n2313 ;
  assign n2315 = n2314 ^ n2311 ;
  assign n2316 = ~n2310 & ~n2315 ;
  assign n2318 = n2317 ^ n2316 ;
  assign n2319 = n1935 ^ x35 ;
  assign n2320 = n2319 ^ x163 ;
  assign n2321 = n2320 ^ n1935 ;
  assign n2322 = n1161 & n2321 ;
  assign n2323 = n2322 ^ n2319 ;
  assign n2324 = ~n2318 & ~n2323 ;
  assign n1939 = n1938 ^ n1935 ;
  assign n2325 = n2324 ^ n1939 ;
  assign n2326 = n1938 ^ x36 ;
  assign n2327 = n2326 ^ x164 ;
  assign n2328 = n2327 ^ n1938 ;
  assign n2329 = n1161 & n2328 ;
  assign n2330 = n2329 ^ n2326 ;
  assign n2331 = n2325 & ~n2330 ;
  assign n2336 = n2335 ^ n2331 ;
  assign n2337 = n2334 ^ x293 ;
  assign n2338 = n2337 ^ x421 ;
  assign n2339 = n2338 ^ n2334 ;
  assign n2340 = n1829 & n2339 ;
  assign n2341 = n2340 ^ n2337 ;
  assign n2342 = ~n2336 & ~n2341 ;
  assign n2344 = n2343 ^ n2342 ;
  assign n2345 = n1931 ^ x38 ;
  assign n2346 = n2345 ^ x166 ;
  assign n2347 = n2346 ^ n1931 ;
  assign n2348 = n1161 & n2347 ;
  assign n2349 = n2348 ^ n2345 ;
  assign n2350 = ~n2344 & ~n2349 ;
  assign n1927 = n1211 & n1829 ;
  assign n1928 = n1927 ^ x295 ;
  assign n1932 = n1931 ^ n1928 ;
  assign n2351 = n2350 ^ n1932 ;
  assign n2355 = n540 & n1161 ;
  assign n2352 = n1928 ^ x39 ;
  assign n2356 = n2355 ^ n2352 ;
  assign n2357 = n2351 & ~n2356 ;
  assign n1924 = n1214 & n1829 ;
  assign n1925 = n1924 ^ x296 ;
  assign n1929 = n1928 ^ n1925 ;
  assign n2358 = n2357 ^ n1929 ;
  assign n2362 = n538 & n1161 ;
  assign n2359 = n1925 ^ x40 ;
  assign n2363 = n2362 ^ n2359 ;
  assign n2364 = n2358 & ~n2363 ;
  assign n1919 = n1207 & n1829 ;
  assign n1920 = n1919 ^ x297 ;
  assign n1926 = n1925 ^ n1920 ;
  assign n2365 = n2364 ^ n1926 ;
  assign n2366 = n1920 ^ x41 ;
  assign n2367 = n2366 ^ x169 ;
  assign n2368 = n2367 ^ n1920 ;
  assign n2369 = n1161 & n2368 ;
  assign n2370 = n2369 ^ n2366 ;
  assign n2371 = n2365 & ~n2370 ;
  assign n1923 = n1922 ^ n1920 ;
  assign n2372 = n2371 ^ n1923 ;
  assign n2373 = n1922 ^ x42 ;
  assign n2374 = n2373 ^ x170 ;
  assign n2375 = n2374 ^ n1922 ;
  assign n2376 = n1161 & n2375 ;
  assign n2377 = n2376 ^ n2373 ;
  assign n2378 = n2372 & ~n2377 ;
  assign n2382 = n2381 ^ n2378 ;
  assign n2386 = n1206 & n1829 ;
  assign n2383 = n2380 ^ x299 ;
  assign n2387 = n2386 ^ n2383 ;
  assign n2388 = ~n2382 & ~n2387 ;
  assign n2392 = n2391 ^ n2388 ;
  assign n2396 = n1203 & n1829 ;
  assign n2393 = n2390 ^ x300 ;
  assign n2397 = n2396 ^ n2393 ;
  assign n2398 = n2392 & ~n2397 ;
  assign n2400 = n2399 ^ n2398 ;
  assign n2401 = n1917 ^ x45 ;
  assign n2402 = n2401 ^ x173 ;
  assign n2403 = n2402 ^ n1917 ;
  assign n2404 = n1161 & n2403 ;
  assign n2405 = n2404 ^ n2401 ;
  assign n2406 = ~n2400 & ~n2405 ;
  assign n1909 = n1829 & n1908 ;
  assign n1910 = n1909 ^ x302 ;
  assign n1918 = n1917 ^ n1910 ;
  assign n2407 = n2406 ^ n1918 ;
  assign n2408 = n1910 ^ x46 ;
  assign n2409 = n2408 ^ x174 ;
  assign n2410 = n2409 ^ n1910 ;
  assign n2411 = n1161 & n2410 ;
  assign n2412 = n2411 ^ n2408 ;
  assign n2413 = n2407 & ~n2412 ;
  assign n1914 = n1913 ^ n1910 ;
  assign n2414 = n2413 ^ n1914 ;
  assign n2415 = n1913 ^ x47 ;
  assign n2416 = n2415 ^ x175 ;
  assign n2417 = n2416 ^ n1913 ;
  assign n2418 = n1161 & n2417 ;
  assign n2419 = n2418 ^ n2415 ;
  assign n2420 = n2414 & ~n2419 ;
  assign n2425 = n2424 ^ n2420 ;
  assign n2426 = n2423 ^ x304 ;
  assign n2427 = n2426 ^ x432 ;
  assign n2428 = n2427 ^ n2423 ;
  assign n2429 = n1829 & n2428 ;
  assign n2430 = n2429 ^ n2426 ;
  assign n2431 = ~n2425 & ~n2430 ;
  assign n2436 = n2435 ^ n2431 ;
  assign n2437 = n2434 ^ x49 ;
  assign n2438 = n2437 ^ x177 ;
  assign n2439 = n2438 ^ n2434 ;
  assign n2440 = n1161 & n2439 ;
  assign n2441 = n2440 ^ n2437 ;
  assign n2442 = ~n2436 & ~n2441 ;
  assign n2447 = n2446 ^ n2442 ;
  assign n2448 = n2445 ^ x306 ;
  assign n2449 = n2448 ^ x434 ;
  assign n2450 = n2449 ^ n2445 ;
  assign n2451 = n1829 & n2450 ;
  assign n2452 = n2451 ^ n2448 ;
  assign n2453 = ~n2447 & ~n2452 ;
  assign n2458 = n2457 ^ n2453 ;
  assign n2459 = n2456 ^ x307 ;
  assign n2460 = n2459 ^ x435 ;
  assign n2461 = n2460 ^ n2456 ;
  assign n2462 = n1829 & n2461 ;
  assign n2463 = n2462 ^ n2459 ;
  assign n2464 = n2458 & ~n2463 ;
  assign n2469 = n2468 ^ n2464 ;
  assign n2470 = n2467 ^ x52 ;
  assign n2471 = n2470 ^ x180 ;
  assign n2472 = n2471 ^ n2467 ;
  assign n2473 = n1161 & n2472 ;
  assign n2474 = n2473 ^ n2470 ;
  assign n2475 = ~n2469 & ~n2474 ;
  assign n2480 = n2479 ^ n2475 ;
  assign n2481 = n2478 ^ x309 ;
  assign n2482 = n2481 ^ x437 ;
  assign n2483 = n2482 ^ n2478 ;
  assign n2484 = n1829 & n2483 ;
  assign n2485 = n2484 ^ n2481 ;
  assign n2486 = ~n2480 & ~n2485 ;
  assign n2491 = n2490 ^ n2486 ;
  assign n2492 = n2489 ^ x54 ;
  assign n2493 = n2492 ^ x182 ;
  assign n2494 = n2493 ^ n2489 ;
  assign n2495 = n1161 & n2494 ;
  assign n2496 = n2495 ^ n2492 ;
  assign n2497 = ~n2491 & ~n2496 ;
  assign n2502 = n2501 ^ n2497 ;
  assign n2503 = n2500 ^ x311 ;
  assign n2504 = n2503 ^ x439 ;
  assign n2505 = n2504 ^ n2500 ;
  assign n2506 = n1829 & n2505 ;
  assign n2507 = n2506 ^ n2503 ;
  assign n2508 = ~n2502 & ~n2507 ;
  assign n2513 = n2512 ^ n2508 ;
  assign n2514 = n2511 ^ x56 ;
  assign n2515 = n2514 ^ x184 ;
  assign n2516 = n2515 ^ n2511 ;
  assign n2517 = n1161 & n2516 ;
  assign n2518 = n2517 ^ n2514 ;
  assign n2519 = ~n2513 & ~n2518 ;
  assign n2524 = n2523 ^ n2519 ;
  assign n2525 = n2522 ^ x313 ;
  assign n2526 = n2525 ^ x441 ;
  assign n2527 = n2526 ^ n2522 ;
  assign n2528 = n1829 & n2527 ;
  assign n2529 = n2528 ^ n2525 ;
  assign n2530 = ~n2524 & ~n2529 ;
  assign n2534 = n2533 ^ n2530 ;
  assign n2535 = n2532 ^ x314 ;
  assign n2536 = n2535 ^ x442 ;
  assign n2537 = n2536 ^ n2532 ;
  assign n2538 = n1829 & n2537 ;
  assign n2539 = n2538 ^ n2535 ;
  assign n2540 = n2534 & ~n2539 ;
  assign n2544 = n2543 ^ n2540 ;
  assign n2548 = n1202 & n1829 ;
  assign n2545 = n2542 ^ x315 ;
  assign n2549 = n2548 ^ n2545 ;
  assign n2550 = n2544 & ~n2549 ;
  assign n2554 = n2553 ^ n2550 ;
  assign n2555 = n2552 ^ x60 ;
  assign n2556 = n2555 ^ x188 ;
  assign n2557 = n2556 ^ n2552 ;
  assign n2558 = n1161 & n2557 ;
  assign n2559 = n2558 ^ n2555 ;
  assign n2560 = ~n2554 & ~n2559 ;
  assign n2564 = n2563 ^ n2560 ;
  assign n2568 = n1194 & n1829 ;
  assign n2565 = n2562 ^ x317 ;
  assign n2569 = n2568 ^ n2565 ;
  assign n2570 = ~n2564 & ~n2569 ;
  assign n2572 = n2571 ^ n2570 ;
  assign n2573 = n1906 ^ x62 ;
  assign n2574 = n2573 ^ x190 ;
  assign n2575 = n2574 ^ n1906 ;
  assign n2576 = n1161 & n2575 ;
  assign n2577 = n2576 ^ n2573 ;
  assign n2578 = ~n2572 & ~n2577 ;
  assign n1902 = n1509 & n1829 ;
  assign n1903 = n1902 ^ x319 ;
  assign n1907 = n1906 ^ n1903 ;
  assign n2579 = n2578 ^ n1907 ;
  assign n2581 = n518 & n1161 ;
  assign n2580 = n1903 ^ x63 ;
  assign n2582 = n2581 ^ n2580 ;
  assign n2583 = n2579 & ~n2582 ;
  assign n1899 = n1187 & n1829 ;
  assign n1900 = n1899 ^ x320 ;
  assign n1904 = n1903 ^ n1900 ;
  assign n2584 = n2583 ^ n1904 ;
  assign n2585 = n1900 ^ x64 ;
  assign n2586 = n2585 ^ x192 ;
  assign n2587 = n2586 ^ n1900 ;
  assign n2588 = n1161 & n2587 ;
  assign n2589 = n2588 ^ n2585 ;
  assign n2590 = n2584 & ~n2589 ;
  assign n1896 = n1829 & n1895 ;
  assign n1897 = n1896 ^ x321 ;
  assign n1901 = n1900 ^ n1897 ;
  assign n2591 = n2590 ^ n1901 ;
  assign n2592 = n1897 ^ x65 ;
  assign n2593 = n2592 ^ x193 ;
  assign n2594 = n2593 ^ n1897 ;
  assign n2595 = n1161 & n2594 ;
  assign n2596 = n2595 ^ n2592 ;
  assign n2597 = n2591 & ~n2596 ;
  assign n1890 = n1183 & n1829 ;
  assign n1891 = n1890 ^ x322 ;
  assign n1898 = n1897 ^ n1891 ;
  assign n2598 = n2597 ^ n1898 ;
  assign n2599 = n1891 ^ x66 ;
  assign n2600 = n2599 ^ x194 ;
  assign n2601 = n2600 ^ n1891 ;
  assign n2602 = n1161 & n2601 ;
  assign n2603 = n2602 ^ n2599 ;
  assign n2604 = n2598 & ~n2603 ;
  assign n1894 = n1893 ^ n1891 ;
  assign n2605 = n2604 ^ n1894 ;
  assign n2606 = n1893 ^ x67 ;
  assign n2607 = n2606 ^ x195 ;
  assign n2608 = n2607 ^ n1893 ;
  assign n2609 = n1161 & n2608 ;
  assign n2610 = n2609 ^ n2606 ;
  assign n2611 = n2605 & ~n2610 ;
  assign n2615 = n2614 ^ n2611 ;
  assign n2619 = n1178 & n1829 ;
  assign n2616 = n2613 ^ x324 ;
  assign n2620 = n2619 ^ n2616 ;
  assign n2621 = ~n2615 & ~n2620 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2624 = n1888 ^ x69 ;
  assign n2625 = n2624 ^ x197 ;
  assign n2626 = n2625 ^ n1888 ;
  assign n2627 = n1161 & n2626 ;
  assign n2628 = n2627 ^ n2624 ;
  assign n2629 = ~n2623 & ~n2628 ;
  assign n1884 = n1172 & n1829 ;
  assign n1885 = n1884 ^ x326 ;
  assign n1889 = n1888 ^ n1885 ;
  assign n2630 = n2629 ^ n1889 ;
  assign n2631 = n1885 ^ x70 ;
  assign n2632 = n2631 ^ x198 ;
  assign n2633 = n2632 ^ n1885 ;
  assign n2634 = n1161 & n2633 ;
  assign n2635 = n2634 ^ n2631 ;
  assign n2636 = n2630 & ~n2635 ;
  assign n1878 = n1169 & n1829 ;
  assign n1879 = n1878 ^ x327 ;
  assign n1886 = n1885 ^ n1879 ;
  assign n2637 = n2636 ^ n1886 ;
  assign n2638 = n1879 ^ x71 ;
  assign n2639 = n2638 ^ x199 ;
  assign n2640 = n2639 ^ n1879 ;
  assign n2641 = n1161 & n2640 ;
  assign n2642 = n2641 ^ n2638 ;
  assign n2643 = n2637 & ~n2642 ;
  assign n1883 = n1882 ^ n1879 ;
  assign n2644 = n2643 ^ n1883 ;
  assign n2645 = n1882 ^ x72 ;
  assign n2646 = n2645 ^ x200 ;
  assign n2647 = n2646 ^ n1882 ;
  assign n2648 = n1161 & n2647 ;
  assign n2649 = n2648 ^ n2645 ;
  assign n2650 = n2644 & ~n2649 ;
  assign n2655 = n2654 ^ n2650 ;
  assign n2656 = n2653 ^ x329 ;
  assign n2657 = n2656 ^ x457 ;
  assign n2658 = n2657 ^ n2653 ;
  assign n2659 = n1829 & n2658 ;
  assign n2660 = n2659 ^ n2656 ;
  assign n2661 = ~n2655 & ~n2660 ;
  assign n2666 = n2665 ^ n2661 ;
  assign n2667 = n2664 ^ x330 ;
  assign n2668 = n2667 ^ x458 ;
  assign n2669 = n2668 ^ n2664 ;
  assign n2670 = n1829 & n2669 ;
  assign n2671 = n2670 ^ n2667 ;
  assign n2672 = n2666 & ~n2671 ;
  assign n2677 = n2676 ^ n2672 ;
  assign n2678 = n2675 ^ x75 ;
  assign n2679 = n2678 ^ x203 ;
  assign n2680 = n2679 ^ n2675 ;
  assign n2681 = n1161 & n2680 ;
  assign n2682 = n2681 ^ n2678 ;
  assign n2683 = ~n2677 & ~n2682 ;
  assign n2688 = n2687 ^ n2683 ;
  assign n2689 = n2686 ^ x332 ;
  assign n2690 = n2689 ^ x460 ;
  assign n2691 = n2690 ^ n2686 ;
  assign n2692 = n1829 & n2691 ;
  assign n2693 = n2692 ^ n2689 ;
  assign n2694 = ~n2688 & ~n2693 ;
  assign n2699 = n2698 ^ n2694 ;
  assign n2700 = n2697 ^ x333 ;
  assign n2701 = n2700 ^ x461 ;
  assign n2702 = n2701 ^ n2697 ;
  assign n2703 = n1829 & n2702 ;
  assign n2704 = n2703 ^ n2700 ;
  assign n2705 = n2699 & ~n2704 ;
  assign n2710 = n2709 ^ n2705 ;
  assign n2711 = n2708 ^ x334 ;
  assign n2712 = n2711 ^ x462 ;
  assign n2713 = n2712 ^ n2708 ;
  assign n2714 = n1829 & n2713 ;
  assign n2715 = n2714 ^ n2711 ;
  assign n2716 = n2710 & ~n2715 ;
  assign n2721 = n2720 ^ n2716 ;
  assign n2722 = n2719 ^ x335 ;
  assign n2723 = n2722 ^ x463 ;
  assign n2724 = n2723 ^ n2719 ;
  assign n2725 = n1829 & n2724 ;
  assign n2726 = n2725 ^ n2722 ;
  assign n2727 = n2721 & ~n2726 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2730 = n1873 ^ x80 ;
  assign n2731 = n2730 ^ x208 ;
  assign n2732 = n2731 ^ n1873 ;
  assign n2733 = n1161 & n2732 ;
  assign n2734 = n2733 ^ n2730 ;
  assign n2735 = ~n2729 & ~n2734 ;
  assign n1877 = n1876 ^ n1873 ;
  assign n2736 = n2735 ^ n1877 ;
  assign n2737 = n1876 ^ x81 ;
  assign n2738 = n2737 ^ x209 ;
  assign n2739 = n2738 ^ n1876 ;
  assign n2740 = n1161 & n2739 ;
  assign n2741 = n2740 ^ n2737 ;
  assign n2742 = n2736 & ~n2741 ;
  assign n2747 = n2746 ^ n2742 ;
  assign n2748 = n2745 ^ x82 ;
  assign n2749 = n2748 ^ x210 ;
  assign n2750 = n2749 ^ n2745 ;
  assign n2751 = n1161 & n2750 ;
  assign n2752 = n2751 ^ n2748 ;
  assign n2753 = n2747 & ~n2752 ;
  assign n2758 = n2757 ^ n2753 ;
  assign n2759 = n2756 ^ x339 ;
  assign n2760 = n2759 ^ x467 ;
  assign n2761 = n2760 ^ n2756 ;
  assign n2762 = n1829 & n2761 ;
  assign n2763 = n2762 ^ n2759 ;
  assign n2764 = ~n2758 & ~n2763 ;
  assign n2769 = n2768 ^ n2764 ;
  assign n2770 = n2767 ^ x340 ;
  assign n2771 = n2770 ^ x468 ;
  assign n2772 = n2771 ^ n2767 ;
  assign n2773 = n1829 & n2772 ;
  assign n2774 = n2773 ^ n2770 ;
  assign n2775 = n2769 & ~n2774 ;
  assign n2780 = n2779 ^ n2775 ;
  assign n2781 = n2778 ^ x341 ;
  assign n2782 = n2781 ^ x469 ;
  assign n2783 = n2782 ^ n2778 ;
  assign n2784 = n1829 & n2783 ;
  assign n2785 = n2784 ^ n2781 ;
  assign n2786 = n2780 & ~n2785 ;
  assign n2791 = n2790 ^ n2786 ;
  assign n2792 = n2789 ^ x342 ;
  assign n2793 = n2792 ^ x470 ;
  assign n2794 = n2793 ^ n2789 ;
  assign n2795 = n1829 & n2794 ;
  assign n2796 = n2795 ^ n2792 ;
  assign n2797 = n2791 & ~n2796 ;
  assign n2802 = n2801 ^ n2797 ;
  assign n2803 = n2800 ^ x343 ;
  assign n2804 = n2803 ^ x471 ;
  assign n2805 = n2804 ^ n2800 ;
  assign n2806 = n1829 & n2805 ;
  assign n2807 = n2806 ^ n2803 ;
  assign n2808 = n2802 & ~n2807 ;
  assign n2813 = n2812 ^ n2808 ;
  assign n2814 = n2811 ^ x88 ;
  assign n2815 = n2814 ^ x216 ;
  assign n2816 = n2815 ^ n2811 ;
  assign n2817 = n1161 & n2816 ;
  assign n2818 = n2817 ^ n2814 ;
  assign n2819 = ~n2813 & ~n2818 ;
  assign n2824 = n2823 ^ n2819 ;
  assign n2825 = n2822 ^ x89 ;
  assign n2826 = n2825 ^ x217 ;
  assign n2827 = n2826 ^ n2822 ;
  assign n2828 = n1161 & n2827 ;
  assign n2829 = n2828 ^ n2825 ;
  assign n2830 = n2824 & ~n2829 ;
  assign n2835 = n2834 ^ n2830 ;
  assign n2836 = n2833 ^ x90 ;
  assign n2837 = n2836 ^ x218 ;
  assign n2838 = n2837 ^ n2833 ;
  assign n2839 = n1161 & n2838 ;
  assign n2840 = n2839 ^ n2836 ;
  assign n2841 = n2835 & ~n2840 ;
  assign n2846 = n2845 ^ n2841 ;
  assign n2847 = n2844 ^ x347 ;
  assign n2848 = n2847 ^ x475 ;
  assign n2849 = n2848 ^ n2844 ;
  assign n2850 = n1829 & n2849 ;
  assign n2851 = n2850 ^ n2847 ;
  assign n2852 = ~n2846 & ~n2851 ;
  assign n2857 = n2856 ^ n2852 ;
  assign n2858 = n2855 ^ x348 ;
  assign n2859 = n2858 ^ x476 ;
  assign n2860 = n2859 ^ n2855 ;
  assign n2861 = n1829 & n2860 ;
  assign n2862 = n2861 ^ n2858 ;
  assign n2863 = n2857 & ~n2862 ;
  assign n2868 = n2867 ^ n2863 ;
  assign n2869 = n2866 ^ x349 ;
  assign n2870 = n2869 ^ x477 ;
  assign n2871 = n2870 ^ n2866 ;
  assign n2872 = n1829 & n2871 ;
  assign n2873 = n2872 ^ n2869 ;
  assign n2874 = n2868 & ~n2873 ;
  assign n2879 = n2878 ^ n2874 ;
  assign n2880 = n2877 ^ x94 ;
  assign n2881 = n2880 ^ x222 ;
  assign n2882 = n2881 ^ n2877 ;
  assign n2883 = n1161 & n2882 ;
  assign n2884 = n2883 ^ n2880 ;
  assign n2885 = ~n2879 & ~n2884 ;
  assign n2890 = n2889 ^ n2885 ;
  assign n2891 = n2888 ^ x95 ;
  assign n2892 = n2891 ^ x223 ;
  assign n2893 = n2892 ^ n2888 ;
  assign n2894 = n1161 & n2893 ;
  assign n2895 = n2894 ^ n2891 ;
  assign n2896 = n2890 & ~n2895 ;
  assign n2898 = n2897 ^ n2896 ;
  assign n2899 = n1866 ^ x96 ;
  assign n2900 = n2899 ^ x224 ;
  assign n2901 = n2900 ^ n1866 ;
  assign n2902 = n1161 & n2901 ;
  assign n2903 = n2902 ^ n2899 ;
  assign n2904 = n2898 & ~n2903 ;
  assign n1870 = n1869 ^ n1866 ;
  assign n2905 = n2904 ^ n1870 ;
  assign n2906 = n1869 ^ x97 ;
  assign n2907 = n2906 ^ x225 ;
  assign n2908 = n2907 ^ n1869 ;
  assign n2909 = n1161 & n2908 ;
  assign n2910 = n2909 ^ n2906 ;
  assign n2911 = n2905 & ~n2910 ;
  assign n2916 = n2915 ^ n2911 ;
  assign n2917 = n2914 ^ x98 ;
  assign n2918 = n2917 ^ x226 ;
  assign n2919 = n2918 ^ n2914 ;
  assign n2920 = n1161 & n2919 ;
  assign n2921 = n2920 ^ n2917 ;
  assign n2922 = n2916 & ~n2921 ;
  assign n2927 = n2926 ^ n2922 ;
  assign n2928 = n2925 ^ x99 ;
  assign n2929 = n2928 ^ x227 ;
  assign n2930 = n2929 ^ n2925 ;
  assign n2931 = n1161 & n2930 ;
  assign n2932 = n2931 ^ n2928 ;
  assign n2933 = n2927 & ~n2932 ;
  assign n2935 = n2934 ^ n2933 ;
  assign n2936 = n1859 ^ x100 ;
  assign n2937 = n2936 ^ x228 ;
  assign n2938 = n2937 ^ n1859 ;
  assign n2939 = n1161 & n2938 ;
  assign n2940 = n2939 ^ n2936 ;
  assign n2941 = n2935 & ~n2940 ;
  assign n1863 = n1862 ^ n1859 ;
  assign n2942 = n2941 ^ n1863 ;
  assign n2943 = n1862 ^ x101 ;
  assign n2944 = n2943 ^ x229 ;
  assign n2945 = n2944 ^ n1862 ;
  assign n2946 = n1161 & n2945 ;
  assign n2947 = n2946 ^ n2943 ;
  assign n2948 = n2942 & ~n2947 ;
  assign n2953 = n2952 ^ n2948 ;
  assign n2954 = n2951 ^ x102 ;
  assign n2955 = n2954 ^ x230 ;
  assign n2956 = n2955 ^ n2951 ;
  assign n2957 = n1161 & n2956 ;
  assign n2958 = n2957 ^ n2954 ;
  assign n2959 = n2953 & ~n2958 ;
  assign n2964 = n2963 ^ n2959 ;
  assign n2965 = n2962 ^ x359 ;
  assign n2966 = n2965 ^ x487 ;
  assign n2967 = n2966 ^ n2962 ;
  assign n2968 = n1829 & n2967 ;
  assign n2969 = n2968 ^ n2965 ;
  assign n2970 = ~n2964 & ~n2969 ;
  assign n2975 = n2974 ^ n2970 ;
  assign n2976 = n2973 ^ x104 ;
  assign n2977 = n2976 ^ x232 ;
  assign n2978 = n2977 ^ n2973 ;
  assign n2979 = n1161 & n2978 ;
  assign n2980 = n2979 ^ n2976 ;
  assign n2981 = ~n2975 & ~n2980 ;
  assign n2986 = n2985 ^ n2981 ;
  assign n2987 = n2984 ^ x105 ;
  assign n2988 = n2987 ^ x233 ;
  assign n2989 = n2988 ^ n2984 ;
  assign n2990 = n1161 & n2989 ;
  assign n2991 = n2990 ^ n2987 ;
  assign n2992 = n2986 & ~n2991 ;
  assign n2997 = n2996 ^ n2992 ;
  assign n2998 = n2995 ^ x362 ;
  assign n2999 = n2998 ^ x490 ;
  assign n3000 = n2999 ^ n2995 ;
  assign n3001 = n1829 & n3000 ;
  assign n3002 = n3001 ^ n2998 ;
  assign n3003 = ~n2997 & ~n3002 ;
  assign n3008 = n3007 ^ n3003 ;
  assign n3009 = n3006 ^ x363 ;
  assign n3010 = n3009 ^ x491 ;
  assign n3011 = n3010 ^ n3006 ;
  assign n3012 = n1829 & n3011 ;
  assign n3013 = n3012 ^ n3009 ;
  assign n3014 = n3008 & ~n3013 ;
  assign n3016 = n3015 ^ n3014 ;
  assign n3017 = n1855 ^ x108 ;
  assign n3018 = n3017 ^ x236 ;
  assign n3019 = n3018 ^ n1855 ;
  assign n3020 = n1161 & n3019 ;
  assign n3021 = n3020 ^ n3017 ;
  assign n3022 = ~n3016 & ~n3021 ;
  assign n1847 = n1829 & n1846 ;
  assign n1848 = n1847 ^ x365 ;
  assign n1856 = n1855 ^ n1848 ;
  assign n3023 = n3022 ^ n1856 ;
  assign n3024 = n1848 ^ x109 ;
  assign n3025 = n3024 ^ x237 ;
  assign n3026 = n3025 ^ n1848 ;
  assign n3027 = n1161 & n3026 ;
  assign n3028 = n3027 ^ n3024 ;
  assign n3029 = n3023 & ~n3028 ;
  assign n1852 = n1851 ^ n1848 ;
  assign n3030 = n3029 ^ n1852 ;
  assign n3031 = n1851 ^ x110 ;
  assign n3032 = n3031 ^ x238 ;
  assign n3033 = n3032 ^ n1851 ;
  assign n3034 = n1161 & n3033 ;
  assign n3035 = n3034 ^ n3031 ;
  assign n3036 = n3030 & ~n3035 ;
  assign n3041 = n3040 ^ n3036 ;
  assign n3042 = n3039 ^ x111 ;
  assign n3043 = n3042 ^ x239 ;
  assign n3044 = n3043 ^ n3039 ;
  assign n3045 = n1161 & n3044 ;
  assign n3046 = n3045 ^ n3042 ;
  assign n3047 = n3041 & ~n3046 ;
  assign n3052 = n3051 ^ n3047 ;
  assign n3053 = n3050 ^ x112 ;
  assign n3054 = n3053 ^ x240 ;
  assign n3055 = n3054 ^ n3050 ;
  assign n3056 = n1161 & n3055 ;
  assign n3057 = n3056 ^ n3053 ;
  assign n3058 = n3052 & ~n3057 ;
  assign n3063 = n3062 ^ n3058 ;
  assign n3064 = n3061 ^ x369 ;
  assign n3065 = n3064 ^ x497 ;
  assign n3066 = n3065 ^ n3061 ;
  assign n3067 = n1829 & n3066 ;
  assign n3068 = n3067 ^ n3064 ;
  assign n3069 = ~n3063 & ~n3068 ;
  assign n3074 = n3073 ^ n3069 ;
  assign n3075 = n3072 ^ x114 ;
  assign n3076 = n3075 ^ x242 ;
  assign n3077 = n3076 ^ n3072 ;
  assign n3078 = n1161 & n3077 ;
  assign n3079 = n3078 ^ n3075 ;
  assign n3080 = ~n3074 & ~n3079 ;
  assign n3085 = n3084 ^ n3080 ;
  assign n3086 = n3083 ^ x115 ;
  assign n3087 = n3086 ^ x243 ;
  assign n3088 = n3087 ^ n3083 ;
  assign n3089 = n1161 & n3088 ;
  assign n3090 = n3089 ^ n3086 ;
  assign n3091 = n3085 & ~n3090 ;
  assign n3096 = n3095 ^ n3091 ;
  assign n3097 = n3094 ^ x372 ;
  assign n3098 = n3097 ^ x500 ;
  assign n3099 = n3098 ^ n3094 ;
  assign n3100 = n1829 & n3099 ;
  assign n3101 = n3100 ^ n3097 ;
  assign n3102 = ~n3096 & ~n3101 ;
  assign n3107 = n3106 ^ n3102 ;
  assign n3108 = n3105 ^ x373 ;
  assign n3109 = n3108 ^ x501 ;
  assign n3110 = n3109 ^ n3105 ;
  assign n3111 = n1829 & n3110 ;
  assign n3112 = n3111 ^ n3108 ;
  assign n3113 = n3107 & ~n3112 ;
  assign n3118 = n3117 ^ n3113 ;
  assign n3119 = n3116 ^ x374 ;
  assign n3120 = n3119 ^ x502 ;
  assign n3121 = n3120 ^ n3116 ;
  assign n3122 = n1829 & n3121 ;
  assign n3123 = n3122 ^ n3119 ;
  assign n3124 = n3118 & ~n3123 ;
  assign n3129 = n3128 ^ n3124 ;
  assign n3130 = n3127 ^ x375 ;
  assign n3131 = n3130 ^ x503 ;
  assign n3132 = n3131 ^ n3127 ;
  assign n3133 = n1829 & n3132 ;
  assign n3134 = n3133 ^ n3130 ;
  assign n3135 = n3129 & ~n3134 ;
  assign n3137 = n3136 ^ n3135 ;
  assign n3138 = n1841 ^ x120 ;
  assign n3139 = n3138 ^ x248 ;
  assign n3140 = n3139 ^ n1841 ;
  assign n3141 = n1161 & n3140 ;
  assign n3142 = n3141 ^ n3138 ;
  assign n3143 = ~n3137 & ~n3142 ;
  assign n1845 = n1844 ^ n1841 ;
  assign n3144 = n3143 ^ n1845 ;
  assign n3145 = n1844 ^ x121 ;
  assign n3146 = n3145 ^ x249 ;
  assign n3147 = n3146 ^ n1844 ;
  assign n3148 = n1161 & n3147 ;
  assign n3149 = n3148 ^ n3145 ;
  assign n3150 = n3144 & ~n3149 ;
  assign n3154 = n3153 ^ n3150 ;
  assign n3155 = n3152 ^ x378 ;
  assign n3156 = n3155 ^ x506 ;
  assign n3157 = n3156 ^ n3152 ;
  assign n3158 = n1829 & n3157 ;
  assign n3159 = n3158 ^ n3155 ;
  assign n3160 = ~n3154 & ~n3159 ;
  assign n3164 = n3163 ^ n3160 ;
  assign n3165 = n3162 ^ x123 ;
  assign n3166 = n3165 ^ x251 ;
  assign n3167 = n3166 ^ n3162 ;
  assign n3168 = n1161 & n3167 ;
  assign n3169 = n3168 ^ n3165 ;
  assign n3170 = ~n3164 & ~n3169 ;
  assign n3174 = n3173 ^ n3170 ;
  assign n3175 = n3172 ^ x124 ;
  assign n3176 = n3175 ^ x252 ;
  assign n3177 = n3176 ^ n3172 ;
  assign n3178 = n1161 & n3177 ;
  assign n3179 = n3178 ^ n3175 ;
  assign n3180 = n3174 & ~n3179 ;
  assign n3184 = n3183 ^ n3180 ;
  assign n3188 = n1167 & n1829 ;
  assign n3185 = n3182 ^ x381 ;
  assign n3189 = n3188 ^ n3185 ;
  assign n3190 = ~n3184 & ~n3189 ;
  assign n3192 = n3191 ^ n3190 ;
  assign n3193 = n1837 ^ x382 ;
  assign n3194 = n3193 ^ x510 ;
  assign n3195 = n3194 ^ n1837 ;
  assign n3196 = n1829 & n3195 ;
  assign n3197 = n3196 ^ n3193 ;
  assign n3198 = n3192 & ~n3197 ;
  assign n1838 = n1837 ^ n1834 ;
  assign n3199 = n3198 ^ n1838 ;
  assign n3200 = ~n1835 & n3199 ;
  assign n3201 = n3200 ^ n1834 ;
  assign n3202 = n1832 & n3201 ;
  assign n3203 = n3202 ^ n1831 ;
  assign n3204 = n2000 & ~n3201 ;
  assign n3205 = n3204 ^ n1999 ;
  assign n3206 = n2017 & ~n3201 ;
  assign n3207 = n3206 ^ n2010 ;
  assign n3208 = n2028 & ~n3201 ;
  assign n3209 = n3208 ^ n2021 ;
  assign n3210 = n2036 & n3201 ;
  assign n3211 = n3210 ^ n1989 ;
  assign n3212 = n2043 & n3201 ;
  assign n3213 = n3212 ^ n1992 ;
  assign n3214 = n2054 & ~n3201 ;
  assign n3215 = n3214 ^ n2047 ;
  assign n3216 = n2065 & n3201 ;
  assign n3217 = n3216 ^ n2058 ;
  assign n3218 = n2076 & ~n3201 ;
  assign n3219 = n3218 ^ n2069 ;
  assign n3220 = n2087 & ~n3201 ;
  assign n3221 = n3220 ^ n2080 ;
  assign n3222 = n2095 & n3201 ;
  assign n3223 = n3222 ^ n1985 ;
  assign n3224 = n2102 & n3201 ;
  assign n3225 = n3224 ^ n1978 ;
  assign n3226 = n2109 & n3201 ;
  assign n3227 = n3226 ^ n1981 ;
  assign n3228 = n2120 & ~n3201 ;
  assign n3229 = n3228 ^ n2113 ;
  assign n3230 = n2131 & ~n3201 ;
  assign n3231 = n3230 ^ n2124 ;
  assign n3232 = n2142 & n3201 ;
  assign n3233 = n3232 ^ n2135 ;
  assign n3234 = n2153 & ~n3201 ;
  assign n3235 = n3234 ^ n2146 ;
  assign n3236 = n2161 & n3201 ;
  assign n3237 = n3236 ^ n1971 ;
  assign n3238 = n2168 & n3201 ;
  assign n3239 = n3238 ^ n1974 ;
  assign n3240 = n2179 & ~n3201 ;
  assign n3241 = n3240 ^ n2172 ;
  assign n3242 = n2190 & n3201 ;
  assign n3243 = n3242 ^ n2183 ;
  assign n3244 = n2201 & ~n3201 ;
  assign n3245 = n3244 ^ n2194 ;
  assign n3246 = n2212 & ~n3201 ;
  assign n3247 = n3246 ^ n2205 ;
  assign n3248 = n2223 & ~n3201 ;
  assign n3249 = n3248 ^ n2216 ;
  assign n3250 = n2231 & n3201 ;
  assign n3251 = n3250 ^ n1967 ;
  assign n3252 = n2238 & n3201 ;
  assign n3253 = n3252 ^ n1960 ;
  assign n3254 = n2245 & n3201 ;
  assign n3255 = n3254 ^ n1963 ;
  assign n3256 = n2256 & ~n3201 ;
  assign n3257 = n3256 ^ n2249 ;
  assign n3258 = n2264 & n3201 ;
  assign n3259 = n3258 ^ n1953 ;
  assign n3260 = n2271 & n3201 ;
  assign n3261 = n3260 ^ n1956 ;
  assign n3262 = n2282 & ~n3201 ;
  assign n3263 = n3262 ^ n2275 ;
  assign n3264 = n2290 & n3201 ;
  assign n3265 = n3264 ^ n1949 ;
  assign n3266 = n2297 & n3201 ;
  assign n3267 = n3266 ^ n1942 ;
  assign n3268 = n2304 & n3201 ;
  assign n3269 = n3268 ^ n1945 ;
  assign n3270 = n2315 & ~n3201 ;
  assign n3271 = n3270 ^ n2308 ;
  assign n3272 = n2323 & n3201 ;
  assign n3273 = n3272 ^ n1935 ;
  assign n3274 = n2330 & n3201 ;
  assign n3275 = n3274 ^ n1938 ;
  assign n3276 = n2341 & ~n3201 ;
  assign n3277 = n3276 ^ n2334 ;
  assign n3278 = n2349 & n3201 ;
  assign n3279 = n3278 ^ n1931 ;
  assign n3280 = n2356 & n3201 ;
  assign n3281 = n3280 ^ n1928 ;
  assign n3282 = n2363 & n3201 ;
  assign n3283 = n3282 ^ n1925 ;
  assign n3284 = n2370 & n3201 ;
  assign n3285 = n3284 ^ n1920 ;
  assign n3286 = n2377 & n3201 ;
  assign n3287 = n3286 ^ n1922 ;
  assign n3288 = n2387 & ~n3201 ;
  assign n3289 = n3288 ^ n2380 ;
  assign n3290 = n2397 & ~n3201 ;
  assign n3291 = n3290 ^ n2390 ;
  assign n3292 = n2405 & n3201 ;
  assign n3293 = n3292 ^ n1917 ;
  assign n3294 = n2412 & n3201 ;
  assign n3295 = n3294 ^ n1910 ;
  assign n3296 = n2419 & n3201 ;
  assign n3297 = n3296 ^ n1913 ;
  assign n3298 = n2430 & ~n3201 ;
  assign n3299 = n3298 ^ n2423 ;
  assign n3300 = n2441 & n3201 ;
  assign n3301 = n3300 ^ n2434 ;
  assign n3302 = n2452 & ~n3201 ;
  assign n3303 = n3302 ^ n2445 ;
  assign n3304 = n2463 & ~n3201 ;
  assign n3305 = n3304 ^ n2456 ;
  assign n3306 = n2474 & n3201 ;
  assign n3307 = n3306 ^ n2467 ;
  assign n3308 = n2485 & ~n3201 ;
  assign n3309 = n3308 ^ n2478 ;
  assign n3310 = n2496 & n3201 ;
  assign n3311 = n3310 ^ n2489 ;
  assign n3312 = n2507 & ~n3201 ;
  assign n3313 = n3312 ^ n2500 ;
  assign n3314 = n2518 & n3201 ;
  assign n3315 = n3314 ^ n2511 ;
  assign n3316 = n2529 & ~n3201 ;
  assign n3317 = n3316 ^ n2522 ;
  assign n3318 = n2539 & ~n3201 ;
  assign n3319 = n3318 ^ n2532 ;
  assign n3320 = n2549 & ~n3201 ;
  assign n3321 = n3320 ^ n2542 ;
  assign n3322 = n2559 & n3201 ;
  assign n3323 = n3322 ^ n2552 ;
  assign n3324 = n2569 & ~n3201 ;
  assign n3325 = n3324 ^ n2562 ;
  assign n3326 = n2577 & n3201 ;
  assign n3327 = n3326 ^ n1906 ;
  assign n3328 = n2582 & n3201 ;
  assign n3329 = n3328 ^ n1903 ;
  assign n3330 = n2589 & n3201 ;
  assign n3331 = n3330 ^ n1900 ;
  assign n3332 = n2596 & n3201 ;
  assign n3333 = n3332 ^ n1897 ;
  assign n3334 = n2603 & n3201 ;
  assign n3335 = n3334 ^ n1891 ;
  assign n3336 = n2610 & n3201 ;
  assign n3337 = n3336 ^ n1893 ;
  assign n3338 = n2620 & ~n3201 ;
  assign n3339 = n3338 ^ n2613 ;
  assign n3340 = n2628 & n3201 ;
  assign n3341 = n3340 ^ n1888 ;
  assign n3342 = n2635 & n3201 ;
  assign n3343 = n3342 ^ n1885 ;
  assign n3344 = n2642 & n3201 ;
  assign n3345 = n3344 ^ n1879 ;
  assign n3346 = n2649 & n3201 ;
  assign n3347 = n3346 ^ n1882 ;
  assign n3348 = n2660 & ~n3201 ;
  assign n3349 = n3348 ^ n2653 ;
  assign n3350 = n2671 & ~n3201 ;
  assign n3351 = n3350 ^ n2664 ;
  assign n3352 = n2682 & n3201 ;
  assign n3353 = n3352 ^ n2675 ;
  assign n3354 = n2693 & ~n3201 ;
  assign n3355 = n3354 ^ n2686 ;
  assign n3356 = n2704 & ~n3201 ;
  assign n3357 = n3356 ^ n2697 ;
  assign n3358 = n2715 & ~n3201 ;
  assign n3359 = n3358 ^ n2708 ;
  assign n3360 = n2726 & ~n3201 ;
  assign n3361 = n3360 ^ n2719 ;
  assign n3362 = n2734 & n3201 ;
  assign n3363 = n3362 ^ n1873 ;
  assign n3364 = n2741 & n3201 ;
  assign n3365 = n3364 ^ n1876 ;
  assign n3366 = n2752 & n3201 ;
  assign n3367 = n3366 ^ n2745 ;
  assign n3368 = n2763 & ~n3201 ;
  assign n3369 = n3368 ^ n2756 ;
  assign n3370 = n2774 & ~n3201 ;
  assign n3371 = n3370 ^ n2767 ;
  assign n3372 = n2785 & ~n3201 ;
  assign n3373 = n3372 ^ n2778 ;
  assign n3374 = n2796 & ~n3201 ;
  assign n3375 = n3374 ^ n2789 ;
  assign n3376 = n2807 & ~n3201 ;
  assign n3377 = n3376 ^ n2800 ;
  assign n3378 = n2818 & n3201 ;
  assign n3379 = n3378 ^ n2811 ;
  assign n3380 = n2829 & n3201 ;
  assign n3381 = n3380 ^ n2822 ;
  assign n3382 = n2840 & n3201 ;
  assign n3383 = n3382 ^ n2833 ;
  assign n3384 = n2851 & ~n3201 ;
  assign n3385 = n3384 ^ n2844 ;
  assign n3386 = n2862 & ~n3201 ;
  assign n3387 = n3386 ^ n2855 ;
  assign n3388 = n2873 & ~n3201 ;
  assign n3389 = n3388 ^ n2866 ;
  assign n3390 = n2884 & n3201 ;
  assign n3391 = n3390 ^ n2877 ;
  assign n3392 = n2895 & n3201 ;
  assign n3393 = n3392 ^ n2888 ;
  assign n3394 = n2903 & n3201 ;
  assign n3395 = n3394 ^ n1866 ;
  assign n3396 = n2910 & n3201 ;
  assign n3397 = n3396 ^ n1869 ;
  assign n3398 = n2921 & n3201 ;
  assign n3399 = n3398 ^ n2914 ;
  assign n3400 = n2932 & n3201 ;
  assign n3401 = n3400 ^ n2925 ;
  assign n3402 = n2940 & n3201 ;
  assign n3403 = n3402 ^ n1859 ;
  assign n3404 = n2947 & n3201 ;
  assign n3405 = n3404 ^ n1862 ;
  assign n3406 = n2958 & n3201 ;
  assign n3407 = n3406 ^ n2951 ;
  assign n3408 = n2969 & ~n3201 ;
  assign n3409 = n3408 ^ n2962 ;
  assign n3410 = n2980 & n3201 ;
  assign n3411 = n3410 ^ n2973 ;
  assign n3412 = n2991 & n3201 ;
  assign n3413 = n3412 ^ n2984 ;
  assign n3414 = n3002 & ~n3201 ;
  assign n3415 = n3414 ^ n2995 ;
  assign n3416 = n3013 & ~n3201 ;
  assign n3417 = n3416 ^ n3006 ;
  assign n3418 = n3021 & n3201 ;
  assign n3419 = n3418 ^ n1855 ;
  assign n3420 = n3028 & n3201 ;
  assign n3421 = n3420 ^ n1848 ;
  assign n3422 = n3035 & n3201 ;
  assign n3423 = n3422 ^ n1851 ;
  assign n3424 = n3046 & n3201 ;
  assign n3425 = n3424 ^ n3039 ;
  assign n3426 = n3057 & n3201 ;
  assign n3427 = n3426 ^ n3050 ;
  assign n3428 = n3068 & ~n3201 ;
  assign n3429 = n3428 ^ n3061 ;
  assign n3430 = n3079 & n3201 ;
  assign n3431 = n3430 ^ n3072 ;
  assign n3432 = n3090 & n3201 ;
  assign n3433 = n3432 ^ n3083 ;
  assign n3434 = n3101 & ~n3201 ;
  assign n3435 = n3434 ^ n3094 ;
  assign n3436 = n3112 & ~n3201 ;
  assign n3437 = n3436 ^ n3105 ;
  assign n3438 = n3123 & ~n3201 ;
  assign n3439 = n3438 ^ n3116 ;
  assign n3440 = n3134 & ~n3201 ;
  assign n3441 = n3440 ^ n3127 ;
  assign n3442 = n3142 & n3201 ;
  assign n3443 = n3442 ^ n1841 ;
  assign n3444 = n3149 & n3201 ;
  assign n3445 = n3444 ^ n1844 ;
  assign n3446 = n3159 & ~n3201 ;
  assign n3447 = n3446 ^ n3152 ;
  assign n3448 = n3169 & n3201 ;
  assign n3449 = n3448 ^ n3162 ;
  assign n3450 = n3179 & n3201 ;
  assign n3451 = n3450 ^ n3172 ;
  assign n3452 = n3189 & ~n3201 ;
  assign n3453 = n3452 ^ n3182 ;
  assign n3454 = n3197 & ~n3201 ;
  assign n3455 = n3454 ^ n1837 ;
  assign n3456 = n1833 & n1834 ;
  assign n3457 = n1829 ^ n1161 ;
  assign n3458 = n3201 & n3457 ;
  assign n3459 = n3458 ^ n1829 ;
  assign y0 = n3203 ;
  assign y1 = n3205 ;
  assign y2 = n3207 ;
  assign y3 = n3209 ;
  assign y4 = n3211 ;
  assign y5 = n3213 ;
  assign y6 = n3215 ;
  assign y7 = n3217 ;
  assign y8 = n3219 ;
  assign y9 = n3221 ;
  assign y10 = n3223 ;
  assign y11 = n3225 ;
  assign y12 = n3227 ;
  assign y13 = n3229 ;
  assign y14 = n3231 ;
  assign y15 = n3233 ;
  assign y16 = n3235 ;
  assign y17 = n3237 ;
  assign y18 = n3239 ;
  assign y19 = n3241 ;
  assign y20 = n3243 ;
  assign y21 = n3245 ;
  assign y22 = n3247 ;
  assign y23 = n3249 ;
  assign y24 = n3251 ;
  assign y25 = n3253 ;
  assign y26 = n3255 ;
  assign y27 = n3257 ;
  assign y28 = n3259 ;
  assign y29 = n3261 ;
  assign y30 = n3263 ;
  assign y31 = n3265 ;
  assign y32 = n3267 ;
  assign y33 = n3269 ;
  assign y34 = n3271 ;
  assign y35 = n3273 ;
  assign y36 = n3275 ;
  assign y37 = n3277 ;
  assign y38 = n3279 ;
  assign y39 = n3281 ;
  assign y40 = n3283 ;
  assign y41 = n3285 ;
  assign y42 = n3287 ;
  assign y43 = n3289 ;
  assign y44 = n3291 ;
  assign y45 = n3293 ;
  assign y46 = n3295 ;
  assign y47 = n3297 ;
  assign y48 = n3299 ;
  assign y49 = n3301 ;
  assign y50 = n3303 ;
  assign y51 = n3305 ;
  assign y52 = n3307 ;
  assign y53 = n3309 ;
  assign y54 = n3311 ;
  assign y55 = n3313 ;
  assign y56 = n3315 ;
  assign y57 = n3317 ;
  assign y58 = n3319 ;
  assign y59 = n3321 ;
  assign y60 = n3323 ;
  assign y61 = n3325 ;
  assign y62 = n3327 ;
  assign y63 = n3329 ;
  assign y64 = n3331 ;
  assign y65 = n3333 ;
  assign y66 = n3335 ;
  assign y67 = n3337 ;
  assign y68 = n3339 ;
  assign y69 = n3341 ;
  assign y70 = n3343 ;
  assign y71 = n3345 ;
  assign y72 = n3347 ;
  assign y73 = n3349 ;
  assign y74 = n3351 ;
  assign y75 = n3353 ;
  assign y76 = n3355 ;
  assign y77 = n3357 ;
  assign y78 = n3359 ;
  assign y79 = n3361 ;
  assign y80 = n3363 ;
  assign y81 = n3365 ;
  assign y82 = n3367 ;
  assign y83 = n3369 ;
  assign y84 = n3371 ;
  assign y85 = n3373 ;
  assign y86 = n3375 ;
  assign y87 = n3377 ;
  assign y88 = n3379 ;
  assign y89 = n3381 ;
  assign y90 = n3383 ;
  assign y91 = n3385 ;
  assign y92 = n3387 ;
  assign y93 = n3389 ;
  assign y94 = n3391 ;
  assign y95 = n3393 ;
  assign y96 = n3395 ;
  assign y97 = n3397 ;
  assign y98 = n3399 ;
  assign y99 = n3401 ;
  assign y100 = n3403 ;
  assign y101 = n3405 ;
  assign y102 = n3407 ;
  assign y103 = n3409 ;
  assign y104 = n3411 ;
  assign y105 = n3413 ;
  assign y106 = n3415 ;
  assign y107 = n3417 ;
  assign y108 = n3419 ;
  assign y109 = n3421 ;
  assign y110 = n3423 ;
  assign y111 = n3425 ;
  assign y112 = n3427 ;
  assign y113 = n3429 ;
  assign y114 = n3431 ;
  assign y115 = n3433 ;
  assign y116 = n3435 ;
  assign y117 = n3437 ;
  assign y118 = n3439 ;
  assign y119 = n3441 ;
  assign y120 = n3443 ;
  assign y121 = n3445 ;
  assign y122 = n3447 ;
  assign y123 = n3449 ;
  assign y124 = n3451 ;
  assign y125 = n3453 ;
  assign y126 = n3455 ;
  assign y127 = n3456 ;
  assign y128 = n3459 ;
  assign y129 = ~n3201 ;
endmodule
