module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n467 , n468 , n469 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n610 , n611 , n612 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 ;
  assign n129 = ~x126 & ~x127 ;
  assign n130 = x127 ^ x125 ;
  assign n131 = ~x122 & ~x123 ;
  assign n132 = x123 ^ x121 ;
  assign n133 = ~x118 & ~x119 ;
  assign n134 = x119 ^ x117 ;
  assign n135 = ~x114 & ~x115 ;
  assign n136 = x115 ^ x113 ;
  assign n137 = ~x110 & ~x111 ;
  assign n138 = x111 ^ x109 ;
  assign n139 = ~x106 & ~x107 ;
  assign n140 = x107 ^ x105 ;
  assign n141 = ~x102 & ~x103 ;
  assign n142 = x103 ^ x101 ;
  assign n143 = ~x98 & ~x99 ;
  assign n144 = x99 ^ x97 ;
  assign n145 = ~x94 & ~x95 ;
  assign n146 = x95 ^ x93 ;
  assign n147 = ~x90 & ~x91 ;
  assign n148 = x91 ^ x89 ;
  assign n149 = ~x86 & ~x87 ;
  assign n150 = x87 ^ x85 ;
  assign n151 = ~x82 & ~x83 ;
  assign n152 = x83 ^ x81 ;
  assign n153 = ~x78 & ~x79 ;
  assign n154 = x79 ^ x77 ;
  assign n155 = ~x74 & ~x75 ;
  assign n156 = x75 ^ x73 ;
  assign n157 = ~x70 & ~x71 ;
  assign n158 = x71 ^ x69 ;
  assign n159 = ~x66 & ~x67 ;
  assign n160 = x67 ^ x65 ;
  assign n161 = ~x62 & ~x63 ;
  assign n162 = x63 ^ x61 ;
  assign n163 = ~x58 & ~x59 ;
  assign n164 = x59 ^ x57 ;
  assign n165 = ~x54 & ~x55 ;
  assign n166 = x55 ^ x53 ;
  assign n167 = ~x50 & ~x51 ;
  assign n168 = x51 ^ x49 ;
  assign n169 = ~x46 & ~x47 ;
  assign n170 = x47 ^ x45 ;
  assign n171 = ~x42 & ~x43 ;
  assign n172 = x43 ^ x41 ;
  assign n173 = ~x38 & ~x39 ;
  assign n174 = x39 ^ x37 ;
  assign n175 = ~x34 & ~x35 ;
  assign n176 = x35 ^ x33 ;
  assign n177 = ~x30 & ~x31 ;
  assign n178 = x31 ^ x29 ;
  assign n179 = ~x26 & ~x27 ;
  assign n180 = x27 ^ x25 ;
  assign n181 = ~x22 & ~x23 ;
  assign n182 = x23 ^ x21 ;
  assign n183 = ~x18 & ~x19 ;
  assign n184 = x19 ^ x17 ;
  assign n185 = ~x14 & ~x15 ;
  assign n186 = x15 ^ x13 ;
  assign n187 = ~x10 & ~x11 ;
  assign n188 = x11 ^ x9 ;
  assign n189 = ~x6 & ~x7 ;
  assign n190 = x7 ^ x5 ;
  assign n191 = ~x2 & ~x3 ;
  assign n196 = x1 & n191 ;
  assign n197 = n196 ^ x3 ;
  assign n198 = ~x4 & n197 ;
  assign n199 = n198 ^ n189 ;
  assign n200 = ~n190 & n199 ;
  assign n201 = n189 & ~n200 ;
  assign n202 = n201 ^ x7 ;
  assign n203 = ~x8 & n202 ;
  assign n204 = n203 ^ n187 ;
  assign n205 = ~n188 & n204 ;
  assign n206 = n187 & ~n205 ;
  assign n207 = n206 ^ x11 ;
  assign n208 = ~x12 & n207 ;
  assign n209 = n208 ^ n185 ;
  assign n210 = ~n186 & n209 ;
  assign n211 = n185 & ~n210 ;
  assign n212 = n211 ^ x15 ;
  assign n213 = ~x16 & n212 ;
  assign n214 = n213 ^ n183 ;
  assign n215 = ~n184 & n214 ;
  assign n216 = n183 & ~n215 ;
  assign n217 = n216 ^ x19 ;
  assign n218 = ~x20 & n217 ;
  assign n219 = n218 ^ n181 ;
  assign n220 = ~n182 & n219 ;
  assign n221 = n181 & ~n220 ;
  assign n222 = n221 ^ x23 ;
  assign n223 = ~x24 & n222 ;
  assign n224 = n223 ^ n179 ;
  assign n225 = ~n180 & n224 ;
  assign n226 = n179 & ~n225 ;
  assign n227 = n226 ^ x27 ;
  assign n228 = ~x28 & n227 ;
  assign n229 = n228 ^ n177 ;
  assign n230 = ~n178 & n229 ;
  assign n231 = n177 & ~n230 ;
  assign n232 = n231 ^ x31 ;
  assign n233 = ~x32 & n232 ;
  assign n234 = n233 ^ n175 ;
  assign n235 = ~n176 & n234 ;
  assign n236 = n175 & ~n235 ;
  assign n237 = n236 ^ x35 ;
  assign n238 = ~x36 & n237 ;
  assign n239 = n238 ^ n173 ;
  assign n240 = ~n174 & n239 ;
  assign n241 = n173 & ~n240 ;
  assign n242 = n241 ^ x39 ;
  assign n243 = ~x40 & n242 ;
  assign n244 = n243 ^ n171 ;
  assign n245 = ~n172 & n244 ;
  assign n246 = n171 & ~n245 ;
  assign n247 = n246 ^ x43 ;
  assign n248 = ~x44 & n247 ;
  assign n249 = n248 ^ n169 ;
  assign n250 = ~n170 & n249 ;
  assign n251 = n169 & ~n250 ;
  assign n252 = n251 ^ x47 ;
  assign n253 = ~x48 & n252 ;
  assign n254 = n253 ^ n167 ;
  assign n255 = ~n168 & n254 ;
  assign n256 = n167 & ~n255 ;
  assign n257 = n256 ^ x51 ;
  assign n258 = ~x52 & n257 ;
  assign n259 = n258 ^ n165 ;
  assign n260 = ~n166 & n259 ;
  assign n261 = n165 & ~n260 ;
  assign n262 = n261 ^ x55 ;
  assign n263 = ~x56 & n262 ;
  assign n264 = n263 ^ n163 ;
  assign n265 = ~n164 & n264 ;
  assign n266 = n163 & ~n265 ;
  assign n267 = n266 ^ x59 ;
  assign n268 = ~x60 & n267 ;
  assign n269 = n268 ^ n161 ;
  assign n270 = ~n162 & n269 ;
  assign n271 = n161 & ~n270 ;
  assign n272 = n271 ^ x63 ;
  assign n273 = ~x64 & n272 ;
  assign n274 = n273 ^ n159 ;
  assign n275 = ~n160 & n274 ;
  assign n276 = n159 & ~n275 ;
  assign n277 = n276 ^ x67 ;
  assign n278 = ~x68 & n277 ;
  assign n279 = n278 ^ n157 ;
  assign n280 = ~n158 & n279 ;
  assign n281 = n157 & ~n280 ;
  assign n282 = n281 ^ x71 ;
  assign n283 = ~x72 & n282 ;
  assign n284 = n283 ^ n155 ;
  assign n285 = ~n156 & n284 ;
  assign n286 = n155 & ~n285 ;
  assign n287 = n286 ^ x75 ;
  assign n288 = ~x76 & n287 ;
  assign n289 = n288 ^ n153 ;
  assign n290 = ~n154 & n289 ;
  assign n291 = n153 & ~n290 ;
  assign n292 = n291 ^ x79 ;
  assign n293 = ~x80 & n292 ;
  assign n294 = n293 ^ n151 ;
  assign n295 = ~n152 & n294 ;
  assign n296 = n151 & ~n295 ;
  assign n297 = n296 ^ x83 ;
  assign n298 = ~x84 & n297 ;
  assign n299 = n298 ^ n149 ;
  assign n300 = ~n150 & n299 ;
  assign n301 = n149 & ~n300 ;
  assign n302 = n301 ^ x87 ;
  assign n303 = ~x88 & n302 ;
  assign n304 = n303 ^ n147 ;
  assign n305 = ~n148 & n304 ;
  assign n306 = n147 & ~n305 ;
  assign n307 = n306 ^ x91 ;
  assign n308 = ~x92 & n307 ;
  assign n309 = n308 ^ n145 ;
  assign n310 = ~n146 & n309 ;
  assign n311 = n145 & ~n310 ;
  assign n312 = n311 ^ x95 ;
  assign n313 = ~x96 & n312 ;
  assign n314 = n313 ^ n143 ;
  assign n315 = ~n144 & n314 ;
  assign n316 = n143 & ~n315 ;
  assign n317 = n316 ^ x99 ;
  assign n318 = ~x100 & n317 ;
  assign n319 = n318 ^ n141 ;
  assign n320 = ~n142 & n319 ;
  assign n321 = n141 & ~n320 ;
  assign n322 = n321 ^ x103 ;
  assign n323 = ~x104 & n322 ;
  assign n324 = n323 ^ n139 ;
  assign n325 = ~n140 & n324 ;
  assign n326 = n139 & ~n325 ;
  assign n327 = n326 ^ x107 ;
  assign n328 = ~x108 & n327 ;
  assign n329 = n328 ^ n137 ;
  assign n330 = ~n138 & n329 ;
  assign n331 = n137 & ~n330 ;
  assign n332 = n331 ^ x111 ;
  assign n333 = ~x112 & n332 ;
  assign n334 = n333 ^ n135 ;
  assign n335 = ~n136 & n334 ;
  assign n336 = n135 & ~n335 ;
  assign n337 = n336 ^ x115 ;
  assign n338 = ~x116 & n337 ;
  assign n339 = n338 ^ n133 ;
  assign n340 = ~n134 & n339 ;
  assign n341 = n133 & ~n340 ;
  assign n342 = n341 ^ x119 ;
  assign n343 = ~x120 & n342 ;
  assign n344 = n343 ^ n131 ;
  assign n345 = ~n132 & n344 ;
  assign n346 = n131 & ~n345 ;
  assign n347 = n346 ^ x123 ;
  assign n348 = ~x124 & n347 ;
  assign n349 = n348 ^ n129 ;
  assign n350 = ~n130 & n349 ;
  assign n351 = n129 & ~n350 ;
  assign n352 = n351 ^ x127 ;
  assign n353 = ~x124 & ~x125 ;
  assign n354 = n129 & n353 ;
  assign n355 = ~x120 & ~x121 ;
  assign n356 = n131 & n355 ;
  assign n357 = ~x116 & ~x117 ;
  assign n358 = n133 & n357 ;
  assign n359 = n356 & n358 ;
  assign n360 = ~x112 & ~x113 ;
  assign n361 = n135 & n359 ;
  assign n362 = n360 & n361 ;
  assign n363 = n354 & n362 ;
  assign n364 = ~x108 & ~x109 ;
  assign n365 = n137 & n364 ;
  assign n366 = n364 ^ n139 ;
  assign n367 = ~x104 & ~x105 ;
  assign n368 = ~x100 & ~x101 ;
  assign n369 = n141 & n368 ;
  assign n370 = n368 ^ n143 ;
  assign n371 = ~x96 & ~x97 ;
  assign n372 = ~x92 & ~x93 ;
  assign n373 = n145 & n372 ;
  assign n374 = n372 ^ n147 ;
  assign n375 = ~x88 & ~x89 ;
  assign n429 = ~x80 & ~x81 ;
  assign n430 = n151 & n429 ;
  assign n431 = n147 & n373 ;
  assign n432 = n375 & n431 ;
  assign n433 = ~x84 & ~x85 ;
  assign n434 = n149 & n433 ;
  assign n435 = n432 & n434 ;
  assign n436 = n430 & n435 ;
  assign n377 = ~x76 & ~x77 ;
  assign n378 = n153 & n377 ;
  assign n379 = n377 ^ n155 ;
  assign n380 = ~x72 & ~x73 ;
  assign n381 = ~x68 & ~x69 ;
  assign n382 = n157 & n381 ;
  assign n383 = n381 ^ n159 ;
  assign n384 = n155 & n380 ;
  assign n385 = n378 & n384 ;
  assign n386 = ~x64 & ~x65 ;
  assign n387 = n159 & n386 ;
  assign n388 = n382 & n387 ;
  assign n389 = n385 & n388 ;
  assign n397 = ~x52 & ~x53 ;
  assign n390 = ~x60 & ~x61 ;
  assign n391 = n161 & n390 ;
  assign n392 = ~x56 & ~x57 ;
  assign n393 = n163 & n392 ;
  assign n394 = n391 & n393 ;
  assign n395 = ~x48 & ~x49 ;
  assign n396 = n167 & n395 ;
  assign n398 = n165 & n397 ;
  assign n399 = n394 & n398 ;
  assign n400 = n396 & n399 ;
  assign n401 = ~x44 & ~x45 ;
  assign n402 = n169 & n401 ;
  assign n403 = ~x40 & ~x41 ;
  assign n404 = n171 & n403 ;
  assign n405 = n402 & n404 ;
  assign n406 = ~x36 & ~x37 ;
  assign n407 = n173 & n406 ;
  assign n408 = ~x32 & ~x33 ;
  assign n409 = n175 & n408 ;
  assign n410 = n405 & n407 ;
  assign n411 = n409 & n410 ;
  assign n412 = n400 & n411 ;
  assign n413 = ~x16 & ~x17 ;
  assign n414 = n183 & n413 ;
  assign n415 = ~x20 & ~x21 ;
  assign n416 = ~x28 & ~x29 ;
  assign n417 = n177 & n416 ;
  assign n418 = ~x24 & ~x25 ;
  assign n419 = n179 & n418 ;
  assign n420 = n417 & n419 ;
  assign n421 = n181 & n420 ;
  assign n422 = n415 & n421 ;
  assign n423 = n414 & n422 ;
  assign n446 = ~x12 & ~x13 ;
  assign n447 = n185 & n446 ;
  assign n460 = n447 ^ n185 ;
  assign n424 = n139 & n367 ;
  assign n425 = n365 & n424 ;
  assign n426 = n143 & n371 ;
  assign n427 = n369 & n426 ;
  assign n428 = n425 & n427 ;
  assign n437 = n428 & n436 ;
  assign n438 = n389 & n400 ;
  assign n439 = n411 & n438 ;
  assign n440 = ~n423 & n439 ;
  assign n441 = n440 ^ n438 ;
  assign n442 = n441 ^ n389 ;
  assign n443 = n437 & ~n442 ;
  assign n444 = n443 ^ n428 ;
  assign n445 = ~x8 & ~x9 ;
  assign n457 = n446 ^ n187 ;
  assign n458 = n447 & ~n457 ;
  assign n449 = n445 & n458 ;
  assign n450 = ~n444 & ~n449 ;
  assign n451 = n189 & ~n450 ;
  assign n455 = n451 ^ n450 ;
  assign n452 = ~x4 & ~x5 ;
  assign n453 = ~n191 & n452 ;
  assign n454 = n451 & n453 ;
  assign n456 = n455 ^ n454 ;
  assign n459 = n456 & n458 ;
  assign n461 = n460 ^ n459 ;
  assign n462 = n423 & ~n461 ;
  assign n467 = ~n181 & n419 ;
  assign n468 = n467 ^ n179 ;
  assign n469 = n417 & ~n468 ;
  assign n474 = ~n183 & n422 ;
  assign n475 = n474 ^ n177 ;
  assign n476 = ~n469 & n475 ;
  assign n477 = ~n462 & n476 ;
  assign n478 = n412 & ~n477 ;
  assign n479 = n175 & ~n478 ;
  assign n480 = n407 & ~n479 ;
  assign n481 = n173 & ~n480 ;
  assign n482 = n405 & ~n481 ;
  assign n483 = n169 & ~n482 ;
  assign n484 = n400 & n483 ;
  assign n491 = ~n171 & n401 ;
  assign n492 = n484 & n491 ;
  assign n493 = n492 ^ n484 ;
  assign n494 = n493 ^ n400 ;
  assign n495 = n165 & ~n494 ;
  assign n496 = n394 & n495 ;
  assign n504 = ~n167 & n496 ;
  assign n505 = n397 & n504 ;
  assign n506 = n505 ^ n397 ;
  assign n497 = n496 ^ n394 ;
  assign n498 = n497 ^ n397 ;
  assign n507 = n506 ^ n498 ;
  assign n508 = n161 & ~n507 ;
  assign n509 = n389 & n508 ;
  assign n512 = ~n163 & n390 ;
  assign n514 = n509 & n512 ;
  assign n510 = n509 ^ n389 ;
  assign n511 = n510 ^ n382 ;
  assign n515 = n514 ^ n511 ;
  assign n516 = ~n383 & n515 ;
  assign n517 = n382 & ~n516 ;
  assign n518 = n517 ^ n157 ;
  assign n519 = n380 & ~n518 ;
  assign n520 = n519 ^ n378 ;
  assign n521 = ~n379 & n520 ;
  assign n522 = n378 & ~n521 ;
  assign n523 = n522 ^ n153 ;
  assign n524 = n436 & ~n523 ;
  assign n525 = n149 & ~n524 ;
  assign n526 = n375 & n525 ;
  assign n528 = ~n151 & n433 ;
  assign n529 = n526 & n528 ;
  assign n376 = n375 ^ n373 ;
  assign n527 = n526 ^ n376 ;
  assign n530 = n529 ^ n527 ;
  assign n531 = ~n374 & n530 ;
  assign n532 = n373 & ~n531 ;
  assign n533 = n532 ^ n145 ;
  assign n534 = n371 & ~n533 ;
  assign n535 = n534 ^ n369 ;
  assign n536 = ~n370 & n535 ;
  assign n537 = n369 & ~n536 ;
  assign n538 = n537 ^ n141 ;
  assign n539 = n367 & ~n538 ;
  assign n540 = n539 ^ n365 ;
  assign n541 = ~n366 & n540 ;
  assign n542 = n365 & ~n541 ;
  assign n543 = n542 ^ n137 ;
  assign n544 = n363 & ~n543 ;
  assign n545 = n135 & ~n544 ;
  assign n546 = n359 & ~n545 ;
  assign n547 = n546 ^ n354 ;
  assign n556 = ~n133 & n356 ;
  assign n557 = n556 ^ n133 ;
  assign n548 = n353 ^ n131 ;
  assign n549 = n548 ^ n133 ;
  assign n558 = n557 ^ n549 ;
  assign n559 = n547 & ~n558 ;
  assign n560 = n354 & ~n559 ;
  assign n561 = n560 ^ n129 ;
  assign n571 = n420 ^ n417 ;
  assign n562 = n414 & n447 ;
  assign n566 = n451 & n452 ;
  assign n567 = n566 ^ n450 ;
  assign n568 = n562 & n567 ;
  assign n569 = n568 ^ n414 ;
  assign n570 = n422 & ~n569 ;
  assign n572 = n571 ^ n570 ;
  assign n573 = n407 & n409 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = n574 ^ n407 ;
  assign n576 = n404 & ~n575 ;
  assign n577 = n402 & ~n576 ;
  assign n578 = n396 & ~n577 ;
  assign n579 = n398 & ~n578 ;
  assign n580 = n393 & ~n579 ;
  assign n581 = n391 & ~n580 ;
  assign n582 = n387 & ~n581 ;
  assign n583 = n382 & ~n582 ;
  assign n584 = n384 & ~n583 ;
  assign n585 = n378 & ~n584 ;
  assign n586 = n430 & ~n585 ;
  assign n587 = n432 & ~n586 ;
  assign n588 = n432 ^ n373 ;
  assign n589 = n588 ^ n434 ;
  assign n590 = n587 & n589 ;
  assign n591 = n590 ^ n588 ;
  assign n592 = n426 & ~n591 ;
  assign n593 = n369 & ~n592 ;
  assign n594 = n424 & ~n593 ;
  assign n595 = n365 & ~n594 ;
  assign n596 = n362 & ~n595 ;
  assign n597 = n358 & ~n596 ;
  assign n598 = n356 & ~n597 ;
  assign n599 = n354 & ~n598 ;
  assign n600 = n354 & n356 ;
  assign n601 = n389 & n436 ;
  assign n610 = n400 & ~n405 ;
  assign n602 = n412 & n420 ;
  assign n603 = ~n450 & n602 ;
  assign n604 = n603 ^ n412 ;
  assign n605 = n604 ^ n394 ;
  assign n611 = n610 ^ n605 ;
  assign n612 = n601 & ~n611 ;
  assign n617 = ~n385 & n436 ;
  assign n618 = n617 ^ n432 ;
  assign n619 = ~n612 & n618 ;
  assign n620 = n427 & ~n619 ;
  assign n621 = n425 & ~n620 ;
  assign n622 = n362 & ~n621 ;
  assign n623 = n600 & ~n622 ;
  assign n624 = n363 & ~n444 ;
  assign n625 = n363 & n428 ;
  assign n626 = n601 & n625 ;
  assign n627 = ~n412 & n626 ;
  assign n628 = n627 ^ n625 ;
  assign n629 = ~x0 & ~x1 ;
  assign n630 = n412 & n629 ;
  assign n631 = n626 & n630 ;
  assign n632 = ~n442 & n631 ;
  assign n633 = n456 & n632 ;
  assign n634 = ~n604 & n633 ;
  assign n635 = ~n569 & n634 ;
  assign y0 = n352 ;
  assign y1 = ~n561 ;
  assign y2 = ~n599 ;
  assign y3 = ~n623 ;
  assign y4 = ~n624 ;
  assign y5 = ~n628 ;
  assign y6 = ~n626 ;
  assign y7 = ~n635 ;
endmodule
