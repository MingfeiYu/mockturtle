module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 ;
  assign n65 = x63 ^ x31 ;
  assign n68 = ~x28 & x60 ;
  assign n67 = x60 ^ x28 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ x62 ;
  assign n66 = x62 ^ x29 ;
  assign n71 = n70 ^ n66 ;
  assign n72 = x61 ^ x29 ;
  assign n75 = n71 & n72 ;
  assign n76 = n75 ^ n70 ;
  assign n78 = x63 ^ x30 ;
  assign n77 = x63 ^ x62 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n76 & ~n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = ~n65 & ~n81 ;
  assign n83 = n82 ^ x31 ;
  assign n84 = ~x27 & x59 ;
  assign n85 = ~x25 & ~x57 ;
  assign n86 = n85 ^ x25 ;
  assign n87 = ~n84 & n86 ;
  assign n88 = ~x26 & x58 ;
  assign n89 = n87 & n88 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = ~x56 & n90 ;
  assign n92 = x24 & n90 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = x31 & ~n68 ;
  assign n95 = ~x63 & n94 ;
  assign n96 = n95 ^ n68 ;
  assign n97 = x61 & ~n96 ;
  assign n98 = n95 ^ x29 ;
  assign n99 = n97 & ~n98 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = ~x30 & x62 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = ~n93 & ~n103 ;
  assign n105 = x49 ^ x17 ;
  assign n106 = x50 ^ x18 ;
  assign n107 = x51 ^ x19 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = ~x16 & x48 ;
  assign n110 = x47 ^ x15 ;
  assign n114 = ~x13 & ~x45 ;
  assign n112 = ~x15 & x47 ;
  assign n111 = x46 ^ x45 ;
  assign n113 = n112 ^ n111 ;
  assign n115 = n114 ^ n113 ;
  assign n118 = x47 ^ x14 ;
  assign n116 = x47 ^ x46 ;
  assign n117 = n116 ^ n112 ;
  assign n119 = n118 ^ n117 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = ~n110 & n121 ;
  assign n123 = n122 ^ x15 ;
  assign n124 = n114 ^ x13 ;
  assign n125 = ~n112 & n124 ;
  assign n126 = ~x14 & x46 ;
  assign n127 = n125 & n126 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = n123 ^ x44 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = x44 ^ x12 ;
  assign n133 = x39 ^ x38 ;
  assign n132 = x39 ^ x6 ;
  assign n134 = n133 ^ n132 ;
  assign n157 = x39 ^ x5 ;
  assign n161 = n157 ^ n132 ;
  assign n136 = x34 ^ x2 ;
  assign n137 = x33 ^ x1 ;
  assign n138 = n137 ^ n136 ;
  assign n141 = ~x0 & x32 ;
  assign n142 = n141 ^ x1 ;
  assign n143 = ~n138 & ~n142 ;
  assign n139 = x34 ^ x1 ;
  assign n144 = n143 ^ n139 ;
  assign n145 = ~n136 & ~n144 ;
  assign n135 = x35 ^ x34 ;
  assign n146 = n145 ^ n135 ;
  assign n148 = x36 ^ x3 ;
  assign n147 = x36 ^ x35 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = ~n146 & ~n149 ;
  assign n151 = n150 ^ n148 ;
  assign n153 = x37 ^ x4 ;
  assign n152 = x37 ^ x36 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n151 & ~n154 ;
  assign n156 = n155 ^ n153 ;
  assign n159 = x37 ^ x5 ;
  assign n160 = n156 & ~n159 ;
  assign n162 = n161 ^ n160 ;
  assign n163 = ~n134 & ~n162 ;
  assign n164 = n163 ^ n133 ;
  assign n175 = x39 ^ x7 ;
  assign n176 = ~n164 & ~n175 ;
  assign n165 = x43 ^ x11 ;
  assign n166 = x42 ^ x10 ;
  assign n167 = ~n165 & ~n166 ;
  assign n169 = x41 ^ x9 ;
  assign n168 = x9 & ~x41 ;
  assign n170 = n169 ^ n168 ;
  assign n171 = x8 & ~n170 ;
  assign n172 = n167 & n171 ;
  assign n173 = n172 ^ x7 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = ~x40 & n167 ;
  assign n179 = ~n170 & n178 ;
  assign n180 = n179 ^ n172 ;
  assign n181 = n177 & n180 ;
  assign n182 = n181 ^ n172 ;
  assign n183 = ~n131 & ~n182 ;
  assign n187 = n168 ^ x43 ;
  assign n184 = x43 ^ x42 ;
  assign n188 = n187 ^ n184 ;
  assign n189 = ~n166 & ~n188 ;
  assign n190 = n189 ^ n184 ;
  assign n191 = ~n165 & n190 ;
  assign n192 = n191 ^ x43 ;
  assign n193 = n183 & n192 ;
  assign n194 = n193 ^ n131 ;
  assign n195 = n194 ^ x44 ;
  assign n196 = n195 ^ n128 ;
  assign n198 = n131 ^ n123 ;
  assign n199 = ~n196 & n198 ;
  assign n200 = n130 & n199 ;
  assign n201 = n200 ^ n194 ;
  assign n202 = n201 ^ n123 ;
  assign n203 = n128 & ~n202 ;
  assign n204 = ~n123 & n203 ;
  assign n205 = n204 ^ n123 ;
  assign n206 = ~n109 & n205 ;
  assign n207 = n108 & n206 ;
  assign n208 = ~n105 & n207 ;
  assign n209 = ~x20 & x52 ;
  assign n210 = ~x22 & x54 ;
  assign n211 = ~x23 & x55 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n212 ^ n210 ;
  assign n214 = ~n209 & ~n213 ;
  assign n215 = ~x21 & x53 ;
  assign n216 = n214 & n215 ;
  assign n217 = n216 ^ n214 ;
  assign n218 = n208 & n217 ;
  assign n219 = n104 & n218 ;
  assign n220 = n83 & ~n219 ;
  assign n221 = n93 ^ n91 ;
  assign n222 = n221 ^ n92 ;
  assign n223 = x59 ^ x27 ;
  assign n224 = x58 ^ x57 ;
  assign n225 = n224 ^ n84 ;
  assign n226 = n225 ^ n85 ;
  assign n229 = x59 ^ x26 ;
  assign n227 = x59 ^ x58 ;
  assign n228 = n227 ^ n84 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = ~n226 & ~n230 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = ~n223 & n232 ;
  assign n234 = n233 ^ x27 ;
  assign n235 = ~n103 & ~n234 ;
  assign n236 = n222 & n235 ;
  assign n237 = n236 ^ n103 ;
  assign n263 = x52 ^ x20 ;
  assign n264 = n263 ^ n209 ;
  assign n265 = n264 ^ x53 ;
  assign n266 = x53 ^ x21 ;
  assign n267 = n265 & ~n266 ;
  assign n268 = n267 ^ x21 ;
  assign n238 = x55 ^ x23 ;
  assign n239 = x54 ^ x22 ;
  assign n240 = n239 ^ n210 ;
  assign n241 = n240 ^ x55 ;
  assign n242 = ~n238 & n241 ;
  assign n243 = n242 ^ x23 ;
  assign n244 = n217 & ~n243 ;
  assign n248 = x50 ^ x49 ;
  assign n249 = n248 ^ x17 ;
  assign n246 = x48 ^ x16 ;
  assign n247 = n246 ^ n109 ;
  assign n250 = n249 ^ n247 ;
  assign n251 = n250 ^ n248 ;
  assign n252 = ~n105 & ~n251 ;
  assign n253 = n252 ^ n248 ;
  assign n254 = ~n106 & n253 ;
  assign n245 = x51 ^ x50 ;
  assign n255 = n254 ^ n245 ;
  assign n256 = ~n107 & ~n255 ;
  assign n257 = n256 ^ x19 ;
  assign n258 = n244 & n257 ;
  assign n259 = n258 ^ n243 ;
  assign n260 = n104 & n259 ;
  assign n261 = n260 ^ n104 ;
  assign n269 = ~n213 & n261 ;
  assign n270 = n268 & n269 ;
  assign n271 = n270 ^ n260 ;
  assign n272 = n237 & ~n271 ;
  assign n273 = n220 & n272 ;
  assign y0 = n273 ;
endmodule
