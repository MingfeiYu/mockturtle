module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n29 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n43 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n107 , n108 , n110 , n111 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n181 , n182 , n183 , n184 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n241 , n242 , n247 , n249 , n250 , n251 , n252 , n255 , n256 , n260 , n261 , n262 , n263 , n265 , n266 , n267 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n362 , n363 , n364 , n365 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n435 , n436 , n437 , n438 , n439 , n440 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n476 , n479 , n480 , n481 , n482 , n483 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n695 , n696 , n697 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n880 , n881 , n882 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n901 , n902 , n903 , n904 , n905 , n906 , n908 , n909 , n910 , n911 , n912 ;
  assign n12 = x9 ^ x8 ;
  assign n11 = x8 & ~x9 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ x8 ;
  assign n15 = x2 & x3 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = x0 & ~x1 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = ~n17 & ~n19 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = x6 ^ x5 ;
  assign n23 = n20 ^ x4 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = x5 & x6 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ x5 ;
  assign n61 = ~x7 & ~x9 ;
  assign n62 = ~n17 & ~n61 ;
  assign n207 = ~x7 & x8 ;
  assign n31 = n207 ^ x7 ;
  assign n63 = n13 ^ x0 ;
  assign n64 = n31 & n63 ;
  assign n65 = n62 & n64 ;
  assign n50 = x3 ^ x2 ;
  assign n51 = x0 & ~n50 ;
  assign n43 = n17 ^ x2 ;
  assign n46 = ~n14 & n43 ;
  assign n38 = n14 ^ n12 ;
  assign n39 = ~n16 & n38 ;
  assign n40 = n39 ^ n38 ;
  assign n47 = n46 ^ n40 ;
  assign n48 = ~x0 & n47 ;
  assign n52 = ~x3 & x9 ;
  assign n53 = n52 ^ n11 ;
  assign n54 = ~n48 & n53 ;
  assign n55 = n51 & n54 ;
  assign n33 = x8 ^ x0 ;
  assign n34 = n33 ^ n11 ;
  assign n35 = n11 ^ x2 ;
  assign n36 = ~x3 & ~n35 ;
  assign n37 = ~n34 & n36 ;
  assign n49 = n48 ^ n37 ;
  assign n56 = n55 ^ n49 ;
  assign n57 = ~x7 & n56 ;
  assign n58 = n57 ^ n37 ;
  assign n59 = ~x1 & ~n58 ;
  assign n32 = n31 ^ x1 ;
  assign n60 = n59 ^ n32 ;
  assign n66 = n65 ^ n60 ;
  assign n71 = ~n27 & n66 ;
  assign n88 = x6 & ~x7 ;
  assign n122 = n43 ^ x8 ;
  assign n125 = ~x5 & n122 ;
  assign n126 = n125 ^ x8 ;
  assign n127 = ~n19 & n126 ;
  assign n128 = x5 & x8 ;
  assign n129 = n128 ^ x8 ;
  assign n80 = x0 & ~x8 ;
  assign n81 = n80 ^ n33 ;
  assign n82 = x1 & ~n81 ;
  assign n73 = ~x1 & x8 ;
  assign n74 = n73 ^ x1 ;
  assign n130 = n82 ^ n74 ;
  assign n131 = n130 ^ x8 ;
  assign n132 = x1 & ~x2 ;
  assign n133 = n132 ^ x2 ;
  assign n134 = n133 ^ x8 ;
  assign n135 = ~x5 & n134 ;
  assign n136 = n135 ^ x8 ;
  assign n137 = n17 & n136 ;
  assign n138 = ~n131 & ~n137 ;
  assign n139 = ~n129 & ~n138 ;
  assign n140 = x5 & x9 ;
  assign n142 = x9 ^ x0 ;
  assign n141 = ~x0 & ~x9 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = ~n140 & n143 ;
  assign n145 = ~n39 & n144 ;
  assign n146 = n145 ^ n139 ;
  assign n147 = ~n139 & ~n146 ;
  assign n148 = ~n127 & n147 ;
  assign n149 = n88 & ~n148 ;
  assign n92 = ~x2 & x8 ;
  assign n93 = n92 ^ x8 ;
  assign n150 = n18 & n93 ;
  assign n151 = n150 ^ n80 ;
  assign n152 = x9 ^ x5 ;
  assign n153 = n152 ^ n140 ;
  assign n154 = x8 ^ x3 ;
  assign n67 = x8 ^ x2 ;
  assign n155 = x8 ^ x1 ;
  assign n158 = n67 & ~n155 ;
  assign n159 = n154 & n158 ;
  assign n160 = n159 ^ n154 ;
  assign n161 = n160 ^ x3 ;
  assign n162 = ~x0 & ~n161 ;
  assign n163 = ~n153 & ~n162 ;
  assign n164 = n151 & n163 ;
  assign n172 = n74 & n164 ;
  assign n173 = ~x3 & n172 ;
  assign n174 = n173 ^ x3 ;
  assign n165 = n164 ^ n163 ;
  assign n166 = n165 ^ x3 ;
  assign n175 = n174 ^ n166 ;
  assign n176 = n149 & ~n175 ;
  assign n183 = n140 ^ n11 ;
  assign n181 = ~x5 & ~n38 ;
  assign n182 = n181 ^ n129 ;
  assign n184 = n183 ^ n182 ;
  assign n189 = n176 & ~n184 ;
  assign n190 = ~n20 & n189 ;
  assign n191 = n190 ^ n20 ;
  assign n84 = x9 ^ x1 ;
  assign n78 = x1 & ~x9 ;
  assign n79 = n78 ^ x1 ;
  assign n83 = n82 ^ n79 ;
  assign n85 = n84 ^ n83 ;
  assign n72 = ~x1 & n14 ;
  assign n75 = n74 ^ n72 ;
  assign n76 = n75 ^ x1 ;
  assign n77 = n76 ^ n38 ;
  assign n86 = n85 ^ n77 ;
  assign n87 = n86 ^ x8 ;
  assign n90 = ~x7 & ~n27 ;
  assign n89 = n88 ^ x7 ;
  assign n91 = n90 ^ n89 ;
  assign n94 = ~x3 & ~n93 ;
  assign n110 = n79 ^ x9 ;
  assign n111 = n110 ^ x2 ;
  assign n116 = n94 & n111 ;
  assign n117 = n18 & n116 ;
  assign n118 = n117 ^ n18 ;
  assign n98 = ~x0 & x2 ;
  assign n97 = x2 ^ x0 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = ~x9 & n99 ;
  assign n95 = x2 & n14 ;
  assign n96 = n95 ^ n93 ;
  assign n101 = n100 ^ n96 ;
  assign n102 = x3 & ~n92 ;
  assign n103 = x1 & n102 ;
  assign n104 = n101 & n103 ;
  assign n105 = n104 ^ n102 ;
  assign n107 = n105 ^ n94 ;
  assign n108 = n107 ^ n18 ;
  assign n119 = n118 ^ n108 ;
  assign n120 = ~n91 & n119 ;
  assign n121 = ~n87 & n120 ;
  assign n178 = n176 ^ n121 ;
  assign n179 = n178 ^ n20 ;
  assign n192 = n191 ^ n179 ;
  assign n193 = ~n71 & ~n192 ;
  assign n194 = n24 & ~n193 ;
  assign n195 = n22 & n194 ;
  assign n196 = n21 & n195 ;
  assign n197 = n196 ^ n194 ;
  assign n198 = n197 ^ n193 ;
  assign n203 = n52 ^ x3 ;
  assign n204 = x1 ^ x0 ;
  assign n208 = n207 ^ x2 ;
  assign n209 = n155 & ~n208 ;
  assign n210 = n209 ^ x2 ;
  assign n211 = n204 & ~n210 ;
  assign n212 = ~n203 & n211 ;
  assign n213 = n38 ^ x7 ;
  assign n214 = ~x3 & ~n133 ;
  assign n215 = n214 ^ x3 ;
  assign n216 = n213 & ~n215 ;
  assign n217 = n99 ^ n19 ;
  assign n218 = n216 & ~n217 ;
  assign n219 = ~n212 & ~n218 ;
  assign n200 = n61 & ~n150 ;
  assign n220 = n219 ^ n200 ;
  assign n199 = n92 ^ x2 ;
  assign n201 = ~n19 & n200 ;
  assign n202 = ~n199 & n201 ;
  assign n221 = n220 ^ n202 ;
  assign n222 = ~n27 & ~n221 ;
  assign n223 = ~x1 & ~x5 ;
  assign n225 = n142 ^ n52 ;
  assign n224 = ~x0 & x3 ;
  assign n226 = n225 ^ n224 ;
  assign n227 = n12 & n226 ;
  assign n228 = n227 ^ x3 ;
  assign n229 = n223 & ~n228 ;
  assign n230 = n182 ^ n152 ;
  assign n231 = x3 ^ x1 ;
  assign n232 = x1 & n231 ;
  assign n233 = n232 ^ n79 ;
  assign n234 = ~n230 & n233 ;
  assign n235 = x2 & ~n140 ;
  assign n236 = ~n234 & n235 ;
  assign n237 = ~n229 & n236 ;
  assign n272 = ~x3 & n19 ;
  assign n262 = x0 & n13 ;
  assign n249 = n231 ^ n13 ;
  assign n250 = x3 & ~n140 ;
  assign n251 = n250 ^ n63 ;
  assign n252 = n251 ^ n249 ;
  assign n263 = n252 ^ x3 ;
  assign n265 = ~n249 & ~n263 ;
  assign n266 = n262 & n265 ;
  assign n238 = n140 ^ x3 ;
  assign n239 = n238 ^ n204 ;
  assign n260 = n239 ^ x3 ;
  assign n261 = n260 ^ n252 ;
  assign n267 = n266 ^ n261 ;
  assign n269 = n267 ^ n63 ;
  assign n270 = n269 ^ n231 ;
  assign n241 = n13 ^ x1 ;
  assign n242 = n241 ^ n238 ;
  assign n255 = n242 ^ x0 ;
  assign n256 = n255 ^ n238 ;
  assign n247 = n256 ^ n140 ;
  assign n271 = n270 ^ n247 ;
  assign n273 = n272 ^ n271 ;
  assign n274 = ~x2 & n153 ;
  assign n275 = n18 ^ x0 ;
  assign n282 = ~n17 & n275 ;
  assign n276 = n274 ^ n140 ;
  assign n277 = n276 ^ n82 ;
  assign n283 = n282 ^ n277 ;
  assign n284 = ~n274 & ~n283 ;
  assign n285 = n284 ^ n277 ;
  assign n287 = n285 ^ n274 ;
  assign n288 = n285 ^ n140 ;
  assign n289 = ~n287 & n288 ;
  assign n286 = n285 ^ n82 ;
  assign n291 = n289 ^ n286 ;
  assign n292 = n291 ^ n82 ;
  assign n293 = n273 & ~n292 ;
  assign n294 = n88 & ~n293 ;
  assign n295 = ~n237 & n294 ;
  assign n304 = n16 ^ x9 ;
  assign n296 = ~x9 & ~n16 ;
  assign n305 = n304 ^ n296 ;
  assign n302 = n96 ^ n40 ;
  assign n303 = n302 ^ n203 ;
  assign n306 = n305 ^ n303 ;
  assign n297 = n52 ^ n16 ;
  assign n298 = n297 ^ n296 ;
  assign n299 = ~x0 & ~n77 ;
  assign n300 = n298 & n299 ;
  assign n301 = ~n296 & ~n300 ;
  assign n307 = n301 ^ n300 ;
  assign n310 = n92 & ~n307 ;
  assign n311 = n310 ^ n300 ;
  assign n312 = ~n306 & ~n311 ;
  assign n313 = n312 ^ n301 ;
  assign n314 = x1 & n313 ;
  assign n315 = n314 ^ n301 ;
  assign n316 = ~n91 & n315 ;
  assign n324 = ~x3 & n316 ;
  assign n325 = n150 & n324 ;
  assign n326 = n325 ^ n150 ;
  assign n317 = n316 ^ n91 ;
  assign n318 = n317 ^ n150 ;
  assign n327 = n326 ^ n318 ;
  assign n328 = ~n295 & n327 ;
  assign n329 = ~n222 & n328 ;
  assign n335 = n14 & n20 ;
  assign n330 = ~x0 & ~x6 ;
  assign n331 = ~x9 & ~n330 ;
  assign n332 = n214 & ~n331 ;
  assign n336 = n335 ^ n332 ;
  assign n337 = ~x4 & ~n336 ;
  assign n338 = n337 ^ n332 ;
  assign n339 = ~n329 & ~n338 ;
  assign n340 = n339 ^ n329 ;
  assign n362 = ~x6 & x8 ;
  assign n382 = ~x1 & n100 ;
  assign n383 = ~n362 & n382 ;
  assign n380 = n38 & n98 ;
  assign n376 = ~x9 & ~n81 ;
  assign n377 = n376 ^ x0 ;
  assign n375 = n141 ^ n11 ;
  assign n378 = n377 ^ n375 ;
  assign n379 = n132 & n378 ;
  assign n381 = n380 ^ n379 ;
  assign n384 = n383 ^ n381 ;
  assign n395 = x8 ^ x6 ;
  assign n396 = n395 ^ n362 ;
  assign n391 = ~x8 & ~n330 ;
  assign n341 = ~x2 & x6 ;
  assign n342 = n341 ^ x2 ;
  assign n392 = n391 ^ n342 ;
  assign n393 = n342 ^ x0 ;
  assign n394 = ~n392 & ~n393 ;
  assign n397 = n396 ^ n394 ;
  assign n398 = n78 & n397 ;
  assign n385 = ~x6 & n38 ;
  assign n386 = n385 ^ x6 ;
  assign n387 = ~n19 & n386 ;
  assign n388 = x2 & n11 ;
  assign n389 = n388 ^ x9 ;
  assign n390 = n387 & n389 ;
  assign n399 = n398 ^ n390 ;
  assign n400 = ~n384 & ~n399 ;
  assign n401 = ~x5 & ~x7 ;
  assign n402 = ~n13 & ~n27 ;
  assign n403 = ~n401 & n402 ;
  assign n405 = x0 & n78 ;
  assign n406 = n403 & n405 ;
  assign n404 = n403 ^ n401 ;
  assign n407 = n406 ^ n404 ;
  assign n352 = ~x1 & ~x6 ;
  assign n351 = x6 ^ x1 ;
  assign n353 = n352 ^ n351 ;
  assign n354 = n353 ^ x1 ;
  assign n408 = x9 ^ x7 ;
  assign n409 = ~x0 & ~x3 ;
  assign n410 = ~n408 & n409 ;
  assign n418 = ~x9 & n410 ;
  assign n419 = n354 & n418 ;
  assign n420 = n419 ^ n354 ;
  assign n411 = n410 ^ x3 ;
  assign n412 = n411 ^ n354 ;
  assign n421 = n420 ^ n412 ;
  assign n422 = n407 & ~n421 ;
  assign n423 = ~n400 & n422 ;
  assign n343 = n342 ^ x6 ;
  assign n345 = ~x2 & ~n81 ;
  assign n344 = n98 ^ n92 ;
  assign n346 = n345 ^ n344 ;
  assign n347 = n52 & n346 ;
  assign n348 = ~x3 & ~n347 ;
  assign n349 = ~n343 & n348 ;
  assign n355 = ~n11 & ~n354 ;
  assign n356 = n349 & n355 ;
  assign n350 = n349 ^ n347 ;
  assign n357 = n356 ^ n350 ;
  assign n358 = ~x0 & n357 ;
  assign n363 = n362 ^ n342 ;
  assign n364 = n363 ^ n199 ;
  assign n365 = n364 ^ x2 ;
  assign n370 = n358 & ~n365 ;
  assign n371 = n79 & n370 ;
  assign n372 = n371 ^ n79 ;
  assign n359 = n358 ^ n357 ;
  assign n360 = n359 ^ n79 ;
  assign n373 = n372 ^ n360 ;
  assign n374 = ~x7 & ~n373 ;
  assign n424 = n423 ^ n374 ;
  assign n425 = ~x2 & ~n19 ;
  assign n476 = ~x8 & n26 ;
  assign n479 = n425 & ~n476 ;
  assign n426 = n353 ^ x0 ;
  assign n427 = x5 & n78 ;
  assign n428 = n427 ^ x9 ;
  assign n429 = ~x0 & n428 ;
  assign n430 = n429 ^ n427 ;
  assign n431 = x2 & ~x5 ;
  assign n432 = n431 ^ n342 ;
  assign n435 = n432 ^ x8 ;
  assign n436 = ~n430 & ~n435 ;
  assign n437 = n436 ^ x0 ;
  assign n438 = ~x8 & ~n437 ;
  assign n439 = ~n426 & n438 ;
  assign n440 = n431 ^ x9 ;
  assign n442 = ~x0 & n440 ;
  assign n443 = n442 ^ x9 ;
  assign n444 = n439 & n443 ;
  assign n445 = n444 ^ n438 ;
  assign n446 = ~x6 & x9 ;
  assign n447 = n446 ^ n26 ;
  assign n448 = n73 & ~n81 ;
  assign n449 = n447 & n448 ;
  assign n450 = n449 ^ n81 ;
  assign n452 = n129 & ~n388 ;
  assign n453 = ~n450 & n452 ;
  assign n454 = n453 ^ n450 ;
  assign n455 = ~x0 & ~n25 ;
  assign n456 = n78 & n431 ;
  assign n457 = ~n274 & ~n456 ;
  assign n458 = n455 & n457 ;
  assign n459 = n454 & n458 ;
  assign n467 = n432 & n459 ;
  assign n468 = ~x1 & n467 ;
  assign n469 = n468 ^ x1 ;
  assign n460 = n459 ^ n454 ;
  assign n461 = n460 ^ x1 ;
  assign n470 = n469 ^ n461 ;
  assign n471 = ~n445 & ~n470 ;
  assign n472 = ~x4 & ~n471 ;
  assign n473 = n472 ^ x4 ;
  assign n480 = n479 ^ n473 ;
  assign n481 = ~x3 & ~n480 ;
  assign n482 = n481 ^ n472 ;
  assign n483 = n424 & n482 ;
  assign n492 = x0 & ~n446 ;
  assign n493 = n25 ^ x5 ;
  assign n498 = ~x1 & ~n493 ;
  assign n499 = n498 ^ n182 ;
  assign n500 = n492 & n499 ;
  assign n501 = n500 ^ n385 ;
  assign n486 = n385 ^ n362 ;
  assign n487 = ~x0 & ~n486 ;
  assign n488 = n487 ^ n385 ;
  assign n489 = x5 & n488 ;
  assign n490 = n489 ^ n385 ;
  assign n491 = x1 & n490 ;
  assign n502 = n501 ^ n491 ;
  assign n503 = x3 & n502 ;
  assign n504 = ~n22 & n214 ;
  assign n505 = n504 ^ x4 ;
  assign n511 = x0 & x5 ;
  assign n512 = n511 ^ x5 ;
  assign n513 = n353 & n512 ;
  assign n507 = x5 ^ x2 ;
  assign n508 = n507 ^ x6 ;
  assign n509 = n25 & ~n508 ;
  assign n506 = n341 ^ n26 ;
  assign n510 = n509 ^ n506 ;
  assign n514 = n513 ^ n510 ;
  assign n515 = ~x3 & ~n81 ;
  assign n516 = n456 & n515 ;
  assign n517 = n516 ^ x3 ;
  assign n518 = n514 & ~n517 ;
  assign n522 = n518 ^ n517 ;
  assign n519 = n79 & n93 ;
  assign n520 = ~x6 & ~n519 ;
  assign n521 = n518 & n520 ;
  assign n523 = n522 ^ n521 ;
  assign n533 = n81 ^ x9 ;
  assign n536 = ~n84 & n533 ;
  assign n537 = n536 ^ x9 ;
  assign n538 = n26 & n537 ;
  assign n539 = n538 ^ x5 ;
  assign n543 = n533 ^ n376 ;
  assign n544 = n543 ^ n19 ;
  assign n540 = x1 & ~n377 ;
  assign n541 = n540 ^ x0 ;
  assign n542 = n541 ^ n83 ;
  assign n545 = n544 ^ n542 ;
  assign n546 = ~x6 & n545 ;
  assign n547 = ~n343 & ~n546 ;
  assign n548 = ~n539 & n547 ;
  assign n524 = n67 ^ x9 ;
  assign n525 = n524 ^ x1 ;
  assign n526 = ~n67 & ~n155 ;
  assign n527 = n526 ^ x1 ;
  assign n528 = ~n525 & n527 ;
  assign n529 = n528 ^ x1 ;
  assign n530 = ~x6 & n529 ;
  assign n531 = n530 ^ x1 ;
  assign n532 = n511 & n531 ;
  assign n549 = n548 ^ n532 ;
  assign n551 = ~n523 & ~n549 ;
  assign n552 = ~x7 & ~n551 ;
  assign n553 = ~n505 & n552 ;
  assign n554 = n503 & n553 ;
  assign n556 = ~n25 & ~n111 ;
  assign n557 = n554 & n556 ;
  assign n555 = n554 ^ n553 ;
  assign n558 = n557 ^ n555 ;
  assign n559 = n19 ^ x2 ;
  assign n560 = n401 ^ x7 ;
  assign n561 = n560 ^ n91 ;
  assign n562 = ~n23 & n561 ;
  assign n563 = ~n559 & n562 ;
  assign n564 = n425 ^ x3 ;
  assign n565 = n425 ^ x4 ;
  assign n566 = n561 & ~n565 ;
  assign n567 = n564 & n566 ;
  assign n678 = ~x2 & ~n561 ;
  assign n668 = x1 & ~n27 ;
  assign n679 = ~x9 & ~n668 ;
  assign n29 = x7 & ~x8 ;
  assign n680 = n476 ^ n29 ;
  assign n569 = n128 ^ x5 ;
  assign n681 = n680 ^ n569 ;
  assign n682 = n679 & ~n681 ;
  assign n683 = n682 ^ x9 ;
  assign n684 = n678 & n683 ;
  assign n688 = ~n31 & ~n353 ;
  assign n689 = n684 & n688 ;
  assign n662 = x2 & n207 ;
  assign n663 = ~n153 & n662 ;
  assign n664 = n353 & n663 ;
  assign n665 = n664 ^ n662 ;
  assign n666 = n665 ^ x2 ;
  assign n673 = ~n207 & n352 ;
  assign n674 = n181 & n673 ;
  assign n667 = n354 ^ x5 ;
  assign n669 = n668 ^ n667 ;
  assign n670 = ~x7 & ~n79 ;
  assign n671 = n669 & n670 ;
  assign n672 = n671 ^ x7 ;
  assign n675 = n674 ^ n672 ;
  assign n677 = n666 & n675 ;
  assign n686 = n684 ^ n677 ;
  assign n615 = ~x2 & n446 ;
  assign n616 = n615 ^ n519 ;
  assign n617 = ~x5 & ~n616 ;
  assign n618 = n617 ^ n519 ;
  assign n619 = ~x7 & ~n618 ;
  assign n620 = n619 ^ x5 ;
  assign n627 = n341 & n401 ;
  assign n628 = n14 & n627 ;
  assign n629 = n628 ^ n14 ;
  assign n621 = n14 ^ x6 ;
  assign n630 = n629 ^ n621 ;
  assign n631 = x0 & ~n630 ;
  assign n632 = ~n620 & n631 ;
  assign n880 = n93 & n110 ;
  assign n658 = x7 & n880 ;
  assign n659 = n658 ^ x7 ;
  assign n640 = ~x2 & ~n13 ;
  assign n641 = n640 ^ n14 ;
  assign n642 = x7 ^ x2 ;
  assign n643 = n642 ^ x1 ;
  assign n644 = n641 & ~n643 ;
  assign n645 = n644 ^ x2 ;
  assign n646 = x1 & ~n645 ;
  assign n648 = n61 & n129 ;
  assign n649 = n646 & n648 ;
  assign n633 = ~x1 & n184 ;
  assign n634 = ~x2 & ~n61 ;
  assign n635 = n633 & n634 ;
  assign n636 = n635 ^ n633 ;
  assign n637 = n636 ^ x7 ;
  assign n647 = n646 ^ n637 ;
  assign n650 = n649 ^ n647 ;
  assign n660 = n659 ^ n650 ;
  assign n661 = n632 & n660 ;
  assign n687 = n686 ^ n661 ;
  assign n690 = n689 ^ n687 ;
  assign n568 = ~n100 & ~n132 ;
  assign n570 = ~n275 & n569 ;
  assign n571 = n568 & n570 ;
  assign n572 = n84 & n128 ;
  assign n580 = ~x1 & n572 ;
  assign n581 = ~n98 & n580 ;
  assign n582 = n581 ^ n98 ;
  assign n573 = n572 ^ n128 ;
  assign n574 = n573 ^ n98 ;
  assign n583 = n582 ^ n574 ;
  assign n584 = ~x4 & ~n583 ;
  assign n585 = ~n571 & n584 ;
  assign n586 = n585 ^ x5 ;
  assign n587 = x1 & n331 ;
  assign n588 = n345 & n587 ;
  assign n601 = n588 ^ n543 ;
  assign n589 = n588 ^ x1 ;
  assign n602 = ~n365 & n589 ;
  assign n603 = ~n601 & n602 ;
  assign n599 = n589 ^ x6 ;
  assign n592 = x0 & ~n93 ;
  assign n593 = ~n446 & n592 ;
  assign n594 = n593 ^ x0 ;
  assign n595 = n594 ^ n81 ;
  assign n590 = n141 ^ n81 ;
  assign n591 = ~n341 & n590 ;
  assign n596 = n595 ^ n591 ;
  assign n597 = ~n75 & ~n596 ;
  assign n600 = n599 ^ n597 ;
  assign n604 = n603 ^ n600 ;
  assign n605 = n585 & ~n604 ;
  assign n606 = n605 ^ x6 ;
  assign n607 = n586 & ~n606 ;
  assign n608 = n607 ^ x5 ;
  assign n609 = x4 & ~n20 ;
  assign n610 = n609 ^ x4 ;
  assign n611 = ~n608 & ~n610 ;
  assign n612 = ~x7 & ~n611 ;
  assign n691 = n690 ^ n612 ;
  assign n692 = ~x3 & ~x4 ;
  assign n693 = ~n691 & n692 ;
  assign n695 = n693 ^ n612 ;
  assign n765 = n12 & n352 ;
  assign n770 = ~x0 & ~n17 ;
  assign n771 = n770 ^ x3 ;
  assign n772 = n765 & ~n771 ;
  assign n736 = n232 ^ n231 ;
  assign n733 = x9 ^ x3 ;
  assign n737 = n736 ^ n733 ;
  assign n734 = n733 ^ x1 ;
  assign n735 = n734 ^ n97 ;
  assign n738 = n737 ^ n735 ;
  assign n722 = n224 ^ n99 ;
  assign n723 = n722 ^ n43 ;
  assign n724 = n723 ^ n231 ;
  assign n725 = n97 ^ x9 ;
  assign n726 = n725 ^ n723 ;
  assign n727 = n723 ^ n97 ;
  assign n728 = n727 ^ x3 ;
  assign n729 = n728 ^ n723 ;
  assign n730 = ~n726 & ~n729 ;
  assign n731 = n730 ^ n723 ;
  assign n732 = n724 & n731 ;
  assign n739 = n738 ^ n732 ;
  assign n740 = n739 ^ n97 ;
  assign n741 = n740 ^ x3 ;
  assign n742 = x8 & n741 ;
  assign n743 = n305 ^ x3 ;
  assign n744 = n743 ^ n141 ;
  assign n745 = n744 ^ n305 ;
  assign n746 = n141 ^ x8 ;
  assign n747 = n50 & n746 ;
  assign n748 = ~n745 & n747 ;
  assign n749 = n748 ^ n743 ;
  assign n750 = ~x1 & n749 ;
  assign n751 = n750 ^ n305 ;
  assign n752 = ~n742 & n751 ;
  assign n753 = ~x6 & ~n752 ;
  assign n696 = n272 ^ x1 ;
  assign n702 = ~x9 & ~n696 ;
  assign n697 = n696 ^ n12 ;
  assign n700 = n697 ^ n272 ;
  assign n701 = n142 & n700 ;
  assign n703 = n702 ^ n701 ;
  assign n704 = x8 & n703 ;
  assign n705 = n704 ^ n702 ;
  assign n706 = n705 ^ x1 ;
  assign n707 = ~x2 & n706 ;
  assign n708 = ~x1 & ~n95 ;
  assign n716 = n224 & n708 ;
  assign n717 = ~n12 & n716 ;
  assign n718 = n717 ^ n12 ;
  assign n709 = n708 ^ x1 ;
  assign n710 = n709 ^ n12 ;
  assign n719 = n718 ^ n710 ;
  assign n720 = ~n40 & n719 ;
  assign n721 = ~n707 & n720 ;
  assign n754 = n753 ^ n721 ;
  assign n755 = ~x4 & ~n754 ;
  assign n756 = n755 ^ x6 ;
  assign n757 = ~x5 & ~n756 ;
  assign n760 = n52 ^ n43 ;
  assign n761 = n80 & ~n760 ;
  assign n758 = n94 ^ x3 ;
  assign n759 = n758 ^ n388 ;
  assign n762 = n761 ^ n759 ;
  assign n763 = x1 & ~n762 ;
  assign n764 = n493 & ~n763 ;
  assign n773 = n764 & ~n772 ;
  assign n774 = n232 ^ n73 ;
  assign n775 = ~x2 & n542 ;
  assign n776 = n77 & n775 ;
  assign n777 = ~n774 & n776 ;
  assign n778 = n777 ^ n775 ;
  assign n786 = ~x3 & n778 ;
  assign n787 = ~n86 & n786 ;
  assign n788 = n787 ^ n86 ;
  assign n779 = n778 ^ x2 ;
  assign n780 = n779 ^ n86 ;
  assign n789 = n788 ^ n780 ;
  assign n790 = n773 & n789 ;
  assign n791 = ~n757 & ~n790 ;
  assign n792 = x0 & n352 ;
  assign n797 = n61 & n92 ;
  assign n798 = n797 ^ n29 ;
  assign n799 = n792 & n798 ;
  assign n800 = ~n609 & ~n799 ;
  assign n801 = ~n791 & n800 ;
  assign n802 = x7 & n801 ;
  assign n803 = ~n772 & n802 ;
  assign n804 = n803 ^ n801 ;
  assign n806 = ~n27 & ~n38 ;
  assign n807 = n806 ^ n386 ;
  assign n808 = n807 ^ n27 ;
  assign n809 = n427 ^ n143 ;
  assign n811 = n376 ^ n78 ;
  assign n810 = ~n72 & n542 ;
  assign n812 = n811 ^ n810 ;
  assign n813 = n809 & n812 ;
  assign n814 = ~x2 & ~n813 ;
  assign n815 = ~x1 & n389 ;
  assign n816 = ~n181 & n815 ;
  assign n817 = n816 ^ n517 ;
  assign n818 = ~n517 & ~n817 ;
  assign n819 = ~n814 & n818 ;
  assign n820 = n808 & n819 ;
  assign n821 = n43 & n493 ;
  assign n826 = n543 ^ n72 ;
  assign n827 = n826 ^ n810 ;
  assign n823 = n110 ^ n74 ;
  assign n824 = n823 ^ x8 ;
  assign n822 = n11 ^ x1 ;
  assign n825 = n824 ^ n822 ;
  assign n828 = n827 ^ n825 ;
  assign n829 = n821 & n828 ;
  assign n830 = ~x9 & ~n391 ;
  assign n831 = x3 & ~x5 ;
  assign n832 = x9 & ~n82 ;
  assign n833 = n832 ^ x2 ;
  assign n834 = n833 ^ x6 ;
  assign n835 = n834 ^ n832 ;
  assign n836 = ~x6 & ~n73 ;
  assign n837 = n836 ^ n832 ;
  assign n838 = ~n835 & n837 ;
  assign n839 = n838 ^ n832 ;
  assign n840 = n831 & n839 ;
  assign n841 = n840 ^ n831 ;
  assign n842 = n830 & n841 ;
  assign n850 = ~n425 & n842 ;
  assign n851 = ~n352 & n850 ;
  assign n852 = n851 ^ n352 ;
  assign n843 = n842 ^ n841 ;
  assign n844 = n843 ^ n352 ;
  assign n853 = n852 ^ n844 ;
  assign n854 = ~n829 & ~n853 ;
  assign n855 = ~n820 & n854 ;
  assign n856 = x7 & n806 ;
  assign n862 = ~x2 & ~n78 ;
  assign n857 = ~n19 & n95 ;
  assign n863 = n862 ^ n857 ;
  assign n864 = n856 & n863 ;
  assign n865 = n864 ^ x7 ;
  assign n866 = ~n855 & ~n865 ;
  assign n805 = n20 & n401 ;
  assign n867 = n866 ^ n805 ;
  assign n868 = x4 & n867 ;
  assign n869 = n868 ^ n866 ;
  assign n870 = n214 ^ x4 ;
  assign n871 = n509 ^ n508 ;
  assign n873 = ~n27 & n810 ;
  assign n872 = n539 & ~n546 ;
  assign n874 = n873 ^ n872 ;
  assign n875 = n871 & n874 ;
  assign n876 = x3 & ~x7 ;
  assign n877 = ~n875 & n876 ;
  assign n881 = ~x3 & n880 ;
  assign n878 = n504 ^ x3 ;
  assign n882 = n881 ^ n878 ;
  assign n885 = ~x2 & n541 ;
  assign n886 = n885 ^ n857 ;
  assign n887 = ~x7 & ~n886 ;
  assign n888 = n887 ^ n857 ;
  assign n889 = ~n882 & ~n888 ;
  assign n890 = n889 ^ n882 ;
  assign n891 = n27 & n133 ;
  assign n892 = ~n890 & n891 ;
  assign n901 = n343 & ~n825 ;
  assign n902 = n892 & n901 ;
  assign n903 = n902 ^ n892 ;
  assign n904 = n903 ^ n890 ;
  assign n905 = ~n877 & n904 ;
  assign n906 = ~n870 & ~n905 ;
  assign n908 = n15 & n810 ;
  assign n909 = n908 ^ n20 ;
  assign n910 = ~x4 & n909 ;
  assign n911 = n910 ^ n20 ;
  assign n912 = n90 & n911 ;
  assign y0 = ~n198 ;
  assign y1 = ~n340 ;
  assign y2 = n483 ;
  assign y3 = n558 ;
  assign y4 = n563 ;
  assign y5 = n567 ;
  assign y6 = ~n695 ;
  assign y7 = ~n804 ;
  assign y8 = ~n869 ;
  assign y9 = n906 ;
  assign y10 = n912 ;
endmodule
