module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n368 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n760 , n761 , n762 , n763 , n764 , n765 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n900 , n903 , n904 , n905 , n906 , n907 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n920 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n954 , n955 , n956 , n957 , n958 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n976 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1241 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1252 , n1256 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1300 , n1301 , n1304 , n1305 , n1306 , n1307 , n1308 , n1311 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1322 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1356 , n1357 , n1358 , n1359 , n1360 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1375 , n1376 , n1377 , n1378 , n1379 , n1382 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1392 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1427 , n1428 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1455 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1501 , n1503 , n1504 , n1505 , n1506 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1539 , n1542 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1555 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1569 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1587 , n1588 , n1589 , n1591 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1606 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1645 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1665 , n1666 , n1667 , n1668 , n1669 , n1672 , n1675 , n1676 , n1677 , n1678 , n1679 , n1682 , n1683 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1699 , n1704 , n1705 , n1706 , n1707 , n1709 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1771 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1816 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1847 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1913 , n1918 , n1919 , n1920 , n1921 , n1923 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1949 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1968 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2003 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2016 , n2020 , n2022 , n2024 , n2025 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2041 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2079 , n2080 , n2081 , n2082 , n2083 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2363 , n2364 , n2365 , n2366 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2773 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2787 , n2788 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3061 , n3066 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3079 , n3080 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3170 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3544 , n3545 , n3546 , n3547 , n3548 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4162 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4268 , n4269 , n4270 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4412 , n4413 , n4414 , n4415 , n4416 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4818 , n4820 , n4821 , n4822 , n4825 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4986 , n4987 , n4988 , n4989 , n4992 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5077 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5120 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5694 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5854 , n5855 , n5856 , n5857 , n5858 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6049 , n6050 , n6053 , n6056 , n6057 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6069 , n6070 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 ;
  assign n58 = x19 & ~x22 ;
  assign n43 = ~x16 & x17 ;
  assign n44 = n43 ^ x16 ;
  assign n45 = x18 & ~x19 ;
  assign n46 = n45 ^ x18 ;
  assign n103 = ~n44 & n46 ;
  assign n84 = x17 ^ x16 ;
  assign n25 = ~x12 & ~x13 ;
  assign n26 = ~x14 & n25 ;
  assign n27 = ~x6 & ~x7 ;
  assign n28 = x2 ^ x1 ;
  assign n29 = ~x0 & x1 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = ~n28 & ~n30 ;
  assign n32 = ~x3 & n31 ;
  assign n33 = ~x4 & n32 ;
  assign n34 = ~x5 & n33 ;
  assign n35 = n27 & n34 ;
  assign n36 = ~x8 & n35 ;
  assign n37 = ~x9 & n36 ;
  assign n38 = ~x10 & n37 ;
  assign n39 = ~x11 & n38 ;
  assign n40 = n26 & n39 ;
  assign n50 = ~x15 & n40 ;
  assign n85 = n50 ^ x17 ;
  assign n86 = ~n84 & n85 ;
  assign n96 = n50 ^ x18 ;
  assign n97 = ~x22 & ~n96 ;
  assign n98 = n86 & n97 ;
  assign n104 = n103 ^ n98 ;
  assign n105 = ~n58 & n104 ;
  assign n41 = ~x22 & ~n40 ;
  assign n42 = n41 ^ x15 ;
  assign n47 = n46 ^ x19 ;
  assign n48 = n47 ^ x18 ;
  assign n49 = ~n44 & ~n48 ;
  assign n51 = ~x22 & ~n50 ;
  assign n52 = n49 & ~n51 ;
  assign n53 = ~x22 & ~n52 ;
  assign n54 = n53 ^ x20 ;
  assign n76 = x22 ^ x21 ;
  assign n77 = n54 & ~n76 ;
  assign n78 = ~n42 & ~n77 ;
  assign n79 = n78 ^ n42 ;
  assign n80 = n79 ^ n77 ;
  assign n55 = n42 & ~n54 ;
  assign n56 = n55 ^ n42 ;
  assign n125 = n80 ^ n56 ;
  assign n124 = n77 ^ n54 ;
  assign n126 = n125 ^ n124 ;
  assign n585 = n105 & ~n126 ;
  assign n65 = n50 ^ x16 ;
  assign n66 = ~x17 & ~n65 ;
  assign n67 = n66 ^ n65 ;
  assign n69 = ~x18 & n58 ;
  assign n70 = n69 ^ n47 ;
  assign n68 = n58 ^ x19 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n46 ;
  assign n73 = ~n67 & n72 ;
  assign n57 = n44 ^ x17 ;
  assign n60 = x22 & n45 ;
  assign n61 = n60 ^ n45 ;
  assign n59 = n58 ^ x22 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n62 ^ n48 ;
  assign n64 = n57 & n63 ;
  assign n74 = n73 ^ n64 ;
  assign n116 = n42 & ~n76 ;
  assign n117 = n116 ^ n80 ;
  assign n90 = x21 ^ x20 ;
  assign n109 = n53 ^ x21 ;
  assign n110 = n90 & n109 ;
  assign n140 = n117 ^ n110 ;
  assign n362 = n74 & ~n140 ;
  assign n2319 = n585 ^ n362 ;
  assign n213 = ~n62 & ~n67 ;
  assign n212 = n57 & n71 ;
  assign n214 = n213 ^ n212 ;
  assign n604 = n110 & n214 ;
  assign n284 = ~n117 & n214 ;
  assign n605 = n604 ^ n284 ;
  assign n91 = n76 & ~n90 ;
  assign n92 = ~n42 & n91 ;
  assign n172 = n61 & n66 ;
  assign n111 = n57 ^ x16 ;
  assign n171 = n70 & n111 ;
  assign n173 = n172 ^ n171 ;
  assign n308 = n92 & n173 ;
  assign n180 = n77 & n173 ;
  assign n175 = n78 & n173 ;
  assign n174 = ~n42 & n173 ;
  assign n176 = n175 ^ n174 ;
  assign n181 = n180 ^ n176 ;
  assign n309 = n308 ^ n181 ;
  assign n306 = n92 ^ n56 ;
  assign n307 = n173 & n306 ;
  assign n310 = n309 ^ n307 ;
  assign n2318 = n605 ^ n310 ;
  assign n2320 = n2319 ^ n2318 ;
  assign n793 = ~n126 & n214 ;
  assign n152 = ~n50 & n111 ;
  assign n153 = n72 & n152 ;
  assign n154 = n153 ^ n52 ;
  assign n262 = n154 ^ n117 ;
  assign n261 = n117 & ~n154 ;
  assign n263 = n262 ^ n261 ;
  assign n1089 = n793 ^ n263 ;
  assign n143 = ~n67 & n69 ;
  assign n142 = n57 & n60 ;
  assign n144 = n143 ^ n142 ;
  assign n288 = ~n126 & n144 ;
  assign n87 = n86 ^ n65 ;
  assign n88 = n72 & n87 ;
  assign n83 = n43 & n63 ;
  assign n89 = n88 ^ n83 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n89 & n93 ;
  assign n289 = n288 ^ n94 ;
  assign n2317 = n1089 ^ n289 ;
  assign n2321 = n2320 ^ n2317 ;
  assign n184 = x19 & n98 ;
  assign n183 = ~n44 & n60 ;
  assign n185 = n184 ^ n183 ;
  assign n337 = n92 & n185 ;
  assign n296 = n89 & n92 ;
  assign n2485 = n337 ^ n296 ;
  assign n240 = n61 & ~n67 ;
  assign n239 = n57 & n70 ;
  assign n241 = n240 ^ n239 ;
  assign n467 = n77 & n241 ;
  assign n242 = ~n42 & n241 ;
  assign n304 = n77 & n242 ;
  assign n468 = n467 ^ n304 ;
  assign n3681 = n2485 ^ n468 ;
  assign n2260 = n105 & ~n125 ;
  assign n3682 = n3681 ^ n2260 ;
  assign n335 = n74 & ~n117 ;
  assign n113 = n66 & n72 ;
  assign n112 = n63 & n111 ;
  assign n114 = n113 ^ n112 ;
  assign n279 = n92 & n114 ;
  assign n783 = n335 ^ n279 ;
  assign n122 = ~n62 & n87 ;
  assign n121 = n43 & n71 ;
  assign n123 = n122 ^ n121 ;
  assign n434 = ~n79 & n123 ;
  assign n3680 = n783 ^ n434 ;
  assign n3683 = n3682 ^ n3680 ;
  assign n349 = n74 & n91 ;
  assign n3675 = n349 ^ n154 ;
  assign n344 = ~n140 & n173 ;
  assign n343 = n308 ^ n175 ;
  assign n345 = n344 ^ n343 ;
  assign n3676 = n3675 ^ n345 ;
  assign n488 = n77 & n214 ;
  assign n3677 = n3676 ^ n488 ;
  assign n158 = n66 & n69 ;
  assign n157 = n60 & n111 ;
  assign n159 = n158 ^ n157 ;
  assign n594 = n185 ^ n159 ;
  assign n595 = n77 & n594 ;
  assign n315 = ~n44 & ~n51 ;
  assign n316 = n47 & n315 ;
  assign n314 = n61 & n152 ;
  assign n317 = n316 ^ n314 ;
  assign n592 = n317 ^ n241 ;
  assign n593 = n110 & n592 ;
  assign n596 = n595 ^ n593 ;
  assign n3678 = n3677 ^ n596 ;
  assign n136 = n69 & n87 ;
  assign n135 = n43 & n60 ;
  assign n137 = n136 ^ n135 ;
  assign n276 = ~n80 & n137 ;
  assign n210 = ~n62 & n66 ;
  assign n209 = n71 & n111 ;
  assign n211 = n210 ^ n209 ;
  assign n260 = ~n117 & n211 ;
  assign n1002 = n276 ^ n260 ;
  assign n446 = n125 & ~n137 ;
  assign n445 = n137 ^ n125 ;
  assign n447 = n446 ^ n445 ;
  assign n278 = n91 & n114 ;
  assign n280 = n279 ^ n278 ;
  assign n862 = n447 ^ n280 ;
  assign n3674 = n1002 ^ n862 ;
  assign n3679 = n3678 ^ n3674 ;
  assign n3684 = n3683 ^ n3679 ;
  assign n3685 = ~n2321 & ~n3684 ;
  assign n548 = n74 & ~n79 ;
  assign n354 = n105 & ~n140 ;
  assign n3687 = n548 ^ n354 ;
  assign n138 = ~n42 & n137 ;
  assign n831 = n124 & n138 ;
  assign n404 = n56 ^ n54 ;
  assign n411 = n159 & n404 ;
  assign n410 = ~n79 & n159 ;
  assign n412 = n411 ^ n410 ;
  assign n2422 = n831 ^ n412 ;
  assign n417 = ~n125 & n144 ;
  assign n2423 = n2422 ^ n417 ;
  assign n230 = ~n92 & ~n159 ;
  assign n293 = n125 & n230 ;
  assign n292 = n230 ^ n125 ;
  assign n294 = n293 ^ n292 ;
  assign n249 = ~n125 & n211 ;
  assign n1225 = n294 ^ n249 ;
  assign n3686 = n2423 ^ n1225 ;
  assign n3688 = n3687 ^ n3686 ;
  assign n607 = n105 & ~n117 ;
  assign n608 = n607 ^ n284 ;
  assign n132 = n61 & n87 ;
  assign n131 = n43 & n70 ;
  assign n133 = n132 ^ n131 ;
  assign n331 = ~n80 & n133 ;
  assign n609 = n608 ^ n331 ;
  assign n168 = n77 & n114 ;
  assign n610 = n609 ^ n168 ;
  assign n170 = ~n79 & n133 ;
  assign n177 = n176 ^ n170 ;
  assign n611 = n610 ^ n177 ;
  assign n3689 = n3688 ^ n611 ;
  assign n251 = ~n79 & n154 ;
  assign n155 = ~n80 & n154 ;
  assign n408 = n251 ^ n155 ;
  assign n405 = ~n77 & n154 ;
  assign n406 = ~n404 & n405 ;
  assign n407 = n406 ^ n154 ;
  assign n409 = n408 ^ n407 ;
  assign n215 = n214 ^ n211 ;
  assign n216 = n215 ^ n123 ;
  assign n217 = n92 & ~n216 ;
  assign n397 = n217 ^ n92 ;
  assign n507 = n409 ^ n397 ;
  assign n502 = n123 ^ n105 ;
  assign n503 = n42 & n502 ;
  assign n504 = n93 & ~n216 ;
  assign n505 = ~n503 & n504 ;
  assign n506 = n505 ^ n93 ;
  assign n508 = n507 ^ n506 ;
  assign n500 = n185 ^ n144 ;
  assign n501 = n110 & n500 ;
  assign n509 = n508 ^ n501 ;
  assign n568 = n417 ^ n144 ;
  assign n524 = n125 & ~n185 ;
  assign n569 = n568 ^ n524 ;
  assign n570 = ~n261 & ~n569 ;
  assign n571 = ~n509 & ~n570 ;
  assign n3690 = n3689 ^ n571 ;
  assign n3691 = n3685 & ~n3690 ;
  assign n472 = n74 & ~n126 ;
  assign n81 = n74 & ~n80 ;
  assign n75 = n56 & n74 ;
  assign n82 = n81 ^ n75 ;
  assign n1163 = n472 ^ n82 ;
  assign n838 = n110 & n137 ;
  assign n267 = ~n117 & n137 ;
  assign n839 = n838 ^ n267 ;
  assign n1164 = n1163 ^ n839 ;
  assign n664 = ~n79 & n105 ;
  assign n225 = ~n80 & n211 ;
  assign n224 = n77 & n211 ;
  assign n226 = n225 ^ n224 ;
  assign n1012 = n664 ^ n226 ;
  assign n1013 = n1012 ^ n434 ;
  assign n2265 = n1164 ^ n1013 ;
  assign n526 = n317 ^ n93 ;
  assign n525 = n93 & n317 ;
  assign n527 = n526 ^ n525 ;
  assign n843 = ~n446 & n527 ;
  assign n229 = n159 ^ n92 ;
  assign n231 = n230 ^ n229 ;
  assign n228 = n91 & n159 ;
  assign n232 = n231 ^ n228 ;
  assign n2264 = n843 ^ n232 ;
  assign n2266 = n2265 ^ n2264 ;
  assign n201 = ~n80 & n144 ;
  assign n200 = n77 & n144 ;
  assign n202 = n201 ^ n200 ;
  assign n2261 = n2260 ^ n202 ;
  assign n2262 = n2261 ^ n407 ;
  assign n829 = n570 ^ n94 ;
  assign n2263 = n2262 ^ n829 ;
  assign n2267 = n2266 ^ n2263 ;
  assign n674 = n92 & n137 ;
  assign n654 = n56 & n214 ;
  assign n245 = ~n80 & n214 ;
  assign n655 = n654 ^ n245 ;
  assign n2258 = n674 ^ n655 ;
  assign n383 = ~n117 & n123 ;
  assign n574 = n383 ^ n123 ;
  assign n127 = n126 ^ n117 ;
  assign n128 = n123 & ~n127 ;
  assign n575 = n574 ^ n128 ;
  assign n478 = n110 & n317 ;
  assign n473 = ~n117 & n317 ;
  assign n479 = n478 ^ n473 ;
  assign n850 = n575 ^ n479 ;
  assign n2256 = n850 ^ n383 ;
  assign n2257 = n2256 ^ n417 ;
  assign n2259 = n2258 ^ n2257 ;
  assign n2268 = n2267 ^ n2259 ;
  assign n1032 = ~n140 & n159 ;
  assign n391 = n93 & n211 ;
  assign n390 = n91 & n211 ;
  assign n392 = n391 ^ n390 ;
  assign n2252 = n1032 ^ n392 ;
  assign n452 = ~n110 & ~n185 ;
  assign n451 = n185 ^ n110 ;
  assign n453 = n452 ^ n451 ;
  assign n399 = n93 & n185 ;
  assign n851 = n453 ^ n399 ;
  assign n553 = ~n117 & n185 ;
  assign n852 = n851 ^ n553 ;
  assign n2253 = n2252 ^ n852 ;
  assign n511 = n56 & n317 ;
  assign n444 = ~n125 & n317 ;
  assign n512 = n511 ^ n444 ;
  assign n429 = n77 & n89 ;
  assign n179 = ~n80 & n89 ;
  assign n430 = n429 ^ n179 ;
  assign n2250 = n512 ^ n430 ;
  assign n2251 = n2250 ^ n294 ;
  assign n2254 = n2253 ^ n2251 ;
  assign n107 = ~n93 & ~n105 ;
  assign n106 = n105 ^ n93 ;
  assign n108 = n107 ^ n106 ;
  assign n363 = n362 ^ n108 ;
  assign n359 = n140 ^ n92 ;
  assign n360 = n144 & ~n359 ;
  assign n358 = n89 & ~n126 ;
  assign n361 = n360 ^ n358 ;
  assign n364 = n363 ^ n361 ;
  assign n323 = n92 & n214 ;
  assign n353 = n323 ^ n279 ;
  assign n355 = n354 ^ n353 ;
  assign n348 = n74 & n92 ;
  assign n350 = n349 ^ n348 ;
  assign n265 = n89 & ~n125 ;
  assign n351 = n350 ^ n265 ;
  assign n352 = n351 ^ n249 ;
  assign n356 = n355 ^ n352 ;
  assign n341 = ~n117 & n173 ;
  assign n342 = n341 ^ n310 ;
  assign n346 = n345 ^ n342 ;
  assign n286 = n123 & ~n140 ;
  assign n347 = n346 ^ n286 ;
  assign n357 = n356 ^ n347 ;
  assign n365 = n364 ^ n357 ;
  assign n2255 = n2254 ^ n365 ;
  assign n2269 = n2268 ^ n2255 ;
  assign n2281 = n267 ^ n177 ;
  assign n881 = n391 ^ n310 ;
  assign n162 = n116 & n159 ;
  assign n882 = n881 ^ n162 ;
  assign n877 = ~n92 & ~n124 ;
  assign n876 = n124 ^ n92 ;
  assign n878 = n877 ^ n876 ;
  assign n270 = ~n42 & ~n114 ;
  assign n271 = ~n124 & n270 ;
  assign n272 = n271 ^ n270 ;
  assign n273 = n272 ^ n126 ;
  assign n879 = n878 ^ n273 ;
  assign n880 = n879 ^ n308 ;
  assign n883 = n882 ^ n880 ;
  assign n2282 = n2281 ^ n883 ;
  assign n543 = ~n125 & n241 ;
  assign n2278 = n607 ^ n543 ;
  assign n1483 = n335 ^ n296 ;
  assign n2279 = n2278 ^ n1483 ;
  assign n312 = ~n126 & n211 ;
  assign n303 = n77 & n138 ;
  assign n2275 = n312 ^ n303 ;
  assign n2276 = n2275 ^ n412 ;
  assign n334 = n93 & n241 ;
  assign n283 = n110 & n242 ;
  assign n2273 = n334 ^ n283 ;
  assign n2274 = n2273 ^ n288 ;
  assign n2277 = n2276 ^ n2274 ;
  assign n2280 = n2279 ^ n2277 ;
  assign n2283 = n2282 ^ n2280 ;
  assign n167 = ~n80 & n114 ;
  assign n2270 = n468 ^ n167 ;
  assign n2271 = n2270 ^ n525 ;
  assign n489 = n488 ^ n245 ;
  assign n799 = n489 ^ n473 ;
  assign n2272 = n2271 ^ n799 ;
  assign n2284 = n2283 ^ n2272 ;
  assign n2285 = ~n2269 & ~n2284 ;
  assign n588 = n260 ^ n77 ;
  assign n597 = n596 ^ n267 ;
  assign n589 = n173 ^ n159 ;
  assign n590 = n589 ^ n133 ;
  assign n591 = n110 & n590 ;
  assign n598 = n597 ^ n591 ;
  assign n599 = ~n588 & ~n598 ;
  assign n606 = n605 ^ n354 ;
  assign n612 = n611 ^ n606 ;
  assign n515 = ~n105 & ~n110 ;
  assign n600 = n515 ^ n181 ;
  assign n601 = n123 ^ n77 ;
  assign n247 = n140 ^ n125 ;
  assign n248 = n211 & n247 ;
  assign n250 = n249 ^ n248 ;
  assign n602 = n601 ^ n250 ;
  assign n603 = ~n600 & n602 ;
  assign n613 = n612 ^ n603 ;
  assign n614 = n599 & ~n613 ;
  assign n481 = n92 & n144 ;
  assign n455 = n144 ^ n93 ;
  assign n190 = ~n93 & ~n144 ;
  assign n456 = n455 ^ n190 ;
  assign n650 = n481 ^ n456 ;
  assign n651 = n650 ^ n360 ;
  assign n118 = n114 & ~n117 ;
  assign n115 = n110 & n114 ;
  assign n119 = n118 ^ n115 ;
  assign n649 = n456 ^ n119 ;
  assign n652 = n651 ^ n649 ;
  assign n653 = n652 ^ n354 ;
  assign n656 = n655 ^ n653 ;
  assign n318 = n92 & n317 ;
  assign n421 = n318 ^ n286 ;
  assign n134 = ~n42 & ~n133 ;
  assign n145 = n144 ^ n133 ;
  assign n146 = ~n134 & n145 ;
  assign n147 = n127 & n146 ;
  assign n422 = n421 ^ n147 ;
  assign n657 = n656 ^ n422 ;
  assign n547 = n317 & n404 ;
  assign n319 = n92 ^ n79 ;
  assign n320 = n317 & ~n319 ;
  assign n321 = n320 ^ n318 ;
  assign n646 = n547 ^ n321 ;
  assign n644 = n185 ^ n125 ;
  assign n645 = n644 ^ n524 ;
  assign n647 = n646 ^ n645 ;
  assign n642 = n93 & n133 ;
  assign n243 = n124 & n242 ;
  assign n641 = n243 ^ n226 ;
  assign n643 = n642 ^ n641 ;
  assign n648 = n647 ^ n643 ;
  assign n658 = n657 ^ n648 ;
  assign n566 = n92 & n105 ;
  assign n637 = n566 ^ n249 ;
  assign n638 = n637 ^ n276 ;
  assign n639 = n638 ^ n118 ;
  assign n635 = n341 ^ n321 ;
  assign n636 = n635 ^ n553 ;
  assign n640 = n639 ^ n636 ;
  assign n659 = n658 ^ n640 ;
  assign n385 = n123 & ~n125 ;
  assign n386 = n385 ^ n288 ;
  assign n305 = n304 ^ n303 ;
  assign n387 = n386 ^ n305 ;
  assign n384 = n383 ^ n177 ;
  assign n388 = n387 ^ n384 ;
  assign n161 = ~n117 & n159 ;
  assign n163 = n162 ^ n161 ;
  assign n160 = n159 ^ n80 ;
  assign n164 = n163 ^ n160 ;
  assign n379 = n93 & n123 ;
  assign n378 = n123 ^ n93 ;
  assign n380 = n379 ^ n378 ;
  assign n381 = ~n164 & n380 ;
  assign n624 = n388 ^ n381 ;
  assign n623 = n575 ^ n489 ;
  assign n625 = n624 ^ n623 ;
  assign n534 = ~n77 & ~n137 ;
  assign n619 = n468 ^ n230 ;
  assign n620 = n619 ^ n228 ;
  assign n621 = n620 ^ n91 ;
  assign n622 = ~n534 & ~n621 ;
  assign n626 = n625 ^ n622 ;
  assign n631 = n312 ^ n231 ;
  assign n632 = n631 ^ n279 ;
  assign n628 = n607 ^ n575 ;
  assign n414 = ~n126 & n185 ;
  assign n629 = n628 ^ n414 ;
  assign n627 = n511 ^ n409 ;
  assign n630 = n629 ^ n627 ;
  assign n633 = n632 ^ n630 ;
  assign n634 = ~n626 & n633 ;
  assign n660 = n659 ^ n634 ;
  assign n683 = n434 ^ n296 ;
  assign n681 = n225 ^ n181 ;
  assign n682 = n681 ^ n331 ;
  assign n684 = n683 ^ n682 ;
  assign n678 = n114 & ~n125 ;
  assign n679 = n678 ^ n391 ;
  assign n680 = n679 ^ n280 ;
  assign n685 = n684 ^ n680 ;
  assign n675 = n674 ^ n200 ;
  assign n676 = n675 ^ n94 ;
  assign n449 = n93 & n173 ;
  assign n673 = n449 ^ n392 ;
  assign n677 = n676 ^ n673 ;
  assign n686 = n685 ^ n677 ;
  assign n668 = ~n125 & n154 ;
  assign n254 = n80 & ~n105 ;
  assign n255 = n254 ^ n77 ;
  assign n253 = n105 ^ n79 ;
  assign n256 = n255 ^ n253 ;
  assign n669 = n668 ^ n256 ;
  assign n670 = n669 ^ n308 ;
  assign n666 = n553 ^ n344 ;
  assign n667 = n666 ^ n453 ;
  assign n671 = n670 ^ n667 ;
  assign n663 = n543 ^ n245 ;
  assign n665 = n664 ^ n663 ;
  assign n672 = n671 ^ n665 ;
  assign n687 = n686 ^ n672 ;
  assign n661 = n214 ^ n138 ;
  assign n662 = n110 & n661 ;
  assign n688 = n687 ^ n662 ;
  assign n689 = n660 & n688 ;
  assign n495 = n362 ^ n260 ;
  assign n496 = n495 ^ n391 ;
  assign n494 = n331 ^ n201 ;
  assign n497 = n496 ^ n494 ;
  assign n394 = n89 & ~n140 ;
  assign n492 = n430 ^ n394 ;
  assign n192 = n93 & n137 ;
  assign n493 = n492 ^ n192 ;
  assign n498 = n497 ^ n493 ;
  assign n490 = n489 ^ n335 ;
  assign n491 = n490 ^ n167 ;
  assign n499 = n498 ^ n491 ;
  assign n252 = n251 ^ n250 ;
  assign n257 = n256 ^ n252 ;
  assign n237 = n42 & n89 ;
  assign n238 = n110 & n237 ;
  assign n244 = n243 ^ n238 ;
  assign n246 = n245 ^ n244 ;
  assign n258 = n257 ^ n246 ;
  assign n234 = n159 ^ n137 ;
  assign n235 = ~n125 & n234 ;
  assign n227 = n226 ^ n176 ;
  assign n233 = n232 ^ n227 ;
  assign n236 = n235 ^ n233 ;
  assign n259 = n258 ^ n236 ;
  assign n510 = n509 ^ n259 ;
  assign n516 = n154 ^ n79 ;
  assign n517 = n516 ^ n251 ;
  assign n518 = ~n515 & ~n517 ;
  assign n519 = n518 ^ n323 ;
  assign n418 = n417 ^ n118 ;
  assign n520 = n519 ^ n418 ;
  assign n513 = n512 ^ n410 ;
  assign n514 = n513 ^ n231 ;
  assign n521 = n520 ^ n514 ;
  assign n522 = n510 & n521 ;
  assign n523 = ~n499 & n522 ;
  assign n120 = n119 ^ n108 ;
  assign n552 = n337 ^ n120 ;
  assign n554 = n553 ^ n552 ;
  assign n550 = n456 ^ n263 ;
  assign n549 = n548 ^ n547 ;
  assign n551 = n550 ^ n549 ;
  assign n555 = n554 ^ n551 ;
  assign n541 = n410 ^ n251 ;
  assign n542 = n541 ^ n202 ;
  assign n544 = n543 ^ n542 ;
  assign n539 = n159 ^ n154 ;
  assign n540 = n77 & n539 ;
  assign n545 = n544 ^ n540 ;
  assign n396 = n392 ^ n323 ;
  assign n398 = n397 ^ n396 ;
  assign n530 = n398 ^ n138 ;
  assign n532 = n241 ^ n77 ;
  assign n533 = n532 ^ n467 ;
  assign n535 = n534 ^ n533 ;
  assign n531 = n241 ^ n137 ;
  assign n536 = n535 ^ n531 ;
  assign n537 = ~n530 & n536 ;
  assign n528 = n527 ^ n154 ;
  assign n529 = ~n524 & n528 ;
  assign n538 = n537 ^ n529 ;
  assign n546 = n545 ^ n538 ;
  assign n556 = n555 ^ n546 ;
  assign n558 = n318 ^ n294 ;
  assign n291 = ~n126 & n133 ;
  assign n557 = n291 ^ n225 ;
  assign n559 = n558 ^ n557 ;
  assign n188 = n159 ^ n123 ;
  assign n189 = n188 ^ n140 ;
  assign n191 = n190 ^ n137 ;
  assign n193 = n192 ^ n191 ;
  assign n194 = ~n189 & ~n193 ;
  assign n186 = ~n80 & n185 ;
  assign n182 = n181 ^ n179 ;
  assign n187 = n186 ^ n182 ;
  assign n195 = n194 ^ n187 ;
  assign n169 = n168 ^ n167 ;
  assign n178 = n177 ^ n169 ;
  assign n196 = n195 ^ n178 ;
  assign n199 = n144 ^ n79 ;
  assign n203 = n202 ^ n199 ;
  assign n219 = n185 ^ n123 ;
  assign n205 = n114 ^ n89 ;
  assign n204 = n154 ^ n74 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n110 & n206 ;
  assign n208 = n207 ^ n110 ;
  assign n218 = n217 ^ n208 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = ~n203 & n220 ;
  assign n222 = ~n196 & n221 ;
  assign n139 = n138 ^ n134 ;
  assign n141 = n140 ^ n81 ;
  assign n148 = n147 ^ n141 ;
  assign n149 = ~n139 & ~n148 ;
  assign n129 = n128 ^ n120 ;
  assign n95 = n94 ^ n82 ;
  assign n130 = n129 ^ n95 ;
  assign n150 = n149 ^ n130 ;
  assign n151 = n150 ^ n126 ;
  assign n156 = n155 ^ n154 ;
  assign n165 = n164 ^ n156 ;
  assign n166 = n151 & ~n165 ;
  assign n197 = n196 ^ n166 ;
  assign n223 = n222 ^ n197 ;
  assign n560 = n559 ^ n223 ;
  assign n561 = n556 & n560 ;
  assign n562 = n523 & n561 ;
  assign n746 = n689 ^ n562 ;
  assign n701 = ~x12 & ~x22 ;
  assign n702 = n39 & n701 ;
  assign n703 = n702 ^ x22 ;
  assign n705 = x13 & ~x22 ;
  assign n706 = n703 & n705 ;
  assign n704 = n703 ^ x14 ;
  assign n707 = n706 ^ n704 ;
  assign n567 = n566 ^ n525 ;
  assign n572 = n571 ^ n567 ;
  assign n563 = n241 ^ n173 ;
  assign n564 = n563 ^ n133 ;
  assign n565 = n91 & n564 ;
  assign n573 = n572 ^ n565 ;
  assign n581 = n214 ^ n173 ;
  assign n582 = n581 ^ n503 ;
  assign n583 = n124 & n582 ;
  assign n584 = n583 ^ n312 ;
  assign n586 = n585 ^ n584 ;
  assign n579 = ~n140 & n206 ;
  assign n577 = ~n125 & n133 ;
  assign n576 = n575 ^ n249 ;
  assign n578 = n577 ^ n576 ;
  assign n580 = n579 ^ n578 ;
  assign n587 = n586 ^ n580 ;
  assign n615 = n110 & n614 ;
  assign n616 = ~n587 & n615 ;
  assign n617 = n616 ^ n587 ;
  assign n618 = n573 & ~n617 ;
  assign n747 = n707 ^ n618 ;
  assign n748 = n618 ^ n562 ;
  assign n749 = n747 & n748 ;
  assign n750 = n749 ^ n618 ;
  assign n751 = ~n746 & ~n750 ;
  assign n752 = n751 ^ n618 ;
  assign n690 = ~n618 & ~n689 ;
  assign n691 = ~n562 & n690 ;
  assign n692 = n691 ^ n618 ;
  assign n695 = ~x22 & ~n39 ;
  assign n696 = n695 ^ x12 ;
  assign n693 = ~x22 & ~n38 ;
  assign n694 = n693 ^ x11 ;
  assign n697 = n696 ^ n694 ;
  assign n698 = ~n614 & n697 ;
  assign n699 = n692 & n698 ;
  assign n700 = n699 ^ n692 ;
  assign n708 = n703 ^ x13 ;
  assign n760 = ~n700 & n708 ;
  assign n710 = ~n124 & n618 ;
  assign n713 = n710 ^ n614 ;
  assign n714 = ~n708 & n713 ;
  assign n709 = n708 ^ n707 ;
  assign n711 = n709 & ~n710 ;
  assign n712 = ~n617 & n711 ;
  assign n715 = n714 ^ n712 ;
  assign n716 = n715 ^ n614 ;
  assign n737 = n713 ^ n617 ;
  assign n738 = ~n708 & n737 ;
  assign n721 = n710 ^ n696 ;
  assign n739 = n738 ^ n721 ;
  assign n1252 = n617 ^ n614 ;
  assign n740 = n739 & n1252 ;
  assign n741 = n740 ^ n721 ;
  assign n757 = n716 & ~n741 ;
  assign n761 = n760 ^ n757 ;
  assign n762 = n752 & n761 ;
  assign n763 = n762 ^ n757 ;
  assign n764 = ~n614 & n763 ;
  assign n718 = n716 ^ n700 ;
  assign n753 = ~n741 & n752 ;
  assign n754 = ~n718 & n753 ;
  assign n717 = ~n700 & n716 ;
  assign n2245 = n754 ^ n717 ;
  assign n2246 = ~n764 & ~n2245 ;
  assign n2243 = ~n617 & ~n707 ;
  assign n2244 = n2243 ^ n707 ;
  assign n2247 = n2246 ^ n2244 ;
  assign n2239 = n694 & n696 ;
  assign n2240 = n2239 ^ n697 ;
  assign n2241 = n2240 ^ n709 ;
  assign n2242 = ~n614 & ~n2241 ;
  assign n2248 = n2247 ^ n2242 ;
  assign n939 = n752 ^ n741 ;
  assign n779 = ~x22 & ~n37 ;
  assign n780 = n779 ^ x10 ;
  assign n777 = ~x22 & ~n36 ;
  assign n778 = n777 ^ x9 ;
  assign n781 = n780 ^ n778 ;
  assign n817 = n398 ^ n331 ;
  assign n818 = n817 ^ n637 ;
  assign n274 = n133 & ~n140 ;
  assign n377 = n312 ^ n274 ;
  assign n816 = n492 ^ n377 ;
  assign n819 = n818 ^ n816 ;
  assign n809 = n665 ^ n605 ;
  assign n808 = n383 ^ n334 ;
  assign n810 = n809 ^ n808 ;
  assign n807 = n273 ^ n254 ;
  assign n811 = n810 ^ n807 ;
  assign n820 = n819 ^ n811 ;
  assign n813 = n241 ^ n114 ;
  assign n814 = ~n127 & ~n813 ;
  assign n815 = n807 & n814 ;
  assign n821 = n820 ^ n815 ;
  assign n802 = n358 ^ n350 ;
  assign n803 = n802 ^ n669 ;
  assign n427 = ~n117 & n241 ;
  assign n800 = n799 ^ n427 ;
  assign n450 = n449 ^ n283 ;
  assign n801 = n800 ^ n450 ;
  assign n804 = n803 ^ n801 ;
  assign n796 = n284 ^ n224 ;
  assign n797 = n796 ^ n645 ;
  assign n794 = n793 ^ n286 ;
  assign n791 = n93 & n214 ;
  assign n792 = n791 ^ n280 ;
  assign n795 = n794 ^ n792 ;
  assign n798 = n797 ^ n795 ;
  assign n805 = n804 ^ n798 ;
  assign n787 = n159 ^ n105 ;
  assign n788 = n787 ^ n89 ;
  assign n789 = ~n125 & n788 ;
  assign n785 = n386 ^ n348 ;
  assign n457 = n456 ^ n238 ;
  assign n330 = n92 & n133 ;
  assign n782 = n457 ^ n330 ;
  assign n784 = n783 ^ n782 ;
  assign n786 = n785 ^ n784 ;
  assign n790 = n789 ^ n786 ;
  assign n806 = n805 ^ n790 ;
  assign n822 = n821 ^ n806 ;
  assign n823 = n560 & n822 ;
  assign n832 = n831 ^ n243 ;
  assign n833 = n832 ^ n379 ;
  assign n834 = n833 ^ n320 ;
  assign n835 = n834 ^ n82 ;
  assign n828 = n789 ^ n304 ;
  assign n830 = n829 ^ n828 ;
  assign n836 = n835 ^ n830 ;
  assign n825 = n427 ^ n341 ;
  assign n826 = n825 ^ n291 ;
  assign n824 = n398 ^ n350 ;
  assign n827 = n826 ^ n824 ;
  assign n837 = n836 ^ n827 ;
  assign n853 = n852 ^ n850 ;
  assign n849 = n456 ^ n249 ;
  assign n854 = n853 ^ n849 ;
  assign n845 = n92 & n241 ;
  assign n846 = n845 ^ n288 ;
  assign n847 = n846 ^ n169 ;
  assign n844 = n843 ^ n323 ;
  assign n848 = n847 ^ n844 ;
  assign n855 = n854 ^ n848 ;
  assign n840 = n839 ^ n354 ;
  assign n841 = n840 ^ n274 ;
  assign n842 = n841 ^ n514 ;
  assign n856 = n855 ^ n842 ;
  assign n865 = n237 ^ n123 ;
  assign n864 = n362 ^ n284 ;
  assign n866 = n865 ^ n864 ;
  assign n867 = n110 & n866 ;
  assign n858 = ~n79 & n185 ;
  assign n859 = n858 ^ n548 ;
  assign n860 = n859 ^ n155 ;
  assign n857 = n288 ^ n186 ;
  assign n861 = n860 ^ n857 ;
  assign n863 = n862 ^ n861 ;
  assign n868 = n867 ^ n863 ;
  assign n872 = n566 ^ n330 ;
  assign n873 = n872 ^ n793 ;
  assign n871 = n414 ^ n167 ;
  assign n874 = n873 ^ n871 ;
  assign n869 = n93 ^ n79 ;
  assign n870 = n204 & ~n869 ;
  assign n875 = n874 ^ n870 ;
  assign n884 = n883 ^ n875 ;
  assign n885 = ~n868 & ~n884 ;
  assign n886 = n856 & n885 ;
  assign n887 = ~n837 & n886 ;
  assign n889 = n823 & n887 ;
  assign n888 = n887 ^ n823 ;
  assign n890 = n889 ^ n888 ;
  assign n892 = n689 & ~n890 ;
  assign n891 = n890 ^ n689 ;
  assign n893 = n892 ^ n891 ;
  assign n894 = n893 ^ n778 ;
  assign n895 = n781 & n894 ;
  assign n896 = n895 ^ n780 ;
  assign n941 = n896 ^ n694 ;
  assign n942 = ~n614 & n941 ;
  assign n897 = n689 ^ n618 ;
  assign n900 = n708 ^ n689 ;
  assign n903 = n897 & ~n900 ;
  assign n904 = n903 ^ n747 ;
  assign n905 = ~n746 & n904 ;
  assign n906 = n905 ^ n747 ;
  assign n940 = n939 ^ n906 ;
  assign n943 = n942 ^ n940 ;
  assign n912 = n710 ^ n617 ;
  assign n913 = n696 & ~n912 ;
  assign n910 = n694 & ~n1252 ;
  assign n907 = n906 ^ n614 ;
  assign n911 = n910 ^ n907 ;
  assign n914 = n913 ^ n911 ;
  assign n920 = n696 ^ n562 ;
  assign n923 = n748 & n920 ;
  assign n917 = n708 ^ n618 ;
  assign n924 = n923 ^ n917 ;
  assign n925 = ~n746 & n924 ;
  assign n926 = n925 ^ n917 ;
  assign n915 = ~n614 & ~n778 ;
  assign n916 = n915 ^ n614 ;
  assign n927 = n926 ^ n916 ;
  assign n928 = n707 ^ n689 ;
  assign n929 = n823 ^ n689 ;
  assign n930 = n928 & n929 ;
  assign n931 = n930 ^ n689 ;
  assign n932 = ~n888 & ~n931 ;
  assign n933 = n932 ^ n689 ;
  assign n934 = n933 ^ n916 ;
  assign n935 = n927 & n934 ;
  assign n936 = n935 ^ n926 ;
  assign n937 = n936 ^ n906 ;
  assign n938 = ~n914 & n937 ;
  assign n944 = n943 ^ n938 ;
  assign n950 = ~n939 & ~n944 ;
  assign n945 = n944 ^ n896 ;
  assign n946 = n939 ^ n614 ;
  assign n947 = n946 ^ n944 ;
  assign n948 = n947 ^ n694 ;
  assign n949 = ~n945 & ~n948 ;
  assign n951 = n950 ^ n949 ;
  assign n954 = ~n614 & n951 ;
  assign n955 = n954 ^ n950 ;
  assign n956 = n955 ^ n944 ;
  assign n755 = n754 ^ n741 ;
  assign n719 = n718 ^ n717 ;
  assign n720 = n614 & n718 ;
  assign n742 = ~n720 & n741 ;
  assign n743 = ~n694 & n742 ;
  assign n744 = n719 & n743 ;
  assign n745 = n744 ^ n742 ;
  assign n756 = n755 ^ n745 ;
  assign n765 = ~n752 & ~n764 ;
  assign n772 = ~n717 & ~n720 ;
  assign n773 = n765 & n772 ;
  assign n774 = n773 ^ n765 ;
  assign n775 = n774 ^ n764 ;
  assign n776 = ~n756 & ~n775 ;
  assign n957 = n956 ^ n776 ;
  assign n998 = x22 ^ x7 ;
  assign n996 = ~x6 & ~x22 ;
  assign n997 = n34 & n996 ;
  assign n999 = n998 ^ n997 ;
  assign n994 = ~x22 & ~n35 ;
  assign n995 = n994 ^ x8 ;
  assign n1000 = n999 ^ n995 ;
  assign n1026 = n409 ^ n392 ;
  assign n1027 = n1026 ^ n283 ;
  assign n1025 = n305 ^ n243 ;
  assign n1028 = n1027 ^ n1025 ;
  assign n1029 = n1028 ^ n195 ;
  assign n1023 = n553 ^ n447 ;
  assign n1024 = n1023 ^ n175 ;
  assign n1030 = n1029 ^ n1024 ;
  assign n1044 = ~n80 & n123 ;
  assign n1045 = n1044 ^ n841 ;
  assign n1041 = ~n126 & n594 ;
  assign n1042 = n1041 ^ n678 ;
  assign n1043 = n1042 ^ n118 ;
  assign n1046 = n1045 ^ n1043 ;
  assign n1040 = ~n125 & n563 ;
  assign n1047 = n1046 ^ n1040 ;
  assign n1037 = n479 ^ n273 ;
  assign n1035 = n642 ^ n391 ;
  assign n1036 = n1035 ^ n489 ;
  assign n1038 = n1037 ^ n1036 ;
  assign n1033 = n1032 ^ n263 ;
  assign n1031 = n383 ^ n330 ;
  assign n1034 = n1033 ^ n1031 ;
  assign n1039 = n1038 ^ n1034 ;
  assign n1048 = n1047 ^ n1039 ;
  assign n1049 = ~n1030 & n1048 ;
  assign n1017 = n845 ^ n394 ;
  assign n1018 = n1017 ^ n525 ;
  assign n1019 = n1018 ^ n312 ;
  assign n1016 = n320 ^ n256 ;
  assign n1020 = n1019 ^ n1016 ;
  assign n1014 = n1013 ^ n654 ;
  assign n1015 = n1014 ^ n231 ;
  assign n1021 = n1020 ^ n1015 ;
  assign n1009 = n859 ^ n512 ;
  assign n1008 = n605 ^ n225 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1004 = n430 ^ n362 ;
  assign n1005 = n1004 ^ n668 ;
  assign n1006 = n1005 ^ n793 ;
  assign n1001 = n334 ^ n286 ;
  assign n1003 = n1002 ^ n1001 ;
  assign n1007 = n1006 ^ n1003 ;
  assign n1011 = n1010 ^ n1007 ;
  assign n1022 = n1021 ^ n1011 ;
  assign n1050 = n1049 ^ n1022 ;
  assign n1051 = n1019 ^ n680 ;
  assign n1058 = n291 ^ n163 ;
  assign n1057 = n478 ^ n331 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1056 = n392 ^ n279 ;
  assign n1060 = n1059 ^ n1056 ;
  assign n1053 = n288 ^ n245 ;
  assign n1052 = n242 ^ n167 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n1055 = n1054 ^ n1032 ;
  assign n1061 = n1060 ^ n1055 ;
  assign n1062 = ~n1051 & ~n1061 ;
  assign n327 = n123 ^ n80 ;
  assign n328 = n327 ^ n133 ;
  assign n329 = ~n261 & ~n328 ;
  assign n1063 = n1062 ^ n329 ;
  assign n370 = ~n107 & n365 ;
  assign n371 = n370 ^ n185 ;
  assign n372 = n140 & n371 ;
  assign n368 = n185 ^ n107 ;
  assign n373 = n372 ^ n368 ;
  assign n1064 = n1063 ^ n373 ;
  assign n1088 = n231 ^ n94 ;
  assign n1090 = n1089 ^ n1088 ;
  assign n1091 = n1090 ^ n623 ;
  assign n1086 = n607 ^ n585 ;
  assign n1085 = n449 ^ n236 ;
  assign n1087 = n1086 ^ n1085 ;
  assign n1092 = n1091 ^ n1087 ;
  assign n437 = n201 ^ n161 ;
  assign n438 = n437 ^ n267 ;
  assign n435 = n434 ^ n179 ;
  assign n436 = n435 ^ n248 ;
  assign n439 = n438 ^ n436 ;
  assign n432 = n317 ^ n114 ;
  assign n433 = ~n126 & n432 ;
  assign n440 = n439 ^ n433 ;
  assign n1093 = n1092 ^ n440 ;
  assign n1079 = n566 ^ n344 ;
  assign n1080 = n1079 ^ n82 ;
  assign n1082 = n566 ^ n274 ;
  assign n298 = n93 & n154 ;
  assign n1081 = n548 ^ n298 ;
  assign n1083 = n1082 ^ n1081 ;
  assign n1084 = ~n1080 & ~n1083 ;
  assign n1094 = n1093 ^ n1084 ;
  assign n1075 = n645 ^ n472 ;
  assign n1073 = n1044 ^ n186 ;
  assign n1074 = n1073 ^ n318 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1077 = n1076 ^ n1002 ;
  assign n1070 = n379 ^ n225 ;
  assign n1071 = n1070 ^ n345 ;
  assign n426 = n92 & n154 ;
  assign n428 = n427 ^ n426 ;
  assign n1069 = n428 ^ n348 ;
  assign n1072 = n1071 ^ n1069 ;
  assign n1078 = n1077 ^ n1072 ;
  assign n1095 = n1094 ^ n1078 ;
  assign n1065 = n296 ^ n117 ;
  assign n1066 = n185 ^ n173 ;
  assign n1067 = n1066 ^ n89 ;
  assign n1068 = ~n1065 & n1067 ;
  assign n1096 = n1095 ^ n1068 ;
  assign n1097 = ~n1064 & n1096 ;
  assign n1098 = ~n887 & ~n1097 ;
  assign n1099 = n1050 & n1098 ;
  assign n1100 = n1099 ^ n887 ;
  assign n1101 = n1100 ^ n999 ;
  assign n1102 = ~n1000 & ~n1101 ;
  assign n1103 = n1102 ^ n999 ;
  assign n1104 = ~n614 & ~n1103 ;
  assign n989 = ~n617 & n694 ;
  assign n986 = n780 ^ n710 ;
  assign n990 = n989 ^ n986 ;
  assign n991 = ~n912 & n990 ;
  assign n992 = n991 ^ n986 ;
  assign n993 = n713 & n992 ;
  assign n1105 = n1104 ^ n993 ;
  assign n967 = ~n689 & n889 ;
  assign n968 = n967 ^ n892 ;
  assign n969 = n900 & n968 ;
  assign n966 = n888 & n928 ;
  assign n970 = n969 ^ n966 ;
  assign n971 = n970 ^ n915 ;
  assign n963 = n617 & n781 ;
  assign n964 = n963 ^ n780 ;
  assign n965 = ~n710 & n964 ;
  assign n972 = n971 ^ n965 ;
  assign n976 = n694 ^ n562 ;
  assign n979 = n748 & n976 ;
  assign n973 = n696 ^ n618 ;
  assign n980 = n979 ^ n973 ;
  assign n981 = ~n746 & ~n980 ;
  assign n982 = n981 ^ n973 ;
  assign n983 = n982 ^ n970 ;
  assign n984 = ~n972 & ~n983 ;
  assign n985 = n984 ^ n982 ;
  assign n1106 = n1105 ^ n985 ;
  assign n958 = n933 ^ n927 ;
  assign n1107 = n1106 ^ n958 ;
  assign n1113 = ~n614 & ~n999 ;
  assign n1110 = n696 ^ n689 ;
  assign n1111 = n968 & ~n1110 ;
  assign n1109 = n888 & n900 ;
  assign n1112 = n1111 ^ n1109 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1115 = n1097 ^ n1050 ;
  assign n1119 = n1050 ^ n707 ;
  assign n1308 = n887 ^ n707 ;
  assign n1120 = ~n1119 & n1308 ;
  assign n1121 = n1120 ^ n707 ;
  assign n1122 = n1115 & ~n1121 ;
  assign n1116 = n1113 ^ n887 ;
  assign n1123 = n1122 ^ n1116 ;
  assign n1124 = ~n1114 & n1123 ;
  assign n1125 = n1124 ^ n1113 ;
  assign n1126 = n1125 ^ n1100 ;
  assign n1108 = ~n614 & ~n1000 ;
  assign n1127 = n1126 ^ n1108 ;
  assign n1241 = n780 ^ n562 ;
  assign n1244 = n748 & n1241 ;
  assign n1238 = n694 ^ n618 ;
  assign n1245 = n1244 ^ n1238 ;
  assign n1246 = ~n746 & ~n1245 ;
  assign n1247 = n1246 ^ n1238 ;
  assign n1128 = ~x22 & ~n34 ;
  assign n1129 = n1128 ^ x6 ;
  assign n1130 = ~n614 & n1129 ;
  assign n1144 = n149 ^ n124 ;
  assign n1145 = n185 ^ n133 ;
  assign n1150 = ~n404 & n1145 ;
  assign n1151 = n1150 ^ n173 ;
  assign n1152 = n1144 & n1151 ;
  assign n1153 = n1152 ^ n379 ;
  assign n1134 = n294 ^ n155 ;
  assign n1133 = n525 ^ n298 ;
  assign n1135 = n1134 ^ n1133 ;
  assign n1136 = n1135 ^ n245 ;
  assign n1131 = n207 ^ n126 ;
  assign n1132 = n89 & ~n1131 ;
  assign n1137 = n1136 ^ n1132 ;
  assign n1138 = n334 ^ n303 ;
  assign n1139 = n1138 ^ n237 ;
  assign n1140 = n1139 ^ n354 ;
  assign n1141 = n1140 ^ n677 ;
  assign n1142 = n1141 ^ n1090 ;
  assign n1143 = n1137 & n1142 ;
  assign n1154 = n1153 ^ n1143 ;
  assign n1157 = n123 ^ n114 ;
  assign n1158 = n1157 ^ n592 ;
  assign n1159 = ~n117 & n1158 ;
  assign n1155 = n337 ^ n186 ;
  assign n1156 = n1155 ^ n169 ;
  assign n1160 = n1159 ^ n1156 ;
  assign n1161 = ~n428 & ~n1160 ;
  assign n454 = n453 ^ n450 ;
  assign n458 = n457 ^ n454 ;
  assign n448 = n447 ^ n444 ;
  assign n459 = n458 ^ n448 ;
  assign n442 = n162 ^ n105 ;
  assign n443 = n54 & n442 ;
  assign n460 = n459 ^ n443 ;
  assign n1162 = n1161 ^ n460 ;
  assign n1171 = n323 ^ n256 ;
  assign n1172 = n1171 ^ n1033 ;
  assign n1168 = n286 ^ n119 ;
  assign n1169 = n1168 ^ n296 ;
  assign n1170 = n1169 ^ n249 ;
  assign n1173 = n1172 ^ n1170 ;
  assign n1165 = n1164 ^ n386 ;
  assign n1166 = n1165 ^ n643 ;
  assign n1167 = n1166 ^ n1010 ;
  assign n1174 = n1173 ^ n1167 ;
  assign n1175 = n1162 & ~n1174 ;
  assign n1176 = n1154 & n1175 ;
  assign n1177 = n1097 & n1176 ;
  assign n1178 = ~n1130 & ~n1177 ;
  assign n1208 = n155 ^ n81 ;
  assign n1209 = n1208 ^ n350 ;
  assign n1210 = n1209 ^ n252 ;
  assign n1211 = n1210 ^ n1079 ;
  assign n1207 = ~n140 & n531 ;
  assign n1212 = n1211 ^ n1207 ;
  assign n1201 = n1066 ^ n539 ;
  assign n1202 = n117 & ~n1201 ;
  assign n1203 = n190 & ~n1066 ;
  assign n1204 = n55 & ~n1203 ;
  assign n1205 = ~n1202 & n1204 ;
  assign n1197 = n604 ^ n478 ;
  assign n1198 = n1197 ^ n231 ;
  assign n1196 = n426 ^ n348 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1200 = n1199 ^ n1031 ;
  assign n1206 = n1205 ^ n1200 ;
  assign n1213 = n1212 ^ n1206 ;
  assign n1215 = n575 ^ n291 ;
  assign n1216 = n1215 ^ n472 ;
  assign n1217 = n1216 ^ n305 ;
  assign n1218 = n1217 ^ n167 ;
  assign n415 = n414 ^ n358 ;
  assign n413 = n412 ^ n409 ;
  assign n416 = n415 ^ n413 ;
  assign n419 = n418 ^ n416 ;
  assign n1219 = n1218 ^ n419 ;
  assign n1214 = ~n79 & ~n1203 ;
  assign n1220 = n1219 ^ n1214 ;
  assign n1221 = n1213 & ~n1220 ;
  assign n1224 = n214 ^ n105 ;
  assign n1226 = n1225 ^ n1224 ;
  assign n1227 = ~n877 & ~n1226 ;
  assign n1228 = n1221 & n1227 ;
  assign n1186 = n791 ^ n170 ;
  assign n1185 = n1074 ^ n513 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1182 = n543 ^ n273 ;
  assign n322 = ~n140 & n154 ;
  assign n1181 = n481 ^ n322 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1179 = n437 ^ n224 ;
  assign n1180 = n1179 ^ n434 ;
  assign n1184 = n1183 ^ n1180 ;
  assign n1188 = n1187 ^ n1184 ;
  assign n1190 = n276 ^ n225 ;
  assign n1191 = n1190 ^ n256 ;
  assign n1189 = n427 ^ n238 ;
  assign n1192 = n1191 ^ n1189 ;
  assign n336 = n335 ^ n334 ;
  assign n338 = n337 ^ n336 ;
  assign n1193 = n1192 ^ n338 ;
  assign n1194 = n1188 & ~n1193 ;
  assign n1195 = n1194 ^ n1153 ;
  assign n1222 = n1221 ^ n1195 ;
  assign n1229 = n1228 ^ n1222 ;
  assign n1232 = ~n1176 & n1229 ;
  assign n1231 = n1229 ^ n1176 ;
  assign n1233 = n1232 ^ n1231 ;
  assign n1234 = ~n1097 & n1233 ;
  assign n1230 = ~n1097 & ~n1229 ;
  assign n1235 = n1234 ^ n1230 ;
  assign n1236 = n1178 & ~n1235 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1248 = n1247 ^ n1237 ;
  assign n1249 = n995 ^ n710 ;
  assign n1262 = n1249 ^ n1237 ;
  assign n1259 = n737 & ~n778 ;
  assign n1260 = n1259 ^ n995 ;
  assign n1261 = n1252 & ~n1260 ;
  assign n1263 = n1262 ^ n1261 ;
  assign n1264 = n1248 & n1263 ;
  assign n1265 = n1264 ^ n1247 ;
  assign n1266 = n1265 ^ n1125 ;
  assign n1267 = ~n1127 & n1266 ;
  assign n1268 = n1267 ^ n1125 ;
  assign n1269 = n1268 ^ n1106 ;
  assign n1270 = n1107 & n1269 ;
  assign n1271 = n1270 ^ n1106 ;
  assign n1272 = n936 ^ n914 ;
  assign n1273 = n1104 ^ n985 ;
  assign n1274 = n1105 & ~n1273 ;
  assign n1275 = n1274 ^ n1104 ;
  assign n1276 = n1275 ^ n1272 ;
  assign n1277 = ~n614 & n781 ;
  assign n1278 = n1277 ^ n893 ;
  assign n1279 = n1278 ^ n1275 ;
  assign n1280 = ~n1276 & n1279 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n1282 = ~n1272 & n1281 ;
  assign n1283 = n1271 & ~n1282 ;
  assign n1284 = n1280 ^ n1272 ;
  assign n1285 = ~n1283 & ~n1284 ;
  assign n1292 = n1282 ^ n1271 ;
  assign n1293 = n1292 ^ n1283 ;
  assign n1294 = n944 & ~n1293 ;
  assign n1289 = n1278 ^ n1276 ;
  assign n1290 = n1289 ^ n1271 ;
  assign n1286 = n1282 ^ n1281 ;
  assign n1287 = n1271 & n1286 ;
  assign n1288 = n1287 ^ n1285 ;
  assign n1291 = n1290 ^ n1288 ;
  assign n1295 = n1294 ^ n1291 ;
  assign n2221 = n1295 ^ n1285 ;
  assign n1297 = n1123 ^ n1112 ;
  assign n1296 = n1263 ^ n1247 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1307 = n887 ^ n708 ;
  assign n1311 = n1097 ^ n887 ;
  assign n1314 = n1307 & n1311 ;
  assign n1315 = n1314 ^ n1308 ;
  assign n1316 = n1115 & n1315 ;
  assign n1317 = n1316 ^ n1308 ;
  assign n1300 = n999 ^ n617 ;
  assign n1301 = n1300 ^ n995 ;
  assign n1304 = ~n1252 & n1301 ;
  assign n1305 = n1304 ^ n995 ;
  assign n1306 = n713 & n1305 ;
  assign n1318 = n1317 ^ n1306 ;
  assign n1322 = n778 ^ n562 ;
  assign n1325 = n748 & n1322 ;
  assign n1319 = n780 ^ n618 ;
  assign n1326 = n1325 ^ n1319 ;
  assign n1327 = ~n746 & ~n1326 ;
  assign n1328 = n1327 ^ n1319 ;
  assign n1329 = n1328 ^ n1317 ;
  assign n1330 = n1318 & ~n1329 ;
  assign n1331 = n1330 ^ n1317 ;
  assign n1332 = n1331 ^ n1296 ;
  assign n1333 = n1298 & ~n1332 ;
  assign n1334 = n1333 ^ n1297 ;
  assign n1335 = n982 ^ n972 ;
  assign n1337 = ~n1334 & n1335 ;
  assign n1336 = n1335 ^ n1334 ;
  assign n1338 = n1337 ^ n1336 ;
  assign n1339 = n1268 ^ n1107 ;
  assign n1340 = n1339 ^ n1337 ;
  assign n1435 = n1129 & ~n1252 ;
  assign n1434 = ~n912 & ~n999 ;
  assign n1436 = n1435 ^ n1434 ;
  assign n1437 = n1436 ^ n614 ;
  assign n1405 = ~x22 & ~n32 ;
  assign n1406 = n1405 ^ x4 ;
  assign n1407 = ~n614 & ~n1406 ;
  assign n1408 = n1407 ^ n614 ;
  assign n1409 = n1408 ^ n1176 ;
  assign n1346 = n1176 ^ n1097 ;
  assign n1417 = n1346 ^ n707 ;
  assign n1418 = n1417 ^ n1229 ;
  assign n1419 = n1418 ^ n709 ;
  assign n1420 = ~n1346 & ~n1419 ;
  assign n1421 = n1420 ^ n709 ;
  assign n1422 = n1231 & n1421 ;
  assign n1423 = n1422 ^ n1417 ;
  assign n1424 = n1423 ^ n1408 ;
  assign n1410 = n1097 ^ n708 ;
  assign n1411 = n1346 & n1410 ;
  assign n1412 = n1231 & n1411 ;
  assign n1413 = n1412 ^ n1176 ;
  assign n1427 = n1413 ^ n1408 ;
  assign n1428 = ~n1424 & n1427 ;
  assign n1414 = n1413 ^ n1229 ;
  assign n1430 = n1428 ^ n1414 ;
  assign n1431 = n1430 ^ n1229 ;
  assign n1432 = n1409 & ~n1431 ;
  assign n1433 = n1432 ^ n1176 ;
  assign n1438 = n1437 ^ n1433 ;
  assign n1448 = n778 ^ n689 ;
  assign n1449 = n968 & ~n1448 ;
  assign n1376 = n780 ^ n689 ;
  assign n1447 = n888 & ~n1376 ;
  assign n1450 = n1449 ^ n1447 ;
  assign n1392 = n887 ^ n696 ;
  assign n1451 = n1450 ^ n1392 ;
  assign n1439 = n887 ^ n694 ;
  assign n1444 = n1311 & ~n1439 ;
  assign n1445 = n1444 ^ n1392 ;
  assign n1446 = n1115 & ~n1445 ;
  assign n1452 = n1451 ^ n1446 ;
  assign n1552 = n999 ^ n618 ;
  assign n1458 = n748 & n1552 ;
  assign n1455 = n995 ^ n618 ;
  assign n1459 = n1458 ^ n1455 ;
  assign n1460 = ~n746 & ~n1459 ;
  assign n1461 = n1460 ^ n1455 ;
  assign n1462 = n1461 ^ n1450 ;
  assign n1463 = ~n1452 & ~n1462 ;
  assign n1453 = n1450 ^ n1437 ;
  assign n1464 = n1463 ^ n1453 ;
  assign n1465 = n1438 & ~n1464 ;
  assign n1466 = n1465 ^ n1437 ;
  assign n1403 = n1328 ^ n1318 ;
  assign n1382 = n995 ^ n562 ;
  assign n1385 = n748 & n1382 ;
  assign n1379 = n778 ^ n618 ;
  assign n1386 = n1385 ^ n1379 ;
  assign n1387 = ~n746 & ~n1386 ;
  assign n1388 = n1387 ^ n1379 ;
  assign n1377 = n968 & ~n1376 ;
  assign n1342 = n694 ^ n689 ;
  assign n1375 = n888 & ~n1342 ;
  assign n1378 = n1377 ^ n1375 ;
  assign n1389 = n1388 ^ n1378 ;
  assign n1397 = n1311 & ~n1392 ;
  assign n1398 = n1397 ^ n1307 ;
  assign n1399 = n1115 & n1398 ;
  assign n1390 = n1378 ^ n1307 ;
  assign n1400 = n1399 ^ n1390 ;
  assign n1401 = ~n1389 & ~n1400 ;
  assign n1402 = n1401 ^ n1388 ;
  assign n1404 = n1403 ^ n1402 ;
  assign n2179 = n1466 ^ n1404 ;
  assign n1522 = n605 ^ n392 ;
  assign n1523 = n1522 ^ n678 ;
  assign n1524 = n1523 ^ n656 ;
  assign n324 = n323 ^ n322 ;
  assign n325 = n324 ^ n321 ;
  assign n275 = n274 ^ n273 ;
  assign n277 = n276 ^ n275 ;
  assign n1521 = n325 ^ n277 ;
  assign n1525 = n1524 ^ n1521 ;
  assign n1518 = n1044 ^ n383 ;
  assign n1519 = n1518 ^ n1208 ;
  assign n1520 = n1519 ^ n479 ;
  assign n1526 = n1525 ^ n1520 ;
  assign n1527 = n1526 ^ n348 ;
  assign n1493 = n877 ^ n117 ;
  assign n1494 = n154 & n1493 ;
  assign n1491 = n93 & n787 ;
  assign n1489 = n243 ^ n118 ;
  assign n1490 = n1489 ^ n291 ;
  assign n1492 = n1491 ^ n1490 ;
  assign n1495 = n1494 ^ n1492 ;
  assign n1485 = n344 ^ n249 ;
  assign n1486 = n1485 ^ n201 ;
  assign n1484 = n1483 ^ n1189 ;
  assign n1487 = n1486 ^ n1484 ;
  assign n1488 = n1487 ^ n632 ;
  assign n1496 = n1495 ^ n1488 ;
  assign n1513 = n645 ^ n417 ;
  assign n1514 = n1513 ^ n398 ;
  assign n1515 = n1514 ^ n611 ;
  assign n1503 = ~n77 & ~n91 ;
  assign n1497 = n144 ^ n105 ;
  assign n1498 = n1497 ^ n185 ;
  assign n1504 = n1503 ^ n1498 ;
  assign n1510 = ~n42 & ~n1497 ;
  assign n1505 = n1498 ^ n42 ;
  assign n1501 = n1498 ^ n91 ;
  assign n1506 = n1505 ^ n1501 ;
  assign n1511 = n1510 ^ n1506 ;
  assign n1512 = n1504 & ~n1511 ;
  assign n1516 = n1515 ^ n1512 ;
  assign n1517 = n1496 & ~n1516 ;
  assign n1528 = n1527 ^ n1517 ;
  assign n1593 = ~n708 & ~n1176 ;
  assign n1594 = n1593 ^ n707 ;
  assign n1595 = ~n1528 & ~n1594 ;
  assign n1591 = n1176 ^ n707 ;
  assign n1596 = n1595 ^ n1591 ;
  assign n1597 = ~n614 & n1596 ;
  assign n1583 = n1407 ^ n710 ;
  assign n1356 = ~x22 & ~n33 ;
  assign n1357 = n1356 ^ x5 ;
  assign n1359 = n614 & ~n1357 ;
  assign n1584 = n1406 ^ n1359 ;
  assign n1587 = ~n617 & ~n1584 ;
  assign n1588 = n1587 ^ n1406 ;
  assign n1589 = ~n1583 & n1588 ;
  assign n1598 = n1597 ^ n1589 ;
  assign n1606 = n1357 ^ n562 ;
  assign n1609 = n748 & n1606 ;
  assign n1603 = n1129 ^ n618 ;
  assign n1610 = n1609 ^ n1603 ;
  assign n1611 = ~n746 & ~n1610 ;
  assign n1612 = n1611 ^ n1603 ;
  assign n1600 = n999 ^ n689 ;
  assign n1601 = n968 & n1600 ;
  assign n1563 = n995 ^ n689 ;
  assign n1599 = n888 & ~n1563 ;
  assign n1602 = n1601 ^ n1599 ;
  assign n1613 = n1612 ^ n1602 ;
  assign n1569 = n887 ^ n780 ;
  assign n1622 = n1602 ^ n1569 ;
  assign n1614 = n887 ^ n778 ;
  assign n1619 = n1311 & ~n1614 ;
  assign n1620 = n1619 ^ n1569 ;
  assign n1621 = n1115 & ~n1620 ;
  assign n1623 = n1622 ^ n1621 ;
  assign n1624 = ~n1613 & n1623 ;
  assign n1625 = n1624 ^ n1612 ;
  assign n1626 = n1625 ^ n1597 ;
  assign n1627 = n1598 & ~n1626 ;
  assign n1628 = n1627 ^ n1597 ;
  assign n1581 = n1461 ^ n1452 ;
  assign n1582 = n1581 ^ n1424 ;
  assign n1629 = n1628 ^ n1582 ;
  assign n1564 = n968 & ~n1563 ;
  assign n1562 = n888 & ~n1448 ;
  assign n1565 = n1564 ^ n1562 ;
  assign n1555 = n1129 ^ n689 ;
  assign n1558 = n897 & n1555 ;
  assign n1559 = n1558 ^ n1552 ;
  assign n1560 = ~n746 & n1559 ;
  assign n1561 = n1560 ^ n1552 ;
  assign n1566 = n1565 ^ n1561 ;
  assign n1574 = n1311 & ~n1569 ;
  assign n1575 = n1574 ^ n1439 ;
  assign n1576 = n1115 & ~n1575 ;
  assign n1567 = n1565 ^ n1439 ;
  assign n1577 = n1576 ^ n1567 ;
  assign n1578 = n1566 & ~n1577 ;
  assign n1579 = n1578 ^ n1565 ;
  assign n1529 = ~n707 & ~n1176 ;
  assign n1530 = ~n1528 & n1529 ;
  assign n1531 = n1530 ^ n1176 ;
  assign n1473 = x22 ^ x2 ;
  assign n1474 = ~x1 & ~x22 ;
  assign n1475 = n1473 & n1474 ;
  assign n1476 = n1475 ^ n1473 ;
  assign n1478 = n30 & n1476 ;
  assign n1479 = n1478 ^ n31 ;
  assign n1477 = n1476 ^ x22 ;
  assign n1480 = n1479 ^ n1477 ;
  assign n1481 = n1480 ^ x3 ;
  assign n1482 = ~n614 & ~n1481 ;
  assign n1532 = n1531 ^ n1482 ;
  assign n1539 = n1229 ^ n1097 ;
  assign n1542 = n1097 ^ n696 ;
  assign n1545 = ~n1539 & ~n1542 ;
  assign n1546 = n1545 ^ n1410 ;
  assign n1547 = n1231 & n1546 ;
  assign n1548 = n1547 ^ n1410 ;
  assign n1549 = n1548 ^ n1531 ;
  assign n1550 = ~n1532 & ~n1549 ;
  assign n1534 = ~n1252 & n1357 ;
  assign n1533 = ~n912 & n1129 ;
  assign n1535 = n1534 ^ n1533 ;
  assign n1536 = n1535 ^ n614 ;
  assign n1537 = n1536 ^ n1531 ;
  assign n1551 = n1550 ^ n1537 ;
  assign n1580 = n1579 ^ n1551 ;
  assign n1630 = n1629 ^ n1580 ;
  assign n1657 = n1577 ^ n1561 ;
  assign n1640 = n1596 ^ n614 ;
  assign n1632 = n1481 ^ n1406 ;
  assign n1637 = ~n1252 & n1632 ;
  assign n1585 = n1406 ^ n617 ;
  assign n1638 = n1637 ^ n1585 ;
  assign n1639 = n713 & n1638 ;
  assign n1641 = n1640 ^ n1639 ;
  assign n1645 = n1097 ^ n694 ;
  assign n1650 = ~n1539 & ~n1645 ;
  assign n1651 = n1650 ^ n1542 ;
  assign n1652 = n1231 & ~n1651 ;
  assign n1653 = n1652 ^ n1542 ;
  assign n1654 = n1653 ^ n1640 ;
  assign n1655 = ~n1641 & n1654 ;
  assign n1642 = n1548 ^ n1532 ;
  assign n1643 = n1642 ^ n1640 ;
  assign n1656 = n1655 ^ n1643 ;
  assign n1658 = n1657 ^ n1656 ;
  assign n1631 = n1625 ^ n1598 ;
  assign n1659 = n1658 ^ n1631 ;
  assign n1692 = n1623 ^ n1612 ;
  assign n1672 = n1406 ^ n562 ;
  assign n1675 = n748 & n1672 ;
  assign n1669 = n1357 ^ n618 ;
  assign n1676 = n1675 ^ n1669 ;
  assign n1677 = ~n746 & ~n1676 ;
  assign n1678 = n1677 ^ n1669 ;
  assign n1660 = n1097 ^ n780 ;
  assign n1665 = ~n1539 & ~n1660 ;
  assign n1666 = n1665 ^ n1645 ;
  assign n1667 = n1231 & ~n1666 ;
  assign n1668 = n1667 ^ n1645 ;
  assign n1679 = n1678 ^ n1668 ;
  assign n1686 = n696 & ~n1176 ;
  assign n1687 = n1686 ^ n708 ;
  assign n1688 = ~n1528 & ~n1687 ;
  assign n1682 = n1176 ^ n708 ;
  assign n1683 = n1682 ^ n1668 ;
  assign n1689 = n1688 ^ n1683 ;
  assign n1690 = n1679 & n1689 ;
  assign n1691 = n1690 ^ n1678 ;
  assign n1693 = n1692 ^ n1691 ;
  assign n1695 = n968 & ~n1555 ;
  assign n1694 = n888 & n1600 ;
  assign n1696 = n1695 ^ n1694 ;
  assign n1720 = n1696 ^ n1692 ;
  assign n1699 = n995 ^ n887 ;
  assign n1704 = n1311 & ~n1699 ;
  assign n1705 = n1704 ^ n1614 ;
  assign n1706 = n1115 & ~n1705 ;
  assign n1697 = n1696 ^ n1614 ;
  assign n1707 = n1706 ^ n1697 ;
  assign n1711 = n694 & ~n1176 ;
  assign n1712 = n1711 ^ n696 ;
  assign n1713 = ~n1528 & n1712 ;
  assign n1709 = n1176 ^ n696 ;
  assign n1714 = n1713 ^ n1709 ;
  assign n1715 = n746 & ~n1481 ;
  assign n1716 = ~n692 & ~n1715 ;
  assign n1717 = ~n1714 & n1716 ;
  assign n1718 = n1717 ^ n1696 ;
  assign n1719 = ~n1707 & n1718 ;
  assign n1721 = n1720 ^ n1719 ;
  assign n1722 = ~n1693 & n1721 ;
  assign n1723 = n1722 ^ n1692 ;
  assign n1724 = n1723 ^ n1631 ;
  assign n1725 = n1659 & ~n1724 ;
  assign n1726 = n1725 ^ n1631 ;
  assign n1727 = n1726 ^ n1629 ;
  assign n1728 = ~n1630 & n1727 ;
  assign n1744 = n1728 ^ n1630 ;
  assign n1745 = n1744 ^ n1726 ;
  assign n1738 = n1579 ^ n1536 ;
  assign n1739 = n1551 & ~n1738 ;
  assign n1740 = n1739 ^ n1536 ;
  assign n1735 = n1400 ^ n1388 ;
  assign n1358 = n1357 ^ n614 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1736 = n1735 ^ n1360 ;
  assign n1348 = n1235 ^ n1177 ;
  assign n1347 = n1346 ^ n1232 ;
  assign n1349 = n1348 ^ n1347 ;
  assign n1350 = n1349 ^ n1233 ;
  assign n1351 = ~n707 & ~n1350 ;
  assign n1734 = ~n1348 & ~n1351 ;
  assign n1737 = n1736 ^ n1734 ;
  assign n1741 = n1740 ^ n1737 ;
  assign n1733 = n1464 ^ n1433 ;
  assign n1742 = n1741 ^ n1733 ;
  assign n1729 = n1628 ^ n1424 ;
  assign n1730 = n1628 ^ n1581 ;
  assign n1731 = n1729 & ~n1730 ;
  assign n1732 = n1731 ^ n1424 ;
  assign n1743 = n1742 ^ n1732 ;
  assign n1746 = n1745 ^ n1743 ;
  assign n1747 = n1657 ^ n1642 ;
  assign n1748 = n1656 & n1747 ;
  assign n1749 = n1748 ^ n1642 ;
  assign n1753 = n1717 ^ n1707 ;
  assign n1752 = ~n912 & ~n1481 ;
  assign n1754 = n1753 ^ n1752 ;
  assign n1765 = n1357 ^ n689 ;
  assign n1766 = n968 & ~n1765 ;
  assign n1764 = n888 & ~n1555 ;
  assign n1767 = n1766 ^ n1764 ;
  assign n1755 = n999 ^ n887 ;
  assign n1760 = n1311 & n1755 ;
  assign n1761 = n1760 ^ n1699 ;
  assign n1762 = n1115 & ~n1761 ;
  assign n1763 = n1762 ^ n1699 ;
  assign n1768 = n1767 ^ n1763 ;
  assign n1771 = n1097 ^ n778 ;
  assign n1776 = ~n1539 & ~n1771 ;
  assign n1777 = n1776 ^ n1660 ;
  assign n1778 = n1231 & ~n1777 ;
  assign n1769 = n1763 ^ n1660 ;
  assign n1779 = n1778 ^ n1769 ;
  assign n1780 = ~n1768 & ~n1779 ;
  assign n1781 = n1780 ^ n1767 ;
  assign n1782 = n1781 ^ n1752 ;
  assign n1783 = ~n1754 & ~n1782 ;
  assign n1784 = n1783 ^ n1753 ;
  assign n1751 = n1721 ^ n1691 ;
  assign n2154 = n1784 ^ n1751 ;
  assign n1785 = ~n1751 & ~n1784 ;
  assign n2155 = n2154 ^ n1785 ;
  assign n1788 = n1781 ^ n1754 ;
  assign n1787 = n1689 ^ n1678 ;
  assign n1789 = n1788 ^ n1787 ;
  assign n1790 = n1406 ^ n618 ;
  assign n1791 = n1790 ^ n1632 ;
  assign n1793 = n748 & n1791 ;
  assign n1794 = n1793 ^ n1790 ;
  assign n1795 = ~n746 & ~n1794 ;
  assign n1796 = n1795 ^ n1790 ;
  assign n1827 = n1796 ^ n1787 ;
  assign n1797 = n1716 ^ n1714 ;
  assign n1798 = n1797 ^ n1796 ;
  assign n1804 = n1129 ^ n887 ;
  assign n1809 = n1311 & ~n1804 ;
  assign n1810 = n1809 ^ n1755 ;
  assign n1811 = n1115 & n1810 ;
  assign n1812 = n1811 ^ n1755 ;
  assign n1800 = n1349 ^ n1234 ;
  assign n1801 = n1097 ^ n995 ;
  assign n1802 = ~n1800 & ~n1801 ;
  assign n1799 = ~n1231 & ~n1771 ;
  assign n1803 = n1802 ^ n1799 ;
  assign n1813 = n1812 ^ n1803 ;
  assign n1816 = n1176 ^ n694 ;
  assign n1821 = n1816 ^ n1803 ;
  assign n1818 = n780 & ~n1176 ;
  assign n1819 = n1818 ^ n694 ;
  assign n1820 = ~n1528 & n1819 ;
  assign n1822 = n1821 ^ n1820 ;
  assign n1823 = n1813 & n1822 ;
  assign n1824 = n1823 ^ n1812 ;
  assign n1825 = n1824 ^ n1796 ;
  assign n1826 = n1798 & ~n1825 ;
  assign n1828 = n1827 ^ n1826 ;
  assign n1829 = ~n1789 & n1828 ;
  assign n1830 = n1829 ^ n1788 ;
  assign n1831 = n1653 ^ n1641 ;
  assign n2156 = ~n1830 & n1831 ;
  assign n1832 = n1831 ^ n1830 ;
  assign n2157 = n2156 ^ n1832 ;
  assign n1750 = n1723 ^ n1659 ;
  assign n2158 = n2157 ^ n1750 ;
  assign n1834 = n1828 ^ n1788 ;
  assign n1858 = n893 & ~n967 ;
  assign n1859 = n1481 & n1858 ;
  assign n1860 = n1859 ^ n967 ;
  assign n1863 = n778 & ~n1176 ;
  assign n1864 = n1863 ^ n780 ;
  assign n1865 = ~n1528 & n1864 ;
  assign n1861 = n1176 ^ n780 ;
  assign n1866 = n1865 ^ n1861 ;
  assign n1867 = n1860 & ~n1866 ;
  assign n1836 = n1406 ^ n689 ;
  assign n1869 = n968 & ~n1836 ;
  assign n1868 = n888 & ~n1765 ;
  assign n1870 = n1869 ^ n1868 ;
  assign n1873 = n1870 ^ n1715 ;
  assign n1871 = n1715 & n1870 ;
  assign n1875 = n1873 ^ n1871 ;
  assign n1876 = ~n1867 & ~n1875 ;
  assign n1872 = n1867 & n1871 ;
  assign n1874 = n1873 ^ n1872 ;
  assign n1877 = n1876 ^ n1874 ;
  assign n1878 = n1877 ^ n1867 ;
  assign n1879 = n1822 ^ n1812 ;
  assign n1887 = n1879 ^ n1872 ;
  assign n1841 = n1097 ^ n999 ;
  assign n1842 = ~n1800 & n1841 ;
  assign n1840 = ~n1231 & ~n1801 ;
  assign n1843 = n1842 ^ n1840 ;
  assign n1837 = n888 & ~n1836 ;
  assign n1835 = n968 & n1481 ;
  assign n1838 = n1837 ^ n1835 ;
  assign n1839 = n1838 ^ n892 ;
  assign n1844 = n1843 ^ n1839 ;
  assign n1847 = n1357 ^ n887 ;
  assign n1852 = n1311 & ~n1847 ;
  assign n1853 = n1852 ^ n1804 ;
  assign n1854 = n1115 & ~n1853 ;
  assign n1845 = n1843 ^ n1804 ;
  assign n1855 = n1854 ^ n1845 ;
  assign n1856 = n1844 & ~n1855 ;
  assign n1857 = n1856 ^ n1843 ;
  assign n1888 = n1872 ^ n1857 ;
  assign n1889 = ~n1887 & n1888 ;
  assign n1890 = n1878 & n1889 ;
  assign n1892 = n1890 ^ n1889 ;
  assign n1893 = n1892 ^ n1872 ;
  assign n1880 = n1879 ^ n1876 ;
  assign n1881 = n1876 ^ n1857 ;
  assign n1882 = n1880 & ~n1881 ;
  assign n1883 = ~n1878 & n1882 ;
  assign n1885 = n1883 ^ n1882 ;
  assign n1886 = n1885 ^ n1876 ;
  assign n1894 = n1893 ^ n1886 ;
  assign n1895 = n1834 & n1894 ;
  assign n1896 = n1895 ^ n1893 ;
  assign n1899 = n1779 ^ n1767 ;
  assign n1904 = n1855 ^ n1839 ;
  assign n1903 = n1866 ^ n1860 ;
  assign n2113 = n1904 ^ n1903 ;
  assign n1905 = ~n1903 & ~n1904 ;
  assign n2114 = n2113 ^ n1905 ;
  assign n1913 = n1406 ^ n887 ;
  assign n1932 = n1913 ^ n1481 ;
  assign n1933 = n1932 ^ n1050 ;
  assign n1934 = n1933 ^ n1913 ;
  assign n1935 = n1913 ^ n1632 ;
  assign n1936 = n1934 & n1935 ;
  assign n1937 = n1936 ^ n1913 ;
  assign n1938 = n1115 & ~n1937 ;
  assign n1939 = n1938 ^ n1913 ;
  assign n1930 = ~n1115 & ~n1481 ;
  assign n1931 = ~n1100 & ~n1930 ;
  assign n1941 = n1939 ^ n1931 ;
  assign n1940 = ~n1931 & n1939 ;
  assign n1942 = n1941 ^ n1940 ;
  assign n1960 = n888 & ~n1481 ;
  assign n1944 = n1357 ^ n1097 ;
  assign n1945 = ~n1800 & ~n1944 ;
  assign n1908 = n1129 ^ n1097 ;
  assign n1943 = ~n1231 & ~n1908 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1956 = n1946 ^ n1940 ;
  assign n1968 = n1176 ^ n999 ;
  assign n1951 = n1176 & n1968 ;
  assign n1952 = n1951 ^ n1000 ;
  assign n1953 = ~n1528 & ~n1952 ;
  assign n1949 = n1176 ^ n995 ;
  assign n1954 = n1953 ^ n1949 ;
  assign n1957 = n1954 ^ n1946 ;
  assign n1958 = ~n1956 & n1957 ;
  assign n1959 = n1958 ^ n1940 ;
  assign n1961 = n1960 ^ n1959 ;
  assign n1955 = n1946 & ~n1954 ;
  assign n1962 = n1961 ^ n1955 ;
  assign n1963 = ~n1942 & n1962 ;
  assign n1964 = n1963 ^ n1955 ;
  assign n2099 = ~n1959 & ~n1960 ;
  assign n2100 = ~n1964 & n2099 ;
  assign n2101 = n2100 ^ n1959 ;
  assign n1918 = n1311 & ~n1913 ;
  assign n1919 = n1918 ^ n1847 ;
  assign n1920 = n1115 & ~n1919 ;
  assign n1909 = ~n1800 & ~n1908 ;
  assign n1907 = ~n1231 & n1841 ;
  assign n1910 = n1909 ^ n1907 ;
  assign n1911 = n1910 ^ n1847 ;
  assign n1921 = n1920 ^ n1911 ;
  assign n1925 = n995 & ~n1176 ;
  assign n1926 = n1925 ^ n778 ;
  assign n1927 = ~n1528 & n1926 ;
  assign n1923 = n1176 ^ n778 ;
  assign n1928 = n1927 ^ n1923 ;
  assign n2104 = n1928 ^ n1910 ;
  assign n2105 = n1921 & ~n2104 ;
  assign n2106 = n2105 ^ n1928 ;
  assign n2116 = ~n2101 & ~n2106 ;
  assign n2115 = n2106 ^ n2101 ;
  assign n2117 = n2116 ^ n2115 ;
  assign n1900 = n1879 ^ n1867 ;
  assign n1901 = n1900 ^ n1873 ;
  assign n1902 = n1901 ^ n1857 ;
  assign n2118 = n2117 ^ n1902 ;
  assign n1929 = n1928 ^ n1921 ;
  assign n1965 = n1964 ^ n1929 ;
  assign n1975 = n1406 ^ n1097 ;
  assign n1976 = ~n1800 & ~n1975 ;
  assign n1974 = ~n1231 & ~n1944 ;
  assign n1977 = n1976 ^ n1974 ;
  assign n1970 = n1129 & ~n1176 ;
  assign n1971 = n1970 ^ n999 ;
  assign n1972 = ~n1528 & ~n1971 ;
  assign n1973 = n1972 ^ n1968 ;
  assign n1978 = n1977 ^ n1973 ;
  assign n1993 = n1481 ^ n1176 ;
  assign n1994 = ~n1231 & n1993 ;
  assign n1995 = n1994 ^ n1176 ;
  assign n1996 = ~n1097 & n1995 ;
  assign n2013 = n1357 ^ n1176 ;
  assign n2005 = ~n1176 & ~n2013 ;
  assign n2000 = n1176 ^ n1129 ;
  assign n2006 = n2005 ^ n2000 ;
  assign n2007 = ~n1528 & ~n2006 ;
  assign n2008 = n2007 ^ n2000 ;
  assign n2079 = n1996 & ~n2008 ;
  assign n2080 = n2079 ^ n1973 ;
  assign n2081 = n1978 & n2080 ;
  assign n1980 = n1357 & n1528 ;
  assign n1979 = n1229 & ~n1481 ;
  assign n1981 = n1980 ^ n1979 ;
  assign n1982 = n1975 ^ n1632 ;
  assign n1984 = n1406 ^ n1229 ;
  assign n1985 = n1984 ^ n1632 ;
  assign n1986 = n1982 & ~n1985 ;
  assign n1987 = n1986 ^ n1632 ;
  assign n1988 = n1231 & ~n1987 ;
  assign n1989 = n1988 ^ n1975 ;
  assign n1991 = n1978 & ~n1989 ;
  assign n2010 = ~n1930 & ~n1991 ;
  assign n1998 = ~n1930 & ~n1996 ;
  assign n1999 = n1998 ^ n1978 ;
  assign n2009 = ~n1999 & n2008 ;
  assign n2011 = n2010 ^ n2009 ;
  assign n1990 = n1989 ^ n1978 ;
  assign n1992 = n1991 ^ n1990 ;
  assign n1997 = n1992 & ~n1996 ;
  assign n2012 = n2011 ^ n1997 ;
  assign n2016 = n1406 ^ n1176 ;
  assign n2028 = n2016 ^ n1528 ;
  assign n2041 = n1528 ^ n1176 ;
  assign n2029 = n2041 ^ n2016 ;
  assign n2030 = n2028 & n2029 ;
  assign n2020 = n2041 ^ n1632 ;
  assign n2022 = n2013 ^ n1632 ;
  assign n2024 = n2022 ^ n1176 ;
  assign n2025 = ~n2020 & n2024 ;
  assign n2031 = n2030 ^ n2025 ;
  assign n2032 = n2031 ^ n1176 ;
  assign n2033 = n2030 ^ n2013 ;
  assign n2034 = n2033 ^ n1176 ;
  assign n2035 = n2032 & ~n2034 ;
  assign n2036 = n1528 & n2035 ;
  assign n2037 = n2036 ^ n2030 ;
  assign n2014 = n1528 ^ n1357 ;
  assign n2050 = n2037 ^ n2014 ;
  assign n2051 = n2050 ^ n2013 ;
  assign n2052 = n2012 & ~n2051 ;
  assign n2053 = ~n1981 & n2052 ;
  assign n2054 = n2053 ^ n2012 ;
  assign n2055 = n1957 ^ n1941 ;
  assign n2056 = n2055 ^ n1998 ;
  assign n2057 = ~n1978 & ~n2056 ;
  assign n2058 = n2057 ^ n2055 ;
  assign n2059 = n2008 & n2058 ;
  assign n2067 = ~n2010 & n2059 ;
  assign n2068 = ~n1992 & n2067 ;
  assign n2069 = n2068 ^ n1992 ;
  assign n2060 = n2059 ^ n2058 ;
  assign n2061 = n2060 ^ n1992 ;
  assign n2070 = n2069 ^ n2061 ;
  assign n2071 = ~n2054 & n2070 ;
  assign n2072 = n2071 ^ n2055 ;
  assign n2073 = n2072 ^ n1973 ;
  assign n2082 = n2081 ^ n2073 ;
  assign n2093 = n2082 ^ n1929 ;
  assign n2088 = ~n1973 & n2057 ;
  assign n2089 = n2088 ^ n2082 ;
  assign n2090 = n2071 & n2089 ;
  assign n2094 = n2093 ^ n2090 ;
  assign n2083 = n2082 ^ n2071 ;
  assign n2091 = ~n2072 & ~n2090 ;
  assign n2092 = ~n2083 & n2091 ;
  assign n2095 = n2094 ^ n2092 ;
  assign n2096 = ~n1965 & n2095 ;
  assign n2097 = n2096 ^ n1964 ;
  assign n2119 = n2118 ^ n2097 ;
  assign n2120 = n2114 & ~n2119 ;
  assign n1906 = n1905 ^ n1902 ;
  assign n2102 = n2101 ^ n1902 ;
  assign n2098 = n2097 ^ n1902 ;
  assign n2103 = n2102 ^ n2098 ;
  assign n2107 = n2106 ^ n1902 ;
  assign n2108 = n2107 ^ n2102 ;
  assign n2109 = n2103 & n2108 ;
  assign n2110 = n2109 ^ n2102 ;
  assign n2111 = ~n1906 & ~n2110 ;
  assign n2112 = n2111 ^ n1905 ;
  assign n2121 = n2116 ^ n1902 ;
  assign n2122 = ~n2112 & ~n2121 ;
  assign n2123 = n2120 & n2122 ;
  assign n2124 = n2123 ^ n2112 ;
  assign n2125 = ~n1899 & ~n2124 ;
  assign n1897 = n1824 ^ n1798 ;
  assign n1898 = n1897 ^ n1834 ;
  assign n2126 = n2125 ^ n1898 ;
  assign n2127 = n1896 & n2126 ;
  assign n2128 = n2127 ^ n1834 ;
  assign n2129 = n2124 ^ n1899 ;
  assign n2130 = n2129 ^ n2125 ;
  assign n2131 = n2130 ^ n1834 ;
  assign n2132 = n1893 ^ n1834 ;
  assign n2133 = n2132 ^ n1897 ;
  assign n2134 = n2133 ^ n2132 ;
  assign n2135 = n2132 ^ n1886 ;
  assign n2136 = n2135 ^ n2132 ;
  assign n2139 = ~n1893 & ~n2136 ;
  assign n2140 = n2134 & n2139 ;
  assign n2141 = n2140 ^ n2134 ;
  assign n2142 = n2141 ^ n2133 ;
  assign n2143 = ~n2131 & ~n2142 ;
  assign n2144 = n2143 ^ n2130 ;
  assign n2145 = ~n2125 & n2144 ;
  assign n2146 = n2128 & n2145 ;
  assign n2147 = n2146 ^ n2144 ;
  assign n2159 = n2158 ^ n2147 ;
  assign n2160 = n2155 & ~n2159 ;
  assign n1786 = n1785 ^ n1750 ;
  assign n2149 = n2147 ^ n1830 ;
  assign n2150 = n1832 & ~n2149 ;
  assign n1833 = n1832 ^ n1750 ;
  assign n2148 = n2147 ^ n1833 ;
  assign n2151 = n2150 ^ n2148 ;
  assign n2152 = n1786 & n2151 ;
  assign n2153 = n2152 ^ n1785 ;
  assign n2161 = n2156 ^ n1750 ;
  assign n2162 = ~n2153 & n2161 ;
  assign n2163 = n2160 & n2162 ;
  assign n2164 = n2163 ^ n2153 ;
  assign n2165 = n1749 & ~n2164 ;
  assign n2166 = n2165 ^ n1745 ;
  assign n2167 = n1746 & n2166 ;
  assign n2168 = n2167 ^ n1629 ;
  assign n2169 = ~n1728 & ~n2168 ;
  assign n2170 = n2169 ^ n1629 ;
  assign n2171 = n2164 ^ n1749 ;
  assign n2172 = n2171 ^ n1746 ;
  assign n2173 = n2172 ^ n2166 ;
  assign n2174 = n2173 ^ n2167 ;
  assign n2175 = n2167 ^ n1743 ;
  assign n2176 = n2174 & n2175 ;
  assign n2177 = ~n2170 & n2176 ;
  assign n2178 = n2177 ^ n2175 ;
  assign n2180 = n2179 ^ n2178 ;
  assign n1467 = n1466 ^ n1402 ;
  assign n1468 = ~n1404 & n1467 ;
  assign n1469 = n1468 ^ n1466 ;
  assign n1370 = n1331 ^ n1298 ;
  assign n1343 = n968 & ~n1342 ;
  assign n1341 = n888 & ~n1110 ;
  assign n1344 = n1343 ^ n1341 ;
  assign n1345 = n1344 ^ n1130 ;
  assign n1363 = ~n1348 & n1360 ;
  assign n1364 = n1363 ^ n1176 ;
  assign n1365 = ~n1351 & ~n1364 ;
  assign n1352 = n1177 ^ n1176 ;
  assign n1366 = n1365 ^ n1352 ;
  assign n1367 = n1366 ^ n1344 ;
  assign n1368 = ~n1345 & n1367 ;
  assign n1369 = n1368 ^ n1237 ;
  assign n1371 = n1370 ^ n1369 ;
  assign n2192 = n1469 ^ n1371 ;
  assign n2184 = n1366 ^ n1345 ;
  assign n2181 = n1740 ^ n1735 ;
  assign n2182 = n1737 & n2181 ;
  assign n2183 = n2182 ^ n1740 ;
  assign n2185 = n2184 ^ n2183 ;
  assign n2186 = n1741 ^ n1732 ;
  assign n2187 = n1742 & n2186 ;
  assign n2188 = n2187 ^ n1741 ;
  assign n2189 = n2188 ^ n2183 ;
  assign n2190 = n2185 & ~n2189 ;
  assign n2191 = n2190 ^ n2185 ;
  assign n2193 = n2192 ^ n2191 ;
  assign n2194 = n2193 ^ n2183 ;
  assign n2195 = n2193 ^ n2192 ;
  assign n2196 = ~n2194 & n2195 ;
  assign n2197 = n2196 ^ n2192 ;
  assign n2198 = n2197 ^ n2178 ;
  assign n2199 = n2180 & ~n2198 ;
  assign n2200 = n2190 ^ n2188 ;
  assign n2201 = n2200 ^ n2196 ;
  assign n2202 = n2201 ^ n2197 ;
  assign n2203 = n2199 & ~n2202 ;
  assign n2204 = n2203 ^ n2197 ;
  assign n2205 = n2204 ^ n1339 ;
  assign n1470 = n1469 ^ n1369 ;
  assign n1471 = n1371 & ~n1470 ;
  assign n1372 = n1265 ^ n1127 ;
  assign n1373 = n1372 ^ n1369 ;
  assign n1472 = n1471 ^ n1373 ;
  assign n2206 = n2205 ^ n1472 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2208 = n1372 ^ n1339 ;
  assign n2209 = n2208 ^ n2206 ;
  assign n2210 = ~n2207 & n2209 ;
  assign n2211 = n2210 ^ n2206 ;
  assign n2212 = n1340 & n2211 ;
  assign n2213 = n2212 ^ n1337 ;
  assign n2214 = ~n1338 & ~n2213 ;
  assign n2215 = ~n1372 & ~n1472 ;
  assign n2216 = n2215 ^ n2206 ;
  assign n2217 = n2215 ^ n1339 ;
  assign n2218 = ~n2216 & n2217 ;
  assign n2219 = n2214 & n2218 ;
  assign n2220 = n2219 ^ n2213 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2223 = n2222 ^ n1287 ;
  assign n2224 = n2223 ^ n2222 ;
  assign n2225 = n2222 ^ n944 ;
  assign n2226 = n2225 ^ n2222 ;
  assign n2227 = ~n2224 & n2226 ;
  assign n2228 = n2227 ^ n2222 ;
  assign n2229 = ~n1285 & ~n2228 ;
  assign n2230 = n2229 ^ n2222 ;
  assign n2231 = n2230 ^ n1295 ;
  assign n2232 = n2220 ^ n1295 ;
  assign n2233 = ~n2229 & ~n2232 ;
  assign n2234 = n2231 & n2233 ;
  assign n2235 = n2234 ^ n2230 ;
  assign n2236 = n2235 ^ n956 ;
  assign n2237 = n957 & n2236 ;
  assign n2238 = n2237 ^ n956 ;
  assign n2249 = n2248 ^ n2238 ;
  assign n2286 = n2285 ^ n2249 ;
  assign n2297 = n379 ^ n308 ;
  assign n2298 = n2297 ^ n252 ;
  assign n2294 = n280 ^ n267 ;
  assign n2295 = n2294 ^ n409 ;
  assign n2293 = n435 ^ n335 ;
  assign n2296 = n2295 ^ n2293 ;
  assign n2299 = n2298 ^ n2296 ;
  assign n2290 = n802 ^ n623 ;
  assign n2291 = n2290 ^ n826 ;
  assign n2292 = n2291 ^ n538 ;
  assign n2300 = n2299 ^ n2292 ;
  assign n2301 = n2300 ^ n1174 ;
  assign n2289 = n1047 ^ n245 ;
  assign n2302 = n2301 ^ n2289 ;
  assign n2288 = n105 & ~n877 ;
  assign n2303 = n2302 ^ n2288 ;
  assign n2287 = n2235 ^ n957 ;
  assign n2304 = n2303 ^ n2287 ;
  assign n281 = n280 ^ n277 ;
  assign n2378 = n281 ^ n115 ;
  assign n2377 = n428 ^ n245 ;
  assign n2379 = n2378 ^ n2377 ;
  assign n2380 = n2379 ^ n859 ;
  assign n2372 = n344 ^ n79 ;
  assign n2373 = n2372 ^ n390 ;
  assign n2366 = n1158 ^ n125 ;
  assign n2369 = ~n105 & n2366 ;
  assign n2370 = n2369 ^ n125 ;
  assign n2371 = ~n253 & ~n2370 ;
  assign n2374 = n2373 ^ n2371 ;
  assign n2357 = n337 ^ n124 ;
  assign n2358 = n185 ^ n74 ;
  assign n2363 = ~n42 & n2358 ;
  assign n2364 = n2363 ^ n661 ;
  assign n2365 = n2357 & n2364 ;
  assign n2375 = n2374 ^ n2365 ;
  assign n2376 = n2375 ^ n2280 ;
  assign n2381 = n2380 ^ n2376 ;
  assign n2354 = n449 ^ n399 ;
  assign n2355 = n2354 ^ n176 ;
  assign n2313 = n2257 ^ n201 ;
  assign n2314 = n2313 ^ n651 ;
  assign n2309 = n284 ^ n265 ;
  assign n2310 = n2309 ^ n2271 ;
  assign n2308 = n678 ^ n260 ;
  assign n2311 = n2310 ^ n2308 ;
  assign n2312 = n2311 ^ n422 ;
  assign n2315 = n2314 ^ n2312 ;
  assign n2306 = n252 ^ n238 ;
  assign n2305 = n1070 ^ n430 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2316 = n2315 ^ n2307 ;
  assign n2356 = n2355 ^ n2316 ;
  assign n2382 = n2381 ^ n2356 ;
  assign n2353 = n2220 ^ n1290 ;
  assign n2383 = n2382 ^ n2353 ;
  assign n2350 = n310 ^ n231 ;
  assign n2351 = n2350 ^ n117 ;
  assign n2352 = n589 & n2351 ;
  assign n2384 = n2383 ^ n2352 ;
  assign n2409 = n2204 ^ n1472 ;
  assign n2410 = n2204 ^ n1336 ;
  assign n2411 = ~n2409 & ~n2410 ;
  assign n2407 = n2215 ^ n1338 ;
  assign n2408 = n2407 ^ n1339 ;
  assign n2412 = n2411 ^ n2408 ;
  assign n332 = n331 ^ n330 ;
  assign n333 = n332 ^ n329 ;
  assign n339 = n338 ^ n333 ;
  assign n311 = n310 ^ n305 ;
  assign n313 = n312 ^ n311 ;
  assign n326 = n325 ^ n313 ;
  assign n340 = n339 ^ n326 ;
  assign n374 = n373 ^ n340 ;
  assign n2399 = n481 ^ n398 ;
  assign n2398 = n845 ^ n655 ;
  assign n2400 = n2399 ^ n2398 ;
  assign n2396 = n430 ^ n167 ;
  assign n2397 = n2396 ^ n81 ;
  assign n2401 = n2400 ^ n2397 ;
  assign n2393 = n678 ^ n291 ;
  assign n2394 = n2393 ^ n668 ;
  assign n2391 = n427 ^ n307 ;
  assign n2392 = n2391 ^ n411 ;
  assign n2395 = n2394 ^ n2392 ;
  assign n2402 = n2401 ^ n2395 ;
  assign n2389 = n512 ^ n385 ;
  assign n2388 = n55 & n145 ;
  assign n2390 = n2389 ^ n2388 ;
  assign n2403 = n2402 ^ n2390 ;
  assign n2404 = n2403 ^ n1094 ;
  assign n2385 = n317 ^ n79 ;
  assign n2386 = n2385 ^ n105 ;
  assign n2387 = ~n524 & ~n2386 ;
  assign n2405 = n2404 ^ n2387 ;
  assign n2406 = n374 & n2405 ;
  assign n2413 = n2412 ^ n2406 ;
  assign n2438 = n1472 ^ n1336 ;
  assign n2439 = n2438 ^ n2204 ;
  assign n2414 = n150 & ~n1011 ;
  assign n2431 = n1032 ^ n585 ;
  assign n2432 = n2431 ^ n852 ;
  assign n2429 = n646 ^ n481 ;
  assign n2428 = n642 ^ n543 ;
  assign n2430 = n2429 ^ n2428 ;
  assign n2433 = n2432 ^ n2430 ;
  assign n2426 = n456 ^ n304 ;
  assign n2427 = n2426 ^ n447 ;
  assign n2434 = n2433 ^ n2427 ;
  assign n2420 = n350 ^ n298 ;
  assign n2421 = n2420 ^ n322 ;
  assign n2424 = n2423 ^ n2421 ;
  assign n2425 = n2424 ^ n1019 ;
  assign n2435 = n2434 ^ n2425 ;
  assign n2415 = n410 ^ n176 ;
  assign n2416 = n2415 ^ n437 ;
  assign n2417 = n2416 ^ n645 ;
  assign n2418 = n2417 ^ n1060 ;
  assign n2419 = n2418 ^ n1014 ;
  assign n2436 = n2435 ^ n2419 ;
  assign n2437 = n2414 & ~n2436 ;
  assign n2440 = n2439 ^ n2437 ;
  assign n2441 = n2188 ^ n2185 ;
  assign n2476 = n2441 ^ n2180 ;
  assign n2460 = n645 ^ n577 ;
  assign n2459 = n260 ^ n118 ;
  assign n2461 = n2460 ^ n2459 ;
  assign n2462 = n2461 ^ n392 ;
  assign n2463 = n2462 ^ n444 ;
  assign n2455 = n154 ^ n140 ;
  assign n2456 = n203 ^ n185 ;
  assign n2457 = n2456 ^ n858 ;
  assign n2458 = ~n2455 & ~n2457 ;
  assign n2464 = n2463 ^ n2458 ;
  assign n2453 = n398 ^ n286 ;
  assign n2454 = n2453 ^ n1013 ;
  assign n2465 = n2464 ^ n2454 ;
  assign n2452 = n55 & n105 ;
  assign n2466 = n2465 ^ n2452 ;
  assign n2471 = n306 & n432 ;
  assign n2468 = n655 ^ n449 ;
  assign n2469 = n2468 ^ n674 ;
  assign n2467 = n785 ^ n473 ;
  assign n2470 = n2469 ^ n2467 ;
  assign n2472 = n2471 ^ n2470 ;
  assign n2473 = ~n2466 & ~n2472 ;
  assign n2448 = n858 ^ n410 ;
  assign n2449 = n2448 ^ n2429 ;
  assign n2447 = n682 ^ n276 ;
  assign n2450 = n2449 ^ n2447 ;
  assign n2445 = n2273 ^ n1089 ;
  assign n2332 = n845 ^ n447 ;
  assign n2333 = n2332 ^ n161 ;
  assign n2446 = n2445 ^ n2333 ;
  assign n2451 = n2450 ^ n2446 ;
  assign n2474 = n2473 ^ n2451 ;
  assign n2475 = ~n837 & n2474 ;
  assign n2477 = n2476 ^ n2475 ;
  assign n2489 = n1035 ^ n280 ;
  assign n2490 = n2489 ^ n323 ;
  assign n2491 = n2490 ^ n415 ;
  assign n2488 = n2468 ^ n2350 ;
  assign n2492 = n2491 ^ n2488 ;
  assign n2486 = n2485 ^ n472 ;
  assign n2484 = n791 ^ n585 ;
  assign n2487 = n2486 ^ n2484 ;
  assign n2493 = n2492 ^ n2487 ;
  assign n400 = n399 ^ n398 ;
  assign n401 = n400 ^ n334 ;
  assign n2483 = n2425 ^ n401 ;
  assign n2494 = n2493 ^ n2483 ;
  assign n285 = n284 ^ n283 ;
  assign n2501 = n1010 ^ n285 ;
  assign n2497 = n479 ^ n94 ;
  assign n2498 = n2497 ^ n321 ;
  assign n2499 = n2498 ^ n155 ;
  assign n2496 = n558 ^ n344 ;
  assign n2500 = n2499 ^ n2496 ;
  assign n2502 = n2501 ^ n2500 ;
  assign n2503 = n2502 ^ n2464 ;
  assign n431 = n430 ^ n428 ;
  assign n441 = n440 ^ n431 ;
  assign n2495 = n626 ^ n441 ;
  assign n2504 = n2503 ^ n2495 ;
  assign n2505 = n2494 & n2504 ;
  assign n2479 = n1749 ^ n1726 ;
  assign n2480 = n2479 ^ n1630 ;
  assign n2481 = n2171 & n2480 ;
  assign n2478 = n1743 ^ n1728 ;
  assign n2482 = n2481 ^ n2478 ;
  assign n2506 = n2505 ^ n2482 ;
  assign n2533 = n1726 ^ n1630 ;
  assign n2534 = n2533 ^ n2171 ;
  assign n2527 = n845 ^ n413 ;
  assign n469 = n468 ^ n202 ;
  assign n2526 = n469 ^ n379 ;
  assign n2528 = n2527 ^ n2526 ;
  assign n2524 = n362 ^ n321 ;
  assign n2525 = n2524 ^ n2468 ;
  assign n2529 = n2528 ^ n2525 ;
  assign n2519 = n211 ^ n133 ;
  assign n2520 = ~n117 & n2519 ;
  assign n2521 = n2520 ^ n427 ;
  assign n2522 = n2521 ^ n577 ;
  assign n2523 = n2522 ^ n795 ;
  assign n2530 = n2529 ^ n2523 ;
  assign n2515 = n74 ^ n42 ;
  assign n2516 = ~n271 & ~n452 ;
  assign n2517 = ~n2515 & n2516 ;
  assign n2511 = n417 ^ n245 ;
  assign n2509 = n394 ^ n250 ;
  assign n2510 = n2509 ^ n192 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2513 = n2512 ^ n228 ;
  assign n2328 = n674 ^ n473 ;
  assign n2507 = n2328 ^ n2275 ;
  assign n2508 = n2507 ^ n180 ;
  assign n2514 = n2513 ^ n2508 ;
  assign n2518 = n2517 ^ n2514 ;
  assign n2531 = n2530 ^ n2518 ;
  assign n2532 = n2531 ^ n2434 ;
  assign n2535 = n2534 ^ n2532 ;
  assign n2536 = n127 & ~n1154 ;
  assign n2542 = n1083 ^ n827 ;
  assign n2543 = n2542 ^ n244 ;
  assign n2544 = n2543 ^ n1171 ;
  assign n2545 = n2544 ^ n2451 ;
  assign n2546 = n2545 ^ n2268 ;
  assign n2539 = n91 & n185 ;
  assign n2537 = n604 ^ n344 ;
  assign n2538 = n2537 ^ n115 ;
  assign n2540 = n2539 ^ n2538 ;
  assign n2541 = ~n864 & ~n2540 ;
  assign n2547 = n2546 ^ n2541 ;
  assign n2548 = n2536 & ~n2547 ;
  assign n2549 = n2548 ^ n2547 ;
  assign n2553 = n2150 ^ n1750 ;
  assign n2550 = n1832 ^ n1784 ;
  assign n2551 = n2550 ^ n2147 ;
  assign n2552 = ~n2154 & ~n2551 ;
  assign n2554 = n2553 ^ n2552 ;
  assign n2555 = ~n2549 & ~n2554 ;
  assign n2556 = n2555 ^ n2532 ;
  assign n2557 = ~n2535 & n2556 ;
  assign n2558 = n2557 ^ n2534 ;
  assign n2559 = n2558 ^ n2482 ;
  assign n2560 = ~n2506 & ~n2559 ;
  assign n2561 = n2560 ^ n2482 ;
  assign n2562 = n2561 ^ n2476 ;
  assign n2563 = n2477 & ~n2562 ;
  assign n2564 = n2563 ^ n2476 ;
  assign n2442 = n2441 ^ n2178 ;
  assign n2443 = n2180 & ~n2442 ;
  assign n2444 = n2443 ^ n2193 ;
  assign n2565 = n2564 ^ n2444 ;
  assign n402 = n401 ^ n344 ;
  assign n393 = n392 ^ n332 ;
  assign n395 = n394 ^ n393 ;
  assign n403 = n402 ^ n395 ;
  assign n420 = n419 ^ n403 ;
  assign n423 = n422 ^ n420 ;
  assign n389 = n123 & n388 ;
  assign n424 = n423 ^ n389 ;
  assign n382 = n381 ^ n377 ;
  assign n425 = n424 ^ n382 ;
  assign n2578 = n379 ^ n250 ;
  assign n2579 = n2578 ^ n296 ;
  assign n2577 = n605 ^ n161 ;
  assign n2580 = n2579 ^ n2577 ;
  assign n2576 = n577 ^ n305 ;
  assign n2581 = n2580 ^ n2576 ;
  assign n2573 = n224 ^ n201 ;
  assign n2574 = n2573 ^ n346 ;
  assign n2575 = n2574 ^ n844 ;
  assign n2582 = n2581 ^ n2575 ;
  assign n463 = n234 ^ n144 ;
  assign n464 = ~n140 & n463 ;
  assign n465 = n464 ^ n260 ;
  assign n2568 = n553 ^ n465 ;
  assign n2569 = n2568 ^ n169 ;
  assign n2566 = n280 ^ n81 ;
  assign n2567 = n2566 ^ n243 ;
  assign n2570 = n2569 ^ n2567 ;
  assign n2571 = n2570 ^ n2469 ;
  assign n2572 = n2571 ^ n1091 ;
  assign n2583 = n2582 ^ n2572 ;
  assign n2584 = ~n425 & n2583 ;
  assign n2585 = n2584 ^ n2444 ;
  assign n2586 = n2565 & ~n2585 ;
  assign n2587 = n2586 ^ n2564 ;
  assign n2588 = n2587 ^ n2439 ;
  assign n2589 = n2440 & n2588 ;
  assign n2590 = n2589 ^ n2439 ;
  assign n2591 = n2590 ^ n2412 ;
  assign n2592 = n2413 & n2591 ;
  assign n2593 = n2592 ^ n2412 ;
  assign n2594 = n2593 ^ n2353 ;
  assign n2595 = n2384 & n2594 ;
  assign n2596 = n2595 ^ n2353 ;
  assign n2599 = n2596 ^ n2287 ;
  assign n2343 = n1278 ^ n1272 ;
  assign n2341 = n2220 ^ n1271 ;
  assign n2344 = n2341 ^ n1278 ;
  assign n2345 = n2344 ^ n1275 ;
  assign n2346 = ~n2343 & ~n2345 ;
  assign n2347 = n2346 ^ n944 ;
  assign n2340 = n2220 ^ n1275 ;
  assign n2342 = n2340 & ~n2341 ;
  assign n2348 = n2347 ^ n2342 ;
  assign n2324 = n647 ^ n427 ;
  assign n2323 = n350 ^ n181 ;
  assign n2325 = n2324 ^ n2323 ;
  assign n2326 = n2325 ^ n643 ;
  assign n2322 = n2321 ^ n545 ;
  assign n2327 = n2326 ^ n2322 ;
  assign n2335 = n519 ^ n506 ;
  assign n2330 = n381 ^ n179 ;
  assign n2329 = n2328 ^ n831 ;
  assign n2331 = n2330 ^ n2329 ;
  assign n2334 = n2333 ^ n2331 ;
  assign n2336 = n2335 ^ n2334 ;
  assign n2337 = n2336 ^ n640 ;
  assign n2338 = ~n2327 & ~n2337 ;
  assign n2339 = n2316 & n2338 ;
  assign n2349 = n2348 ^ n2339 ;
  assign n2597 = n2596 ^ n2348 ;
  assign n2598 = n2349 & ~n2597 ;
  assign n2600 = n2599 ^ n2598 ;
  assign n2601 = ~n2304 & n2600 ;
  assign n2602 = n2601 ^ n2303 ;
  assign n2603 = n2602 ^ n2249 ;
  assign n2604 = ~n2286 & ~n2603 ;
  assign n2605 = n2604 ^ n2249 ;
  assign n461 = n460 ^ n441 ;
  assign n480 = n479 ^ n348 ;
  assign n482 = n481 ^ n480 ;
  assign n483 = n482 ^ n308 ;
  assign n476 = ~n79 & n432 ;
  assign n474 = n473 ^ n472 ;
  assign n475 = n474 ^ n256 ;
  assign n477 = n476 ^ n475 ;
  assign n484 = n483 ^ n477 ;
  assign n470 = n469 ^ n120 ;
  assign n462 = n298 ^ n170 ;
  assign n466 = n465 ^ n462 ;
  assign n471 = n470 ^ n466 ;
  assign n485 = n484 ^ n471 ;
  assign n486 = ~n461 & n485 ;
  assign n487 = ~n425 & n486 ;
  assign n2606 = n2605 ^ n487 ;
  assign n2608 = ~n708 & ~n2240 ;
  assign n2609 = n2608 ^ n2240 ;
  assign n2610 = ~n707 & n2609 ;
  assign n2611 = ~n614 & n2610 ;
  assign n2612 = n2611 ^ n2244 ;
  assign n2613 = ~n2238 & n2246 ;
  assign n2614 = ~n2612 & n2613 ;
  assign n2615 = n2614 ^ n2238 ;
  assign n5665 = ~n708 & n2240 ;
  assign n2618 = ~n614 & n5665 ;
  assign n2619 = n2243 & n2618 ;
  assign n2620 = ~n2615 & n2619 ;
  assign n2607 = n2238 ^ n487 ;
  assign n2616 = n2615 ^ n2607 ;
  assign n2621 = n2620 ^ n2616 ;
  assign n2622 = ~n2606 & ~n2621 ;
  assign n2623 = n2622 ^ n2605 ;
  assign n2627 = n205 ^ n185 ;
  assign n2628 = n2627 ^ n1224 ;
  assign n2629 = ~n79 & n2628 ;
  assign n2625 = n1485 ^ n330 ;
  assign n2624 = n468 ^ n181 ;
  assign n2626 = n2625 ^ n2624 ;
  assign n2630 = n2629 ^ n2626 ;
  assign n2631 = n2630 ^ n2434 ;
  assign n2635 = n791 ^ n606 ;
  assign n2636 = n2635 ^ n108 ;
  assign n2633 = n674 ^ n345 ;
  assign n2632 = n231 ^ n225 ;
  assign n2634 = n2633 ^ n2632 ;
  assign n2637 = n2636 ^ n2634 ;
  assign n2638 = n2637 ^ n2273 ;
  assign n2639 = n2638 ^ n1165 ;
  assign n2640 = n2639 ^ n498 ;
  assign n2641 = ~n2631 & ~n2640 ;
  assign n2642 = n1526 & n2641 ;
  assign n2742 = ~n2623 & n2642 ;
  assign n2700 = n472 ^ n108 ;
  assign n2701 = n2700 ^ n251 ;
  assign n2697 = n2399 ^ n310 ;
  assign n2698 = n2697 ^ n286 ;
  assign n2699 = n2698 ^ n322 ;
  assign n2702 = n2701 ^ n2699 ;
  assign n2703 = n2702 ^ n2272 ;
  assign n2695 = ~n117 & n1145 ;
  assign n2693 = n345 ^ n81 ;
  assign n2694 = n2693 ^ n226 ;
  assign n2696 = n2695 ^ n2694 ;
  assign n2704 = n2703 ^ n2696 ;
  assign n2691 = n317 ^ n89 ;
  assign n2692 = ~n1131 & n2691 ;
  assign n2705 = n2704 ^ n2692 ;
  assign n2706 = n2705 ^ n835 ;
  assign n2710 = n2258 ^ n381 ;
  assign n2709 = n2511 ^ n1186 ;
  assign n2711 = n2710 ^ n2709 ;
  assign n2707 = n276 ^ n181 ;
  assign n2708 = n2707 ^ n607 ;
  assign n2712 = n2711 ^ n2708 ;
  assign n266 = n265 ^ n202 ;
  assign n268 = n267 ^ n266 ;
  assign n264 = n263 ^ n260 ;
  assign n269 = n268 ^ n264 ;
  assign n2713 = n2712 ^ n269 ;
  assign n2714 = n2713 ^ n856 ;
  assign n2715 = n2706 & n2714 ;
  assign n2787 = n2742 ^ n2715 ;
  assign n2743 = ~n2715 & ~n2742 ;
  assign n3673 = n2787 ^ n2743 ;
  assign n3692 = n3691 ^ n3673 ;
  assign n3805 = n3692 ^ n1473 ;
  assign n3802 = x22 ^ x1 ;
  assign n3735 = ~n3673 & n3691 ;
  assign n3720 = n2627 ^ n74 ;
  assign n3721 = n124 & n3720 ;
  assign n3722 = n3721 ^ n571 ;
  assign n3728 = ~n126 & n502 ;
  assign n3727 = n1032 ^ n437 ;
  assign n3729 = n3728 ^ n3727 ;
  assign n3726 = n468 ^ n186 ;
  assign n3730 = n3729 ^ n3726 ;
  assign n3731 = n3730 ^ n584 ;
  assign n3732 = n3731 ^ n613 ;
  assign n3723 = n110 ^ n79 ;
  assign n3724 = n500 ^ n137 ;
  assign n3725 = ~n3723 & n3724 ;
  assign n3733 = n3732 ^ n3725 ;
  assign n3734 = n3722 & ~n3733 ;
  assign n3763 = n3735 ^ n3734 ;
  assign n3803 = n3802 ^ n3763 ;
  assign n2673 = n487 & ~n2605 ;
  assign n2674 = n2673 ^ n2606 ;
  assign n2679 = n2612 & ~n2618 ;
  assign n2680 = n2679 ^ n2238 ;
  assign n2681 = n2248 & ~n2680 ;
  assign n2682 = n2674 & ~n2681 ;
  assign n2717 = n2602 ^ n2286 ;
  assign n2718 = n2600 ^ n2303 ;
  assign n2719 = n2596 ^ n2349 ;
  assign n2720 = n2593 ^ n2384 ;
  assign n2721 = n2590 ^ n2413 ;
  assign n2722 = n2587 ^ n2440 ;
  assign n2723 = n2585 ^ n2564 ;
  assign n2724 = n2561 ^ n2477 ;
  assign n2725 = n2558 ^ n2506 ;
  assign n2744 = n2554 ^ n2549 ;
  assign n2745 = ~n2535 & n2744 ;
  assign n2746 = n2745 ^ n2744 ;
  assign n2726 = n2555 ^ n2535 ;
  assign n2747 = n2746 ^ n2726 ;
  assign n2748 = ~n2725 & ~n2747 ;
  assign n2749 = n2724 & ~n2748 ;
  assign n2750 = n2723 & ~n2749 ;
  assign n2751 = ~n2722 & ~n2750 ;
  assign n2752 = n2721 & ~n2751 ;
  assign n2753 = ~n2720 & ~n2752 ;
  assign n2754 = ~n2719 & ~n2753 ;
  assign n2755 = n2718 & ~n2754 ;
  assign n2756 = ~n2717 & ~n2755 ;
  assign n2761 = n2682 & ~n2756 ;
  assign n2683 = n2673 & n2681 ;
  assign n2757 = ~n2683 & n2756 ;
  assign n2758 = ~n2623 & n2757 ;
  assign n2759 = n2758 ^ n2683 ;
  assign n2760 = n2759 ^ n2623 ;
  assign n2762 = n2761 ^ n2760 ;
  assign n2763 = n2642 & n2762 ;
  assign n2764 = n2763 ^ n2759 ;
  assign n2765 = n2743 & ~n2764 ;
  assign n3751 = ~n2765 & n3691 ;
  assign n2716 = n2715 ^ n2642 ;
  assign n2684 = n2683 ^ n2682 ;
  assign n2685 = n2684 ^ n2623 ;
  assign n2727 = n2725 & n2726 ;
  assign n2728 = ~n2724 & ~n2727 ;
  assign n2729 = ~n2723 & ~n2728 ;
  assign n2730 = n2722 & ~n2729 ;
  assign n2731 = ~n2721 & ~n2730 ;
  assign n2732 = n2720 & ~n2731 ;
  assign n2733 = n2719 & ~n2732 ;
  assign n2734 = ~n2718 & ~n2733 ;
  assign n2735 = n2717 & ~n2734 ;
  assign n2736 = n2685 & ~n2735 ;
  assign n2737 = n2736 ^ n2715 ;
  assign n2738 = n2716 & n2737 ;
  assign n2739 = n2736 ^ n2623 ;
  assign n2740 = n2738 & n2739 ;
  assign n2741 = n2740 ^ n2715 ;
  assign n3719 = ~n2741 & ~n3691 ;
  assign n3800 = n3751 ^ n3719 ;
  assign n3801 = n28 & n3800 ;
  assign n3804 = n3803 ^ n3801 ;
  assign n3806 = n3805 ^ n3804 ;
  assign n3797 = x2 & ~n2787 ;
  assign n3792 = n3692 ^ x22 ;
  assign n3798 = n3797 ^ n3792 ;
  assign n3799 = ~x1 & ~n3798 ;
  assign n3807 = n3806 ^ n3799 ;
  assign n3808 = ~x0 & ~n3807 ;
  assign n3809 = n3808 ^ n3804 ;
  assign n2648 = x22 & n29 ;
  assign n2649 = n2648 ^ n28 ;
  assign n4656 = ~n29 & n2649 ;
  assign n4663 = n4656 ^ n2649 ;
  assign n3821 = n28 & ~n30 ;
  assign n2645 = x0 & ~x22 ;
  assign n2644 = x0 & x2 ;
  assign n2646 = n2645 ^ n2644 ;
  assign n3776 = ~n3821 ^ n2646 ;
  assign n4664 = n4663 ^ n3776 ;
  assign n2667 = ~n4664 ^ n1481 ;
  assign n2781 = n2762 ^ n2735 ;
  assign n2782 = n2781 ^ n2736 ;
  assign n2783 = n2782 ^ n2735 ;
  assign n3626 = ~n2667 & n2783 ;
  assign n2643 = n2642 ^ n2623 ;
  assign n3627 = n2643 ^ n1406 ;
  assign n2668 = ~n1406 & ~n2667 ;
  assign n2669 = n2668 ^ n1406 ;
  assign n2663 = ~n1481 & n4664 ;
  assign n2664 = ~n4664 ^ n2663 ;
  assign n2665 = ~n1406 & ~n2664 ;
  assign n2670 = n2669 ^ n2665 ;
  assign n3635 = ~n2670 & ~n2685 ;
  assign n2666 = n2665 ^ n2664 ;
  assign n2671 = n2670 ^ n2666 ;
  assign n3386 = n2671 ^ n2667 ;
  assign n2773 = n2665 ^ n1357 ;
  assign n3387 = n3386 ^ n2773 ;
  assign n3384 = n1357 & ~n2671 ;
  assign n2688 = n1357 & n2667 ;
  assign n3385 = n3384 ^ n2688 ;
  assign n3388 = n3387 ^ n3385 ;
  assign n3389 = n3388 ^ n2665 ;
  assign n3380 = ~n1357 & n2665 ;
  assign n3422 = n3389 ^ n3380 ;
  assign n3634 = n2717 & n3422 ;
  assign n3636 = n3635 ^ n3634 ;
  assign n3398 = n2685 ^ n1406 ;
  assign n3628 = n3398 ^ n2685 ;
  assign n3629 = n1357 & n2717 ;
  assign n3630 = n3629 ^ n2685 ;
  assign n3631 = ~n3628 & ~n3630 ;
  assign n3632 = n3631 ^ n2685 ;
  assign n3633 = ~n2664 & ~n3632 ;
  assign n3637 = n3636 ^ n3633 ;
  assign n3639 = ~n1357 & ~n3637 ;
  assign n3638 = n3637 ^ n1357 ;
  assign n3640 = n3639 ^ n3638 ;
  assign n3641 = ~n3627 & n3640 ;
  assign n3642 = n3626 & n3641 ;
  assign n3643 = n3642 ^ n3640 ;
  assign n3464 = n1357 & ~n2667 ;
  assign n2780 = n2684 ^ n2642 ;
  assign n2784 = ~n2780 & ~n2783 ;
  assign n3623 = n2784 ^ n2736 ;
  assign n3624 = n3623 ^ n2783 ;
  assign n3625 = n3464 & ~n3624 ;
  assign n3645 = n3643 ^ n3625 ;
  assign n3646 = n3645 ^ n3639 ;
  assign n3647 = n3646 ^ n3645 ;
  assign n3648 = ~n2667 & ~n3623 ;
  assign n3649 = n3647 & n3648 ;
  assign n3650 = n3649 ^ n3646 ;
  assign n2003 = n1357 ^ n1129 ;
  assign n3282 = n2003 & n2718 ;
  assign n2801 = n2754 ^ n2733 ;
  assign n2797 = n1357 ^ n999 ;
  assign n2798 = n1129 ^ n995 ;
  assign n2799 = ~n2003 & n2798 ;
  assign n2800 = n2797 & n2799 ;
  assign n3274 = n2801 ^ n2800 ;
  assign n3276 = n2800 ^ n2720 ;
  assign n3280 = ~n3274 & n3276 ;
  assign n2809 = n1129 & n1357 ;
  assign n2810 = n2809 ^ n2003 ;
  assign n2808 = n999 & ~n2003 ;
  assign n2811 = n2810 ^ n2808 ;
  assign n3273 = ~n2801 & n2811 ;
  assign n3275 = n3274 ^ n995 ;
  assign n3277 = n3276 ^ n3275 ;
  assign n3278 = n3273 & ~n3277 ;
  assign n3272 = n2733 ^ n995 ;
  assign n3279 = n3278 ^ n3272 ;
  assign n3281 = n3280 ^ n3279 ;
  assign n3283 = n3282 ^ n3281 ;
  assign n3269 = ~n999 & ~n2801 ;
  assign n3270 = n3269 ^ n2754 ;
  assign n3271 = n2811 & ~n3270 ;
  assign n3284 = n3283 ^ n3271 ;
  assign n2842 = n708 & n2239 ;
  assign n2843 = n2842 ^ n2608 ;
  assign n2844 = n2726 & n2843 ;
  assign n2837 = n707 & ~n2240 ;
  assign n2838 = n2837 ^ n2240 ;
  assign n2835 = ~n707 & n2239 ;
  assign n2836 = n2835 ^ n2239 ;
  assign n2839 = n2838 ^ n2836 ;
  assign n2840 = n709 & ~n2839 ;
  assign n2841 = ~n2744 & n2840 ;
  assign n2845 = n2844 ^ n2841 ;
  assign n2828 = n2746 ^ n2725 ;
  assign n2829 = n2828 ^ n2725 ;
  assign n2830 = n2725 ^ n709 ;
  assign n2831 = n2830 ^ n2725 ;
  assign n2832 = n2829 & n2831 ;
  assign n2833 = n2832 ^ n2725 ;
  assign n2834 = n697 & n2833 ;
  assign n2846 = n2845 ^ n2834 ;
  assign n2847 = n2838 ^ n2239 ;
  assign n2848 = n2239 ^ n708 ;
  assign n2849 = ~n2744 & ~n2848 ;
  assign n2850 = n2849 ^ n2239 ;
  assign n2851 = ~n2847 & ~n2850 ;
  assign n2852 = n2851 ^ n2239 ;
  assign n2853 = ~n2745 & ~n2852 ;
  assign n2854 = ~n2846 & ~n2853 ;
  assign n3092 = n2854 ^ n2744 ;
  assign n2855 = n2748 ^ n2727 ;
  assign n2856 = n2855 ^ n2724 ;
  assign n2857 = n2856 ^ n2724 ;
  assign n2858 = n2724 ^ n709 ;
  assign n2859 = n2858 ^ n2724 ;
  assign n2860 = ~n2857 & n2859 ;
  assign n2861 = n2860 ^ n2724 ;
  assign n2862 = n697 & ~n2861 ;
  assign n2868 = n2862 ^ n2239 ;
  assign n2869 = n2868 ^ n2862 ;
  assign n2864 = ~n707 & n708 ;
  assign n2870 = n2864 ^ n709 ;
  assign n2871 = n2726 & n2870 ;
  assign n2872 = n2869 & n2871 ;
  assign n2873 = n2872 ^ n2868 ;
  assign n2865 = ~n2240 & n2864 ;
  assign n2866 = n2726 & n2865 ;
  assign n2863 = n2862 ^ n2240 ;
  assign n2867 = n2866 ^ n2863 ;
  assign n2874 = n2873 ^ n2867 ;
  assign n2875 = n2867 ^ n2862 ;
  assign n2876 = n2875 ^ n708 ;
  assign n2879 = ~n2725 & ~n2876 ;
  assign n2880 = n2879 ^ n708 ;
  assign n2881 = ~n2874 & n2880 ;
  assign n2882 = n2881 ^ n2873 ;
  assign n3093 = n2882 ^ n707 ;
  assign n3094 = n2854 ^ n707 ;
  assign n3095 = n3094 ^ n707 ;
  assign n3096 = ~n3093 & n3095 ;
  assign n3097 = n3096 ^ n707 ;
  assign n3098 = n3092 & ~n3097 ;
  assign n1256 = n995 ^ n778 ;
  assign n2972 = n2751 ^ n2730 ;
  assign n3086 = n1256 & ~n2972 ;
  assign n3087 = n2721 ^ n780 ;
  assign n3088 = n3086 & n3087 ;
  assign n2914 = n780 & n1256 ;
  assign n2922 = n2914 ^ n1256 ;
  assign n2923 = n2922 ^ n780 ;
  assign n2916 = n778 & n995 ;
  assign n2917 = n2916 ^ n1256 ;
  assign n2924 = n2923 ^ n2917 ;
  assign n3074 = ~n2722 & n2924 ;
  assign n1814 = n780 ^ n694 ;
  assign n2918 = n2917 ^ n694 ;
  assign n2919 = n1814 & n2918 ;
  assign n2915 = ~n694 & n2914 ;
  assign n2920 = n2919 ^ n2915 ;
  assign n3073 = ~n2723 & n2920 ;
  assign n3075 = n3074 ^ n3073 ;
  assign n3076 = n3075 ^ n694 ;
  assign n3079 = n3076 ^ n2721 ;
  assign n3082 = ~n2972 & n3079 ;
  assign n3083 = n3082 ^ n2721 ;
  assign n3084 = n1256 & ~n3083 ;
  assign n3085 = n3084 ^ n3076 ;
  assign n3089 = n3088 ^ n3085 ;
  assign n3091 = n3089 ^ n2882 ;
  assign n3099 = n3098 ^ n3091 ;
  assign n3001 = ~n707 & n2853 ;
  assign n3002 = n3001 ^ n2846 ;
  assign n2967 = n2750 ^ n2729 ;
  assign n2968 = n2722 & n2922 ;
  assign n2969 = ~n2967 & n2968 ;
  assign n2970 = n2969 ^ n1256 ;
  assign n2971 = n2970 ^ n2969 ;
  assign n2973 = n2972 ^ n2750 ;
  assign n2976 = n2971 & n2973 ;
  assign n2977 = n2976 ^ n2969 ;
  assign n2979 = ~n2723 & n2924 ;
  assign n2978 = n2724 & n2920 ;
  assign n2980 = n2979 ^ n2978 ;
  assign n2981 = n2980 ^ n694 ;
  assign n2982 = n2981 ^ n2969 ;
  assign n2983 = n2982 ^ n2980 ;
  assign n2984 = n2977 & ~n2983 ;
  assign n2985 = n2984 ^ n2981 ;
  assign n2988 = ~n2967 & ~n2980 ;
  assign n2989 = n2988 ^ n1256 ;
  assign n2990 = ~n694 & n2989 ;
  assign n2991 = n2990 ^ n1256 ;
  assign n2992 = n2985 & n2991 ;
  assign n2997 = n780 & ~n2967 ;
  assign n2993 = n2967 ^ n2722 ;
  assign n2998 = n2997 ^ n2993 ;
  assign n2999 = n2992 & n2998 ;
  assign n3000 = n2999 ^ n2985 ;
  assign n3003 = n3002 ^ n3000 ;
  assign n3045 = ~n708 & ~n2744 ;
  assign n3037 = n2744 ^ n2726 ;
  assign n3038 = n3037 ^ n2726 ;
  assign n3041 = n694 & ~n3038 ;
  assign n3042 = n3041 ^ n2726 ;
  assign n3043 = ~n697 & n3042 ;
  assign n3044 = n3043 ^ n2726 ;
  assign n3046 = n3045 ^ n3044 ;
  assign n3004 = n697 & ~n2744 ;
  assign n3011 = n2726 & n2924 ;
  assign n3010 = ~n2744 & n2920 ;
  assign n3012 = n3011 ^ n3010 ;
  assign n3005 = n2725 ^ n1814 ;
  assign n3006 = n3005 ^ n2725 ;
  assign n3007 = n2829 & n3006 ;
  assign n3008 = n3007 ^ n2725 ;
  assign n3009 = n1256 & n3008 ;
  assign n3013 = n3012 ^ n3009 ;
  assign n3014 = n2535 ^ n781 ;
  assign n3015 = n1256 & ~n3014 ;
  assign n3016 = n3015 ^ n781 ;
  assign n3017 = n2744 ^ n1256 ;
  assign n3018 = n3017 ^ n694 ;
  assign n3019 = n3016 & n3018 ;
  assign n3020 = n3019 ^ n1256 ;
  assign n3021 = n694 & n3020 ;
  assign n3022 = n3021 ^ n694 ;
  assign n3023 = ~n3013 & n3022 ;
  assign n3024 = ~n3004 & ~n3023 ;
  assign n3031 = n2725 & n2924 ;
  assign n3030 = n2726 & n2920 ;
  assign n3032 = n3031 ^ n3030 ;
  assign n3033 = n3032 ^ n694 ;
  assign n3025 = n2724 ^ n1814 ;
  assign n3026 = n3025 ^ n2724 ;
  assign n3027 = ~n2857 & n3026 ;
  assign n3028 = n3027 ^ n2724 ;
  assign n3029 = n1256 & n3028 ;
  assign n3034 = n3033 ^ n3029 ;
  assign n3035 = n3024 & n3034 ;
  assign n3036 = n3035 ^ n3034 ;
  assign n3047 = n3046 ^ n3036 ;
  assign n3055 = n1256 & ~n2723 ;
  assign n3052 = n2723 ^ n780 ;
  assign n3049 = n2724 & n2924 ;
  assign n3048 = n2725 & n2920 ;
  assign n3050 = n3049 ^ n3048 ;
  assign n3051 = n3050 ^ n694 ;
  assign n3053 = n3052 ^ n3051 ;
  assign n3054 = n3053 ^ n3052 ;
  assign n3056 = n3055 ^ n3054 ;
  assign n3057 = n3056 ^ n3052 ;
  assign n2888 = n2749 ^ n2728 ;
  assign n3058 = n1256 & ~n2888 ;
  assign n3059 = ~n3057 & n3058 ;
  assign n3061 = n3059 ^ n3056 ;
  assign n3066 = n3061 ^ n3046 ;
  assign n3068 = n3047 & n3066 ;
  assign n3069 = n3068 ^ n3046 ;
  assign n3070 = n3069 ^ n3002 ;
  assign n3071 = ~n3003 & n3070 ;
  assign n3072 = n3071 ^ n3069 ;
  assign n3265 = n3099 ^ n3072 ;
  assign n3620 = n3284 ^ n3265 ;
  assign n3116 = n3069 ^ n3003 ;
  assign n3113 = ~n2720 & ~n2811 ;
  assign n2909 = n2753 ^ n2732 ;
  assign n3105 = n2811 & ~n2909 ;
  assign n3111 = n999 & n3105 ;
  assign n3108 = n2909 ^ n2721 ;
  assign n3109 = n2800 & n3108 ;
  assign n3110 = n3109 ^ n2811 ;
  assign n3112 = n3111 ^ n3110 ;
  assign n3114 = n3113 ^ n3112 ;
  assign n2819 = n2811 ^ n995 ;
  assign n3106 = n2819 & ~n3105 ;
  assign n3104 = n2003 & n2719 ;
  assign n3107 = n3106 ^ n3104 ;
  assign n3115 = n3114 ^ n3107 ;
  assign n3117 = n3116 ^ n3115 ;
  assign n2910 = n2909 ^ n2752 ;
  assign n3120 = n2003 & n2910 ;
  assign n3119 = n2720 ^ n999 ;
  assign n3121 = n3120 ^ n3119 ;
  assign n2928 = n2752 ^ n2731 ;
  assign n3124 = n2003 & ~n2928 ;
  assign n3131 = ~n3121 & ~n3124 ;
  assign n3139 = n3131 ^ n3120 ;
  assign n3129 = ~n2722 & n2800 ;
  assign n3127 = ~n2721 & ~n2811 ;
  assign n3125 = n3124 ^ n995 ;
  assign n3126 = n3125 ^ n3120 ;
  assign n3128 = n3127 ^ n3126 ;
  assign n3130 = n3129 ^ n3128 ;
  assign n3132 = n3131 ^ n3121 ;
  assign n3133 = n3132 ^ n3120 ;
  assign n3134 = n3120 ^ n995 ;
  assign n3135 = n3134 ^ n3120 ;
  assign n3136 = ~n3133 & ~n3135 ;
  assign n3137 = n3136 ^ n3120 ;
  assign n3138 = n3130 & ~n3137 ;
  assign n3140 = n3139 ^ n3138 ;
  assign n3123 = n3121 ^ n3120 ;
  assign n3141 = n3140 ^ n3123 ;
  assign n3118 = n3066 ^ n3036 ;
  assign n3142 = n3141 ^ n3118 ;
  assign n3162 = n2972 ^ n2723 ;
  assign n3163 = ~n2800 & n3162 ;
  assign n3159 = n2003 & ~n2721 ;
  assign n3153 = n2972 ^ n2819 ;
  assign n3156 = n2811 & ~n2972 ;
  assign n3157 = n3153 & n3156 ;
  assign n3152 = n2723 ^ n2722 ;
  assign n3154 = n3153 ^ n3152 ;
  assign n3158 = n3157 ^ n3154 ;
  assign n3160 = n3159 ^ n3158 ;
  assign n3147 = n2722 ^ n999 ;
  assign n3148 = n3147 ^ n2722 ;
  assign n3149 = ~n2972 & n3148 ;
  assign n3150 = n3149 ^ n2722 ;
  assign n3151 = n2811 & n3150 ;
  assign n3161 = n3160 ^ n3151 ;
  assign n3164 = n3163 ^ n3161 ;
  assign n3143 = n3023 ^ n3004 ;
  assign n3144 = n3143 ^ n3034 ;
  assign n3165 = n3164 ^ n3144 ;
  assign n3191 = n2967 ^ n2724 ;
  assign n3192 = ~n2800 & ~n3191 ;
  assign n3188 = n2003 & ~n2722 ;
  assign n3178 = n2811 & ~n2967 ;
  assign n3181 = n2973 ^ n995 ;
  assign n3182 = n3181 ^ n2811 ;
  assign n3180 = n2972 ^ n2729 ;
  assign n3183 = n3182 ^ n3180 ;
  assign n3186 = n3178 & ~n3183 ;
  assign n3179 = n2724 ^ n2723 ;
  assign n3184 = n3183 ^ n3179 ;
  assign n3187 = n3186 ^ n3184 ;
  assign n3189 = n3188 ^ n3187 ;
  assign n3175 = ~n999 & ~n2967 ;
  assign n3176 = n3175 ^ n2723 ;
  assign n3177 = n2811 & n3176 ;
  assign n3190 = n3189 ^ n3177 ;
  assign n3193 = n3192 ^ n3190 ;
  assign n3170 = n3021 ^ n3013 ;
  assign n3194 = n3193 ^ n3170 ;
  assign n3211 = n2724 & ~n2811 ;
  assign n3210 = n2725 & n2800 ;
  assign n3212 = n3211 ^ n3210 ;
  assign n3203 = n2723 ^ n995 ;
  assign n3204 = n3203 ^ n999 ;
  assign n3205 = n3204 ^ n2723 ;
  assign n3206 = ~n2888 & ~n3205 ;
  assign n3207 = n3206 ^ n2723 ;
  assign n3208 = n2003 & ~n3207 ;
  assign n3209 = n3208 ^ n995 ;
  assign n3213 = n3212 ^ n3209 ;
  assign n3252 = n3213 ^ n3170 ;
  assign n3196 = n2726 ^ n995 ;
  assign n3197 = n3196 ^ n2726 ;
  assign n3198 = ~n3038 & n3197 ;
  assign n3199 = n3198 ^ n2726 ;
  assign n3200 = ~n1256 & n3199 ;
  assign n3201 = n3200 ^ n2726 ;
  assign n3195 = n780 & ~n2744 ;
  assign n3202 = n3201 ^ n3195 ;
  assign n3214 = n3213 ^ n3202 ;
  assign n3215 = n1256 & ~n2744 ;
  assign n3216 = n2809 ^ n2808 ;
  assign n3217 = n995 & ~n3216 ;
  assign n3218 = n2003 & n2726 ;
  assign n3219 = n2744 & ~n3218 ;
  assign n3220 = n3217 & n3219 ;
  assign n3221 = n3220 ^ n3217 ;
  assign n3222 = n3221 ^ n995 ;
  assign n3229 = n2726 & ~n2811 ;
  assign n3228 = ~n2744 & n2800 ;
  assign n3230 = n3229 ^ n3228 ;
  assign n3223 = n2725 ^ n1000 ;
  assign n3224 = n3223 ^ n2725 ;
  assign n3225 = n2829 & ~n3224 ;
  assign n3226 = n3225 ^ n2725 ;
  assign n3227 = n2003 & n3226 ;
  assign n3231 = n3230 ^ n3227 ;
  assign n3232 = n3222 & ~n3231 ;
  assign n3234 = n3215 & n3232 ;
  assign n3233 = n3232 ^ n3215 ;
  assign n3235 = n3234 ^ n3233 ;
  assign n3242 = n2855 ^ n2726 ;
  assign n3243 = ~n2800 & ~n3242 ;
  assign n3237 = n2811 & ~n2855 ;
  assign n3241 = n999 & n3237 ;
  assign n3244 = n3243 ^ n3241 ;
  assign n3245 = n3244 ^ n2726 ;
  assign n3240 = n2725 & ~n2811 ;
  assign n3246 = n3245 ^ n3240 ;
  assign n3238 = n2855 ^ n995 ;
  assign n3239 = ~n3237 & ~n3238 ;
  assign n3247 = n3246 ^ n3239 ;
  assign n3236 = n2003 & n2724 ;
  assign n3248 = n3247 ^ n3236 ;
  assign n3249 = n3235 & n3248 ;
  assign n3250 = n3249 ^ n3202 ;
  assign n3251 = n3214 & ~n3250 ;
  assign n3253 = n3252 ^ n3251 ;
  assign n3254 = n3194 & ~n3253 ;
  assign n3255 = n3254 ^ n3193 ;
  assign n3256 = n3255 ^ n3164 ;
  assign n3257 = ~n3165 & ~n3256 ;
  assign n3258 = n3257 ^ n3164 ;
  assign n3259 = n3258 ^ n3141 ;
  assign n3260 = ~n3142 & n3259 ;
  assign n3261 = n3260 ^ n3141 ;
  assign n3262 = n3261 ^ n3116 ;
  assign n3263 = ~n3117 & ~n3262 ;
  assign n3264 = n3263 ^ n3261 ;
  assign n3621 = n3620 ^ n3264 ;
  assign n2785 = n1406 ^ n1357 ;
  assign n3399 = n3398 ^ n2785 ;
  assign n3400 = n3399 ^ n3398 ;
  assign n3362 = n2756 ^ n2735 ;
  assign n3401 = n3398 ^ n3362 ;
  assign n3402 = n3401 ^ n3398 ;
  assign n3403 = n3400 & n3402 ;
  assign n3404 = n3403 ^ n3398 ;
  assign n3405 = ~n2667 & n3404 ;
  assign n3379 = n2717 ^ n1357 ;
  assign n3382 = n2671 & ~n3379 ;
  assign n3383 = n3382 ^ n3380 ;
  assign n3395 = ~n2718 & n3388 ;
  assign n3396 = n3395 ^ n2665 ;
  assign n3397 = ~n3383 & ~n3396 ;
  assign n3406 = n3405 ^ n3397 ;
  assign n3378 = n3261 ^ n3117 ;
  assign n3407 = n3406 ^ n3378 ;
  assign n3433 = n3258 ^ n3142 ;
  assign n3411 = n2717 ^ n1406 ;
  assign n2802 = n2734 ^ n2733 ;
  assign n2803 = n2802 ^ n2755 ;
  assign n2804 = n2803 ^ n2801 ;
  assign n2805 = n2804 ^ n2754 ;
  assign n3412 = ~n2667 & ~n2805 ;
  assign n3413 = n3411 & n3412 ;
  assign n2690 = n3464 ^ n2667 ;
  assign n3408 = n3362 ^ n2755 ;
  assign n3410 = ~n2690 & ~n3408 ;
  assign n3414 = n3413 ^ n3410 ;
  assign n3424 = ~n2670 & n2718 ;
  assign n3423 = n2719 & n3422 ;
  assign n3425 = n3424 ^ n3423 ;
  assign n3426 = n3425 ^ n1357 ;
  assign n3415 = n2718 ^ n1406 ;
  assign n3416 = n3415 ^ n2718 ;
  assign n3417 = n1357 & n2719 ;
  assign n3418 = n3417 ^ n2718 ;
  assign n3419 = ~n3416 & n3418 ;
  assign n3420 = n3419 ^ n2718 ;
  assign n3421 = ~n2664 & n3420 ;
  assign n3427 = n3426 ^ n3421 ;
  assign n3428 = ~n3414 & n3427 ;
  assign n3431 = n3428 ^ n3414 ;
  assign n3409 = n3408 ^ n2805 ;
  assign n3429 = n3428 & n3464 ;
  assign n3430 = n3409 & n3429 ;
  assign n3432 = n3431 ^ n3430 ;
  assign n3434 = n3433 ^ n3432 ;
  assign n3444 = ~n2803 & n3464 ;
  assign n3439 = n2671 & n2719 ;
  assign n3438 = ~n2720 & n3388 ;
  assign n3440 = n3439 ^ n3438 ;
  assign n3442 = ~n1357 & ~n3440 ;
  assign n3441 = n3440 ^ n1357 ;
  assign n3443 = n3442 ^ n3441 ;
  assign n3445 = n3444 ^ n3443 ;
  assign n3436 = ~n2667 & ~n2801 ;
  assign n3437 = ~n3415 & n3436 ;
  assign n3446 = n3445 ^ n3437 ;
  assign n3447 = n3446 ^ n3442 ;
  assign n3448 = n3447 ^ n3446 ;
  assign n3449 = ~n2667 & n2804 ;
  assign n3450 = n3448 & n3449 ;
  assign n3451 = n3450 ^ n3447 ;
  assign n3435 = n3255 ^ n3165 ;
  assign n3452 = n3451 ^ n3435 ;
  assign n3314 = n2801 ^ n2732 ;
  assign n3457 = n2671 & ~n2720 ;
  assign n3456 = ~n2721 & n3388 ;
  assign n3458 = n3457 ^ n3456 ;
  assign n3465 = n3314 & ~n3458 ;
  assign n3466 = n3464 & n3465 ;
  assign n3460 = ~n2667 & ~n2909 ;
  assign n3461 = n2719 ^ n1406 ;
  assign n3462 = n3460 & n3461 ;
  assign n3459 = n3458 ^ n1357 ;
  assign n3463 = n3462 ^ n3459 ;
  assign n3467 = n3466 ^ n3463 ;
  assign n3454 = n2801 ^ n2753 ;
  assign n3455 = ~n2690 & ~n3454 ;
  assign n3468 = n3467 ^ n3455 ;
  assign n3453 = n3253 ^ n3193 ;
  assign n3469 = n3468 ^ n3453 ;
  assign n3489 = n3250 ^ n3213 ;
  assign n3485 = ~n2667 & ~n2928 ;
  assign n3486 = n2720 ^ n1406 ;
  assign n3487 = n3485 & n3486 ;
  assign n3473 = n2671 & ~n2721 ;
  assign n3472 = ~n2722 & n3388 ;
  assign n3474 = n3473 ^ n3472 ;
  assign n3470 = n2909 ^ n2731 ;
  assign n3471 = n3464 & ~n3470 ;
  assign n3475 = n3474 ^ n3471 ;
  assign n3476 = ~n2667 & n2910 ;
  assign n3477 = n3476 ^ n3474 ;
  assign n3478 = ~n3475 & ~n3477 ;
  assign n3479 = n3478 ^ n3474 ;
  assign n3480 = n3474 ^ n1357 ;
  assign n3483 = ~n3479 & ~n3480 ;
  assign n3481 = n3480 ^ n3471 ;
  assign n3484 = n3483 ^ n3481 ;
  assign n3488 = n3487 ^ n3484 ;
  assign n3490 = n3489 ^ n3488 ;
  assign n3575 = n3248 ^ n3235 ;
  assign n3576 = n3575 ^ n3234 ;
  assign n3508 = n3231 ^ n3221 ;
  assign n3500 = ~n2690 & ~n3180 ;
  assign n3495 = n2671 & ~n2723 ;
  assign n3494 = n2724 & n3388 ;
  assign n3496 = n3495 ^ n3494 ;
  assign n3498 = n1357 & ~n3496 ;
  assign n3497 = n3496 ^ n1357 ;
  assign n3499 = n3498 ^ n3497 ;
  assign n3501 = n3500 ^ n3499 ;
  assign n3491 = ~n2667 & ~n2967 ;
  assign n3492 = n2722 ^ n1406 ;
  assign n3493 = n3491 & ~n3492 ;
  assign n3502 = n3501 ^ n3493 ;
  assign n3503 = n3502 ^ n3498 ;
  assign n3504 = n3503 ^ n3502 ;
  assign n3505 = ~n2667 & n2973 ;
  assign n3506 = n3504 & n3505 ;
  assign n3507 = n3506 ^ n3503 ;
  assign n3509 = n3508 ^ n3507 ;
  assign n3526 = n2724 ^ n1357 ;
  assign n3514 = n2723 ^ n1357 ;
  assign n3513 = n2723 ^ n1406 ;
  assign n3515 = n3514 ^ n3513 ;
  assign n3516 = n2888 & n3515 ;
  assign n3517 = n3516 ^ n3513 ;
  assign n3527 = n3526 ^ n3517 ;
  assign n3518 = n2724 ^ n1481 ;
  assign n3519 = n3518 ^ n1357 ;
  assign n3520 = n3519 ^ n2724 ;
  assign n3523 = n2725 & ~n3520 ;
  assign n3524 = n3523 ^ n2724 ;
  assign n3525 = n1632 & n3524 ;
  assign n3528 = n3527 ^ n3525 ;
  assign n3529 = n2667 & ~n3528 ;
  assign n3530 = n3529 ^ n3517 ;
  assign n3510 = n2809 ^ n999 ;
  assign n3511 = ~n2744 & ~n3510 ;
  assign n3512 = n3511 ^ n3218 ;
  assign n3531 = n3530 ^ n3512 ;
  assign n3538 = n2671 & n2725 ;
  assign n3537 = n2726 & n3388 ;
  assign n3539 = n3538 ^ n3537 ;
  assign n3534 = n2785 & ~n2857 ;
  assign n3535 = n3534 ^ n2724 ;
  assign n3536 = ~n2667 & n3535 ;
  assign n3540 = n3539 ^ n3536 ;
  assign n3544 = n2785 & ~n3038 ;
  assign n3545 = n3544 ^ n2726 ;
  assign n3546 = n1632 & n3545 ;
  assign n3547 = n3546 ^ n2726 ;
  assign n3548 = n3547 ^ n2725 ;
  assign n3551 = n3548 ^ n2746 ;
  assign n3552 = n3551 ^ n3548 ;
  assign n3553 = n2785 & n3552 ;
  assign n3554 = n3553 ^ n3548 ;
  assign n3555 = ~n2667 & n3554 ;
  assign n3556 = n3555 ^ n3547 ;
  assign n3557 = n1357 & ~n3556 ;
  assign n3558 = ~n2745 & ~n3386 ;
  assign n3559 = n3557 & n3558 ;
  assign n3560 = n3559 ^ n3557 ;
  assign n3561 = ~n3540 & ~n3560 ;
  assign n3562 = n3561 ^ n1357 ;
  assign n3541 = n3540 ^ n1357 ;
  assign n3563 = n3562 ^ n3541 ;
  assign n3568 = n3563 ^ n3512 ;
  assign n3565 = n3561 ^ n1129 ;
  assign n3566 = ~n2744 & n3565 ;
  assign n3567 = ~n3562 & n3566 ;
  assign n3569 = n3568 ^ n3567 ;
  assign n3570 = ~n3531 & n3569 ;
  assign n3571 = n3570 ^ n3530 ;
  assign n3572 = n3571 ^ n3507 ;
  assign n3573 = n3509 & n3572 ;
  assign n3574 = n3573 ^ n3508 ;
  assign n3577 = n3576 ^ n3574 ;
  assign n3593 = n2928 ^ n2730 ;
  assign n3583 = n2671 & ~n2722 ;
  assign n3582 = ~n2723 & n3388 ;
  assign n3584 = n3583 ^ n3582 ;
  assign n3594 = n3584 ^ n1357 ;
  assign n3595 = n3594 ^ n2688 ;
  assign n3596 = n3595 ^ n3584 ;
  assign n3597 = n3593 & n3596 ;
  assign n3598 = n3597 ^ n3594 ;
  assign n3601 = n3598 ^ n3576 ;
  assign n3578 = n2721 ^ n1406 ;
  assign n3579 = n3578 ^ n2721 ;
  assign n3580 = ~n2972 & n3579 ;
  assign n3581 = n3580 ^ n2721 ;
  assign n3589 = ~n2972 & ~n3584 ;
  assign n3590 = n3589 ^ n2667 ;
  assign n3591 = n1357 & ~n3590 ;
  assign n3592 = n3591 ^ n2667 ;
  assign n3599 = ~n3592 & ~n3598 ;
  assign n3600 = ~n3581 & n3599 ;
  assign n3602 = n3601 ^ n3600 ;
  assign n3603 = n3577 & n3602 ;
  assign n3604 = n3603 ^ n3576 ;
  assign n3605 = n3604 ^ n3488 ;
  assign n3606 = n3490 & ~n3605 ;
  assign n3607 = n3606 ^ n3489 ;
  assign n3608 = n3607 ^ n3453 ;
  assign n3609 = n3469 & ~n3608 ;
  assign n3610 = n3609 ^ n3468 ;
  assign n3611 = n3610 ^ n3435 ;
  assign n3612 = ~n3452 & n3611 ;
  assign n3613 = n3612 ^ n3451 ;
  assign n3614 = n3613 ^ n3432 ;
  assign n3615 = n3434 & n3614 ;
  assign n3616 = n3615 ^ n3432 ;
  assign n3617 = n3616 ^ n3378 ;
  assign n3618 = ~n3407 & n3617 ;
  assign n3619 = n3618 ^ n3406 ;
  assign n3622 = n3621 ^ n3619 ;
  assign n3791 = n3650 ^ n3622 ;
  assign n3810 = n3809 ^ n3791 ;
  assign n4039 = n3616 ^ n3407 ;
  assign n4040 = n4039 ^ n3791 ;
  assign n2766 = n2765 ^ n2741 ;
  assign n4026 = n28 & ~n2766 ;
  assign n4027 = n4026 ^ n3692 ;
  assign n4036 = ~n4664 ^ n4027 ;
  assign n4028 = n4027 ^ n2787 ;
  assign n4029 = n4028 ^ n4027 ;
  assign n4023 = n2787 ^ n2643 ;
  assign n4030 = n4029 ^ n4023 ;
  assign n4031 = ~x2 & n4030 ;
  assign n4032 = n4031 ^ n4023 ;
  assign n4033 = ~x1 & ~n4032 ;
  assign n4034 = n4033 ^ n4028 ;
  assign n4035 = ~x0 & ~n4034 ;
  assign n4037 = n4036 ^ n4035 ;
  assign n3840 = n3607 ^ n3469 ;
  assign n3855 = ~n4664 ^ n3840 ;
  assign n3842 = n28 & ~n3362 ;
  assign n3843 = n3842 ^ n2685 ;
  assign n3856 = n3855 ^ n3843 ;
  assign n3848 = n2717 ^ x2 ;
  assign n3849 = n3848 ^ n2717 ;
  assign n3850 = n2718 & n3849 ;
  assign n3851 = n3850 ^ n2717 ;
  assign n3852 = ~x1 & n3851 ;
  assign n3844 = n3843 ^ n2717 ;
  assign n3853 = n3852 ^ n3844 ;
  assign n3854 = ~x0 & ~n3853 ;
  assign n3857 = n3856 ^ n3854 ;
  assign n3867 = n3571 ^ n3509 ;
  assign n3877 = n3569 ^ n3530 ;
  assign n3878 = ~n4664 ^ n3877 ;
  assign n3876 = n29 & ~n2721 ;
  assign n3879 = n3878 ^ n3876 ;
  assign n3875 = ~n2722 & n3821 ;
  assign n3880 = n3879 ^ n3875 ;
  assign n3872 = n28 & ~n2928 ;
  assign n3873 = n3872 ^ n2720 ;
  assign n3874 = x0 & ~n3873 ;
  assign n3881 = n3880 ^ n3874 ;
  assign n3897 = n3560 ^ n3541 ;
  assign n3898 = n3897 ^ n3565 ;
  assign n3899 = n2744 & ~n3898 ;
  assign n3900 = n3899 ^ n3565 ;
  assign n3958 = n3900 ^ n3877 ;
  assign n2650 = x0 & n28 ;
  assign n3895 = n2650 & n2993 ;
  assign n3885 = n3556 ^ n3385 ;
  assign n3886 = n3885 ^ n3556 ;
  assign n3887 = ~n2667 & n2726 ;
  assign n3888 = n2744 & ~n3887 ;
  assign n3889 = n3886 & n3888 ;
  assign n3890 = n3889 ^ n3885 ;
  assign n3891 = ~n4664 ^ n3890 ;
  assign n3779 = n2650 ^ x0 ;
  assign n3884 = ~n2722 & n3779 ;
  assign n3892 = n3891 ^ n3884 ;
  assign n3883 = n2724 & n3821 ;
  assign n3893 = n3892 ^ n3883 ;
  assign n3882 = n29 & ~n2723 ;
  assign n3894 = n3893 ^ n3882 ;
  assign n3896 = n3895 ^ n3894 ;
  assign n2889 = n2888 ^ n2723 ;
  assign n3916 = n2650 & n2889 ;
  assign n3912 = n31 ^ x0 ;
  assign n3913 = ~n2725 & ~n3912 ;
  assign n3521 = n2725 ^ n2724 ;
  assign n3910 = n29 & n3521 ;
  assign n2654 = x2 & n2645 ;
  assign n2651 = n2645 ^ x0 ;
  assign n2652 = n2651 ^ x1 ;
  assign n2653 = n2652 ^ n29 ;
  assign n2655 = n2654 ^ n2653 ;
  assign n2656 = ~n1479 & n2655 ;
  assign n2657 = n2656 ^ n2650 ;
  assign n2658 = n2657 ^ n1479 ;
  assign n2659 = n2658 ^ n2649 ;
  assign n2647 = n2646 ^ n1478 ;
  assign n2660 = n2659 ^ n2647 ;
  assign n2661 = n2660 ^ n2656 ;
  assign n3908 = n2661 ^ x0 ;
  assign n3902 = n2663 ^ n1481 ;
  assign n3903 = n3902 ^ n1406 ;
  assign n3904 = ~n2744 & ~n3903 ;
  assign n3905 = n3904 ^ n3887 ;
  assign n3909 = n3908 ^ n3905 ;
  assign n3911 = n3910 ^ n3909 ;
  assign n3914 = n3913 ^ n3911 ;
  assign n3907 = ~n2723 & n3779 ;
  assign n3915 = n3914 ^ n3907 ;
  assign n3917 = n3916 ^ n3915 ;
  assign n3927 = n2744 ^ n1481 ;
  assign n3928 = n3927 ^ n1481 ;
  assign n3929 = ~n2535 & ~n2725 ;
  assign n3930 = n3929 ^ n1481 ;
  assign n3931 = n3928 & n3930 ;
  assign n3932 = n3931 ^ n1481 ;
  assign n3933 = n3932 & ~n4664 ;
  assign n3941 = n3933 ^ n3905 ;
  assign n3924 = n29 & n2725 ;
  assign n3923 = n2726 & n3821 ;
  assign n3925 = n3924 ^ n3923 ;
  assign n3920 = n28 & ~n2857 ;
  assign n3921 = n3920 ^ n2724 ;
  assign n3922 = x0 & n3921 ;
  assign n3926 = n3925 ^ n3922 ;
  assign n3934 = n3933 ^ n2663 ;
  assign n3935 = n3934 ^ n3933 ;
  assign n3938 = ~n3928 & n3935 ;
  assign n3939 = n3938 ^ n3933 ;
  assign n3940 = n3926 & n3939 ;
  assign n3942 = n3941 ^ n3940 ;
  assign n3943 = ~n3917 & n3942 ;
  assign n3906 = n3905 ^ n3900 ;
  assign n3944 = n3943 ^ n3906 ;
  assign n3901 = n3900 ^ n3890 ;
  assign n3945 = n3944 ^ n3901 ;
  assign n3946 = ~n3896 & n3945 ;
  assign n3947 = n3946 ^ n3944 ;
  assign n3080 = n2972 ^ n2721 ;
  assign n3955 = n2650 & n3080 ;
  assign n3950 = ~n2721 & n3779 ;
  assign n3949 = ~n2723 & n3821 ;
  assign n3951 = n3950 ^ n3949 ;
  assign n3952 = ~n4664 ^ n3951 ;
  assign n3948 = n29 & ~n2722 ;
  assign n3953 = n3952 ^ n3948 ;
  assign n3954 = n3953 ^ n3900 ;
  assign n3956 = n3955 ^ n3954 ;
  assign n3957 = ~n3947 & ~n3956 ;
  assign n3959 = n3958 ^ n3957 ;
  assign n3960 = n3881 & ~n3959 ;
  assign n3961 = n3960 ^ n3877 ;
  assign n3963 = n3867 & ~n3961 ;
  assign n3962 = n3961 ^ n3867 ;
  assign n3964 = n3963 ^ n3962 ;
  assign n3973 = x2 & ~n2721 ;
  assign n3974 = n3973 ^ n2720 ;
  assign n3975 = ~x1 & ~n3974 ;
  assign n3965 = n28 & ~n2909 ;
  assign n3966 = n3965 ^ n2719 ;
  assign n3967 = n3966 ^ n2720 ;
  assign n3976 = n3975 ^ n3967 ;
  assign n3977 = ~x0 & ~n3976 ;
  assign n3978 = n3977 ^ n3966 ;
  assign n3979 = ~n4664 ^ n3978 ;
  assign n3989 = n29 & n2719 ;
  assign n3988 = ~n2720 & n3821 ;
  assign n3990 = n3989 ^ n3988 ;
  assign n3985 = n28 & ~n2801 ;
  assign n3986 = n3985 ^ n2718 ;
  assign n3987 = x0 & n3986 ;
  assign n3991 = n3990 ^ n3987 ;
  assign n3992 = n3991 ^ n3978 ;
  assign n3980 = n3602 ^ n3574 ;
  assign n3993 = n3992 ^ n3980 ;
  assign n3994 = ~n3979 & n3993 ;
  assign n3995 = ~n3964 & n3994 ;
  assign n3996 = n3980 ^ n3963 ;
  assign n3997 = ~n4664 ^ n3991 ;
  assign n3998 = n3997 ^ n3980 ;
  assign n3999 = ~n3996 & ~n3998 ;
  assign n4000 = n3999 ^ n3963 ;
  assign n4001 = ~n3995 & ~n4000 ;
  assign n4002 = ~n4664 ^ n4001 ;
  assign n3866 = n29 & n2718 ;
  assign n4003 = n4002 ^ n3866 ;
  assign n3865 = n2719 & n3821 ;
  assign n4004 = n4003 ^ n3865 ;
  assign n3862 = n28 & ~n2805 ;
  assign n3863 = n3862 ^ n2717 ;
  assign n3864 = x0 & n3863 ;
  assign n4005 = n4004 ^ n3864 ;
  assign n4006 = n4001 ^ n3840 ;
  assign n4007 = n4006 ^ n3604 ;
  assign n4008 = n4007 ^ n3490 ;
  assign n4009 = n4008 ^ n3840 ;
  assign n4010 = n4005 & n4009 ;
  assign n4011 = n4010 ^ n4006 ;
  assign n4012 = ~n3857 & n4011 ;
  assign n3834 = n28 & n2783 ;
  assign n3833 = ~n4664 ^ n2643 ;
  assign n3835 = n3834 ^ n3833 ;
  assign n3832 = n2685 ^ n1473 ;
  assign n3836 = n3835 ^ n3832 ;
  assign n3824 = n2685 ^ x22 ;
  assign n3825 = n3824 ^ n2717 ;
  assign n3826 = n3825 ^ n3824 ;
  assign n3829 = x2 & n3826 ;
  assign n3830 = n3829 ^ n3824 ;
  assign n3831 = ~x1 & n3830 ;
  assign n3837 = n3836 ^ n3831 ;
  assign n3838 = ~x0 & n3837 ;
  assign n3839 = n3838 ^ n3835 ;
  assign n3841 = n3840 ^ n3839 ;
  assign n4013 = n4012 ^ n3841 ;
  assign n4014 = n3839 ^ n3452 ;
  assign n4015 = n4014 ^ n3610 ;
  assign n4016 = n4013 & ~n4015 ;
  assign n4017 = n4016 ^ n3839 ;
  assign n3822 = n2685 & n3821 ;
  assign n3819 = n29 & n2643 ;
  assign n3817 = n2660 ^ n30 ;
  assign n3813 = n2787 ^ n2657 ;
  assign n3814 = n2784 ^ x0 ;
  assign n3815 = ~n3813 & ~n3814 ;
  assign n3811 = n2787 ^ n2656 ;
  assign n3812 = ~n2784 & ~n3811 ;
  assign n3816 = n3815 ^ n3812 ;
  assign n3818 = n3817 ^ n3816 ;
  assign n3820 = n3819 ^ n3818 ;
  assign n3823 = n3822 ^ n3820 ;
  assign n4018 = n4017 ^ n3823 ;
  assign n4019 = n3823 ^ n3434 ;
  assign n4020 = n4019 ^ n3613 ;
  assign n4021 = ~n4018 & n4020 ;
  assign n4022 = n4021 ^ n4017 ;
  assign n4038 = n4037 ^ n4022 ;
  assign n4041 = n4040 ^ n4038 ;
  assign n4042 = n4041 ^ n4040 ;
  assign n4043 = n4022 ^ n3791 ;
  assign n4044 = n4043 ^ n4040 ;
  assign n4045 = ~n4042 & ~n4044 ;
  assign n4046 = n4045 ^ n4040 ;
  assign n4047 = n3810 & n4046 ;
  assign n4048 = n4047 ^ n3809 ;
  assign n3752 = n3751 ^ n3735 ;
  assign n3753 = ~n3734 & ~n3752 ;
  assign n3754 = n3753 ^ n3735 ;
  assign n3736 = n3734 & ~n3735 ;
  assign n3737 = ~n3719 & n3736 ;
  assign n3786 = n3754 ^ n3737 ;
  assign n3738 = n3736 ^ n3734 ;
  assign n3714 = n592 ^ n146 ;
  assign n3715 = n3714 ^ n234 ;
  assign n3746 = n124 & n3715 ;
  assign n3747 = ~n2576 & ~n3746 ;
  assign n3743 = n432 ^ n144 ;
  assign n3744 = n77 & n3743 ;
  assign n3741 = n3722 ^ n288 ;
  assign n3739 = n839 ^ n276 ;
  assign n3740 = n3739 ^ n598 ;
  assign n3742 = n3741 ^ n3740 ;
  assign n3745 = n3744 ^ n3742 ;
  assign n3748 = n3747 ^ n3745 ;
  assign n3749 = ~n3738 & n3748 ;
  assign n3787 = n3786 ^ n3749 ;
  assign n3788 = n2650 & n3787 ;
  assign n3784 = n29 & ~n3763 ;
  assign n3780 = n3749 & n3779 ;
  assign n3778 = ~n3692 & n3821 ;
  assign n3781 = n3780 ^ n3778 ;
  assign n3782 = n3781 ^ n2659 ;
  assign n3777 = n3776 ^ n2658 ;
  assign n3783 = n3782 ^ n3777 ;
  assign n3785 = n3784 ^ n3783 ;
  assign n3789 = n3788 ^ n3785 ;
  assign n3651 = n3650 ^ n3619 ;
  assign n3652 = ~n3622 & n3651 ;
  assign n3653 = n3652 ^ n3650 ;
  assign n3266 = n3265 ^ n3264 ;
  assign n3285 = n3284 ^ n3264 ;
  assign n3286 = n3266 & n3285 ;
  assign n3287 = n3286 ^ n3265 ;
  assign n3090 = n3089 ^ n3072 ;
  assign n3100 = n3090 & ~n3099 ;
  assign n3101 = n3100 ^ n3089 ;
  assign n2929 = n1256 & ~n2928 ;
  assign n2936 = n2929 ^ n694 ;
  assign n2925 = ~n2721 & n2924 ;
  assign n2921 = ~n2722 & n2920 ;
  assign n2926 = n2925 ^ n2921 ;
  assign n2927 = n2926 ^ n694 ;
  assign n2930 = n2929 ^ n2927 ;
  assign n2911 = n1256 & n2910 ;
  assign n2931 = n2930 ^ n2911 ;
  assign n2937 = n2936 ^ n2931 ;
  assign n2938 = n2937 ^ n2926 ;
  assign n2908 = n2720 ^ n780 ;
  assign n2912 = n2911 ^ n2908 ;
  assign n2913 = n2912 ^ n2911 ;
  assign n2939 = n2938 ^ n2913 ;
  assign n2962 = n2939 ^ n2938 ;
  assign n2942 = n2936 ^ n2911 ;
  assign n2943 = n2942 ^ n2931 ;
  assign n2944 = n2943 ^ n2939 ;
  assign n2935 = n2931 ^ n2929 ;
  assign n2940 = n2939 ^ n2935 ;
  assign n2941 = n2940 ^ n2911 ;
  assign n2945 = n2944 ^ n2941 ;
  assign n2946 = n2944 ^ n2940 ;
  assign n2947 = n2946 ^ n2939 ;
  assign n2948 = n2947 ^ n2946 ;
  assign n2949 = ~n2929 & n2948 ;
  assign n2951 = n2949 ^ n2947 ;
  assign n2952 = ~n2945 & ~n2951 ;
  assign n2957 = n2952 ^ n2949 ;
  assign n2953 = n2952 ^ n2946 ;
  assign n2954 = n2940 ^ n2939 ;
  assign n2955 = n2954 ^ n2929 ;
  assign n2956 = ~n2953 & ~n2955 ;
  assign n2958 = n2957 ^ n2956 ;
  assign n2959 = n2958 ^ n2944 ;
  assign n2960 = n2959 ^ n2947 ;
  assign n2963 = n2962 ^ n2960 ;
  assign n2932 = n2931 ^ n2913 ;
  assign n2933 = n2932 ^ n2911 ;
  assign n2934 = n2933 ^ n2926 ;
  assign n2964 = n2963 ^ n2934 ;
  assign n2965 = n2964 ^ n2913 ;
  assign n2899 = n2724 & n2843 ;
  assign n2898 = n2725 & n2840 ;
  assign n2900 = n2899 ^ n2898 ;
  assign n2895 = n709 & ~n2888 ;
  assign n2896 = n2895 ^ n2723 ;
  assign n2897 = n697 & ~n2896 ;
  assign n2901 = n2900 ^ n2897 ;
  assign n2902 = n2901 ^ n2726 ;
  assign n2883 = ~n2854 & n2882 ;
  assign n2884 = ~n707 & n2883 ;
  assign n2885 = ~n2744 & n2884 ;
  assign n2886 = n2885 ^ n2883 ;
  assign n2887 = n2886 ^ n2882 ;
  assign n2903 = n2902 ^ n2887 ;
  assign n2904 = n2903 ^ n2901 ;
  assign n2905 = n707 & ~n2887 ;
  assign n2906 = ~n2904 & n2905 ;
  assign n2907 = n2906 ^ n2903 ;
  assign n2966 = n2965 ^ n2907 ;
  assign n3102 = n3101 ^ n2966 ;
  assign n2822 = n2003 & n2717 ;
  assign n2820 = n2811 & n2819 ;
  assign n2821 = ~n2805 & n2820 ;
  assign n2823 = n2822 ^ n2821 ;
  assign n2824 = n2823 ^ n2819 ;
  assign n2825 = n2824 ^ n2718 ;
  assign n2816 = n999 & ~n2805 ;
  assign n2817 = n2816 ^ n2718 ;
  assign n2818 = n2811 & ~n2817 ;
  assign n2826 = n2825 ^ n2818 ;
  assign n2806 = n2805 ^ n2719 ;
  assign n2807 = n2800 & ~n2806 ;
  assign n2827 = n2826 ^ n2807 ;
  assign n3103 = n3102 ^ n2827 ;
  assign n3288 = n3287 ^ n3103 ;
  assign n2775 = ~n1357 & ~n2671 ;
  assign n2776 = n2775 ^ n2665 ;
  assign n2777 = ~n2685 & ~n2776 ;
  assign n2767 = n2766 ^ n2764 ;
  assign n2768 = n2767 ^ n2685 ;
  assign n2769 = ~n2690 & ~n2768 ;
  assign n2686 = n2685 ^ n1357 ;
  assign n2687 = n2686 ^ n2671 ;
  assign n2770 = n2769 ^ n2687 ;
  assign n2778 = n2777 ^ n2770 ;
  assign n2672 = ~n2643 & n2671 ;
  assign n2779 = n2778 ^ n2672 ;
  assign n2790 = ~n1357 & ~n2787 ;
  assign n2791 = n2790 ^ n1406 ;
  assign n2792 = ~n2784 & ~n2791 ;
  assign n2788 = n2787 ^ n1406 ;
  assign n2793 = n2792 ^ n2788 ;
  assign n2794 = ~n2667 & n2793 ;
  assign n2795 = ~n2779 & n2794 ;
  assign n2796 = n2795 ^ n2779 ;
  assign n3289 = n3288 ^ n2796 ;
  assign n3774 = n3653 ^ n3289 ;
  assign n3790 = n3789 ^ n3774 ;
  assign n4084 = n4048 ^ n3790 ;
  assign n4068 = n154 & ~n374 ;
  assign n4060 = n116 & n144 ;
  assign n4061 = n4060 ^ n379 ;
  assign n4062 = n4061 ^ n276 ;
  assign n4063 = n4062 ^ n167 ;
  assign n4059 = n3687 ^ n2393 ;
  assign n4064 = n4063 ^ n4059 ;
  assign n4056 = n512 ^ n181 ;
  assign n4055 = n577 ^ n284 ;
  assign n4057 = n4056 ^ n4055 ;
  assign n4058 = n4057 ^ n1001 ;
  assign n4065 = n4064 ^ n4058 ;
  assign n4054 = n93 & n2627 ;
  assign n4066 = n4065 ^ n4054 ;
  assign n4067 = n4066 ^ n849 ;
  assign n4069 = n4068 ^ n4067 ;
  assign n4076 = n607 ^ n169 ;
  assign n4077 = n4076 ^ n341 ;
  assign n4078 = n4077 ^ n793 ;
  assign n4079 = n4078 ^ n2696 ;
  assign n4080 = n4079 ^ n672 ;
  assign n4072 = n817 ^ n434 ;
  assign n4073 = n4072 ^ n495 ;
  assign n4074 = n4073 ^ n2324 ;
  assign n4071 = n480 ^ n268 ;
  assign n4075 = n4074 ^ n4071 ;
  assign n4081 = n4080 ^ n4075 ;
  assign n4070 = n626 ^ n585 ;
  assign n4082 = n4081 ^ n4070 ;
  assign n4083 = n4069 & n4082 ;
  assign n4085 = n4084 ^ n4083 ;
  assign n4093 = n1044 ^ n163 ;
  assign n4094 = n4093 ^ n477 ;
  assign n4095 = n4094 ^ n786 ;
  assign n4099 = n447 ^ n170 ;
  assign n4100 = n4099 ^ n394 ;
  assign n4101 = n4100 ^ n2468 ;
  assign n4102 = n4101 ^ n2581 ;
  assign n4097 = n354 ^ n120 ;
  assign n4098 = n4097 ^ n2496 ;
  assign n4103 = n4102 ^ n4098 ;
  assign n4096 = n116 & n205 ;
  assign n4104 = n4103 ^ n4096 ;
  assign n4105 = n4095 & ~n4104 ;
  assign n4087 = n1032 ^ n489 ;
  assign n4088 = n4087 ^ n231 ;
  assign n4089 = n4088 ^ n2295 ;
  assign n4090 = n4089 ^ n2395 ;
  assign n4086 = n791 ^ n243 ;
  assign n4091 = n4090 ^ n4086 ;
  assign n4092 = n4091 ^ n251 ;
  assign n4106 = n4105 ^ n4092 ;
  assign n4107 = n4039 ^ n4037 ;
  assign n4137 = n795 ^ n444 ;
  assign n4138 = n4137 ^ n605 ;
  assign n4131 = n211 ^ n190 ;
  assign n4132 = n4131 ^ n391 ;
  assign n4133 = n399 ^ n117 ;
  assign n4134 = n4133 ^ n4131 ;
  assign n4135 = ~n4132 & ~n4134 ;
  assign n4127 = n845 ^ n82 ;
  assign n295 = n294 ^ n291 ;
  assign n297 = n296 ^ n295 ;
  assign n4128 = n4127 ^ n297 ;
  assign n4129 = n4128 ^ n395 ;
  assign n4130 = n4129 ^ n1193 ;
  assign n4136 = n4135 ^ n4130 ;
  assign n4139 = n4138 ^ n4136 ;
  assign n4121 = n385 ^ n362 ;
  assign n4122 = n4121 ^ n2700 ;
  assign n4123 = n4122 ^ n1033 ;
  assign n4119 = ~n254 & ~n293 ;
  assign n4120 = n4119 ^ n859 ;
  assign n4124 = n4123 ^ n4120 ;
  assign n4125 = n4124 ^ n2508 ;
  assign n4116 = n629 ^ n285 ;
  assign n4113 = n383 ^ n161 ;
  assign n4114 = n4113 ^ n304 ;
  assign n4112 = n398 ^ n170 ;
  assign n4115 = n4114 ^ n4112 ;
  assign n4117 = n4116 ^ n4115 ;
  assign n4110 = n646 ^ n350 ;
  assign n4108 = n449 ^ n232 ;
  assign n4109 = n4108 ^ n831 ;
  assign n4111 = n4110 ^ n4109 ;
  assign n4118 = n4117 ^ n4111 ;
  assign n4126 = n4125 ^ n4118 ;
  assign n4140 = n4139 ^ n4126 ;
  assign n4141 = n4022 & n4106 ;
  assign n4142 = n4140 & ~n4141 ;
  assign n4143 = n4141 ^ n4140 ;
  assign n4144 = n4143 ^ n4022 ;
  assign n4145 = n4144 ^ n4142 ;
  assign n4146 = n4145 ^ n4022 ;
  assign n4147 = n4039 ^ n4022 ;
  assign n4148 = n4147 ^ n4022 ;
  assign n4149 = ~n4146 & ~n4148 ;
  assign n4150 = n4149 ^ n4022 ;
  assign n4151 = n4107 & n4150 ;
  assign n4152 = n4151 ^ n4022 ;
  assign n4153 = n3810 & ~n4152 ;
  assign n4154 = n4140 ^ n3810 ;
  assign n4162 = n3810 & n4154 ;
  assign n4155 = n4154 ^ n4141 ;
  assign n4164 = n4162 ^ n4155 ;
  assign n4165 = ~n4039 & ~n4164 ;
  assign n4173 = n4165 ^ n4162 ;
  assign n4166 = n4165 ^ n4141 ;
  assign n4167 = n4037 ^ n3810 ;
  assign n4168 = n4167 ^ n4154 ;
  assign n4169 = n4168 ^ n4039 ;
  assign n4170 = n4169 ^ n4154 ;
  assign n4171 = n4170 ^ n3810 ;
  assign n4172 = ~n4166 & ~n4171 ;
  assign n4174 = n4173 ^ n4172 ;
  assign n4175 = n4174 ^ n3810 ;
  assign n4176 = n4175 ^ n4155 ;
  assign n4177 = ~n4153 & n4176 ;
  assign n4182 = n4177 ^ n4153 ;
  assign n4178 = ~n4106 & n4177 ;
  assign n4179 = ~n4022 & n4178 ;
  assign n4183 = n4182 ^ n4179 ;
  assign n4180 = n4037 & ~n4039 ;
  assign n4181 = n4179 & n4180 ;
  assign n4184 = n4183 ^ n4181 ;
  assign n4185 = n4142 & n4184 ;
  assign n4186 = ~n4107 & n4185 ;
  assign n4187 = n4106 & n4186 ;
  assign n4188 = n4187 ^ n4185 ;
  assign n4189 = n4188 ^ n4184 ;
  assign n4190 = n4189 ^ n4083 ;
  assign n4191 = ~n4085 & ~n4190 ;
  assign n4192 = n4191 ^ n4085 ;
  assign n4049 = n4048 ^ n3789 ;
  assign n4050 = ~n3790 & ~n4049 ;
  assign n4051 = n4050 ^ n3789 ;
  assign n3755 = ~n3748 & ~n3754 ;
  assign n3750 = ~n3737 & n3749 ;
  assign n3756 = n3755 ^ n3750 ;
  assign n3757 = n28 & ~n3756 ;
  assign n3707 = n845 ^ n274 ;
  assign n3705 = n278 ^ n94 ;
  assign n3706 = n3705 ^ n642 ;
  assign n3708 = n3707 ^ n3706 ;
  assign n3703 = n787 ^ n531 ;
  assign n3704 = ~n117 & n3703 ;
  assign n3709 = n3708 ^ n3704 ;
  assign n3710 = n429 ^ n218 ;
  assign n3711 = n3710 ^ n548 ;
  assign n3712 = ~n3709 & ~n3711 ;
  assign n3713 = n1213 & n3712 ;
  assign n3716 = n91 & n3715 ;
  assign n3717 = n3713 & n3716 ;
  assign n3718 = n3717 ^ n3713 ;
  assign n3758 = n3757 ^ n3718 ;
  assign n3771 = ~n4664 ^ n3758 ;
  assign n3759 = n3758 ^ n3749 ;
  assign n3760 = n3759 ^ n3758 ;
  assign n3761 = n3760 ^ x2 ;
  assign n3762 = n3761 ^ n3760 ;
  assign n3766 = n3762 & ~n3763 ;
  assign n3767 = n3766 ^ n3760 ;
  assign n3768 = ~x1 & n3767 ;
  assign n3769 = n3768 ^ n3759 ;
  assign n3770 = ~x0 & ~n3769 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3694 = n3692 ^ n1406 ;
  assign n3693 = n3692 ^ n1357 ;
  assign n3695 = n3694 ^ n3693 ;
  assign n3696 = n3693 ^ n2766 ;
  assign n3697 = n3696 ^ n3693 ;
  assign n3698 = n3695 & ~n3697 ;
  assign n3699 = n3698 ^ n3693 ;
  assign n3700 = ~n2667 & ~n3699 ;
  assign n3661 = n2690 ^ n1357 ;
  assign n3662 = n3661 ^ n3422 ;
  assign n3659 = n3380 ^ n2671 ;
  assign n3660 = ~n2787 & n3659 ;
  assign n3663 = n3662 ^ n3660 ;
  assign n3668 = ~n2643 & ~n3380 ;
  assign n3669 = n3388 & n3668 ;
  assign n3670 = n3669 ^ n3388 ;
  assign n3671 = n3670 ^ n3389 ;
  assign n3672 = ~n3663 & ~n3671 ;
  assign n3701 = n3700 ^ n3672 ;
  assign n3656 = n3653 ^ n2796 ;
  assign n3657 = ~n3289 & ~n3656 ;
  assign n3375 = n2717 & ~n2811 ;
  assign n3366 = n2811 & n3362 ;
  assign n3372 = ~n999 & n2811 ;
  assign n3373 = ~n3366 & ~n3372 ;
  assign n3367 = n3366 ^ n2811 ;
  assign n3368 = ~n995 & ~n3367 ;
  assign n3365 = n2003 & ~n2685 ;
  assign n3369 = n3368 ^ n3365 ;
  assign n3370 = n3369 ^ n2811 ;
  assign n3363 = n3362 ^ n2718 ;
  assign n3364 = n2800 & ~n3363 ;
  assign n3371 = n3370 ^ n3364 ;
  assign n3374 = n3373 ^ n3371 ;
  assign n3376 = n3375 ^ n3374 ;
  assign n3322 = n1256 & ~n2909 ;
  assign n3329 = n3322 ^ n694 ;
  assign n3319 = ~n2720 & n2924 ;
  assign n3318 = ~n2721 & n2920 ;
  assign n3320 = n3319 ^ n3318 ;
  assign n3321 = n3320 ^ n694 ;
  assign n3323 = n3322 ^ n3321 ;
  assign n3315 = n1256 & n3314 ;
  assign n3324 = n3323 ^ n3315 ;
  assign n3330 = n3329 ^ n3324 ;
  assign n3331 = n3330 ^ n3320 ;
  assign n3313 = n2719 ^ n780 ;
  assign n3316 = n3315 ^ n3313 ;
  assign n3317 = n3316 ^ n3315 ;
  assign n3332 = n3331 ^ n3317 ;
  assign n3355 = n3332 ^ n3331 ;
  assign n3335 = n3329 ^ n3315 ;
  assign n3336 = n3335 ^ n3324 ;
  assign n3337 = n3336 ^ n3332 ;
  assign n3328 = n3324 ^ n3322 ;
  assign n3333 = n3332 ^ n3328 ;
  assign n3334 = n3333 ^ n3315 ;
  assign n3338 = n3337 ^ n3334 ;
  assign n3339 = n3337 ^ n3333 ;
  assign n3340 = n3339 ^ n3332 ;
  assign n3341 = n3340 ^ n3339 ;
  assign n3342 = ~n3322 & ~n3341 ;
  assign n3344 = n3342 ^ n3340 ;
  assign n3345 = ~n3338 & n3344 ;
  assign n3350 = n3345 ^ n3342 ;
  assign n3346 = n3345 ^ n3339 ;
  assign n3347 = n3333 ^ n3332 ;
  assign n3348 = n3347 ^ n3322 ;
  assign n3349 = ~n3346 & ~n3348 ;
  assign n3351 = n3350 ^ n3349 ;
  assign n3352 = n3351 ^ n3337 ;
  assign n3353 = n3352 ^ n3340 ;
  assign n3356 = n3355 ^ n3353 ;
  assign n3325 = n3324 ^ n3317 ;
  assign n3326 = n3325 ^ n3315 ;
  assign n3327 = n3326 ^ n3320 ;
  assign n3357 = n3356 ^ n3327 ;
  assign n3358 = n3357 ^ n3317 ;
  assign n3309 = n2726 ^ n2725 ;
  assign n3307 = n2901 ^ n2887 ;
  assign n3308 = ~n2902 & n3307 ;
  assign n3310 = n3309 ^ n3308 ;
  assign n3311 = ~n707 & ~n3310 ;
  assign n3304 = ~n2723 & n2843 ;
  assign n3303 = n2724 & n2840 ;
  assign n3305 = n3304 ^ n3303 ;
  assign n3298 = n2722 ^ n709 ;
  assign n3299 = n3298 ^ n2722 ;
  assign n3300 = ~n2967 & n3299 ;
  assign n3301 = n3300 ^ n2722 ;
  assign n3302 = n697 & ~n3301 ;
  assign n3306 = n3305 ^ n3302 ;
  assign n3312 = n3311 ^ n3306 ;
  assign n3359 = n3358 ^ n3312 ;
  assign n3293 = n3101 ^ n2965 ;
  assign n3294 = ~n2966 & ~n3293 ;
  assign n3295 = n3294 ^ n3101 ;
  assign n3360 = n3359 ^ n3295 ;
  assign n3290 = n3287 ^ n2827 ;
  assign n3291 = ~n3103 & ~n3290 ;
  assign n3292 = n3291 ^ n3287 ;
  assign n3361 = n3360 ^ n3292 ;
  assign n3377 = n3376 ^ n3361 ;
  assign n3654 = n3653 ^ n3377 ;
  assign n3658 = n3657 ^ n3654 ;
  assign n3702 = n3701 ^ n3658 ;
  assign n3773 = n3772 ^ n3702 ;
  assign n4052 = n4051 ^ n3773 ;
  assign n299 = n298 ^ n297 ;
  assign n287 = n286 ^ n285 ;
  assign n290 = n289 ^ n287 ;
  assign n300 = n299 ^ n290 ;
  assign n282 = n281 ^ n269 ;
  assign n301 = n300 ^ n282 ;
  assign n302 = n259 & ~n301 ;
  assign n375 = n374 ^ n302 ;
  assign n376 = ~n223 & ~n375 ;
  assign n4053 = n4052 ^ n376 ;
  assign n4193 = n4192 ^ n4053 ;
  assign n4360 = ~n4084 & ~n4192 ;
  assign n4361 = n4360 ^ n4192 ;
  assign n4357 = n376 & n4052 ;
  assign n4358 = n4357 ^ n4053 ;
  assign n4337 = ~n3718 & ~n3755 ;
  assign n4336 = n3718 & ~n3750 ;
  assign n4338 = n4337 ^ n4336 ;
  assign n4339 = n28 & ~n4338 ;
  assign n4198 = n447 ^ n345 ;
  assign n4199 = n4198 ^ n273 ;
  assign n4331 = n4199 ^ n1495 ;
  assign n4328 = n211 ^ n105 ;
  assign n4329 = n4328 ^ n137 ;
  assign n4330 = n92 & n4329 ;
  assign n4332 = n4331 ^ n4330 ;
  assign n4327 = n2429 ^ n95 ;
  assign n4333 = n4332 ^ n4327 ;
  assign n4321 = n2297 ^ n318 ;
  assign n4322 = n4321 ^ n793 ;
  assign n4323 = n4322 ^ n843 ;
  assign n4324 = n4323 ^ n580 ;
  assign n4319 = n813 ^ n594 ;
  assign n4320 = ~n125 & n4319 ;
  assign n4325 = n4324 ^ n4320 ;
  assign n4326 = n790 & ~n4325 ;
  assign n4334 = n4333 ^ n4326 ;
  assign n4335 = n2494 & ~n4334 ;
  assign n4340 = n4339 ^ n4335 ;
  assign n4352 = ~n4664 ^ n4340 ;
  assign n4347 = x2 & n3749 ;
  assign n4348 = n4347 ^ n3718 ;
  assign n4349 = ~x1 & ~n4348 ;
  assign n4341 = n4340 ^ n3718 ;
  assign n4350 = n4349 ^ n4341 ;
  assign n4351 = ~x0 & n4350 ;
  assign n4353 = n4352 ^ n4351 ;
  assign n4313 = n3692 ^ n2688 ;
  assign n4309 = n3752 ^ n3692 ;
  assign n4310 = n4309 ^ n3786 ;
  assign n4308 = ~n1357 & n3800 ;
  assign n4311 = n4310 ^ n4308 ;
  assign n4312 = ~n2671 & ~n4311 ;
  assign n4314 = n4313 ^ n4312 ;
  assign n4301 = n3763 ^ n1406 ;
  assign n4302 = n3800 ^ n2667 ;
  assign n4303 = n4302 ^ n2667 ;
  assign n4305 = ~n2671 & n4303 ;
  assign n4306 = n4305 ^ n2667 ;
  assign n4307 = ~n4301 & ~n4306 ;
  assign n4315 = n4314 ^ n4307 ;
  assign n4299 = n3800 ^ n2787 ;
  assign n4300 = n3388 & ~n4299 ;
  assign n4316 = n4315 ^ n4300 ;
  assign n4233 = n2643 ^ n999 ;
  assign n4234 = n2003 & ~n4233 ;
  assign n4235 = n2783 & n4234 ;
  assign n4230 = ~n2685 & ~n2811 ;
  assign n4229 = n2717 & n2800 ;
  assign n4231 = n4230 ^ n4229 ;
  assign n4232 = n4231 ^ n995 ;
  assign n4236 = n4235 ^ n4232 ;
  assign n4284 = n4236 ^ n4235 ;
  assign n4285 = n2003 & ~n3623 ;
  assign n4286 = n4284 & n4285 ;
  assign n4263 = n708 ^ n694 ;
  assign n4268 = n2722 ^ n707 ;
  assign n4269 = n4268 ^ n694 ;
  assign n4270 = n4269 ^ n2722 ;
  assign n4272 = ~n2723 & ~n4270 ;
  assign n4273 = n4272 ^ n2722 ;
  assign n4274 = n4263 & ~n4273 ;
  assign n4264 = n709 & ~n2972 ;
  assign n4265 = n4264 ^ n2721 ;
  assign n4266 = n4265 ^ n2722 ;
  assign n4275 = n4274 ^ n4266 ;
  assign n4276 = ~n697 & n4275 ;
  assign n4277 = n4276 ^ n4265 ;
  assign n4255 = n3306 ^ n2725 ;
  assign n4258 = n3310 & ~n4255 ;
  assign n4259 = n4258 ^ n2725 ;
  assign n4260 = ~n707 & n4259 ;
  assign n4261 = n4260 ^ n2724 ;
  assign n4262 = ~n707 & ~n4261 ;
  assign n4278 = n4277 ^ n4262 ;
  assign n4244 = n694 & n1256 ;
  assign n4245 = ~n2803 & n4244 ;
  assign n4279 = n4278 ^ n4245 ;
  assign n4252 = n1256 & ~n2801 ;
  assign n4253 = n2718 ^ n780 ;
  assign n4254 = n4252 & ~n4253 ;
  assign n4280 = n4279 ^ n4254 ;
  assign n4241 = n2719 & n2924 ;
  assign n4240 = ~n2720 & n2920 ;
  assign n4242 = n4241 ^ n4240 ;
  assign n4243 = n4242 ^ n694 ;
  assign n4246 = n4245 ^ n4242 ;
  assign n4247 = n1256 & n2804 ;
  assign n4248 = n4247 ^ n4245 ;
  assign n4249 = ~n4246 & n4248 ;
  assign n4250 = n4249 ^ n4245 ;
  assign n4251 = ~n4243 & ~n4250 ;
  assign n4281 = n4280 ^ n4251 ;
  assign n4237 = n3312 ^ n3295 ;
  assign n4238 = n3359 & ~n4237 ;
  assign n4239 = n4238 ^ n3358 ;
  assign n4282 = n4281 ^ n4239 ;
  assign n4283 = n4282 ^ n4236 ;
  assign n4287 = n4286 ^ n4283 ;
  assign n4288 = n4287 ^ n4282 ;
  assign n4289 = n4231 ^ n2003 ;
  assign n4290 = n4289 ^ n4231 ;
  assign n4291 = n4231 ^ n3624 ;
  assign n4292 = n4291 ^ n4231 ;
  assign n4293 = n4290 & ~n4292 ;
  assign n4294 = n4293 ^ n4231 ;
  assign n4295 = ~n995 & n4294 ;
  assign n4296 = ~n4288 & n4295 ;
  assign n4297 = n4296 ^ n4287 ;
  assign n4226 = n3376 ^ n3292 ;
  assign n4227 = n3361 & ~n4226 ;
  assign n4228 = n4227 ^ n3376 ;
  assign n4298 = n4297 ^ n4228 ;
  assign n4317 = n4316 ^ n4298 ;
  assign n4223 = n3701 ^ n3377 ;
  assign n4224 = ~n3658 & ~n4223 ;
  assign n4225 = n4224 ^ n3377 ;
  assign n4318 = n4317 ^ n4225 ;
  assign n4354 = n4353 ^ n4318 ;
  assign n4220 = n4051 ^ n3772 ;
  assign n4221 = ~n3773 & n4220 ;
  assign n4222 = n4221 ^ n4051 ;
  assign n4355 = n4354 ^ n4222 ;
  assign n4211 = n1044 ^ n256 ;
  assign n4212 = n4211 ^ n553 ;
  assign n4210 = n845 ^ n645 ;
  assign n4213 = n4212 ^ n4210 ;
  assign n4214 = n4213 ^ n268 ;
  assign n4208 = n4087 ^ n481 ;
  assign n4207 = ~n117 & n2691 ;
  assign n4209 = n4208 ^ n4207 ;
  assign n4215 = n4214 ^ n4209 ;
  assign n4216 = n4215 ^ n2375 ;
  assign n4205 = n843 ^ n252 ;
  assign n4204 = n410 ^ n385 ;
  assign n4206 = n4205 ^ n4204 ;
  assign n4217 = n4216 ^ n4206 ;
  assign n4218 = n4217 ^ n4066 ;
  assign n4200 = n4199 ^ n3726 ;
  assign n4201 = n4200 ^ n4071 ;
  assign n4202 = n2358 & ~n4201 ;
  assign n4197 = n417 ^ n303 ;
  assign n4203 = n4202 ^ n4197 ;
  assign n4219 = n4218 ^ n4203 ;
  assign n4356 = n4355 ^ n4219 ;
  assign n4359 = n4358 ^ n4356 ;
  assign n4362 = n4361 ^ n4359 ;
  assign n4194 = x23 ^ x22 ;
  assign n4195 = n4194 ^ n4053 ;
  assign n4196 = n4193 & ~n4195 ;
  assign n4363 = n4362 ^ n4196 ;
  assign n4524 = n335 ^ n161 ;
  assign n4525 = n4524 ^ n831 ;
  assign n4522 = n549 ^ n260 ;
  assign n4523 = n4522 ^ n481 ;
  assign n4526 = n4525 ^ n4523 ;
  assign n4517 = n434 ^ n170 ;
  assign n4518 = n4517 ^ n858 ;
  assign n4519 = n4518 ^ n512 ;
  assign n4520 = n4519 ^ n298 ;
  assign n4516 = n575 ^ n192 ;
  assign n4521 = n4520 ^ n4516 ;
  assign n4527 = n4526 ^ n4521 ;
  assign n4528 = n4527 ^ n821 ;
  assign n4529 = n4528 ^ n4092 ;
  assign n4512 = n4353 ^ n4222 ;
  assign n4513 = n4354 & n4512 ;
  assign n4514 = n4513 ^ n4353 ;
  assign n4507 = n4316 ^ n4225 ;
  assign n4508 = n4317 & ~n4507 ;
  assign n4509 = n4508 ^ n4316 ;
  assign n4503 = n4282 ^ n4228 ;
  assign n4504 = n4297 & n4503 ;
  assign n4505 = n4504 ^ n4282 ;
  assign n4495 = n2717 ^ n780 ;
  assign n4496 = n1256 & ~n2805 ;
  assign n4497 = ~n4495 & n4496 ;
  assign n4483 = n2718 & n2924 ;
  assign n4482 = n2719 & n2920 ;
  assign n4484 = n4483 ^ n4482 ;
  assign n4485 = n4484 ^ n694 ;
  assign n4490 = n3409 ^ n3408 ;
  assign n4491 = ~n4485 & ~n4490 ;
  assign n4492 = n4491 ^ n3408 ;
  assign n4493 = n1256 & ~n4492 ;
  assign n4494 = n4493 ^ n4485 ;
  assign n4498 = n4497 ^ n4494 ;
  assign n4479 = ~n2721 & n2843 ;
  assign n4478 = ~n2722 & n2840 ;
  assign n4480 = n4479 ^ n4478 ;
  assign n4475 = n709 & ~n2928 ;
  assign n4476 = n4475 ^ n2720 ;
  assign n4477 = n697 & ~n4476 ;
  assign n4481 = n4480 ^ n4477 ;
  assign n4499 = n4498 ^ n4481 ;
  assign n4468 = n4277 ^ n4260 ;
  assign n4469 = n4277 ^ n2724 ;
  assign n4470 = ~n4468 & n4469 ;
  assign n4471 = n4470 ^ n3179 ;
  assign n4472 = ~n707 & n4471 ;
  assign n4500 = n4499 ^ n4472 ;
  assign n4465 = n4278 ^ n4239 ;
  assign n4466 = n4281 & ~n4465 ;
  assign n4467 = n4466 ^ n4278 ;
  assign n4501 = n4500 ^ n4467 ;
  assign n4443 = n999 & ~n2643 ;
  assign n4459 = n2643 ^ n995 ;
  assign n4460 = ~n2811 & n4459 ;
  assign n4463 = n4443 & n4460 ;
  assign n4453 = n995 & ~n2643 ;
  assign n4454 = n999 & n2809 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4452 = n2685 & n2800 ;
  assign n4456 = n4455 ^ n4452 ;
  assign n4457 = n4456 ^ n2809 ;
  assign n4444 = n2787 ^ n995 ;
  assign n4447 = n4444 ^ n2784 ;
  assign n4448 = n4447 ^ n4444 ;
  assign n4449 = ~n1000 & n4448 ;
  assign n4450 = n4449 ^ n4444 ;
  assign n4451 = n2003 & ~n4450 ;
  assign n4458 = n4457 ^ n4451 ;
  assign n4461 = n4460 ^ n4458 ;
  assign n4464 = n4463 ^ n4461 ;
  assign n4502 = n4501 ^ n4464 ;
  assign n4506 = n4505 ^ n4502 ;
  assign n4510 = n4509 ^ n4506 ;
  assign n4433 = n4335 & n4338 ;
  assign n4434 = n4433 ^ n4338 ;
  assign n4435 = n4434 ^ n4337 ;
  assign n4436 = n28 & ~n4435 ;
  assign n4437 = n4436 ^ n3802 ;
  assign n4432 = n4335 ^ n1473 ;
  assign n4438 = n4437 ^ n4432 ;
  assign n4429 = x2 & ~n3718 ;
  assign n4424 = n4335 ^ x22 ;
  assign n4430 = n4429 ^ n4424 ;
  assign n4431 = ~x1 & n4430 ;
  assign n4439 = n4438 ^ n4431 ;
  assign n4440 = ~x0 & ~n4439 ;
  assign n4441 = n4440 ^ n4437 ;
  assign n4405 = n2668 ^ n2667 ;
  assign n4406 = n3756 ^ n3754 ;
  assign n4407 = n4406 ^ n3787 ;
  assign n4408 = ~n4405 & n4407 ;
  assign n4396 = ~n2670 & ~n3763 ;
  assign n4395 = n3422 & n3692 ;
  assign n4397 = n4396 ^ n4395 ;
  assign n4389 = n4301 ^ n3763 ;
  assign n4390 = n1357 & n3692 ;
  assign n4391 = n4390 ^ n3763 ;
  assign n4392 = ~n4389 & ~n4391 ;
  assign n4393 = n4392 ^ n3763 ;
  assign n4394 = ~n2664 & ~n4393 ;
  assign n4398 = n4397 ^ n4394 ;
  assign n4399 = n4398 ^ n1357 ;
  assign n4400 = n4399 ^ n4398 ;
  assign n4401 = n3756 ^ n3737 ;
  assign n4402 = ~n2667 & n4401 ;
  assign n4403 = n4400 & n4402 ;
  assign n4404 = n4403 ^ n4399 ;
  assign n4409 = n4408 ^ n4404 ;
  assign n4412 = ~n3786 & ~n4398 ;
  assign n4413 = n4412 ^ n2667 ;
  assign n4414 = n1357 & ~n4413 ;
  assign n4415 = n4414 ^ n2667 ;
  assign n4416 = ~n4409 & ~n4415 ;
  assign n4418 = n3787 ^ n1406 ;
  assign n4419 = n4418 ^ n3787 ;
  assign n4420 = ~n3786 & ~n4419 ;
  assign n4421 = n4420 ^ n3787 ;
  assign n4422 = n4416 & ~n4421 ;
  assign n4423 = n4422 ^ n4409 ;
  assign n4442 = n4441 ^ n4423 ;
  assign n4511 = n4510 ^ n4442 ;
  assign n4515 = n4514 ^ n4511 ;
  assign n4530 = n4529 ^ n4515 ;
  assign n4387 = n317 ^ n188 ;
  assign n4388 = ~n125 & n4387 ;
  assign n4531 = n4530 ^ n4388 ;
  assign n4367 = n4191 ^ n4189 ;
  assign n4375 = n4053 & n4361 ;
  assign n4376 = ~n4367 & n4375 ;
  assign n4382 = n4376 ^ n4357 ;
  assign n4381 = n4375 ^ n4053 ;
  assign n4383 = n4382 ^ n4381 ;
  assign n4384 = n4383 ^ n4219 ;
  assign n4385 = n4356 & ~n4384 ;
  assign n4386 = n4385 ^ n4355 ;
  assign n4532 = n4531 ^ n4386 ;
  assign n4377 = n4356 & n4376 ;
  assign n4368 = ~n4357 & n4367 ;
  assign n4364 = ~n4053 & ~n4356 ;
  assign n4373 = n4368 ^ n4364 ;
  assign n4374 = n4360 & ~n4373 ;
  assign n4378 = n4377 ^ n4374 ;
  assign n4533 = n4532 ^ n4378 ;
  assign n4369 = ~n4360 & n4368 ;
  assign n4370 = n4356 & n4369 ;
  assign n4371 = n4358 & n4370 ;
  assign n4365 = n4364 ^ n4358 ;
  assign n4366 = ~n4361 & ~n4365 ;
  assign n4372 = n4371 ^ n4366 ;
  assign n4379 = n4378 ^ n4372 ;
  assign n4380 = n4194 & ~n4379 ;
  assign n4534 = n4533 ^ n4380 ;
  assign n4535 = n4378 & ~n4532 ;
  assign n4536 = ~n4194 & ~n4535 ;
  assign n4537 = n4515 ^ n4386 ;
  assign n4538 = n4531 & n4537 ;
  assign n4539 = n4538 ^ n4515 ;
  assign n4689 = n4372 ^ n4194 ;
  assign n4686 = n4539 ^ n4532 ;
  assign n4687 = n4686 ^ n4372 ;
  assign n4688 = n4687 ^ n4539 ;
  assign n4690 = n4689 ^ n4688 ;
  assign n4691 = n4690 ^ n4539 ;
  assign n4692 = n4691 ^ n4690 ;
  assign n4694 = n4689 ^ n4372 ;
  assign n4695 = n4692 & ~n4694 ;
  assign n4696 = n4695 ^ n4690 ;
  assign n4697 = n4695 ^ n4694 ;
  assign n4698 = n4379 & ~n4697 ;
  assign n4699 = n4698 ^ n4378 ;
  assign n4700 = n4699 ^ n4379 ;
  assign n4701 = n4696 & ~n4700 ;
  assign n4702 = n4701 ^ n4698 ;
  assign n4703 = n4702 ^ n4686 ;
  assign n4704 = n4703 ^ n4372 ;
  assign n4680 = n4514 ^ n4506 ;
  assign n4681 = n4510 ^ n4441 ;
  assign n4682 = n4681 ^ n4423 ;
  assign n4683 = ~n4680 & n4682 ;
  assign n4672 = n394 ^ n256 ;
  assign n4673 = n4672 ^ n179 ;
  assign n4674 = n4673 ^ n1071 ;
  assign n4670 = n4204 ^ n2431 ;
  assign n4669 = n267 ^ n94 ;
  assign n4671 = n4670 ^ n4669 ;
  assign n4675 = n4674 ^ n4671 ;
  assign n4676 = n4675 ^ n2280 ;
  assign n4677 = n4676 ^ n1527 ;
  assign n4667 = n4111 ^ n422 ;
  assign n4668 = ~n875 & n4667 ;
  assign n4678 = n4677 ^ n4668 ;
  assign n4657 = n4656 ^ ~n3821 ;
  assign n4660 = ~n4336 & ~n4657 ;
  assign n4661 = n4660 ^ ~n3821 ;
  assign n4662 = ~n4335 & ~n4661 ;
  assign n4665 = n4664 ^ n4662 ;
  assign n4651 = n4505 ^ n4464 ;
  assign n4652 = n4502 & n4651 ;
  assign n4653 = n4652 ^ n4505 ;
  assign n4644 = n4498 ^ n4467 ;
  assign n4645 = n4500 & ~n4644 ;
  assign n4646 = n4645 ^ n4498 ;
  assign n4641 = ~n2720 & n2843 ;
  assign n4640 = ~n2721 & n2840 ;
  assign n4642 = n4641 ^ n4640 ;
  assign n4635 = n2719 ^ n709 ;
  assign n4636 = n4635 ^ n2719 ;
  assign n4637 = ~n2909 & n4636 ;
  assign n4638 = n4637 ^ n2719 ;
  assign n4639 = n697 & n4638 ;
  assign n4643 = n4642 ^ n4639 ;
  assign n4647 = n4646 ^ n4643 ;
  assign n4628 = n4481 ^ n2723 ;
  assign n4629 = ~n4471 & n4628 ;
  assign n4630 = n4629 ^ n2723 ;
  assign n4631 = n4630 ^ n2722 ;
  assign n4632 = ~n707 & ~n4631 ;
  assign n4648 = n4647 ^ n4632 ;
  assign n4610 = n2685 ^ n780 ;
  assign n4611 = n1256 & ~n3362 ;
  assign n4612 = ~n4610 & n4611 ;
  assign n4607 = n2717 & n2924 ;
  assign n4606 = n2718 & n2920 ;
  assign n4608 = n4607 ^ n4606 ;
  assign n4609 = n4608 ^ n694 ;
  assign n4613 = n4612 ^ n4609 ;
  assign n4614 = n4613 ^ n4612 ;
  assign n4615 = n2783 ^ n2756 ;
  assign n4616 = n1256 & ~n4615 ;
  assign n4617 = n4614 & n4616 ;
  assign n4618 = n4617 ^ n4613 ;
  assign n4619 = ~n694 & ~n4618 ;
  assign n4620 = n4608 ^ n1256 ;
  assign n4621 = n4620 ^ n4608 ;
  assign n4622 = n4608 ^ n2782 ;
  assign n4623 = n4622 ^ n4608 ;
  assign n4624 = n4621 & n4623 ;
  assign n4625 = n4624 ^ n4608 ;
  assign n4626 = n4619 & n4625 ;
  assign n4627 = n4626 ^ n4618 ;
  assign n4649 = n4648 ^ n4627 ;
  assign n4577 = ~n995 & n2787 ;
  assign n4592 = n4453 ^ n4444 ;
  assign n4593 = n4444 ^ n1357 ;
  assign n4594 = n4593 ^ n4444 ;
  assign n4595 = ~n4592 & ~n4594 ;
  assign n4596 = n4595 ^ n4444 ;
  assign n4597 = ~n2003 & n4596 ;
  assign n4586 = n2787 ^ n1357 ;
  assign n4587 = n4586 ^ n2787 ;
  assign n4588 = n4023 & n4587 ;
  assign n4589 = n4588 ^ n2787 ;
  assign n4590 = n2799 & ~n4589 ;
  assign n4599 = n4597 ^ n4590 ;
  assign n4600 = n999 & n4599 ;
  assign n4578 = n3692 ^ n995 ;
  assign n4581 = n4578 ^ n2766 ;
  assign n4582 = n4581 ^ n4578 ;
  assign n4583 = ~n1000 & ~n4582 ;
  assign n4584 = n4583 ^ n4578 ;
  assign n4585 = n2003 & ~n4584 ;
  assign n4591 = n4590 ^ n4585 ;
  assign n4601 = n4600 ^ n4591 ;
  assign n4602 = n4601 ^ n4585 ;
  assign n4603 = ~n2810 & ~n4602 ;
  assign n4604 = n4577 & n4603 ;
  assign n4605 = n4604 ^ n4601 ;
  assign n4650 = n4649 ^ n4605 ;
  assign n4654 = n4653 ^ n4650 ;
  assign n4410 = n2667 ^ n1357 ;
  assign n4550 = ~n2670 & n3749 ;
  assign n4549 = n3422 & ~n3763 ;
  assign n4551 = n4550 ^ n4549 ;
  assign n4544 = n3380 ^ n2664 ;
  assign n4545 = n3763 ^ n3749 ;
  assign n4546 = n4389 & ~n4545 ;
  assign n4547 = n4546 ^ n3763 ;
  assign n4548 = ~n4544 & ~n4547 ;
  assign n4552 = n4551 ^ n4548 ;
  assign n4553 = n1357 & n4552 ;
  assign n4542 = ~n3718 & ~n4405 ;
  assign n4543 = ~n3756 & n4542 ;
  assign n4554 = n4553 ^ n4543 ;
  assign n4555 = n4552 ^ n1357 ;
  assign n4556 = n4555 ^ n4552 ;
  assign n4557 = ~n2667 & ~n3756 ;
  assign n4558 = n4557 ^ n4552 ;
  assign n4559 = n4556 & ~n4558 ;
  assign n4560 = n4559 ^ n4552 ;
  assign n4561 = ~n4554 & ~n4560 ;
  assign n4566 = n1406 & ~n3756 ;
  assign n4567 = n4566 ^ n3718 ;
  assign n4568 = n4561 & n4567 ;
  assign n4569 = n4568 ^ n4554 ;
  assign n4570 = n4410 & ~n4569 ;
  assign n4571 = n4338 ^ n3750 ;
  assign n4572 = n4571 ^ n4552 ;
  assign n4573 = n4556 & n4572 ;
  assign n4574 = n4573 ^ n4552 ;
  assign n4575 = n4570 & ~n4574 ;
  assign n4576 = n4575 ^ n4569 ;
  assign n4655 = n4654 ^ n4576 ;
  assign n4666 = n4665 ^ n4655 ;
  assign n4679 = n4678 ^ n4666 ;
  assign n4684 = n4683 ^ n4679 ;
  assign n4540 = n4509 ^ n4441 ;
  assign n4541 = n4442 & n4540 ;
  assign n4685 = n4684 ^ n4541 ;
  assign n4705 = n4704 ^ n4685 ;
  assign n4706 = n4705 ^ n4685 ;
  assign n4707 = n4539 & ~n4706 ;
  assign n4708 = n4536 & n4707 ;
  assign n4709 = n4708 ^ n4705 ;
  assign n4872 = n4685 ^ n4539 ;
  assign n4875 = n4372 & n4532 ;
  assign n4876 = n4872 & n4875 ;
  assign n4877 = n4194 & ~n4876 ;
  assign n4878 = n4877 ^ n4194 ;
  assign n4873 = n4535 & ~n4872 ;
  assign n4874 = ~n4194 & ~n4873 ;
  assign n4879 = n4878 ^ n4874 ;
  assign n4840 = n4665 ^ n4576 ;
  assign n4841 = ~n4655 & n4840 ;
  assign n4842 = n4841 ^ n4665 ;
  assign n4838 = ~n2690 & ~n4338 ;
  assign n4831 = n3422 & n3749 ;
  assign n4830 = ~n2666 & ~n3718 ;
  assign n4832 = n4831 ^ n4830 ;
  assign n4825 = n3718 ^ n1357 ;
  assign n4833 = n4832 ^ n4825 ;
  assign n4827 = n1357 & n3749 ;
  assign n4828 = n4827 ^ n3718 ;
  assign n4829 = n2665 & ~n4828 ;
  assign n4834 = n4833 ^ n4829 ;
  assign n4818 = n3718 ^ n2667 ;
  assign n4835 = n4834 ^ n4818 ;
  assign n4815 = n4338 ^ n3718 ;
  assign n4820 = ~n2667 & n4815 ;
  assign n4821 = n4820 ^ n3718 ;
  assign n4822 = ~n1406 & ~n4821 ;
  assign n4836 = n4835 ^ n4822 ;
  assign n4814 = ~n2667 & n4335 ;
  assign n4837 = n4836 ^ n4814 ;
  assign n4839 = n4838 ^ n4837 ;
  assign n4847 = n4842 ^ n4839 ;
  assign n4843 = ~n4839 & ~n4842 ;
  assign n4848 = n4847 ^ n4843 ;
  assign n4810 = n4653 ^ n4649 ;
  assign n4811 = n4650 & n4810 ;
  assign n4812 = n4811 ^ n4653 ;
  assign n4807 = n2003 & ~n3763 ;
  assign n4803 = ~n995 & ~n3800 ;
  assign n4804 = n4803 ^ n3692 ;
  assign n4805 = n2811 & n4804 ;
  assign n4795 = n999 & ~n2809 ;
  assign n4796 = n4795 ^ n2800 ;
  assign n4797 = ~n3800 & n4796 ;
  assign n4794 = ~n2787 & n2800 ;
  assign n4798 = n4797 ^ n4794 ;
  assign n4799 = n4798 ^ n4578 ;
  assign n4806 = n4805 ^ n4799 ;
  assign n4808 = n4807 ^ n4806 ;
  assign n4777 = n2643 ^ n780 ;
  assign n4778 = n1256 & n2783 ;
  assign n4779 = ~n4777 & n4778 ;
  assign n4772 = ~n2685 & n2924 ;
  assign n4771 = n2717 & n2920 ;
  assign n4773 = n4772 ^ n4771 ;
  assign n4774 = ~n694 & ~n4773 ;
  assign n4775 = n4774 ^ n694 ;
  assign n4776 = n4775 ^ n4773 ;
  assign n4780 = n4779 ^ n4776 ;
  assign n4770 = ~n3624 & n4244 ;
  assign n4781 = n4780 ^ n4770 ;
  assign n4782 = n4781 ^ n4774 ;
  assign n4783 = n4782 ^ n4781 ;
  assign n4784 = n1256 & ~n3623 ;
  assign n4785 = n4783 & n4784 ;
  assign n4786 = n4785 ^ n4782 ;
  assign n4748 = n697 & n2804 ;
  assign n4747 = n2718 ^ n708 ;
  assign n4749 = n4748 ^ n4747 ;
  assign n4754 = n697 & ~n2801 ;
  assign n4758 = ~n4749 & ~n4754 ;
  assign n4766 = n4758 ^ n4748 ;
  assign n4752 = n2719 & n2843 ;
  assign n4751 = ~n2720 & n2840 ;
  assign n4753 = n4752 ^ n4751 ;
  assign n4755 = n4754 ^ n4753 ;
  assign n4756 = n4755 ^ n4748 ;
  assign n4757 = n4756 ^ n707 ;
  assign n4759 = n4758 ^ n4749 ;
  assign n4760 = n4759 ^ n4748 ;
  assign n4763 = ~n707 & ~n4760 ;
  assign n4764 = n4763 ^ n4748 ;
  assign n4765 = n4757 & ~n4764 ;
  assign n4767 = n4766 ^ n4765 ;
  assign n4750 = n4749 ^ n4748 ;
  assign n4768 = n4767 ^ n4750 ;
  assign n4769 = n4768 ^ ~n4664 ;
  assign n4787 = n4786 ^ n4769 ;
  assign n4736 = n4643 ^ n2722 ;
  assign n4737 = n4643 ^ n4630 ;
  assign n4738 = n4737 ^ n4643 ;
  assign n4741 = ~n707 & ~n4738 ;
  assign n4742 = n4741 ^ n4643 ;
  assign n4743 = n4736 & n4742 ;
  assign n4744 = n4743 ^ n2722 ;
  assign n4745 = n4744 ^ n2721 ;
  assign n4746 = ~n707 & n4745 ;
  assign n4788 = n4787 ^ n4746 ;
  assign n4789 = n4788 ^ n4646 ;
  assign n4790 = n4789 ^ n4788 ;
  assign n4791 = n4790 ^ n4627 ;
  assign n4792 = n4648 & n4791 ;
  assign n4793 = n4792 ^ n4789 ;
  assign n4809 = n4808 ^ n4793 ;
  assign n4845 = n4812 ^ n4809 ;
  assign n4813 = ~n4809 & ~n4812 ;
  assign n4846 = n4845 ^ n4813 ;
  assign n4849 = n4848 ^ n4846 ;
  assign n4844 = n4843 ^ n4813 ;
  assign n4850 = n4849 ^ n4844 ;
  assign n4711 = n4423 & ~n4441 ;
  assign n4710 = n4506 ^ n4442 ;
  assign n4712 = n4711 ^ n4710 ;
  assign n4713 = n4712 ^ n4506 ;
  assign n4715 = n4514 & n4713 ;
  assign n4716 = n4715 ^ n4506 ;
  assign n4717 = ~n4510 & ~n4716 ;
  assign n4718 = n4717 ^ n4509 ;
  assign n4719 = n4514 ^ n4441 ;
  assign n4720 = n4442 & n4719 ;
  assign n4721 = n4720 ^ n4514 ;
  assign n4722 = n4666 & ~n4721 ;
  assign n4723 = n4509 & n4722 ;
  assign n4724 = ~n4506 & n4723 ;
  assign n4725 = n4724 ^ n4722 ;
  assign n4726 = n4725 ^ n4721 ;
  assign n4727 = n4718 & n4726 ;
  assign n4730 = n4666 ^ n4514 ;
  assign n4731 = n4730 ^ n4666 ;
  assign n4732 = n4711 & ~n4731 ;
  assign n4733 = n4732 ^ n4666 ;
  assign n4734 = n4727 & ~n4733 ;
  assign n4735 = n4734 ^ n4726 ;
  assign n4851 = n4850 ^ n4735 ;
  assign n4859 = n2518 ^ n837 ;
  assign n4855 = n1075 ^ n457 ;
  assign n4854 = n462 ^ n81 ;
  assign n4856 = n4855 ^ n4854 ;
  assign n4852 = n2485 ^ n279 ;
  assign n4853 = n4852 ^ n519 ;
  assign n4857 = n4856 ^ n4853 ;
  assign n4858 = n1039 & n4857 ;
  assign n4860 = n4859 ^ n4858 ;
  assign n4862 = n4851 & n4860 ;
  assign n4864 = n4678 ^ n4539 ;
  assign n4865 = ~n4685 & ~n4864 ;
  assign n4866 = n4865 ^ n4539 ;
  assign n4868 = n4862 & n4866 ;
  assign n4867 = n4866 ^ n4862 ;
  assign n4869 = n4868 ^ n4867 ;
  assign n4861 = n4860 ^ n4851 ;
  assign n4863 = n4862 ^ n4861 ;
  assign n4870 = n4869 ^ n4863 ;
  assign n4871 = n4870 ^ n4868 ;
  assign n4880 = n4879 ^ n4871 ;
  assign n5011 = n4863 & n4869 ;
  assign n4994 = n995 & ~n3786 ;
  assign n4995 = n4994 ^ n3763 ;
  assign n4996 = n2811 & ~n4995 ;
  assign n4992 = n3763 ^ n995 ;
  assign n4997 = n4996 ^ n4992 ;
  assign n4989 = n2003 & n3749 ;
  assign n4998 = n4997 ^ n4989 ;
  assign n4984 = n3372 ^ n2800 ;
  assign n4987 = ~n3786 & n4984 ;
  assign n4986 = n2800 & n3692 ;
  assign n4988 = n4987 ^ n4986 ;
  assign n4999 = n4998 ^ n4988 ;
  assign n4978 = ~n4769 & n4786 ;
  assign n4975 = n4786 ^ n4744 ;
  assign n4971 = n4786 ^ n707 ;
  assign n4972 = n4971 ^ n4769 ;
  assign n4976 = n4972 ^ n2721 ;
  assign n4977 = ~n4975 & ~n4976 ;
  assign n4979 = n4978 ^ n4977 ;
  assign n4980 = ~n707 & n4979 ;
  assign n4981 = n4980 ^ n4978 ;
  assign n4982 = n4981 ^ n4786 ;
  assign n4959 = ~n2685 & n2920 ;
  assign n4958 = n2643 & n2924 ;
  assign n4960 = n4959 ^ n4958 ;
  assign n4968 = n4960 ^ n694 ;
  assign n4964 = n1814 & n2784 ;
  assign n4961 = n4960 ^ n2787 ;
  assign n4962 = ~n694 & n4960 ;
  assign n4963 = ~n4961 & n4962 ;
  assign n4965 = n4964 ^ n4963 ;
  assign n4966 = n4965 ^ n4961 ;
  assign n4967 = n1256 & ~n4966 ;
  assign n4969 = n4968 ^ n4967 ;
  assign n4946 = ~n707 & ~n2721 ;
  assign n4948 = n4664 & n4768 ;
  assign n4951 = n4948 ^ n4769 ;
  assign n4949 = ~n2721 & n4948 ;
  assign n4947 = ~n707 & ~n2720 ;
  assign n4950 = n4949 ^ n4947 ;
  assign n4952 = n4951 ^ n4950 ;
  assign n4953 = n4952 ^ n4947 ;
  assign n4954 = ~n4946 & n4953 ;
  assign n4955 = n4954 ^ n4950 ;
  assign n4936 = n2240 ^ n707 ;
  assign n4937 = n4936 ^ n2839 ;
  assign n4938 = ~n3408 & n4937 ;
  assign n4932 = n2717 ^ n708 ;
  assign n4933 = n697 & ~n2805 ;
  assign n4934 = ~n4932 & n4933 ;
  assign n4917 = ~n708 & ~n2718 ;
  assign n4928 = n4917 ^ n707 ;
  assign n4918 = ~n2608 & ~n4917 ;
  assign n4929 = n4928 ^ n4918 ;
  assign n4921 = ~n707 & n2719 ;
  assign n4922 = n4921 ^ n2719 ;
  assign n4923 = n4922 ^ n2718 ;
  assign n4925 = ~n708 & n4923 ;
  assign n4926 = n4925 ^ n2718 ;
  assign n4927 = n2239 & n4926 ;
  assign n4930 = n4929 ^ n4927 ;
  assign n4919 = n2719 & ~n2838 ;
  assign n4920 = n4918 & n4919 ;
  assign n4931 = n4930 ^ n4920 ;
  assign n4935 = n4934 ^ n4931 ;
  assign n4939 = n4938 ^ n4935 ;
  assign n4956 = n4955 ^ n4939 ;
  assign n4940 = n4939 ^ n707 ;
  assign n4941 = n697 & n3409 ;
  assign n4942 = n4941 ^ n707 ;
  assign n4943 = n4940 & ~n4942 ;
  assign n4944 = n4943 ^ n707 ;
  assign n4945 = n4931 & ~n4944 ;
  assign n4957 = n4956 ^ n4945 ;
  assign n4970 = n4969 ^ n4957 ;
  assign n4983 = n4982 ^ n4970 ;
  assign n5000 = n4999 ^ n4983 ;
  assign n5002 = n5000 ^ n4788 ;
  assign n5001 = n5000 ^ n4808 ;
  assign n5003 = n5002 ^ n5001 ;
  assign n5004 = n4793 & n5003 ;
  assign n5005 = n5004 ^ n5002 ;
  assign n4898 = n2671 & ~n4335 ;
  assign n4899 = n4898 ^ n1357 ;
  assign n4902 = n4899 ^ n1406 ;
  assign n4903 = n4435 & n4902 ;
  assign n4906 = n4903 ^ n4899 ;
  assign n4897 = ~n1406 & n4664 ;
  assign n4900 = ~n3718 & n4899 ;
  assign n4901 = n4897 & n4900 ;
  assign n4904 = n4903 ^ n4901 ;
  assign n4905 = n2667 & n4904 ;
  assign n4907 = n4906 ^ n4905 ;
  assign n4908 = ~n1357 & ~n4907 ;
  assign n4913 = n3388 & ~n3718 ;
  assign n4914 = n4913 ^ n4898 ;
  assign n4915 = n4908 & n4914 ;
  assign n4916 = n4915 ^ n4907 ;
  assign n5006 = n5005 ^ n4916 ;
  assign n5007 = n5006 ^ n4844 ;
  assign n4894 = n4839 ^ n4735 ;
  assign n4895 = n4894 ^ n4842 ;
  assign n4896 = n4850 & n4895 ;
  assign n5008 = n5007 ^ n4896 ;
  assign n4886 = n414 ^ n323 ;
  assign n4887 = n4886 ^ n179 ;
  assign n4888 = n4887 ^ n2390 ;
  assign n4884 = n4076 ^ n332 ;
  assign n4883 = n437 ^ n280 ;
  assign n4885 = n4884 ^ n4883 ;
  assign n4889 = n4888 ^ n4885 ;
  assign n4890 = n4889 ^ n4325 ;
  assign n4891 = n4890 ^ n4203 ;
  assign n4881 = n605 ^ n533 ;
  assign n4882 = ~n515 & n4881 ;
  assign n4892 = n4891 ^ n4882 ;
  assign n4893 = n2705 & ~n4892 ;
  assign n5009 = n5008 ^ n4893 ;
  assign n5010 = n5009 ^ n4877 ;
  assign n5012 = n5011 ^ n5010 ;
  assign n5013 = n5012 ^ n5009 ;
  assign n5014 = n5013 ^ n5011 ;
  assign n5015 = n4866 ^ n4851 ;
  assign n5016 = n5015 ^ n4860 ;
  assign n5017 = ~n4874 & ~n5016 ;
  assign n5018 = ~n5014 & n5017 ;
  assign n5019 = n5018 ^ n5012 ;
  assign n5150 = n5006 ^ n4843 ;
  assign n5151 = ~n4813 & ~n5150 ;
  assign n5152 = n5006 ^ n4848 ;
  assign n5153 = n5152 ^ n5006 ;
  assign n5154 = n5006 ^ n4846 ;
  assign n5155 = n5154 ^ n5006 ;
  assign n5156 = ~n5153 & n5155 ;
  assign n5157 = n5156 ^ n5006 ;
  assign n5158 = n4735 & n5157 ;
  assign n5159 = n5151 & ~n5158 ;
  assign n5160 = n4842 ^ n4735 ;
  assign n5161 = n4894 & ~n5160 ;
  assign n5162 = n5161 ^ n4839 ;
  assign n5163 = n4846 & n5006 ;
  assign n5164 = ~n5162 & n5163 ;
  assign n5165 = n5164 ^ n5162 ;
  assign n5166 = ~n5159 & n5165 ;
  assign n5145 = n5000 ^ n4916 ;
  assign n5146 = ~n5005 & ~n5145 ;
  assign n5147 = n5146 ^ n5000 ;
  assign n5130 = n2664 ^ n1406 ;
  assign n5131 = n2664 ^ n1357 ;
  assign n5132 = ~n4335 & n5131 ;
  assign n5133 = ~n5130 & n5132 ;
  assign n5134 = n5133 ^ n1357 ;
  assign n5138 = ~n1406 & n4335 ;
  assign n5139 = n5138 ^ n2785 ;
  assign n5140 = ~n4336 & n5139 ;
  assign n5141 = n5140 ^ n1357 ;
  assign n5142 = n3902 & ~n5141 ;
  assign n5143 = n5134 & n5142 ;
  assign n5144 = n5143 ^ n5134 ;
  assign n5148 = n5147 ^ n5144 ;
  assign n5122 = n995 & ~n3756 ;
  assign n5123 = n5122 ^ n3749 ;
  assign n5124 = n2811 & n5123 ;
  assign n5120 = n3749 ^ n995 ;
  assign n5125 = n5124 ^ n5120 ;
  assign n5117 = n2003 & ~n3718 ;
  assign n5126 = n5125 ^ n5117 ;
  assign n5115 = ~n3756 & n4984 ;
  assign n5114 = n2800 & ~n3763 ;
  assign n5116 = n5115 ^ n5114 ;
  assign n5127 = n5126 ^ n5116 ;
  assign n5084 = n2842 ^ n2837 ;
  assign n5098 = n4949 ^ n4921 ;
  assign n5091 = n4949 ^ n4946 ;
  assign n5092 = n5091 ^ n4949 ;
  assign n5093 = n4951 ^ n4949 ;
  assign n5094 = n5093 ^ n4949 ;
  assign n5095 = ~n5092 & n5094 ;
  assign n5096 = n5095 ^ n4949 ;
  assign n5097 = ~n4947 & n5096 ;
  assign n5099 = n5098 ^ n5097 ;
  assign n5088 = ~n707 & ~n2718 ;
  assign n5089 = ~n2609 & ~n5088 ;
  assign n5087 = n2836 & n4917 ;
  assign n5090 = n5089 ^ n5087 ;
  assign n5100 = n5099 ^ n5090 ;
  assign n5085 = ~n707 & n2717 ;
  assign n5086 = n2608 & n5085 ;
  assign n5101 = n5100 ^ n5086 ;
  assign n5102 = n5101 ^ n5099 ;
  assign n5103 = n2717 ^ n707 ;
  assign n5104 = ~n5102 & n5103 ;
  assign n5105 = n5084 & n5104 ;
  assign n5106 = n5105 ^ n5101 ;
  assign n5077 = n2685 ^ n707 ;
  assign n5079 = n5077 ^ n3362 ;
  assign n5080 = n5079 ^ n5077 ;
  assign n5081 = n709 & ~n5080 ;
  assign n5082 = n5081 ^ n5077 ;
  assign n5083 = n697 & ~n5082 ;
  assign n5107 = n5106 ^ n5083 ;
  assign n5056 = n1256 & ~n2766 ;
  assign n5062 = n1256 & n3692 ;
  assign n5059 = ~n2787 & n2924 ;
  assign n5058 = n2643 & n2920 ;
  assign n5060 = n5059 ^ n5058 ;
  assign n5061 = n5060 ^ n694 ;
  assign n5063 = n5062 ^ n5061 ;
  assign n5057 = n3692 ^ n780 ;
  assign n5064 = n5063 ^ n5057 ;
  assign n5065 = n5056 & n5064 ;
  assign n5066 = n5065 ^ n5063 ;
  assign n5108 = n5107 ^ n5066 ;
  assign n5109 = n5108 ^ n4969 ;
  assign n5110 = n5109 ^ n5108 ;
  assign n5111 = n5110 ^ n4955 ;
  assign n5112 = ~n4957 & n5111 ;
  assign n5113 = n5112 ^ n5109 ;
  assign n5128 = n5127 ^ n5113 ;
  assign n5053 = n4999 ^ n4982 ;
  assign n5054 = ~n4983 & ~n5053 ;
  assign n5055 = n5054 ^ n4999 ;
  assign n5129 = n5128 ^ n5055 ;
  assign n5149 = n5148 ^ n5129 ;
  assign n5167 = n5166 ^ n5149 ;
  assign n5047 = n4204 ^ n4199 ;
  assign n5044 = n2275 ^ n332 ;
  assign n5045 = n5044 ^ n381 ;
  assign n5046 = n5045 ^ n2487 ;
  assign n5048 = n5047 ^ n5046 ;
  assign n5036 = n124 ^ n117 ;
  assign n5041 = ~n42 & n539 ;
  assign n5042 = n5041 ^ n317 ;
  assign n5043 = ~n5036 & n5042 ;
  assign n5049 = n5048 ^ n5043 ;
  assign n5033 = n3726 ^ n288 ;
  assign n5034 = n5033 ^ n321 ;
  assign n5030 = n2428 ^ n170 ;
  assign n5031 = n5030 ^ n668 ;
  assign n5032 = n5031 ^ n881 ;
  assign n5035 = n5034 ^ n5032 ;
  assign n5050 = n5049 ^ n5035 ;
  assign n5051 = n5050 ^ n2512 ;
  assign n5052 = n4069 & n5051 ;
  assign n5168 = n5167 ^ n5052 ;
  assign n5027 = n5011 ^ n5008 ;
  assign n5028 = ~n5009 & ~n5027 ;
  assign n5029 = n5028 ^ n5008 ;
  assign n5169 = n5168 ^ n5029 ;
  assign n5020 = n5009 ^ n4866 ;
  assign n5021 = n5020 ^ n4863 ;
  assign n5022 = n5021 ^ n4866 ;
  assign n5023 = n5009 ^ n4869 ;
  assign n5024 = ~n4868 & n4873 ;
  assign n5025 = n5023 & n5024 ;
  assign n5026 = n5022 & n5025 ;
  assign n5170 = n5169 ^ n5026 ;
  assign n5171 = n5170 ^ n5169 ;
  assign n5172 = n5009 ^ n4868 ;
  assign n5173 = n5172 ^ n4868 ;
  assign n5176 = n4871 & ~n5173 ;
  assign n5177 = n5176 ^ n4868 ;
  assign n5178 = n4876 & n5177 ;
  assign n5179 = n4194 & ~n5178 ;
  assign n5180 = ~n5171 & n5179 ;
  assign n5181 = n5180 ^ n5170 ;
  assign n5182 = n5026 & ~n5169 ;
  assign n5183 = ~n4194 & ~n5182 ;
  assign n5286 = n5167 ^ n5029 ;
  assign n5287 = ~n5168 & n5286 ;
  assign n5288 = n5287 ^ n5167 ;
  assign n5281 = n5055 & n5128 ;
  assign n5282 = n5281 ^ n5129 ;
  assign n5278 = n5144 & ~n5147 ;
  assign n5279 = n5278 ^ n5148 ;
  assign n5275 = n2003 & ~n4335 ;
  assign n5271 = ~n4338 & n4795 ;
  assign n5269 = n4338 ^ n3749 ;
  assign n5270 = n2800 & ~n5269 ;
  assign n5272 = n5271 ^ n5270 ;
  assign n5264 = n3718 ^ n995 ;
  assign n5273 = n5272 ^ n5264 ;
  assign n5266 = ~n995 & ~n4338 ;
  assign n5267 = n5266 ^ n3718 ;
  assign n5268 = n2811 & ~n5267 ;
  assign n5274 = n5273 ^ n5268 ;
  assign n5276 = n5275 ^ n5274 ;
  assign n5210 = n2719 & n4664 ;
  assign n5211 = ~n2720 & ~n2721 ;
  assign n5212 = n4768 & n5211 ;
  assign n5213 = n5210 & n5212 ;
  assign n5214 = n5213 ^ n2718 ;
  assign n5220 = n2842 ^ n2839 ;
  assign n5221 = n5220 ^ n2840 ;
  assign n5219 = ~n5665 ^ n707 ;
  assign n5222 = n5221 ^ n5219 ;
  assign n5223 = n5222 ^ n2840 ;
  assign n5224 = n2783 & ~n5223 ;
  assign n5218 = ~n2685 & n2843 ;
  assign n5225 = n5224 ^ n5218 ;
  assign n5216 = n697 & n2643 ;
  assign n5215 = n2717 & n2840 ;
  assign n5217 = n5216 ^ n5215 ;
  assign n5226 = n5225 ^ n5217 ;
  assign n5227 = n707 & ~n4951 ;
  assign n5228 = ~n5226 & n5227 ;
  assign n5229 = n5228 ^ n5226 ;
  assign n5240 = n5229 ^ n5214 ;
  assign n5237 = n5088 ^ ~n4664 ;
  assign n5232 = ~n4946 & ~n4947 ;
  assign n5233 = ~n4921 & n5232 ;
  assign n5234 = n4769 & n5233 ;
  assign n5235 = ~n4664 & ~n5234 ;
  assign n5231 = n5229 ^ n5213 ;
  assign n5236 = n5235 ^ n5231 ;
  assign n5238 = n5237 ^ n5236 ;
  assign n5239 = ~n5228 & ~n5238 ;
  assign n5241 = n5240 ^ n5239 ;
  assign n5242 = ~n5213 & ~n5241 ;
  assign n5243 = ~n5214 & ~n5242 ;
  assign n5249 = n5228 ^ n1357 ;
  assign n5250 = n5249 ^ n5214 ;
  assign n5251 = n5250 ^ n5242 ;
  assign n5247 = n5214 ^ n5213 ;
  assign n5248 = n5247 ^ n5240 ;
  assign n5252 = n5251 ^ n5248 ;
  assign n5244 = n5099 ^ n5066 ;
  assign n5245 = ~n5107 & n5244 ;
  assign n5246 = n5245 ^ n5099 ;
  assign n5253 = n5252 ^ n5246 ;
  assign n5254 = n5253 ^ n5251 ;
  assign n5255 = n5254 ^ n5246 ;
  assign n5256 = n5243 & ~n5255 ;
  assign n5257 = n5256 ^ n5253 ;
  assign n5207 = n2922 & ~n3800 ;
  assign n5206 = n2924 & n3692 ;
  assign n5208 = n5207 ^ n5206 ;
  assign n5204 = ~n2787 & n2920 ;
  assign n5200 = ~n694 & ~n3800 ;
  assign n5201 = n5200 ^ n3763 ;
  assign n5202 = n1256 & ~n5201 ;
  assign n5203 = n5202 ^ n694 ;
  assign n5205 = n5204 ^ n5203 ;
  assign n5209 = n5208 ^ n5205 ;
  assign n5258 = n5257 ^ n5209 ;
  assign n5260 = n5258 ^ n5108 ;
  assign n5259 = n5258 ^ n5127 ;
  assign n5261 = n5260 ^ n5259 ;
  assign n5262 = ~n5113 & ~n5261 ;
  assign n5263 = n5262 ^ n5260 ;
  assign n5277 = n5276 ^ n5263 ;
  assign n5280 = n5279 ^ n5277 ;
  assign n5283 = n5282 ^ n5280 ;
  assign n5194 = n5166 ^ n5148 ;
  assign n5195 = ~n5149 & n5194 ;
  assign n5284 = n5283 ^ n5195 ;
  assign n5188 = n840 ^ n75 ;
  assign n5187 = n4887 ^ n3680 ;
  assign n5189 = n5188 ^ n5187 ;
  assign n5190 = n5189 ^ n5049 ;
  assign n5186 = ~n319 & n563 ;
  assign n5191 = n5190 ^ n5186 ;
  assign n5185 = n159 & ~n4124 ;
  assign n5192 = n5191 ^ n5185 ;
  assign n5193 = n2356 & n5192 ;
  assign n5285 = n5284 ^ n5193 ;
  assign n5289 = n5288 ^ n5285 ;
  assign n5184 = n5169 & n5178 ;
  assign n5290 = n5289 ^ n5184 ;
  assign n5291 = n5290 ^ n5289 ;
  assign n5292 = n5183 & ~n5291 ;
  assign n5293 = n5292 ^ n5290 ;
  assign n5422 = n5182 & ~n5289 ;
  assign n5423 = ~n4194 & ~n5422 ;
  assign n5424 = n5423 ^ n4194 ;
  assign n5420 = n5184 & n5289 ;
  assign n5421 = n4194 & ~n5420 ;
  assign n5425 = n5424 ^ n5421 ;
  assign n5416 = n5288 ^ n5284 ;
  assign n5417 = n5285 & n5416 ;
  assign n5418 = n5417 ^ n5288 ;
  assign n5409 = n5276 ^ n5258 ;
  assign n5410 = ~n5263 & ~n5409 ;
  assign n5411 = n5410 ^ n5258 ;
  assign n5396 = n2915 & n4407 ;
  assign n5386 = n2924 & ~n3763 ;
  assign n5385 = n2920 & n3692 ;
  assign n5387 = n5386 ^ n5385 ;
  assign n5388 = n5387 ^ n694 ;
  assign n5389 = n1256 & n5388 ;
  assign n5392 = ~n780 & ~n3786 ;
  assign n5393 = n5392 ^ n3749 ;
  assign n5394 = n5389 & n5393 ;
  assign n5395 = n5394 ^ n5388 ;
  assign n5397 = n5396 ^ n5395 ;
  assign n5398 = ~n694 & ~n5397 ;
  assign n5401 = n1256 & n4406 ;
  assign n5402 = n3749 & n5401 ;
  assign n5403 = ~n780 & n5402 ;
  assign n5404 = n5403 ^ n5401 ;
  assign n5399 = n5387 ^ n1256 ;
  assign n5405 = n5404 ^ n5399 ;
  assign n5406 = n5398 & n5405 ;
  assign n5407 = n5406 ^ n5397 ;
  assign n5377 = n1357 ^ n707 ;
  assign n5378 = n5377 ^ ~n4664 ;
  assign n5372 = n4921 & n5212 ;
  assign n5373 = ~n5235 & n5372 ;
  assign n5374 = n5373 ^ n5235 ;
  assign n5375 = n5374 ^ n5088 ;
  assign n5376 = n5237 & n5375 ;
  assign n5379 = n5378 ^ n5376 ;
  assign n5380 = n5374 ^ n5226 ;
  assign n5381 = n5380 ^ n707 ;
  assign n5382 = ~n5379 & ~n5381 ;
  assign n5383 = n5382 ^ n5374 ;
  assign n5365 = ~n4664 ^ n1357 ;
  assign n5366 = ~n4664 ^ n707 ;
  assign n5367 = n5366 ^ n5088 ;
  assign n5368 = n5365 & ~n5367 ;
  assign n5369 = n5368 ^ n1357 ;
  assign n5370 = n5369 ^ n5085 ;
  assign n5355 = n2787 ^ n708 ;
  assign n5356 = n697 & n2784 ;
  assign n5357 = ~n5355 & n5356 ;
  assign n5342 = ~n2685 & n2840 ;
  assign n5341 = n2643 & n2843 ;
  assign n5343 = n5342 ^ n5341 ;
  assign n5344 = n5343 ^ n2787 ;
  assign n5345 = n5344 ^ n5343 ;
  assign n5348 = n5343 ^ n2784 ;
  assign n5349 = n5348 ^ n5343 ;
  assign n5350 = n697 & ~n5349 ;
  assign n5351 = ~n5345 & n5350 ;
  assign n5352 = n5351 ^ n5345 ;
  assign n5353 = n5352 ^ n5344 ;
  assign n5354 = ~n707 & n5353 ;
  assign n5358 = n5357 ^ n5354 ;
  assign n5359 = n5343 ^ n707 ;
  assign n5360 = ~n5358 & n5359 ;
  assign n5362 = n697 & n2767 ;
  assign n5363 = n5360 & n5362 ;
  assign n5361 = n5360 ^ n5358 ;
  assign n5364 = n5363 ^ n5361 ;
  assign n5371 = n5370 ^ n5364 ;
  assign n5384 = n5383 ^ n5371 ;
  assign n5408 = n5407 ^ n5384 ;
  assign n5412 = n5411 ^ n5408 ;
  assign n5332 = n2003 & n4435 ;
  assign n5334 = ~n2811 & ~n4335 ;
  assign n5333 = n2800 & ~n3718 ;
  assign n5335 = n5334 ^ n5333 ;
  assign n5336 = n5335 ^ n995 ;
  assign n5337 = n5336 ^ n999 ;
  assign n5338 = n5332 & ~n5337 ;
  assign n5339 = n5338 ^ n5336 ;
  assign n5329 = n5246 ^ n5209 ;
  assign n5330 = ~n5257 & n5329 ;
  assign n5331 = n5330 ^ n5209 ;
  assign n5340 = n5339 ^ n5331 ;
  assign n5413 = n5412 ^ n5340 ;
  assign n5310 = n5282 ^ n5277 ;
  assign n5311 = n5281 ^ n5166 ;
  assign n5312 = ~n5278 & ~n5281 ;
  assign n5313 = ~n5277 & n5312 ;
  assign n5314 = n5313 ^ n5281 ;
  assign n5315 = n5311 & ~n5314 ;
  assign n5317 = n5310 ^ n5280 ;
  assign n5318 = n5282 & n5317 ;
  assign n5319 = n5318 ^ n5310 ;
  assign n5320 = n5315 & ~n5319 ;
  assign n5321 = n5320 ^ n5314 ;
  assign n5322 = ~n5310 & n5321 ;
  assign n5323 = n5166 ^ n5147 ;
  assign n5324 = n5166 ^ n5144 ;
  assign n5325 = n5323 & ~n5324 ;
  assign n5326 = n5325 ^ n5166 ;
  assign n5327 = n5322 & ~n5326 ;
  assign n5328 = n5327 ^ n5321 ;
  assign n5414 = n5413 ^ n5328 ;
  assign n5303 = n341 ^ n284 ;
  assign n5304 = n5303 ^ n550 ;
  assign n5305 = n5304 ^ n2262 ;
  assign n5306 = n5305 ^ n4070 ;
  assign n5301 = n2627 ^ n144 ;
  assign n5302 = ~n80 & n5301 ;
  assign n5307 = n5306 ^ n5302 ;
  assign n5298 = n1024 ^ n858 ;
  assign n5297 = n838 ^ n577 ;
  assign n5299 = n5298 ^ n5297 ;
  assign n5295 = n2697 ^ n2497 ;
  assign n5294 = n2428 ^ n418 ;
  assign n5296 = n5295 ^ n5294 ;
  assign n5300 = n5299 ^ n5296 ;
  assign n5308 = n5307 ^ n5300 ;
  assign n5309 = n4139 & n5308 ;
  assign n5415 = n5414 ^ n5309 ;
  assign n5419 = n5418 ^ n5415 ;
  assign n5426 = n5425 ^ n5419 ;
  assign n5529 = n5421 ^ n5418 ;
  assign n5514 = n5331 & n5339 ;
  assign n5515 = n5408 & ~n5411 ;
  assign n5522 = n5515 ^ n5412 ;
  assign n5523 = ~n5514 & ~n5522 ;
  assign n5517 = ~n5514 & n5515 ;
  assign n5516 = n5515 ^ n5514 ;
  assign n5518 = n5517 ^ n5516 ;
  assign n5519 = n5412 & n5518 ;
  assign n5493 = n5407 ^ n5383 ;
  assign n5494 = n5384 & n5493 ;
  assign n5495 = n5494 ^ n5407 ;
  assign n5496 = n5495 ^ n995 ;
  assign n5497 = n5496 ^ n2810 ;
  assign n5498 = n5497 ^ n5495 ;
  assign n5499 = ~n1000 & ~n4335 ;
  assign n5500 = n5498 & n5499 ;
  assign n5501 = n5500 ^ n5496 ;
  assign n5502 = n5501 ^ n5495 ;
  assign n5505 = n999 & ~n4335 ;
  assign n5506 = n5505 ^ n995 ;
  assign n5507 = ~n4336 & ~n5506 ;
  assign n5508 = n5507 ^ n995 ;
  assign n5509 = ~n2809 & ~n5508 ;
  assign n5510 = n5502 & n5509 ;
  assign n5511 = n5510 ^ n5501 ;
  assign n5469 = n3718 ^ n780 ;
  assign n5470 = n1256 & ~n5469 ;
  assign n5471 = ~n3756 & n5470 ;
  assign n5466 = n2924 & n3749 ;
  assign n5465 = n2920 & ~n3763 ;
  assign n5467 = n5466 ^ n5465 ;
  assign n5468 = n5467 ^ n694 ;
  assign n5472 = n5471 ^ n5468 ;
  assign n5477 = n5472 ^ n5471 ;
  assign n5478 = n4338 ^ n3755 ;
  assign n5479 = n1256 & n5478 ;
  assign n5480 = n5477 & n5479 ;
  assign n5473 = n5369 ^ n5364 ;
  assign n5474 = n5370 & ~n5473 ;
  assign n5475 = n5474 ^ n5085 ;
  assign n5476 = n5475 ^ n5472 ;
  assign n5481 = n5480 ^ n5476 ;
  assign n5482 = n5481 ^ n5475 ;
  assign n5485 = n5467 ^ n4571 ;
  assign n5486 = n5485 ^ n5467 ;
  assign n5487 = n1256 & ~n5486 ;
  assign n5488 = n5487 ^ n5467 ;
  assign n5489 = ~n694 & n5488 ;
  assign n5490 = ~n5482 & n5489 ;
  assign n5491 = n5490 ^ n5481 ;
  assign n5451 = n2643 & n2865 ;
  assign n5450 = ~n2787 & n2842 ;
  assign n5452 = n5451 ^ n5450 ;
  assign n5453 = n5452 ^ n697 ;
  assign n5455 = n2717 ^ n2643 ;
  assign n5456 = ~n707 & n5455 ;
  assign n5454 = n5085 ^ n4023 ;
  assign n5457 = n5456 ^ n5454 ;
  assign n5458 = n694 & ~n5457 ;
  assign n5459 = n5458 ^ n2787 ;
  assign n5460 = ~n708 & ~n5459 ;
  assign n5461 = ~n5453 & n5460 ;
  assign n5462 = n5461 ^ n5453 ;
  assign n5443 = n3692 ^ n2766 ;
  assign n5444 = n5443 ^ n3692 ;
  assign n5447 = n709 & ~n5444 ;
  assign n5448 = n5447 ^ n3692 ;
  assign n5449 = n697 & ~n5448 ;
  assign n5463 = n5462 ^ n5449 ;
  assign n5441 = n2717 ^ n2685 ;
  assign n5442 = ~n707 & n5441 ;
  assign n5464 = n5463 ^ n5442 ;
  assign n5492 = n5491 ^ n5464 ;
  assign n5512 = n5511 ^ n5492 ;
  assign n5513 = n5512 ^ n5340 ;
  assign n5520 = n5519 ^ n5513 ;
  assign n5439 = n5340 ^ n5328 ;
  assign n5440 = ~n5413 & ~n5439 ;
  assign n5521 = n5520 ^ n5440 ;
  assign n5524 = n5523 ^ n5521 ;
  assign n5435 = n5034 ^ n842 ;
  assign n5431 = n2393 ^ n284 ;
  assign n5432 = n5431 ^ n409 ;
  assign n5430 = n783 ^ n383 ;
  assign n5433 = n5432 ^ n5430 ;
  assign n5434 = n5433 ^ n4209 ;
  assign n5436 = n5435 ^ n5434 ;
  assign n5437 = n5436 ^ n4080 ;
  assign n5438 = n2494 & ~n5437 ;
  assign n5525 = n5524 ^ n5438 ;
  assign n5427 = n5309 & ~n5414 ;
  assign n5428 = n5427 ^ n5415 ;
  assign n5429 = n5428 ^ n5423 ;
  assign n5526 = n5525 ^ n5429 ;
  assign n5527 = n5526 ^ n5428 ;
  assign n5528 = n5527 ^ n5525 ;
  assign n5530 = n5529 ^ n5528 ;
  assign n5531 = n5419 & ~n5530 ;
  assign n5532 = n5531 ^ n5526 ;
  assign n5639 = n4335 ^ n780 ;
  assign n5640 = n1256 & ~n4338 ;
  assign n5641 = n5639 & n5640 ;
  assign n5633 = n2920 & n3749 ;
  assign n5632 = n2924 & ~n3718 ;
  assign n5634 = n5633 ^ n5632 ;
  assign n5636 = n694 & n5634 ;
  assign n5642 = n5641 ^ n5636 ;
  assign n5638 = n4244 & n4434 ;
  assign n5643 = n5642 ^ n5638 ;
  assign n5635 = n5634 ^ n694 ;
  assign n5637 = n5636 ^ n5635 ;
  assign n5644 = n5643 ^ n5637 ;
  assign n5645 = n5644 ^ n5643 ;
  assign n5646 = n1256 & ~n4433 ;
  assign n5647 = ~n5645 & n5646 ;
  assign n5648 = n5647 ^ n5644 ;
  assign n5629 = n5495 ^ n5492 ;
  assign n5630 = ~n5511 & n5629 ;
  assign n5631 = n5630 ^ n5492 ;
  assign n5649 = n5648 ^ n5631 ;
  assign n5625 = n5456 ^ n995 ;
  assign n5620 = n5463 ^ n707 ;
  assign n5621 = n5620 ^ n2685 ;
  assign n5622 = ~n707 & ~n5441 ;
  assign n5623 = n5621 & n5622 ;
  assign n5624 = n5623 ^ n5620 ;
  assign n5626 = n5625 ^ n5624 ;
  assign n5590 = n2835 & ~n3692 ;
  assign n5614 = n2787 & n2836 ;
  assign n5611 = n3692 ^ n707 ;
  assign n5612 = ~n2240 & n5611 ;
  assign n5591 = n3763 ^ n707 ;
  assign n5594 = n5591 ^ n3800 ;
  assign n5595 = n5594 ^ n5591 ;
  assign n5596 = n709 & ~n5595 ;
  assign n5597 = n5596 ^ n5591 ;
  assign n5598 = n697 & n5597 ;
  assign n5610 = n5598 ^ n697 ;
  assign n5613 = n5612 ^ n5610 ;
  assign n5615 = n5614 ^ n5613 ;
  assign n5599 = n3692 ^ n2787 ;
  assign n5600 = n5599 ^ n694 ;
  assign n5601 = n5600 ^ n707 ;
  assign n5602 = n5601 ^ n5599 ;
  assign n5603 = n707 & ~n3692 ;
  assign n5604 = n5603 ^ n5599 ;
  assign n5605 = n5602 & n5604 ;
  assign n5606 = n5605 ^ n5599 ;
  assign n5607 = ~n697 & n5606 ;
  assign n5608 = n5607 ^ n697 ;
  assign n5609 = n708 & ~n5608 ;
  assign n5616 = n5615 ^ n5609 ;
  assign n5617 = n5616 ^ n5598 ;
  assign n5618 = n5590 & n5617 ;
  assign n5619 = n5618 ^ n5616 ;
  assign n5627 = n5626 ^ n5619 ;
  assign n5587 = n5475 ^ n5464 ;
  assign n5588 = ~n5491 & n5587 ;
  assign n5589 = n5588 ^ n5475 ;
  assign n5628 = n5627 ^ n5589 ;
  assign n5650 = n5649 ^ n5628 ;
  assign n5568 = n5514 ^ n5340 ;
  assign n5563 = n5512 ^ n5408 ;
  assign n5562 = n5514 ^ n5512 ;
  assign n5564 = n5563 ^ n5562 ;
  assign n5565 = n5564 ^ n5512 ;
  assign n5566 = ~n5412 & ~n5565 ;
  assign n5569 = n5566 ^ n5565 ;
  assign n5570 = ~n5568 & ~n5569 ;
  assign n5567 = n5566 ^ n5408 ;
  assign n5571 = n5570 ^ n5567 ;
  assign n5572 = n5412 ^ n5339 ;
  assign n5573 = n5572 ^ n5331 ;
  assign n5574 = n5512 ^ n5331 ;
  assign n5575 = n5574 ^ n5563 ;
  assign n5576 = n5512 ^ n5339 ;
  assign n5577 = n5576 ^ n5563 ;
  assign n5578 = ~n5575 & ~n5577 ;
  assign n5579 = n5578 ^ n5563 ;
  assign n5580 = ~n5573 & ~n5579 ;
  assign n5581 = n5328 & n5580 ;
  assign n5582 = n5581 ^ n5512 ;
  assign n5583 = n5582 ^ n5570 ;
  assign n5584 = n5583 ^ n5581 ;
  assign n5585 = ~n5571 & ~n5584 ;
  assign n5586 = n5585 ^ n5582 ;
  assign n5651 = n5650 ^ n5586 ;
  assign n5556 = n2520 ^ n570 ;
  assign n5554 = n295 ^ n250 ;
  assign n5555 = n5554 ^ n344 ;
  assign n5557 = n5556 ^ n5555 ;
  assign n5558 = n5557 ^ n4201 ;
  assign n5559 = ~n499 & ~n5558 ;
  assign n5560 = n4118 ^ n1174 ;
  assign n5561 = n5559 & n5560 ;
  assign n5652 = n5651 ^ n5561 ;
  assign n5536 = n5427 ^ n5418 ;
  assign n5550 = n5536 ^ n5438 ;
  assign n5533 = n5415 & ~n5418 ;
  assign n5551 = n5550 ^ n5533 ;
  assign n5552 = n5525 & n5551 ;
  assign n5553 = n5552 ^ n5524 ;
  assign n5653 = n5652 ^ n5553 ;
  assign n5535 = n5525 ^ n5427 ;
  assign n5537 = n5535 & n5536 ;
  assign n5538 = n5537 ^ n5428 ;
  assign n5543 = n5538 ^ n5537 ;
  assign n5544 = n5537 ^ n5525 ;
  assign n5545 = n5544 ^ n5537 ;
  assign n5546 = n5543 & n5545 ;
  assign n5547 = n5546 ^ n5537 ;
  assign n5548 = n5420 & n5547 ;
  assign n5654 = n5653 ^ n5548 ;
  assign n5534 = n5422 & ~n5533 ;
  assign n5539 = n5525 & ~n5538 ;
  assign n5540 = n5539 ^ n5428 ;
  assign n5541 = n5534 & n5540 ;
  assign n5542 = ~n4194 & ~n5541 ;
  assign n5549 = n5542 & ~n5548 ;
  assign n5655 = n5654 ^ n5549 ;
  assign n5656 = n5541 & n5653 ;
  assign n5657 = ~n4194 & ~n5656 ;
  assign n5714 = n5651 ^ n5553 ;
  assign n5715 = ~n5652 & ~n5714 ;
  assign n5716 = n5715 ^ n5651 ;
  assign n5710 = n3709 ^ n1080 ;
  assign n5706 = n358 ^ n273 ;
  assign n5707 = n5706 ^ n478 ;
  assign n5708 = n5707 ^ n583 ;
  assign n5705 = n1075 ^ n1031 ;
  assign n5709 = n5708 ^ n5705 ;
  assign n5711 = n5710 ^ n5709 ;
  assign n5712 = n561 & n5711 ;
  assign n5700 = n5631 & n5648 ;
  assign n5701 = n5700 ^ n5649 ;
  assign n5699 = ~n5589 & ~n5627 ;
  assign n5702 = n5701 ^ n5699 ;
  assign n5689 = n1256 & n4435 ;
  assign n5696 = n1814 & n5689 ;
  assign n5691 = n2924 & ~n4335 ;
  assign n5690 = n2920 & ~n3718 ;
  assign n5692 = n5691 ^ n5690 ;
  assign n5694 = n5692 ^ n694 ;
  assign n5697 = n5696 ^ n5694 ;
  assign n5675 = n2717 ^ n995 ;
  assign n5676 = ~n5455 & ~n5675 ;
  assign n5677 = n5676 ^ n995 ;
  assign n5678 = ~n2787 & ~n5677 ;
  assign n5679 = n5677 ^ n2787 ;
  assign n5680 = n5679 ^ n5678 ;
  assign n5681 = ~n707 & n5680 ;
  assign n5682 = ~n5678 & n5681 ;
  assign n5673 = n697 & n3749 ;
  assign n5669 = ~n707 & ~n3786 ;
  assign n5670 = n5669 ^ n3763 ;
  assign n5671 = ~n2843 & ~n5670 ;
  assign n5666 = ~n3786 & n5665 ;
  assign n5661 = n3786 ^ n3692 ;
  assign n5662 = n2840 & ~n5661 ;
  assign n5663 = n5662 ^ n3763 ;
  assign n5664 = n5663 ^ n707 ;
  assign n5667 = n5666 ^ n5664 ;
  assign n5672 = n5671 ^ n5667 ;
  assign n5674 = n5673 ^ n5672 ;
  assign n5683 = n5682 ^ n5674 ;
  assign n5684 = n5683 ^ n5624 ;
  assign n5685 = n5684 ^ n5619 ;
  assign n5686 = n5685 ^ n5683 ;
  assign n5687 = n5626 & n5686 ;
  assign n5688 = n5687 ^ n5684 ;
  assign n5698 = n5697 ^ n5688 ;
  assign n5703 = n5702 ^ n5698 ;
  assign n5659 = n5628 ^ n5586 ;
  assign n5660 = n5650 & ~n5659 ;
  assign n5704 = n5703 ^ n5660 ;
  assign n5713 = n5712 ^ n5704 ;
  assign n5717 = n5716 ^ n5713 ;
  assign n5658 = n5548 & ~n5653 ;
  assign n5718 = n5717 ^ n5658 ;
  assign n5719 = n5718 ^ n5717 ;
  assign n5720 = n5657 & ~n5719 ;
  assign n5721 = n5720 ^ n5718 ;
  assign n5722 = n5656 & ~n5717 ;
  assign n5723 = ~n4194 & ~n5722 ;
  assign n5777 = n5699 ^ n5628 ;
  assign n5778 = n5700 ^ n5698 ;
  assign n5779 = n5777 & n5778 ;
  assign n5784 = ~n5699 & ~n5701 ;
  assign n5785 = n5784 ^ n5698 ;
  assign n5786 = ~n5586 & ~n5785 ;
  assign n5787 = n5779 & ~n5786 ;
  assign n5788 = n5631 ^ n5586 ;
  assign n5789 = n5649 & ~n5788 ;
  assign n5790 = n5789 ^ n5648 ;
  assign n5791 = ~n5698 & ~n5699 ;
  assign n5792 = n5790 & n5791 ;
  assign n5793 = n5792 ^ n5790 ;
  assign n5794 = ~n5787 & ~n5793 ;
  assign n5766 = n3718 ^ n708 ;
  assign n5767 = n697 & ~n3756 ;
  assign n5768 = n5766 & n5767 ;
  assign n5760 = n2843 & n3749 ;
  assign n5759 = n2840 & ~n3763 ;
  assign n5761 = n5760 ^ n5759 ;
  assign n5763 = n707 & n5761 ;
  assign n5769 = n5768 ^ n5763 ;
  assign n5765 = ~n4571 & n4937 ;
  assign n5770 = n5769 ^ n5765 ;
  assign n5762 = n5761 ^ n707 ;
  assign n5764 = n5763 ^ n5762 ;
  assign n5771 = n5770 ^ n5764 ;
  assign n5772 = n5771 ^ n5770 ;
  assign n5773 = n697 & n5478 ;
  assign n5774 = ~n5772 & n5773 ;
  assign n5775 = n5774 ^ n5771 ;
  assign n5748 = n2919 & ~n4335 ;
  assign n5749 = n5748 ^ n694 ;
  assign n5750 = ~n2916 & n5749 ;
  assign n5753 = ~n780 & n4335 ;
  assign n5754 = n5753 ^ n1814 ;
  assign n5755 = ~n4336 & n5754 ;
  assign n5756 = n5755 ^ n5748 ;
  assign n5757 = n5750 & n5756 ;
  assign n5758 = n5757 ^ n5749 ;
  assign n5776 = n5775 ^ n5758 ;
  assign n5795 = n5794 ^ n5776 ;
  assign n5743 = n5674 & n5678 ;
  assign n5744 = n5743 ^ n3692 ;
  assign n5745 = ~n707 & n5744 ;
  assign n5742 = ~n5674 & ~n5681 ;
  assign n5746 = n5745 ^ n5742 ;
  assign n5739 = n5697 ^ n5683 ;
  assign n5740 = n5688 & ~n5739 ;
  assign n5741 = n5740 ^ n5683 ;
  assign n5747 = n5746 ^ n5741 ;
  assign n5796 = n5795 ^ n5747 ;
  assign n5728 = n2566 ^ n456 ;
  assign n5729 = n5728 ^ n467 ;
  assign n5730 = n5729 ^ n1071 ;
  assign n5731 = n5730 ^ n4521 ;
  assign n5732 = n5731 ^ n2327 ;
  assign n5733 = ~n424 & n5732 ;
  assign n5736 = ~n524 & n1064 ;
  assign n5734 = n607 ^ n267 ;
  assign n5735 = n5734 ^ n472 ;
  assign n5737 = n5736 ^ n5735 ;
  assign n5738 = n5733 & ~n5737 ;
  assign n5797 = n5796 ^ n5738 ;
  assign n5725 = n5716 ^ n5704 ;
  assign n5726 = n5713 & n5725 ;
  assign n5727 = n5726 ^ n5716 ;
  assign n5798 = n5797 ^ n5727 ;
  assign n5724 = n5658 & n5717 ;
  assign n5799 = n5798 ^ n5724 ;
  assign n5800 = n5799 ^ n5798 ;
  assign n5801 = n5723 & ~n5800 ;
  assign n5802 = n5801 ^ n5799 ;
  assign n5803 = n5722 & n5798 ;
  assign n5804 = ~n4194 & ~n5803 ;
  assign n5890 = n5796 ^ n5727 ;
  assign n5891 = n5797 & ~n5890 ;
  assign n5892 = n5891 ^ n5796 ;
  assign n5873 = n365 & n4091 ;
  assign n5882 = n543 ^ n444 ;
  assign n5883 = n5882 ^ n1012 ;
  assign n5880 = n447 ^ n381 ;
  assign n5881 = n5880 ^ n3728 ;
  assign n5884 = n5883 ^ n5881 ;
  assign n5878 = n4120 ^ n458 ;
  assign n5876 = n645 ^ n81 ;
  assign n5875 = n2459 ^ n225 ;
  assign n5877 = n5876 ^ n5875 ;
  assign n5879 = n5878 ^ n5877 ;
  assign n5885 = n5884 ^ n5879 ;
  assign n5874 = ~n359 & n432 ;
  assign n5886 = n5885 ^ n5874 ;
  assign n5887 = ~n4203 & ~n5886 ;
  assign n5888 = n5873 & n5887 ;
  assign n5841 = ~n3692 & n3734 ;
  assign n5842 = n5841 ^ n3692 ;
  assign n5843 = n5842 ^ n3763 ;
  assign n5844 = ~n707 & ~n5841 ;
  assign n5845 = ~n5843 & n5844 ;
  assign n5813 = n4335 ^ n708 ;
  assign n5814 = ~n4338 & n5813 ;
  assign n5817 = n5814 ^ n4433 ;
  assign n5819 = ~n707 & ~n3749 ;
  assign n5820 = ~n2610 & ~n5819 ;
  assign n5818 = ~n3718 & ~n5221 ;
  assign n5821 = n5820 ^ n5818 ;
  assign n5822 = n3718 ^ n707 ;
  assign n5834 = n2608 & n5822 ;
  assign n5831 = ~n2838 & ~n3749 ;
  assign n5832 = n708 & n5831 ;
  assign n5826 = n707 & ~n3749 ;
  assign n5827 = n5826 ^ n5822 ;
  assign n5828 = ~n708 & ~n5827 ;
  assign n5829 = n5828 ^ n5822 ;
  assign n5830 = n2239 & n5829 ;
  assign n5833 = n5832 ^ n5830 ;
  assign n5835 = n5834 ^ n5833 ;
  assign n5836 = ~n5821 & ~n5835 ;
  assign n5837 = n5817 & n5836 ;
  assign n5838 = n5837 ^ n5835 ;
  assign n5815 = n5814 ^ n4434 ;
  assign n5816 = n4937 & n5815 ;
  assign n5839 = n5838 ^ n5816 ;
  assign n5840 = n5839 ^ n694 ;
  assign n5846 = n5845 ^ n5840 ;
  assign n5809 = ~n707 & n3692 ;
  assign n5810 = ~n5742 & ~n5743 ;
  assign n5811 = n5809 & n5810 ;
  assign n5812 = n5811 ^ n5742 ;
  assign n5847 = n5846 ^ n5812 ;
  assign n5806 = ~n5741 & n5746 ;
  assign n5867 = n5847 ^ n5806 ;
  assign n5848 = ~n5806 & ~n5847 ;
  assign n5868 = n5867 ^ n5848 ;
  assign n5858 = ~n5747 & n5847 ;
  assign n5869 = n5868 ^ n5858 ;
  assign n5857 = n5794 ^ n5747 ;
  assign n5850 = ~n5758 & n5775 ;
  assign n5861 = n5858 ^ n5850 ;
  assign n5862 = n5861 ^ n5776 ;
  assign n5863 = n5858 & n5862 ;
  assign n5864 = n5863 ^ n5776 ;
  assign n5865 = ~n5857 & ~n5864 ;
  assign n5866 = n5865 ^ n5861 ;
  assign n5870 = n5869 ^ n5866 ;
  assign n5871 = n5870 ^ n5848 ;
  assign n5807 = n5806 ^ n5747 ;
  assign n5808 = ~n5794 & ~n5807 ;
  assign n5849 = n5848 ^ n5806 ;
  assign n5851 = n5850 ^ n5776 ;
  assign n5854 = ~n5849 & ~n5851 ;
  assign n5855 = n5854 ^ n5806 ;
  assign n5856 = n5808 & ~n5855 ;
  assign n5872 = n5871 ^ n5856 ;
  assign n5889 = n5888 ^ n5872 ;
  assign n5893 = n5892 ^ n5889 ;
  assign n5805 = n5724 & ~n5798 ;
  assign n5894 = n5893 ^ n5805 ;
  assign n5895 = n5894 ^ n5893 ;
  assign n5896 = n5804 & ~n5895 ;
  assign n5897 = n5896 ^ n5894 ;
  assign n5898 = n5803 & ~n5893 ;
  assign n5899 = ~n4194 & ~n5898 ;
  assign n5957 = n2268 & ~n2289 ;
  assign n5955 = ~n140 & n5301 ;
  assign n5949 = n473 ^ n410 ;
  assign n5950 = n5949 ^ n2566 ;
  assign n5946 = n831 ^ n331 ;
  assign n5947 = n5946 ^ n558 ;
  assign n5948 = n5947 ^ n3726 ;
  assign n5951 = n5950 ^ n5948 ;
  assign n5952 = n5951 ^ n1010 ;
  assign n5953 = n5952 ^ n1488 ;
  assign n5940 = n5839 ^ n5812 ;
  assign n5941 = ~n5846 & ~n5940 ;
  assign n5942 = n5941 ^ n5839 ;
  assign n5937 = n709 & n4435 ;
  assign n5938 = n697 & n5937 ;
  assign n5928 = n707 & ~n3718 ;
  assign n5929 = n5928 ^ n4335 ;
  assign n5930 = ~n708 & ~n5929 ;
  assign n5931 = n5930 ^ n4335 ;
  assign n5932 = n2239 & ~n5931 ;
  assign n5933 = n5932 ^ n2239 ;
  assign n5921 = ~n707 & n3718 ;
  assign n5922 = n5921 ^ n707 ;
  assign n5923 = n5922 ^ n4335 ;
  assign n5925 = n708 & n5923 ;
  assign n5926 = n5925 ^ n4335 ;
  assign n5927 = ~n2240 & n5926 ;
  assign n5934 = n5933 ^ n5927 ;
  assign n5935 = n5934 ^ n697 ;
  assign n5939 = n5938 ^ n5935 ;
  assign n5943 = n5942 ^ n5939 ;
  assign n5916 = ~n694 & ~n5841 ;
  assign n5917 = ~n5843 & n5916 ;
  assign n5918 = n5917 ^ n5843 ;
  assign n5919 = n5918 ^ n3749 ;
  assign n5920 = ~n707 & ~n5919 ;
  assign n5944 = n5943 ^ n5920 ;
  assign n5904 = n5808 & n5851 ;
  assign n5906 = ~n5850 & ~n5869 ;
  assign n5905 = n5869 ^ n5850 ;
  assign n5907 = n5906 ^ n5905 ;
  assign n5908 = ~n5848 & n5907 ;
  assign n5909 = ~n5794 & n5908 ;
  assign n5910 = n5851 ^ n5847 ;
  assign n5911 = n5867 & n5910 ;
  assign n5912 = n5911 ^ n5847 ;
  assign n5913 = ~n5906 & ~n5912 ;
  assign n5914 = ~n5909 & n5913 ;
  assign n5915 = ~n5904 & n5914 ;
  assign n5945 = n5944 ^ n5915 ;
  assign n5954 = n5953 ^ n5945 ;
  assign n5956 = n5955 ^ n5954 ;
  assign n5958 = n5957 ^ n5956 ;
  assign n5901 = n5892 ^ n5872 ;
  assign n5902 = ~n5889 & n5901 ;
  assign n5903 = n5902 ^ n5892 ;
  assign n5959 = n5958 ^ n5903 ;
  assign n5900 = n5805 & n5893 ;
  assign n5960 = n5959 ^ n5900 ;
  assign n5961 = n5960 ^ n5959 ;
  assign n5962 = n5899 & ~n5961 ;
  assign n5963 = n5962 ^ n5960 ;
  assign n5964 = n5900 & n5959 ;
  assign n5965 = n4194 & ~n5964 ;
  assign n6034 = n5945 ^ n5903 ;
  assign n6035 = n5958 & n6034 ;
  assign n6036 = n6035 ^ n5945 ;
  assign n5981 = ~n4335 & ~n5222 ;
  assign n5982 = n697 & n4336 ;
  assign n5983 = n5981 & ~n5982 ;
  assign n5993 = n3749 & ~n5922 ;
  assign n6026 = ~n5983 & n5993 ;
  assign n6001 = n3718 & ~n3749 ;
  assign n6007 = n6001 ^ n5983 ;
  assign n6008 = n6007 ^ n707 ;
  assign n6009 = n6008 ^ n5983 ;
  assign n6010 = n6009 ^ n5939 ;
  assign n5988 = n5939 ^ n707 ;
  assign n5989 = n5988 ^ n5918 ;
  assign n5990 = ~n707 & n5919 ;
  assign n5991 = n5989 & n5990 ;
  assign n5992 = n5991 ^ n5988 ;
  assign n5994 = n5992 & ~n5993 ;
  assign n6011 = n6010 ^ n5994 ;
  assign n6012 = n6011 ^ n6010 ;
  assign n6015 = ~n6001 & ~n6012 ;
  assign n6016 = n6015 ^ n6010 ;
  assign n6017 = ~n6007 & n6016 ;
  assign n6021 = n6008 & ~n6017 ;
  assign n5995 = n5994 ^ n5992 ;
  assign n6018 = n6010 ^ n5995 ;
  assign n6019 = n6018 ^ n6017 ;
  assign n6022 = n6019 ^ n5995 ;
  assign n6023 = n6022 ^ n707 ;
  assign n6024 = n6021 & ~n6023 ;
  assign n5984 = ~n3749 & ~n5983 ;
  assign n5985 = ~n5918 & ~n5939 ;
  assign n5986 = n5985 ^ n5921 ;
  assign n5987 = n5984 & n5986 ;
  assign n5996 = n5995 ^ n5987 ;
  assign n6002 = n5983 & ~n6001 ;
  assign n6003 = n5992 & n6002 ;
  assign n6004 = n6003 ^ n5992 ;
  assign n5997 = n5922 ^ n5819 ;
  assign n5998 = ~n5983 & ~n5997 ;
  assign n5999 = n5998 ^ n5983 ;
  assign n6000 = ~n5992 & n5999 ;
  assign n6005 = n6004 ^ n6000 ;
  assign n6006 = ~n5996 & n6005 ;
  assign n6020 = n6019 ^ n6006 ;
  assign n6025 = n6024 ^ n6020 ;
  assign n6027 = n6026 ^ n6025 ;
  assign n6028 = n5942 ^ n5915 ;
  assign n6029 = n5944 & ~n6028 ;
  assign n6030 = n6029 ^ n5942 ;
  assign n6031 = n6027 & ~n6030 ;
  assign n6032 = n6031 ^ n6006 ;
  assign n5969 = n4060 ^ n118 ;
  assign n5970 = n5969 ^ n201 ;
  assign n5971 = n5970 ^ n1035 ;
  assign n5972 = n5971 ^ n409 ;
  assign n5967 = n5946 ^ n286 ;
  assign n5968 = n5967 ^ n350 ;
  assign n5973 = n5972 ^ n5968 ;
  assign n5974 = n5973 ^ n4097 ;
  assign n5975 = n5974 ^ n1137 ;
  assign n5976 = n5975 ^ n2572 ;
  assign n5977 = n1004 ^ n321 ;
  assign n5978 = n5977 ^ n1195 ;
  assign n5979 = n5976 & n5978 ;
  assign n5980 = ~n5737 & n5979 ;
  assign n6033 = n6032 ^ n5980 ;
  assign n6037 = n6036 ^ n6033 ;
  assign n5966 = n5898 & ~n5959 ;
  assign n6038 = n6037 ^ n5966 ;
  assign n6039 = n6038 ^ n6037 ;
  assign n6040 = n5965 & ~n6039 ;
  assign n6041 = n6040 ^ n6038 ;
  assign n6042 = n5966 & n6037 ;
  assign n6043 = ~n4194 & ~n6042 ;
  assign n6108 = n6036 ^ n6032 ;
  assign n6109 = n6033 & ~n6108 ;
  assign n6110 = n6109 ^ n6036 ;
  assign n6094 = n391 ^ n245 ;
  assign n6093 = n4086 ^ n831 ;
  assign n6095 = n6094 ^ n6093 ;
  assign n6096 = n6095 ^ n2697 ;
  assign n6097 = n6096 ^ n4058 ;
  assign n6098 = n6097 ^ n5877 ;
  assign n6099 = n6098 ^ n4095 ;
  assign n6100 = n6099 ^ n1094 ;
  assign n6056 = n5832 ^ n3749 ;
  assign n6049 = n4335 ^ n3718 ;
  assign n6050 = n6049 ^ n5832 ;
  assign n6053 = n6050 ^ n3749 ;
  assign n6057 = n6056 ^ n6053 ;
  assign n6069 = n6056 ^ n4335 ;
  assign n6070 = n6069 ^ n6057 ;
  assign n6072 = ~n6056 & n6070 ;
  assign n6062 = n4335 ^ n707 ;
  assign n6065 = n6057 ^ n4335 ;
  assign n6063 = n6057 ^ n3749 ;
  assign n6064 = n6063 ^ n707 ;
  assign n6066 = n6065 ^ n6064 ;
  assign n6067 = n6062 & ~n6066 ;
  assign n6073 = n6072 ^ n6067 ;
  assign n6074 = n6073 ^ n6065 ;
  assign n6075 = n6072 ^ n6063 ;
  assign n6076 = n6075 ^ n6065 ;
  assign n6077 = ~n6074 & ~n6076 ;
  assign n6078 = ~n6057 & n6077 ;
  assign n6079 = n6078 ^ n6072 ;
  assign n6087 = n6079 ^ n3749 ;
  assign n6090 = n707 & ~n5983 ;
  assign n6091 = n6087 & n6090 ;
  assign n6088 = n6087 ^ n6000 ;
  assign n6045 = n6004 ^ n5998 ;
  assign n6046 = ~n6000 & ~n6030 ;
  assign n6047 = ~n6045 & n6046 ;
  assign n6089 = n6088 ^ n6047 ;
  assign n6092 = n6091 ^ n6089 ;
  assign n6101 = n6100 ^ n6092 ;
  assign n6102 = n6101 ^ n6092 ;
  assign n6103 = ~n2457 & ~n6102 ;
  assign n6104 = n2338 & n6103 ;
  assign n6105 = n117 & n6104 ;
  assign n6106 = n6105 ^ n6103 ;
  assign n6107 = n6106 ^ n6101 ;
  assign n6111 = n6110 ^ n6107 ;
  assign n6044 = n5964 & ~n6037 ;
  assign n6112 = n6111 ^ n6044 ;
  assign n6113 = n6112 ^ n6111 ;
  assign n6114 = n6043 & ~n6113 ;
  assign n6115 = n6114 ^ n6112 ;
  assign n6124 = n330 ^ n304 ;
  assign n6125 = n6124 ^ n480 ;
  assign n6126 = n6125 ^ n1089 ;
  assign n6122 = n2281 ^ n861 ;
  assign n6123 = n6122 ^ n5880 ;
  assign n6127 = n6126 ^ n6123 ;
  assign n6128 = n6127 ^ n688 ;
  assign n6129 = n6128 ^ n2705 ;
  assign n6120 = n380 ^ n105 ;
  assign n6121 = ~n524 & n6120 ;
  assign n6130 = n6129 ^ n6121 ;
  assign n6117 = n6110 ^ n6092 ;
  assign n6118 = ~n6107 & ~n6117 ;
  assign n6119 = n6118 ^ n6110 ;
  assign n6131 = n6130 ^ n6119 ;
  assign n6116 = n6042 & ~n6111 ;
  assign n6132 = n6131 ^ n6116 ;
  assign n6133 = n6132 ^ n6131 ;
  assign n6134 = n6044 & n6111 ;
  assign n6135 = n4194 & ~n6134 ;
  assign n6136 = ~n6133 & n6135 ;
  assign n6137 = n6136 ^ n6132 ;
  assign n6149 = n1015 ^ n364 ;
  assign n6146 = n1041 ^ n549 ;
  assign n6145 = n4669 ^ n4056 ;
  assign n6147 = n6146 ^ n6145 ;
  assign n6148 = n6147 ^ n1212 ;
  assign n6150 = n6149 ^ n6148 ;
  assign n6151 = n6150 ^ n626 ;
  assign n6152 = n6151 ^ n1153 ;
  assign n6153 = n4136 & ~n6152 ;
  assign n6144 = n6119 & ~n6130 ;
  assign n6154 = n6153 ^ n6144 ;
  assign n6138 = n6131 ^ n4194 ;
  assign n6139 = n6134 ^ n6116 ;
  assign n6141 = n6131 & n6139 ;
  assign n6142 = n6141 ^ n6116 ;
  assign n6143 = ~n6138 & ~n6142 ;
  assign n6155 = n6154 ^ n6143 ;
  assign n6172 = n6116 & ~n6153 ;
  assign n6173 = n6172 ^ n6153 ;
  assign n6174 = n6173 ^ n6119 ;
  assign n6175 = n6174 ^ n6172 ;
  assign n6176 = n6172 ^ n6134 ;
  assign n6177 = n6176 ^ n6172 ;
  assign n6178 = ~n6175 & n6177 ;
  assign n6179 = n6178 ^ n6172 ;
  assign n6180 = n6131 & n6179 ;
  assign n6181 = n6180 ^ n6172 ;
  assign n6182 = n4194 & ~n6181 ;
  assign n6164 = n444 ^ n265 ;
  assign n6165 = n6164 ^ n400 ;
  assign n6161 = n548 ^ n154 ;
  assign n6162 = n6161 ^ n517 ;
  assign n6163 = n6162 ^ n263 ;
  assign n6166 = n6165 ^ n6163 ;
  assign n6167 = n6166 ^ n4887 ;
  assign n6168 = ~n2630 & n6167 ;
  assign n6169 = n1062 & n6168 ;
  assign n6170 = n5978 & n6169 ;
  assign n6156 = n6130 ^ n6116 ;
  assign n6157 = n6119 ^ n6116 ;
  assign n6158 = n6156 & ~n6157 ;
  assign n6159 = n6158 ^ n6116 ;
  assign n6160 = ~n6153 & n6159 ;
  assign n6171 = n6170 ^ n6160 ;
  assign n6183 = n6182 ^ n6171 ;
  assign n6190 = n4328 ^ n154 ;
  assign n6191 = n247 & n6190 ;
  assign n6188 = n335 ^ n238 ;
  assign n6187 = n674 ^ n80 ;
  assign n6189 = n6188 ^ n6187 ;
  assign n6192 = n6191 ^ n6189 ;
  assign n6193 = ~n4884 & n6192 ;
  assign n6194 = n6193 ^ n3721 ;
  assign n6195 = n1022 & n6194 ;
  assign n6196 = n5307 & n6195 ;
  assign n6197 = n6196 ^ n4194 ;
  assign n6184 = n6182 ^ n4194 ;
  assign n6185 = n6184 ^ n6160 ;
  assign n6186 = n6171 & n6185 ;
  assign n6198 = n6197 ^ n6186 ;
  assign n6201 = n173 ^ n110 ;
  assign n6202 = n642 ^ n566 ;
  assign n6203 = n6202 ^ n614 ;
  assign n6204 = n6203 ^ n3741 ;
  assign n6205 = ~n689 & ~n6204 ;
  assign n6206 = n6201 & n6205 ;
  assign n6207 = n6206 ^ n6204 ;
  assign n6208 = n6207 ^ n4194 ;
  assign n6199 = n6196 ^ n6170 ;
  assign n6200 = n6186 & ~n6199 ;
  assign n6209 = n6208 ^ n6200 ;
  assign n6215 = n6207 ^ n6160 ;
  assign n6216 = n6207 ^ n6196 ;
  assign n6217 = ~n6199 & n6216 ;
  assign n6218 = ~n6215 & n6217 ;
  assign n6219 = n6181 & n6218 ;
  assign n6220 = n4194 & ~n6219 ;
  assign n6211 = ~n6170 & ~n6196 ;
  assign n6212 = n6207 & n6211 ;
  assign n6213 = n6160 & n6212 ;
  assign n6210 = n1252 & ~n3746 ;
  assign n6214 = n6213 ^ n6210 ;
  assign n6221 = n6220 ^ n6214 ;
  assign n6222 = n6210 & ~n6213 ;
  assign n6223 = n6222 ^ n6214 ;
  assign n6224 = ~n6184 & n6223 ;
  assign n6225 = n6224 ^ n4194 ;
  assign n6226 = ~x21 & ~x22 ;
  assign n6227 = n6222 & ~n6226 ;
  assign n6228 = n6219 & n6227 ;
  assign n6231 = n6228 ^ n6226 ;
  assign n6232 = n6231 ^ n6228 ;
  assign n6233 = n1252 & n6232 ;
  assign n6234 = n6233 ^ n6228 ;
  assign n6235 = ~n6225 & ~n6234 ;
  assign n6236 = n6235 ^ n6228 ;
  assign n6237 = n4194 & ~n6228 ;
  assign y0 = n4193 ;
  assign y1 = ~n4363 ;
  assign y2 = ~n4534 ;
  assign y3 = ~n4709 ;
  assign y4 = n4880 ;
  assign y5 = n5019 ;
  assign y6 = ~n5181 ;
  assign y7 = n5293 ;
  assign y8 = n5426 ;
  assign y9 = ~n5532 ;
  assign y10 = ~n5655 ;
  assign y11 = n5721 ;
  assign y12 = ~n5802 ;
  assign y13 = n5897 ;
  assign y14 = n5963 ;
  assign y15 = n6041 ;
  assign y16 = n6115 ;
  assign y17 = ~n6137 ;
  assign y18 = n6155 ;
  assign y19 = ~n6183 ;
  assign y20 = ~n6198 ;
  assign y21 = n6209 ;
  assign y22 = ~n6221 ;
  assign y23 = ~n6236 ;
  assign y24 = n6237 ;
endmodule
