module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n18 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n36 , n37 , n38 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n142 , n150 , n151 , n154 , n155 , n156 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n269 , n271 , n275 , n276 , n277 , n278 , n281 , n282 , n283 , n286 , n287 , n288 , n289 , n290 , n293 , n294 , n295 , n310 , n313 , n317 , n318 , n319 , n320 , n321 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n480 , n481 , n482 , n483 , n484 , n485 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n600 , n601 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n814 , n821 , n822 , n823 , n824 , n826 , n827 , n829 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n840 , n843 , n847 , n848 , n854 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n925 , n926 , n927 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n940 , n941 , n942 , n943 , n945 , n946 , n947 , n948 , n949 ;
  assign n11 = x5 & x6 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ x5 ;
  assign n29 = x3 ^ x2 ;
  assign n30 = x0 & ~n29 ;
  assign n31 = ~x3 & x9 ;
  assign n24 = x8 & ~x9 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n30 & n32 ;
  assign n23 = x9 ^ x8 ;
  assign n25 = n24 ^ n23 ;
  assign n34 = n25 ^ x8 ;
  assign n14 = x2 & x3 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n15 ^ x3 ;
  assign n38 = n16 ^ x2 ;
  assign n43 = ~n34 & n38 ;
  assign n632 = n25 ^ x9 ;
  assign n36 = ~n15 & n632 ;
  assign n37 = n632 ^ n36 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = ~x0 & n44 ;
  assign n46 = ~n33 & ~n45 ;
  assign n47 = ~x7 & ~n46 ;
  assign n48 = n24 ^ x2 ;
  assign n49 = ~x3 & ~n48 ;
  assign n51 = n632 ^ x0 ;
  assign n52 = ~x7 & ~n632 ;
  assign n53 = ~n51 & n52 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n49 & ~n54 ;
  assign n56 = ~n47 & ~n55 ;
  assign n57 = ~x1 & ~n56 ;
  assign n221 = ~x7 & x8 ;
  assign n20 = n221 ^ x7 ;
  assign n58 = n57 ^ n20 ;
  assign n21 = ~n16 & n20 ;
  assign n22 = ~x7 & ~x9 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = n21 & n27 ;
  assign n59 = n58 ^ n28 ;
  assign n60 = ~n13 & ~n59 ;
  assign n66 = ~x0 & x2 ;
  assign n65 = x2 ^ x0 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = ~x9 & n67 ;
  assign n63 = x2 & n34 ;
  assign n61 = ~x2 & x8 ;
  assign n62 = n61 ^ x8 ;
  assign n64 = n63 ^ n62 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = x1 & n69 ;
  assign n71 = x3 & ~n61 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = x1 & ~x9 ;
  assign n74 = n73 ^ x1 ;
  assign n75 = n74 ^ x9 ;
  assign n76 = n75 ^ x2 ;
  assign n77 = x0 & ~x1 ;
  assign n78 = ~x3 & ~n62 ;
  assign n79 = n77 & n78 ;
  assign n80 = n76 & n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = ~n72 & ~n81 ;
  assign n94 = x9 ^ x1 ;
  assign n90 = x8 ^ x0 ;
  assign n89 = x0 & ~x8 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = x1 & ~n91 ;
  assign n93 = n92 ^ n74 ;
  assign n95 = n94 ^ n93 ;
  assign n85 = ~x1 & n34 ;
  assign n83 = ~x1 & x8 ;
  assign n84 = n83 ^ x1 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n86 ^ x1 ;
  assign n88 = n632 ^ n87 ;
  assign n96 = n95 ^ n88 ;
  assign n97 = n96 ^ x8 ;
  assign n100 = ~x7 & ~n13 ;
  assign n98 = x6 & ~x7 ;
  assign n99 = n98 ^ x7 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = ~n97 & ~n101 ;
  assign n103 = ~n82 & n102 ;
  assign n124 = n38 ^ x8 ;
  assign n125 = ~x5 & n124 ;
  assign n126 = n125 ^ x8 ;
  assign n117 = x5 & x9 ;
  assign n135 = n126 ^ n117 ;
  assign n123 = n77 ^ x1 ;
  assign n150 = n135 ^ n123 ;
  assign n119 = x9 ^ x0 ;
  assign n118 = ~x0 & ~x9 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = ~n117 & n120 ;
  assign n122 = n120 ^ n36 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = ~n123 & ~n127 ;
  assign n129 = n128 ^ n117 ;
  assign n130 = n129 ^ n122 ;
  assign n131 = n130 ^ n123 ;
  assign n132 = n122 & ~n131 ;
  assign n133 = n121 & n132 ;
  assign n134 = n133 ^ n130 ;
  assign n151 = n150 ^ n134 ;
  assign n159 = n151 ^ n117 ;
  assign n160 = n159 ^ n123 ;
  assign n136 = n135 ^ n127 ;
  assign n142 = n136 ^ n120 ;
  assign n137 = n136 ^ n36 ;
  assign n138 = n137 ^ n127 ;
  assign n154 = n142 ^ n138 ;
  assign n155 = n154 ^ n135 ;
  assign n156 = n155 ^ n126 ;
  assign n161 = n160 ^ n156 ;
  assign n104 = n84 ^ x8 ;
  assign n105 = n104 ^ n92 ;
  assign n162 = n161 ^ n105 ;
  assign n106 = n16 ^ x8 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = n107 ^ x8 ;
  assign n109 = n105 ^ x5 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = n108 & n110 ;
  assign n116 = n111 ^ n98 ;
  assign n163 = n162 ^ n116 ;
  assign n112 = x1 & ~x2 ;
  assign n113 = n112 ^ x2 ;
  assign n114 = n107 & ~n113 ;
  assign n115 = n111 & n114 ;
  assign n164 = n163 ^ n115 ;
  assign n165 = ~n16 & ~n123 ;
  assign n170 = n117 ^ n24 ;
  assign n168 = ~x5 & ~n632 ;
  assign n166 = x5 & x8 ;
  assign n167 = n166 ^ x8 ;
  assign n169 = n168 ^ n167 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = n98 & ~n171 ;
  assign n173 = ~n165 & n172 ;
  assign n174 = n173 ^ n98 ;
  assign n175 = n161 & n174 ;
  assign n176 = ~n164 & n175 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n62 & n77 ;
  assign n179 = n178 ^ n89 ;
  assign n180 = x9 ^ x5 ;
  assign n181 = n180 ^ n117 ;
  assign n182 = ~x0 & ~n181 ;
  assign n183 = x8 ^ x3 ;
  assign n184 = x2 ^ x1 ;
  assign n185 = ~n29 & n184 ;
  assign n186 = n183 & n185 ;
  assign n187 = n186 ^ x8 ;
  assign n188 = n182 & ~n187 ;
  assign n189 = n188 ^ n181 ;
  assign n190 = n179 & ~n189 ;
  assign n198 = ~x3 & n190 ;
  assign n199 = n84 & n198 ;
  assign n200 = n199 ^ n84 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = n191 ^ n84 ;
  assign n201 = n200 ^ n192 ;
  assign n202 = n177 & n201 ;
  assign n203 = ~n103 & ~n202 ;
  assign n204 = ~n60 & n203 ;
  assign n205 = x6 ^ x5 ;
  assign n206 = ~n34 & n165 ;
  assign n207 = n165 ^ x4 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = n206 & n208 ;
  assign n210 = n205 & n209 ;
  assign n211 = n210 ^ n208 ;
  assign n212 = ~n204 & ~n211 ;
  assign n217 = n31 ^ x3 ;
  assign n218 = x1 ^ x0 ;
  assign n222 = n221 ^ x2 ;
  assign n536 = x8 ^ x1 ;
  assign n223 = ~n222 & n536 ;
  assign n224 = n223 ^ x2 ;
  assign n225 = n218 & ~n224 ;
  assign n226 = ~n217 & n225 ;
  assign n227 = n632 ^ x7 ;
  assign n228 = ~x3 & ~n113 ;
  assign n229 = n228 ^ x3 ;
  assign n230 = n227 & ~n229 ;
  assign n231 = n123 ^ n67 ;
  assign n232 = n230 & ~n231 ;
  assign n233 = ~n226 & ~n232 ;
  assign n214 = n22 & ~n178 ;
  assign n234 = n233 ^ n214 ;
  assign n213 = n61 ^ x2 ;
  assign n215 = ~n123 & n214 ;
  assign n216 = ~n213 & n215 ;
  assign n235 = n234 ^ n216 ;
  assign n236 = ~n13 & ~n235 ;
  assign n237 = ~x1 & ~x5 ;
  assign n239 = n119 ^ n31 ;
  assign n238 = ~x0 & x3 ;
  assign n240 = n239 ^ n238 ;
  assign n241 = n23 & n240 ;
  assign n242 = n241 ^ x3 ;
  assign n243 = n237 & ~n242 ;
  assign n244 = n180 ^ n169 ;
  assign n245 = x3 ^ x1 ;
  assign n246 = x1 & n245 ;
  assign n247 = n246 ^ n74 ;
  assign n248 = ~n244 & n247 ;
  assign n249 = x2 & ~n117 ;
  assign n250 = ~n248 & n249 ;
  assign n251 = ~n243 & n250 ;
  assign n293 = n245 ^ x0 ;
  assign n294 = n293 ^ n117 ;
  assign n295 = n294 ^ x3 ;
  assign n275 = ~n294 & n295 ;
  assign n276 = n275 ^ x1 ;
  assign n277 = n276 ^ n26 ;
  assign n278 = n277 ^ x3 ;
  assign n281 = ~n278 & ~n293 ;
  assign n310 = n117 ^ x3 ;
  assign n282 = n310 ^ n25 ;
  assign n283 = n282 ^ n117 ;
  assign n286 = n245 & ~n283 ;
  assign n287 = n281 & n286 ;
  assign n288 = n287 ^ n275 ;
  assign n271 = n25 ^ x1 ;
  assign n289 = n288 ^ n271 ;
  assign n313 = n310 ^ n26 ;
  assign n269 = n313 ^ n117 ;
  assign n290 = n289 ^ n269 ;
  assign n317 = n98 & n290 ;
  assign n318 = ~x2 & n181 ;
  assign n319 = n77 ^ x0 ;
  assign n326 = ~n16 & n319 ;
  assign n320 = n318 ^ n117 ;
  assign n321 = n320 ^ n92 ;
  assign n327 = n326 ^ n321 ;
  assign n328 = ~n318 & ~n327 ;
  assign n329 = n328 ^ n321 ;
  assign n330 = n329 ^ n318 ;
  assign n331 = n117 ^ n92 ;
  assign n332 = n320 & ~n331 ;
  assign n333 = ~n330 & n332 ;
  assign n334 = n333 ^ n329 ;
  assign n335 = n317 & ~n334 ;
  assign n336 = n335 ^ n98 ;
  assign n337 = ~n251 & n336 ;
  assign n339 = n31 ^ n15 ;
  assign n338 = ~x9 & ~n15 ;
  assign n340 = n339 ^ n338 ;
  assign n341 = ~n88 & n340 ;
  assign n342 = ~x0 & n341 ;
  assign n343 = x1 & ~n61 ;
  assign n344 = n338 & n343 ;
  assign n345 = n344 ^ n338 ;
  assign n346 = ~n342 & ~n345 ;
  assign n350 = n64 ^ n37 ;
  assign n351 = n350 ^ n217 ;
  assign n348 = n15 ^ x9 ;
  assign n349 = n348 ^ n338 ;
  assign n352 = n351 ^ n349 ;
  assign n353 = x1 & n352 ;
  assign n347 = ~x3 & n178 ;
  assign n354 = n353 ^ n347 ;
  assign n355 = n346 & ~n354 ;
  assign n356 = ~n101 & ~n355 ;
  assign n357 = ~n337 & ~n356 ;
  assign n358 = ~n236 & n357 ;
  assign n366 = n34 & n165 ;
  assign n359 = ~x0 & ~x6 ;
  assign n360 = ~x9 & ~n359 ;
  assign n361 = n228 & ~n360 ;
  assign n367 = n366 ^ n361 ;
  assign n368 = ~x4 & ~n367 ;
  assign n369 = n368 ^ n361 ;
  assign n370 = ~n358 & n369 ;
  assign n428 = ~x2 & ~n91 ;
  assign n427 = n66 ^ n61 ;
  assign n429 = n428 ^ n427 ;
  assign n430 = n31 & n429 ;
  assign n412 = ~x1 & ~x6 ;
  assign n411 = x6 ^ x1 ;
  assign n413 = n412 ^ n411 ;
  assign n414 = n413 ^ x1 ;
  assign n431 = ~n24 & ~n414 ;
  assign n389 = ~x2 & x6 ;
  assign n390 = n389 ^ x2 ;
  assign n432 = n390 ^ x6 ;
  assign n433 = ~x3 & ~n432 ;
  assign n434 = ~n431 & n433 ;
  assign n435 = ~n430 & ~n434 ;
  assign n378 = ~x6 & x8 ;
  assign n436 = n390 ^ n378 ;
  assign n437 = n436 ^ n213 ;
  assign n438 = n437 ^ x2 ;
  assign n439 = ~x0 & n74 ;
  assign n440 = ~n438 & n439 ;
  assign n441 = n440 ^ x0 ;
  assign n442 = ~n435 & n441 ;
  assign n443 = ~x7 & ~n442 ;
  assign n379 = ~x1 & n68 ;
  assign n380 = ~n378 & n379 ;
  assign n376 = n66 & n632 ;
  assign n372 = ~x9 & ~n91 ;
  assign n373 = n372 ^ x0 ;
  assign n371 = n118 ^ n24 ;
  assign n374 = n373 ^ n371 ;
  assign n375 = n112 & n374 ;
  assign n377 = n376 ^ n375 ;
  assign n381 = n380 ^ n377 ;
  assign n394 = x8 ^ x6 ;
  assign n395 = n394 ^ n378 ;
  assign n388 = ~x8 & ~n359 ;
  assign n391 = n390 ^ n388 ;
  assign n392 = n390 ^ x0 ;
  assign n393 = ~n391 & ~n392 ;
  assign n396 = n395 ^ n393 ;
  assign n397 = n73 & n396 ;
  assign n382 = ~x6 & n632 ;
  assign n383 = n382 ^ x6 ;
  assign n384 = ~n123 & n383 ;
  assign n385 = x2 & n24 ;
  assign n386 = n385 ^ x9 ;
  assign n387 = n384 & n386 ;
  assign n398 = n397 ^ n387 ;
  assign n399 = ~n381 & ~n398 ;
  assign n400 = ~x5 & ~x7 ;
  assign n401 = ~n13 & ~n25 ;
  assign n402 = ~n400 & n401 ;
  assign n404 = x0 & n73 ;
  assign n405 = n402 & n404 ;
  assign n403 = n402 ^ n400 ;
  assign n406 = n405 ^ n403 ;
  assign n407 = x9 ^ x7 ;
  assign n408 = ~x0 & ~x3 ;
  assign n409 = ~n407 & n408 ;
  assign n421 = ~x9 & n409 ;
  assign n422 = n414 & n421 ;
  assign n423 = n422 ^ n414 ;
  assign n410 = n409 ^ x3 ;
  assign n415 = n414 ^ n410 ;
  assign n424 = n423 ^ n415 ;
  assign n425 = n406 & ~n424 ;
  assign n426 = ~n399 & n425 ;
  assign n444 = n443 ^ n426 ;
  assign n449 = x2 & ~x5 ;
  assign n450 = n449 ^ n390 ;
  assign n451 = ~x1 & n450 ;
  assign n452 = n73 & n449 ;
  assign n453 = ~x0 & ~n11 ;
  assign n454 = ~n318 & n453 ;
  assign n455 = ~n452 & n454 ;
  assign n456 = ~n451 & n455 ;
  assign n457 = ~x6 & x9 ;
  assign n458 = n457 ^ n12 ;
  assign n460 = ~n91 & n167 ;
  assign n461 = ~n385 & n460 ;
  assign n462 = n461 ^ n91 ;
  assign n463 = n83 & ~n462 ;
  assign n464 = n458 & n463 ;
  assign n465 = n464 ^ n462 ;
  assign n466 = ~n456 & n465 ;
  assign n467 = n413 ^ x0 ;
  assign n468 = n449 ^ x9 ;
  assign n471 = ~n413 & n468 ;
  assign n472 = n471 ^ x9 ;
  assign n473 = ~n467 & n472 ;
  assign n474 = x5 & n73 ;
  assign n475 = n474 ^ x9 ;
  assign n476 = ~x0 & n475 ;
  assign n477 = n476 ^ n474 ;
  assign n480 = n450 ^ x8 ;
  assign n481 = ~n477 & ~n480 ;
  assign n482 = n481 ^ x0 ;
  assign n483 = ~x8 & ~n482 ;
  assign n484 = ~n473 & n483 ;
  assign n485 = ~n466 & ~n484 ;
  assign n488 = ~x4 & ~n485 ;
  assign n445 = ~x2 & ~n123 ;
  assign n446 = ~x8 & n12 ;
  assign n447 = n445 & ~n446 ;
  assign n448 = n447 ^ x4 ;
  assign n489 = n488 ^ n448 ;
  assign n490 = x3 & ~n489 ;
  assign n491 = n490 ^ n448 ;
  assign n492 = n444 & ~n491 ;
  assign n493 = ~n205 & n228 ;
  assign n494 = n493 ^ x4 ;
  assign n495 = ~x7 & ~n494 ;
  assign n496 = x0 & x5 ;
  assign n517 = n91 ^ x9 ;
  assign n518 = n517 ^ n372 ;
  assign n519 = n518 ^ n123 ;
  assign n514 = x1 & ~n373 ;
  assign n515 = n514 ^ x0 ;
  assign n516 = n515 ^ n93 ;
  assign n520 = n519 ^ n516 ;
  assign n521 = ~x6 & n520 ;
  assign n522 = ~n432 & ~n521 ;
  assign n502 = n496 ^ x5 ;
  assign n503 = n413 & n502 ;
  assign n498 = x5 ^ x2 ;
  assign n499 = n498 ^ x6 ;
  assign n500 = n11 & ~n499 ;
  assign n497 = n389 ^ n12 ;
  assign n501 = n500 ^ n497 ;
  assign n504 = n503 ^ n501 ;
  assign n505 = ~x3 & ~n91 ;
  assign n506 = n452 & n505 ;
  assign n507 = n506 ^ x3 ;
  assign n508 = n504 & ~n507 ;
  assign n512 = n508 ^ n507 ;
  assign n509 = n62 & n74 ;
  assign n510 = ~x6 & ~n509 ;
  assign n511 = n508 & n510 ;
  assign n513 = n512 ^ n511 ;
  assign n525 = ~n94 & n517 ;
  assign n526 = n525 ^ x9 ;
  assign n527 = n12 & n526 ;
  assign n528 = n527 ^ x5 ;
  assign n529 = ~n513 & ~n528 ;
  assign n530 = n522 & n529 ;
  assign n531 = n530 ^ n513 ;
  assign n532 = n496 & ~n531 ;
  assign n533 = x8 ^ x2 ;
  assign n534 = n533 ^ x9 ;
  assign n535 = n534 ^ x1 ;
  assign n537 = ~n533 & ~n536 ;
  assign n538 = n537 ^ x1 ;
  assign n539 = ~n535 & n538 ;
  assign n540 = n539 ^ x1 ;
  assign n541 = ~x6 & n540 ;
  assign n542 = n541 ^ x1 ;
  assign n543 = n532 & n542 ;
  assign n544 = n543 ^ n531 ;
  assign n545 = n495 & n544 ;
  assign n554 = n11 ^ x5 ;
  assign n555 = ~x1 & ~n554 ;
  assign n556 = n555 ^ n169 ;
  assign n557 = x0 & ~n457 ;
  assign n558 = n556 & n557 ;
  assign n559 = n558 ^ n382 ;
  assign n548 = n382 ^ n378 ;
  assign n549 = ~x0 & ~n548 ;
  assign n550 = n549 ^ n382 ;
  assign n551 = x5 & n550 ;
  assign n552 = n551 ^ n382 ;
  assign n553 = x1 & n552 ;
  assign n560 = n559 ^ n553 ;
  assign n561 = x3 & n560 ;
  assign n562 = ~n11 & ~n76 ;
  assign n563 = n561 & n562 ;
  assign n564 = n563 ^ n561 ;
  assign n565 = n545 & ~n564 ;
  assign n566 = n123 ^ x2 ;
  assign n567 = ~n207 & ~n566 ;
  assign n568 = n400 ^ x7 ;
  assign n569 = n568 ^ n101 ;
  assign n570 = n567 & n569 ;
  assign n571 = x4 ^ x3 ;
  assign n572 = n445 ^ x4 ;
  assign n573 = n571 & ~n572 ;
  assign n574 = n569 & n573 ;
  assign n578 = n166 ^ x5 ;
  assign n644 = ~n319 & n578 ;
  assign n645 = ~n112 & n644 ;
  assign n646 = ~n68 & n645 ;
  assign n647 = ~x4 & n166 ;
  assign n648 = ~n73 & n647 ;
  assign n650 = n66 & n75 ;
  assign n651 = n648 & n650 ;
  assign n649 = n648 ^ x4 ;
  assign n652 = n651 ^ n649 ;
  assign n653 = ~n646 & ~n652 ;
  assign n654 = n653 ^ x5 ;
  assign n660 = x1 & n360 ;
  assign n661 = n428 & n660 ;
  assign n662 = n661 ^ n518 ;
  assign n663 = n661 ^ x1 ;
  assign n664 = ~n438 & n663 ;
  assign n665 = ~n662 & n664 ;
  assign n666 = n665 ^ n663 ;
  assign n674 = n666 ^ x6 ;
  assign n655 = n118 ^ n91 ;
  assign n658 = n389 & n655 ;
  assign n659 = n658 ^ n118 ;
  assign n667 = x0 & ~n86 ;
  assign n668 = ~n62 & n667 ;
  assign n669 = ~n457 & n668 ;
  assign n670 = n669 ^ n667 ;
  assign n671 = n670 ^ n86 ;
  assign n673 = ~n659 & ~n671 ;
  assign n675 = n674 ^ n673 ;
  assign n676 = n653 & ~n675 ;
  assign n677 = n676 ^ x6 ;
  assign n678 = n654 & ~n677 ;
  assign n679 = n678 ^ x5 ;
  assign n680 = x4 & ~n165 ;
  assign n681 = n680 ^ x4 ;
  assign n682 = ~n679 & ~n681 ;
  assign n683 = ~x7 & n682 ;
  assign n604 = ~x2 & n457 ;
  assign n605 = n604 ^ n509 ;
  assign n606 = ~x5 & ~n605 ;
  assign n607 = n606 ^ n509 ;
  assign n608 = ~x7 & ~n607 ;
  assign n609 = n608 ^ x5 ;
  assign n616 = n389 & n400 ;
  assign n617 = n34 & n616 ;
  assign n618 = n617 ^ n34 ;
  assign n610 = n34 ^ x6 ;
  assign n619 = n618 ^ n610 ;
  assign n620 = x0 & ~n619 ;
  assign n621 = ~n609 & n620 ;
  assign n622 = n22 & n167 ;
  assign n18 = x7 & ~x8 ;
  assign n623 = x1 & ~n18 ;
  assign n624 = ~n622 & n623 ;
  assign n625 = x2 & ~x7 ;
  assign n626 = n34 & n625 ;
  assign n627 = n626 ^ x2 ;
  assign n628 = n624 & ~n627 ;
  assign n629 = ~x1 & n171 ;
  assign n630 = x7 ^ x2 ;
  assign n631 = n630 ^ n629 ;
  assign n634 = ~x7 & ~n25 ;
  assign n635 = n634 ^ n632 ;
  assign n636 = n631 & ~n635 ;
  assign n637 = n636 ^ x7 ;
  assign n638 = n629 & ~n637 ;
  assign n639 = ~n628 & ~n638 ;
  assign n640 = n621 & ~n639 ;
  assign n575 = ~n20 & ~n413 ;
  assign n576 = ~x2 & ~n569 ;
  assign n577 = ~n575 & n576 ;
  assign n579 = n578 ^ n446 ;
  assign n580 = n579 ^ n18 ;
  assign n581 = x1 & ~n13 ;
  assign n582 = ~x9 & ~n581 ;
  assign n583 = ~n580 & n582 ;
  assign n584 = n583 ^ x9 ;
  assign n585 = n577 & n584 ;
  assign n586 = x2 & n221 ;
  assign n587 = ~n181 & n586 ;
  assign n588 = n413 & n587 ;
  assign n589 = n588 ^ n586 ;
  assign n590 = n589 ^ x2 ;
  assign n596 = ~n221 & n412 ;
  assign n597 = n168 & n596 ;
  assign n591 = n414 ^ x5 ;
  assign n592 = n591 ^ n581 ;
  assign n593 = ~x7 & ~n74 ;
  assign n594 = n592 & n593 ;
  assign n595 = n594 ^ x7 ;
  assign n598 = n597 ^ n595 ;
  assign n600 = n590 & n598 ;
  assign n601 = ~n585 & ~n600 ;
  assign n641 = n640 ^ n601 ;
  assign n642 = n641 ^ x7 ;
  assign n684 = n683 ^ n642 ;
  assign n687 = n684 ^ n641 ;
  assign n685 = ~x3 & ~x4 ;
  assign n686 = ~n684 & n685 ;
  assign n688 = n687 ^ n686 ;
  assign n691 = n38 ^ n31 ;
  assign n692 = n89 & ~n691 ;
  assign n689 = n78 ^ x3 ;
  assign n690 = n689 ^ n385 ;
  assign n693 = n692 ^ n690 ;
  assign n694 = x1 & ~n693 ;
  assign n695 = n23 & n412 ;
  assign n696 = ~x0 & ~n16 ;
  assign n697 = n696 ^ x3 ;
  assign n698 = n695 & ~n697 ;
  assign n699 = n554 & ~n698 ;
  assign n700 = ~n694 & n699 ;
  assign n706 = n246 ^ n83 ;
  assign n701 = ~x2 & n516 ;
  assign n702 = ~x3 & ~n96 ;
  assign n703 = n701 & n702 ;
  assign n704 = n703 ^ n701 ;
  assign n707 = n88 & n704 ;
  assign n708 = ~n706 & n707 ;
  assign n705 = n704 ^ x2 ;
  assign n709 = n708 ^ n705 ;
  assign n710 = n700 & n709 ;
  assign n753 = n246 ^ n245 ;
  assign n750 = x9 ^ x3 ;
  assign n754 = n753 ^ n750 ;
  assign n751 = n750 ^ x1 ;
  assign n752 = n751 ^ n65 ;
  assign n755 = n754 ^ n752 ;
  assign n739 = n238 ^ n67 ;
  assign n740 = n739 ^ n38 ;
  assign n741 = n740 ^ n245 ;
  assign n742 = n65 ^ x9 ;
  assign n743 = n742 ^ n740 ;
  assign n744 = n740 ^ n65 ;
  assign n745 = n744 ^ x3 ;
  assign n746 = n745 ^ n740 ;
  assign n747 = ~n743 & ~n746 ;
  assign n748 = n747 ^ n740 ;
  assign n749 = n741 & n748 ;
  assign n756 = n755 ^ n749 ;
  assign n757 = n756 ^ n65 ;
  assign n758 = n757 ^ x3 ;
  assign n759 = x8 & n758 ;
  assign n760 = n118 ^ x8 ;
  assign n761 = ~n533 & n760 ;
  assign n765 = n183 & n761 ;
  assign n762 = n349 ^ x3 ;
  assign n766 = n765 ^ n762 ;
  assign n767 = ~x1 & n766 ;
  assign n768 = n767 ^ n349 ;
  assign n769 = n759 & n768 ;
  assign n770 = n769 ^ n768 ;
  assign n771 = ~x6 & ~n770 ;
  assign n711 = n90 ^ x9 ;
  assign n712 = ~n94 & ~n711 ;
  assign n717 = ~n34 & ~n751 ;
  assign n718 = n717 ^ n23 ;
  assign n719 = n718 ^ x9 ;
  assign n720 = n712 & n719 ;
  assign n721 = n720 ^ n717 ;
  assign n722 = n721 ^ ~n34 ;
  assign n723 = n722 ^ x1 ;
  assign n724 = ~x2 & n723 ;
  assign n725 = ~x1 & ~n63 ;
  assign n733 = n238 & n725 ;
  assign n734 = ~n23 & n733 ;
  assign n735 = n734 ^ n23 ;
  assign n726 = n725 ^ x1 ;
  assign n727 = n726 ^ n23 ;
  assign n736 = n735 ^ n727 ;
  assign n737 = ~n37 & n736 ;
  assign n738 = ~n724 & n737 ;
  assign n772 = n771 ^ n738 ;
  assign n773 = ~x4 & ~n772 ;
  assign n774 = n773 ^ x6 ;
  assign n775 = ~x5 & ~n774 ;
  assign n776 = ~n710 & ~n775 ;
  assign n783 = n412 ^ n18 ;
  assign n784 = n783 ^ n698 ;
  assign n782 = n22 & n61 ;
  assign n785 = n784 ^ n782 ;
  assign n778 = n698 ^ x7 ;
  assign n840 = n785 ^ n778 ;
  assign n777 = n698 ^ n412 ;
  assign n779 = n778 ^ n777 ;
  assign n780 = n779 ^ x0 ;
  assign n781 = n780 ^ n778 ;
  assign n856 = n840 ^ n781 ;
  assign n857 = n856 ^ n777 ;
  assign n858 = n857 ^ n698 ;
  assign n802 = n785 ^ n412 ;
  assign n803 = n802 ^ n778 ;
  assign n804 = n803 ^ x0 ;
  assign n805 = n804 ^ n778 ;
  assign n843 = n840 ^ n805 ;
  assign n847 = n858 ^ n843 ;
  assign n821 = n698 & ~n778 ;
  assign n806 = n805 ^ n785 ;
  assign n807 = n806 ^ n777 ;
  assign n808 = n807 ^ n778 ;
  assign n822 = n821 ^ n808 ;
  assign n823 = n822 ^ n779 ;
  assign n824 = n823 ^ x7 ;
  assign n826 = n840 ^ x7 ;
  assign n827 = ~n824 & ~n826 ;
  assign n814 = n785 ^ x7 ;
  assign n829 = n843 ^ n814 ;
  assign n832 = x0 & ~n829 ;
  assign n833 = n827 & n832 ;
  assign n834 = n833 ^ n821 ;
  assign n835 = n847 ^ n834 ;
  assign n836 = n835 ^ n412 ;
  assign n837 = n836 ^ n806 ;
  assign n838 = n837 ^ n814 ;
  assign n848 = n847 ^ n838 ;
  assign n854 = n848 ^ x7 ;
  assign n859 = n858 ^ n854 ;
  assign n860 = ~n680 & ~n859 ;
  assign n861 = ~n776 & n860 ;
  assign n862 = n400 & n681 ;
  assign n863 = ~n13 & ~n632 ;
  assign n864 = n863 ^ n13 ;
  assign n865 = n864 ^ n383 ;
  assign n866 = n474 ^ n120 ;
  assign n868 = n372 ^ n73 ;
  assign n867 = ~n85 & n516 ;
  assign n869 = n868 ^ n867 ;
  assign n870 = ~x2 & n869 ;
  assign n871 = n866 & n870 ;
  assign n872 = n871 ^ x2 ;
  assign n873 = ~x1 & n386 ;
  assign n874 = ~n168 & n873 ;
  assign n875 = n874 ^ n507 ;
  assign n876 = ~n507 & ~n875 ;
  assign n877 = n872 & n876 ;
  assign n878 = n865 & n877 ;
  assign n879 = ~n412 & ~n445 ;
  assign n880 = ~x9 & ~n388 ;
  assign n881 = ~n879 & n880 ;
  assign n882 = x6 ^ x2 ;
  assign n883 = x9 & n882 ;
  assign n884 = ~n92 & n883 ;
  assign n885 = ~n83 & ~n390 ;
  assign n886 = x3 & ~x5 ;
  assign n887 = ~n885 & n886 ;
  assign n888 = ~n884 & n887 ;
  assign n889 = ~n881 & n888 ;
  assign n890 = n38 & n554 ;
  assign n895 = n518 ^ n85 ;
  assign n896 = n895 ^ n867 ;
  assign n892 = n84 ^ n75 ;
  assign n893 = n892 ^ x8 ;
  assign n891 = n24 ^ x1 ;
  assign n894 = n893 ^ n891 ;
  assign n897 = n896 ^ n894 ;
  assign n898 = n890 & n897 ;
  assign n899 = ~n889 & ~n898 ;
  assign n900 = ~n878 & n899 ;
  assign n901 = x7 & n863 ;
  assign n907 = ~x2 & ~n73 ;
  assign n902 = n63 & ~n123 ;
  assign n908 = n907 ^ n902 ;
  assign n909 = n901 & n908 ;
  assign n910 = n909 ^ x7 ;
  assign n911 = ~x4 & ~n910 ;
  assign n912 = ~n900 & n911 ;
  assign n913 = ~n862 & ~n912 ;
  assign n914 = n228 ^ x4 ;
  assign n915 = n500 ^ n499 ;
  assign n917 = ~n13 & n867 ;
  assign n916 = ~n521 & n528 ;
  assign n918 = n917 ^ n916 ;
  assign n919 = n915 & n918 ;
  assign n920 = x3 & ~x7 ;
  assign n921 = ~n919 & n920 ;
  assign n922 = n432 & ~n894 ;
  assign n925 = n62 & n75 ;
  assign n926 = ~x3 & n925 ;
  assign n923 = n493 ^ x3 ;
  assign n927 = n926 ^ n923 ;
  assign n930 = ~x2 & n515 ;
  assign n931 = n930 ^ n902 ;
  assign n932 = ~x7 & ~n931 ;
  assign n933 = n932 ^ n902 ;
  assign n934 = ~n927 & ~n933 ;
  assign n935 = n934 ^ n927 ;
  assign n936 = n13 & n113 ;
  assign n937 = ~n935 & n936 ;
  assign n940 = n922 & n937 ;
  assign n938 = n937 ^ n935 ;
  assign n941 = n940 ^ n938 ;
  assign n942 = ~n921 & n941 ;
  assign n943 = ~n914 & ~n942 ;
  assign n945 = n14 & n867 ;
  assign n946 = n945 ^ n165 ;
  assign n947 = ~x4 & n946 ;
  assign n948 = n947 ^ n165 ;
  assign n949 = n100 & n948 ;
  assign y0 = n212 ;
  assign y1 = n370 ;
  assign y2 = n492 ;
  assign y3 = n565 ;
  assign y4 = n570 ;
  assign y5 = n574 ;
  assign y6 = n688 ;
  assign y7 = ~n861 ;
  assign y8 = n913 ;
  assign y9 = n943 ;
  assign y10 = n949 ;
endmodule
