module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n127 , n128 , n129 , n133 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n146 , n147 , n148 , n151 , n152 , n153 , n154 , n155 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 ;
  assign n35 = x5 ^ x3 ;
  assign n28 = x1 & x4 ;
  assign n26 = x3 ^ x2 ;
  assign n24 = x3 ^ x1 ;
  assign n25 = n24 ^ x0 ;
  assign n27 = n26 ^ n25 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~x5 & n29 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = ~x6 & n31 ;
  assign n23 = x4 ^ x2 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = ~x7 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = ~x8 & n36 ;
  assign n22 = x6 ^ x4 ;
  assign n38 = n37 ^ n22 ;
  assign n39 = ~x9 & n38 ;
  assign n20 = x6 ^ x5 ;
  assign n13 = x6 & x7 ;
  assign n15 = ~x8 & ~n13 ;
  assign n14 = n13 ^ x8 ;
  assign n16 = n15 ^ n14 ;
  assign n18 = ~x9 & ~n16 ;
  assign n12 = x7 ^ x6 ;
  assign n17 = n16 ^ n12 ;
  assign n19 = n18 ^ n17 ;
  assign n21 = n20 ^ n19 ;
  assign n40 = n39 ^ n21 ;
  assign n41 = ~x10 & ~n40 ;
  assign n42 = n41 ^ n19 ;
  assign n44 = ~x7 & ~x8 ;
  assign n59 = ~x2 & ~x3 ;
  assign n60 = n59 ^ n26 ;
  assign n54 = x1 & x2 ;
  assign n47 = ~x0 & n28 ;
  assign n45 = x2 & x4 ;
  assign n46 = n45 ^ x1 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ x3 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = x5 & n55 ;
  assign n57 = n56 ^ n48 ;
  assign n58 = n57 ^ x4 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = n61 ^ n57 ;
  assign n65 = ~x9 & n62 ;
  assign n66 = n65 ^ n57 ;
  assign n67 = x6 & ~n66 ;
  assign n68 = n67 ^ n57 ;
  assign n69 = n44 & ~n68 ;
  assign n82 = ~x5 & ~x6 ;
  assign n83 = n82 ^ n20 ;
  assign n84 = n83 ^ x7 ;
  assign n71 = x4 & x5 ;
  assign n72 = n71 ^ x6 ;
  assign n85 = n84 ^ n72 ;
  assign n70 = x9 ^ x8 ;
  assign n74 = x3 & x4 ;
  assign n73 = n72 ^ x5 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = n75 ^ n72 ;
  assign n79 = x7 & ~n76 ;
  assign n80 = n79 ^ n72 ;
  assign n81 = ~n70 & ~n80 ;
  assign n86 = n85 ^ n81 ;
  assign n87 = ~x9 & ~n86 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = ~n69 & ~n88 ;
  assign n43 = ~n15 & ~n18 ;
  assign n90 = n89 ^ n43 ;
  assign n91 = x10 & n90 ;
  assign n92 = n91 ^ n89 ;
  assign n178 = x5 & n13 ;
  assign n177 = n16 ^ x8 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = ~x10 & n179 ;
  assign n181 = n180 ^ n16 ;
  assign n109 = n72 ^ n12 ;
  assign n93 = x8 ^ x7 ;
  assign n100 = n93 ^ n71 ;
  assign n110 = n100 ^ n12 ;
  assign n111 = n109 & ~n110 ;
  assign n101 = n100 ^ x3 ;
  assign n104 = n100 ^ n72 ;
  assign n102 = n93 ^ n72 ;
  assign n103 = n102 ^ x3 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n101 & ~n105 ;
  assign n112 = n111 ^ n106 ;
  assign n113 = n112 ^ n104 ;
  assign n114 = n111 ^ n102 ;
  assign n115 = n114 ^ n104 ;
  assign n116 = ~n113 & n115 ;
  assign n117 = n72 & n116 ;
  assign n118 = n117 ^ n111 ;
  assign n119 = n118 ^ n109 ;
  assign n127 = x6 & ~n60 ;
  assign n128 = n71 & n127 ;
  assign n129 = ~x7 & ~n128 ;
  assign n133 = x6 ^ x2 ;
  assign n136 = ~x4 & ~n133 ;
  assign n137 = n136 ^ x5 ;
  assign n138 = x6 ^ x3 ;
  assign n139 = n136 ^ n133 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = n140 ^ x6 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = n142 ^ x5 ;
  assign n144 = n129 & n143 ;
  assign n151 = x3 & ~x5 ;
  assign n152 = n151 ^ x6 ;
  assign n153 = x4 & ~n152 ;
  assign n146 = x3 & ~x6 ;
  assign n147 = n45 & n146 ;
  assign n148 = n147 ^ n20 ;
  assign n154 = n153 ^ n148 ;
  assign n155 = x3 ^ x0 ;
  assign n158 = x5 & n155 ;
  assign n159 = n158 ^ x0 ;
  assign n160 = x1 & n159 ;
  assign n161 = n154 & ~n160 ;
  assign n162 = n161 ^ n147 ;
  assign n163 = n144 & ~n162 ;
  assign n164 = ~x8 & ~n163 ;
  assign n172 = ~x3 & n164 ;
  assign n173 = n13 & n172 ;
  assign n174 = n173 ^ n13 ;
  assign n165 = n164 ^ x8 ;
  assign n166 = n165 ^ n13 ;
  assign n175 = n174 ^ n166 ;
  assign n176 = ~n119 & n175 ;
  assign n182 = n181 ^ n176 ;
  assign n183 = n182 ^ n16 ;
  assign n184 = ~x10 & ~n183 ;
  assign n185 = n184 ^ n16 ;
  assign n187 = n181 ^ x9 ;
  assign n186 = n181 ^ x10 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = ~n185 & ~n188 ;
  assign n190 = n189 ^ n187 ;
  assign n191 = ~x9 & ~x10 ;
  assign n192 = ~x3 & n191 ;
  assign n196 = ~x2 & ~n16 ;
  assign n197 = n71 & n196 ;
  assign n193 = x4 & n82 ;
  assign n194 = n193 ^ n82 ;
  assign n195 = n44 & n194 ;
  assign n198 = n197 ^ n195 ;
  assign n199 = n192 & n198 ;
  assign n200 = n13 & ~n59 ;
  assign n201 = n71 & n200 ;
  assign n203 = n193 ^ x6 ;
  assign n202 = n147 & n160 ;
  assign n204 = n203 ^ n202 ;
  assign n224 = n44 & ~n128 ;
  assign n206 = n204 & n224 ;
  assign n207 = n206 ^ x8 ;
  assign n208 = ~x9 & n207 ;
  assign n209 = ~n201 & n208 ;
  assign n210 = ~x10 & ~n70 ;
  assign n211 = n178 & n210 ;
  assign n219 = ~x8 & n211 ;
  assign n220 = ~n74 & n219 ;
  assign n221 = n220 ^ n74 ;
  assign n212 = n211 ^ x10 ;
  assign n213 = n212 ^ n74 ;
  assign n222 = n221 ^ n213 ;
  assign n223 = ~n209 & ~n222 ;
  assign n225 = n191 & n224 ;
  assign n227 = n82 & ~n202 ;
  assign n228 = n225 & n227 ;
  assign n226 = n225 ^ n191 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = x8 & n201 ;
  assign n231 = n229 & n230 ;
  assign n232 = n231 ^ n229 ;
  assign y0 = ~n42 ;
  assign y1 = n92 ;
  assign y2 = ~n190 ;
  assign y3 = ~n199 ;
  assign y4 = ~n223 ;
  assign y5 = ~n232 ;
  assign y6 = ~n225 ;
endmodule
