module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
output y0;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, y0;
assign n_0 = x0 & ~x32;
assign n_1 = x34 ^ x2;
assign n_2 = x34 ^ x33;
assign n_3 = x34 ^ x1;
assign n_4 = x35 ^ x3;
assign n_5 = x37 ^ x5;
assign n_6 = x6 & ~x38;
assign n_7 = x38 ^ x6;
assign n_8 = x7 & ~x39;
assign n_9 = x39 ^ x7;
assign n_10 = x41 ^ x9;
assign n_11 = ~x9 & x41;
assign n_12 = x10 & ~x42;
assign n_13 = x42 ^ x10;
assign n_14 = x11 & ~x43;
assign n_15 = x43 ^ x11;
assign n_16 = x44 ^ x12;
assign n_17 = x12 & ~x44;
assign n_18 = x45 ^ x13;
assign n_19 = x13 ^ ~x45;
assign n_20 = x46 ^ x14;
assign n_21 = x14 & ~x46;
assign n_22 = x47 ^ x15;
assign n_23 = x15 ^ ~x47;
assign n_24 = x48 ^ x16;
assign n_25 = x16 & ~x48;
assign n_26 = x49 ^ x17;
assign n_27 = x17 & ~x49;
assign n_28 = x50 ^ x18;
assign n_29 = x18 & ~x50;
assign n_30 = x51 ^ x19;
assign n_31 = x19 & ~x51;
assign n_32 = x52 ^ x20;
assign n_33 = x20 & ~x52;
assign n_34 = x53 ^ x21;
assign n_35 = x21 & ~x53;
assign n_36 = x54 ^ x22;
assign n_37 = x22 & ~x54;
assign n_38 = x55 ^ x23;
assign n_39 = x23 & ~x55;
assign n_40 = x57 ^ x25;
assign n_41 = x26 & ~x58;
assign n_42 = x58 ^ x26;
assign n_43 = x27 & ~x59;
assign n_44 = x59 ^ x27;
assign n_45 = x28 & ~x60;
assign n_46 = x60 ^ x28;
assign n_47 = x29 & ~x61;
assign n_48 = x61 ^ x29;
assign n_49 = x30 & ~x62;
assign n_50 = x31 & ~x63;
assign n_51 = x63 ^ x31;
assign n_52 = n_0 ^ x34;
assign n_53 = n_2 ^ n_3;
assign n_54 = x37 & ~n_5;
assign n_55 = ~n_6 & ~n_8;
assign n_56 = n_7 ^ n_8;
assign n_57 = n_10 ^ n_11;
assign n_58 = n_11 ^ x42;
assign n_59 = ~n_12 & ~n_14;
assign n_60 = n_16 ^ n_17;
assign n_61 = ~n_17 & n_19;
assign n_62 = n_20 ^ n_21;
assign n_63 = ~n_21 & n_23;
assign n_64 = n_24 ^ n_25;
assign n_65 = n_26 ^ n_27;
assign n_66 = n_28 ^ n_29;
assign n_67 = ~n_27 & ~n_31;
assign n_68 = n_32 ^ n_33;
assign n_69 = n_34 ^ n_35;
assign n_70 = n_36 ^ n_37;
assign n_71 = ~n_35 & ~n_39;
assign n_72 = x57 & ~n_40;
assign n_73 = ~n_41 & ~n_43;
assign n_74 = n_42 ^ n_43;
assign n_75 = n_46 ^ n_45;
assign n_76 = ~n_45 & ~n_47;
assign n_77 = n_49 ^ x30;
assign n_78 = ~n_49 & ~n_50;
assign n_79 = n_52 ^ n_3;
assign n_80 = n_54 ^ x5;
assign n_81 = n_54 ^ x6;
assign n_82 = x40 & ~n_57;
assign n_83 = ~x8 & ~n_57;
assign n_84 = ~n_13 & n_58;
assign n_85 = n_60 ^ x45;
assign n_86 = n_62 ^ x47;
assign n_87 = ~n_64 & ~n_65;
assign n_88 = n_66 ^ x51;
assign n_89 = ~n_29 & n_67;
assign n_90 = ~n_68 & ~n_69;
assign n_91 = n_70 ^ x55;
assign n_92 = ~n_37 & n_71;
assign n_93 = n_72 ^ x25;
assign n_94 = n_72 ^ x26;
assign n_95 = n_75 ^ x61;
assign n_96 = n_77 ^ x62;
assign n_97 = n_76 & n_78;
assign n_98 = ~n_53 & n_79;
assign n_99 = n_55 & ~n_80;
assign n_100 = n_81 ^ x37;
assign n_101 = n_82 & n_59;
assign n_102 = n_59 & n_83;
assign n_103 = n_84 ^ x42;
assign n_104 = ~n_18 & ~n_85;
assign n_105 = ~n_22 & ~n_86;
assign n_106 = ~n_30 & ~n_88;
assign n_107 = ~n_87 & n_89;
assign n_108 = ~n_38 & ~n_91;
assign n_109 = ~n_90 & n_92;
assign n_110 = ~n_33 & n_92;
assign n_111 = n_73 & ~n_93;
assign n_112 = n_94 ^ x57;
assign n_113 = ~n_48 & ~n_95;
assign n_114 = n_98 ^ n_3;
assign n_115 = ~x4 & n_99;
assign n_116 = x36 & n_99;
assign n_117 = n_56 & ~n_100;
assign n_118 = ~x8 & n_101;
assign n_119 = n_102 ^ n_101;
assign n_120 = n_103 ^ x43;
assign n_121 = n_104 ^ x13;
assign n_122 = n_105 ^ x15;
assign n_123 = n_106 ^ x19;
assign n_124 = n_108 ^ x23;
assign n_125 = x56 & n_111;
assign n_126 = ~x24 & n_111;
assign n_127 = n_74 & ~n_112;
assign n_128 = n_113 ^ x29;
assign n_129 = ~n_1 & n_114;
assign n_130 = n_115 ^ n_116;
assign n_131 = ~x4 & n_116;
assign n_132 = n_117 ^ n_54;
assign n_133 = ~n_15 & n_120;
assign n_134 = n_123 & ~n_107;
assign n_135 = n_124 & ~n_109;
assign n_136 = ~n_125 & ~n_126;
assign n_137 = n_127 ^ n_72;
assign n_138 = n_128 ^ x63;
assign n_139 = n_129 ^ x2;
assign n_140 = n_132 ^ x37;
assign n_141 = n_133 ^ x43;
assign n_142 = n_110 & ~n_134;
assign n_143 = n_97 & ~n_136;
assign n_144 = n_136 ^ n_125;
assign n_145 = n_137 ^ x57;
assign n_146 = n_138 ^ x63;
assign n_147 = n_139 ^ x35;
assign n_148 = n_140 ^ x39;
assign n_149 = ~n_118 & ~n_141;
assign n_150 = n_135 & ~n_142;
assign n_151 = n_144 ^ n_126;
assign n_152 = n_145 ^ x59;
assign n_153 = ~n_49 & ~n_146;
assign n_154 = ~n_4 & n_147;
assign n_155 = ~n_9 & n_148;
assign n_156 = n_143 & ~n_150;
assign n_157 = ~n_44 & n_152;
assign n_158 = n_153 ^ x62;
assign n_159 = n_153 ^ x63;
assign n_160 = n_154 ^ x3;
assign n_161 = n_155 ^ x39;
assign n_162 = n_157 ^ x59;
assign n_163 = ~n_158 & n_96;
assign n_164 = n_130 & ~n_160;
assign n_165 = ~n_131 & ~n_161;
assign n_166 = ~n_162 & n_151;
assign n_167 = n_163 ^ n_77;
assign n_168 = ~n_164 & n_165;
assign n_169 = n_97 & ~n_166;
assign n_170 = n_167 ^ n_159;
assign n_171 = n_119 & ~n_168;
assign n_172 = ~n_156 & ~n_169;
assign n_173 = n_170 ^ x62;
assign n_174 = n_149 & ~n_171;
assign n_175 = ~n_51 & ~n_173;
assign n_176 = n_174 ^ n_61;
assign n_177 = n_63 ^ n_174;
assign n_178 = n_175 ^ x31;
assign n_179 = ~n_174 & ~n_177;
assign n_180 = n_179 ^ n_174;
assign n_181 = ~n_176 & ~n_180;
assign n_182 = n_181 ^ n_179;
assign n_183 = n_182 ^ n_174;
assign n_184 = n_183 ^ n_63;
assign n_185 = n_121 & ~n_184;
assign n_186 = n_185 ^ n_63;
assign n_187 = n_122 & ~n_186;
assign n_188 = ~n_25 & ~n_187;
assign n_189 = n_89 & n_188;
assign n_190 = n_110 & n_189;
assign n_191 = n_143 & n_190;
assign n_192 = n_178 & ~n_191;
assign n_193 = n_172 & n_192;
assign y0 = ~n_193;
endmodule