module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n131 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n516 , n518 , n519 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n600 , n601 , n602 , n603 , n604 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 ;
  assign n131 = ~x2 & ~x3 ;
  assign n134 = x1 & n131 ;
  assign n135 = n134 ^ x3 ;
  assign n136 = ~x6 & ~x7 ;
  assign n137 = n136 ^ x7 ;
  assign n138 = n137 ^ x5 ;
  assign n139 = n136 & n138 ;
  assign n140 = ~x4 & n139 ;
  assign n141 = n135 & n140 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = n142 ^ n137 ;
  assign n144 = ~x10 & ~x11 ;
  assign n456 = ~x8 & ~x9 ;
  assign n457 = n144 & n456 ;
  assign n149 = n143 & n457 ;
  assign n145 = n144 ^ x11 ;
  assign n146 = n145 ^ x9 ;
  assign n147 = n144 & n146 ;
  assign n150 = n149 ^ n147 ;
  assign n151 = n150 ^ n145 ;
  assign n152 = ~x14 & ~x15 ;
  assign n451 = ~x12 & ~x13 ;
  assign n452 = n152 & n451 ;
  assign n157 = n151 & n452 ;
  assign n153 = n152 ^ x15 ;
  assign n154 = n153 ^ x13 ;
  assign n155 = n152 & n154 ;
  assign n158 = n157 ^ n155 ;
  assign n159 = n158 ^ n153 ;
  assign n160 = ~x18 & ~x19 ;
  assign n448 = ~x16 & ~x17 ;
  assign n449 = n160 & n448 ;
  assign n165 = n159 & n449 ;
  assign n161 = n160 ^ x19 ;
  assign n162 = n161 ^ x17 ;
  assign n163 = n160 & n162 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = n166 ^ n161 ;
  assign n168 = ~x22 & ~x23 ;
  assign n434 = ~x20 & ~x21 ;
  assign n435 = n168 & n434 ;
  assign n173 = n167 & n435 ;
  assign n169 = n168 ^ x23 ;
  assign n170 = n169 ^ x21 ;
  assign n171 = n168 & n170 ;
  assign n174 = n173 ^ n171 ;
  assign n175 = n174 ^ n169 ;
  assign n176 = ~x26 & ~x27 ;
  assign n431 = ~x24 & ~x25 ;
  assign n432 = n176 & n431 ;
  assign n181 = n175 & n432 ;
  assign n177 = n176 ^ x27 ;
  assign n178 = n177 ^ x25 ;
  assign n179 = n176 & n178 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ n177 ;
  assign n184 = ~x30 & ~x31 ;
  assign n429 = ~x28 & ~x29 ;
  assign n430 = n184 & n429 ;
  assign n189 = n183 & n430 ;
  assign n185 = n184 ^ x31 ;
  assign n186 = n185 ^ x29 ;
  assign n187 = n184 & n186 ;
  assign n190 = n189 ^ n187 ;
  assign n191 = n190 ^ n185 ;
  assign n192 = ~x34 & ~x35 ;
  assign n491 = ~x32 & ~x33 ;
  assign n492 = n192 & n491 ;
  assign n197 = n191 & n492 ;
  assign n193 = n192 ^ x35 ;
  assign n194 = n193 ^ x33 ;
  assign n195 = n192 & n194 ;
  assign n198 = n197 ^ n195 ;
  assign n199 = n198 ^ n193 ;
  assign n200 = ~x38 & ~x39 ;
  assign n489 = ~x36 & ~x37 ;
  assign n490 = n200 & n489 ;
  assign n205 = n199 & n490 ;
  assign n201 = n200 ^ x39 ;
  assign n202 = n201 ^ x37 ;
  assign n203 = n200 & n202 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = n206 ^ n201 ;
  assign n208 = ~x42 & ~x43 ;
  assign n486 = ~x40 & ~x41 ;
  assign n487 = n208 & n486 ;
  assign n213 = n207 & n487 ;
  assign n209 = n208 ^ x43 ;
  assign n210 = n209 ^ x41 ;
  assign n211 = n208 & n210 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ n209 ;
  assign n216 = ~x46 & ~x47 ;
  assign n426 = ~x44 & ~x45 ;
  assign n427 = n216 & n426 ;
  assign n221 = n215 & n427 ;
  assign n217 = n216 ^ x47 ;
  assign n218 = n217 ^ x45 ;
  assign n219 = n216 & n218 ;
  assign n222 = n221 ^ n219 ;
  assign n223 = n222 ^ n217 ;
  assign n224 = ~x50 & ~x51 ;
  assign n420 = ~x48 & ~x49 ;
  assign n421 = n224 & n420 ;
  assign n229 = n223 & n421 ;
  assign n225 = n224 ^ x51 ;
  assign n226 = n225 ^ x49 ;
  assign n227 = n224 & n226 ;
  assign n230 = n229 ^ n227 ;
  assign n231 = n230 ^ n225 ;
  assign n232 = ~x54 & ~x55 ;
  assign n412 = ~x52 & ~x53 ;
  assign n419 = n232 & n412 ;
  assign n237 = n231 & n419 ;
  assign n233 = n232 ^ x55 ;
  assign n234 = n233 ^ x53 ;
  assign n235 = n232 & n234 ;
  assign n238 = n237 ^ n235 ;
  assign n239 = n238 ^ n233 ;
  assign n240 = ~x58 & ~x59 ;
  assign n416 = ~x56 & ~x57 ;
  assign n417 = n240 & n416 ;
  assign n245 = n239 & n417 ;
  assign n241 = n240 ^ x59 ;
  assign n242 = n241 ^ x57 ;
  assign n243 = n240 & n242 ;
  assign n246 = n245 ^ n243 ;
  assign n247 = n246 ^ n241 ;
  assign n248 = ~x62 & ~x63 ;
  assign n409 = ~x60 & ~x61 ;
  assign n410 = n248 & n409 ;
  assign n253 = n247 & n410 ;
  assign n249 = n248 ^ x63 ;
  assign n250 = n249 ^ x61 ;
  assign n251 = n248 & n250 ;
  assign n254 = n253 ^ n251 ;
  assign n255 = n254 ^ n249 ;
  assign n256 = ~x66 & ~x67 ;
  assign n482 = ~x64 & ~x65 ;
  assign n483 = n256 & n482 ;
  assign n261 = n255 & n483 ;
  assign n257 = n256 ^ x67 ;
  assign n258 = n257 ^ x65 ;
  assign n259 = n256 & n258 ;
  assign n262 = n261 ^ n259 ;
  assign n263 = n262 ^ n257 ;
  assign n264 = ~x70 & ~x71 ;
  assign n407 = ~x68 & ~x69 ;
  assign n481 = n264 & n407 ;
  assign n269 = n263 & n481 ;
  assign n265 = n264 ^ x71 ;
  assign n266 = n265 ^ x69 ;
  assign n267 = n264 & n266 ;
  assign n270 = n269 ^ n267 ;
  assign n271 = n270 ^ n265 ;
  assign n272 = ~x74 & ~x75 ;
  assign n478 = ~x72 & ~x73 ;
  assign n479 = n272 & n478 ;
  assign n277 = n271 & n479 ;
  assign n273 = n272 ^ x75 ;
  assign n274 = n273 ^ x73 ;
  assign n275 = n272 & n274 ;
  assign n278 = n277 ^ n275 ;
  assign n279 = n278 ^ n273 ;
  assign n280 = ~x78 & ~x79 ;
  assign n405 = ~x76 & ~x77 ;
  assign n477 = n280 & n405 ;
  assign n285 = n279 & n477 ;
  assign n281 = n280 ^ x79 ;
  assign n282 = n281 ^ x77 ;
  assign n283 = n280 & n282 ;
  assign n286 = n285 ^ n283 ;
  assign n287 = n286 ^ n281 ;
  assign n288 = ~x82 & ~x83 ;
  assign n463 = ~x80 & ~x81 ;
  assign n464 = n288 & n463 ;
  assign n293 = n287 & n464 ;
  assign n289 = n288 ^ x83 ;
  assign n290 = n289 ^ x81 ;
  assign n291 = n288 & n290 ;
  assign n294 = n293 ^ n291 ;
  assign n295 = n294 ^ n289 ;
  assign n296 = ~x86 & ~x87 ;
  assign n459 = ~x84 & ~x85 ;
  assign n460 = n296 & n459 ;
  assign n301 = n295 & n460 ;
  assign n297 = n296 ^ x87 ;
  assign n298 = n297 ^ x85 ;
  assign n299 = n296 & n298 ;
  assign n302 = n301 ^ n299 ;
  assign n303 = n302 ^ n297 ;
  assign n304 = ~x90 & ~x91 ;
  assign n403 = ~x88 & ~x89 ;
  assign n461 = n304 & n403 ;
  assign n309 = n303 & n461 ;
  assign n305 = n304 ^ x91 ;
  assign n306 = n305 ^ x89 ;
  assign n307 = n304 & n306 ;
  assign n310 = n309 ^ n307 ;
  assign n311 = n310 ^ n305 ;
  assign n312 = ~x94 & ~x95 ;
  assign n400 = ~x92 & ~x93 ;
  assign n402 = n312 & n400 ;
  assign n317 = n311 & n402 ;
  assign n313 = n312 ^ x95 ;
  assign n314 = n313 ^ x93 ;
  assign n315 = n312 & n314 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n318 ^ n313 ;
  assign n320 = ~x98 & ~x99 ;
  assign n472 = ~x96 & ~x97 ;
  assign n473 = n320 & n472 ;
  assign n325 = n319 & n473 ;
  assign n321 = n320 ^ x99 ;
  assign n322 = n321 ^ x97 ;
  assign n323 = n320 & n322 ;
  assign n326 = n325 ^ n323 ;
  assign n327 = n326 ^ n321 ;
  assign n328 = ~x102 & ~x103 ;
  assign n398 = ~x100 & ~x101 ;
  assign n471 = n328 & n398 ;
  assign n333 = n327 & n471 ;
  assign n329 = n328 ^ x103 ;
  assign n330 = n329 ^ x101 ;
  assign n331 = n328 & n330 ;
  assign n334 = n333 ^ n331 ;
  assign n335 = n334 ^ n329 ;
  assign n336 = ~x106 & ~x107 ;
  assign n468 = ~x104 & ~x105 ;
  assign n469 = n336 & n468 ;
  assign n341 = n335 & n469 ;
  assign n337 = n336 ^ x107 ;
  assign n338 = n337 ^ x105 ;
  assign n339 = n336 & n338 ;
  assign n342 = n341 ^ n339 ;
  assign n343 = n342 ^ n337 ;
  assign n344 = ~x110 & ~x111 ;
  assign n396 = ~x108 & ~x109 ;
  assign n467 = n344 & n396 ;
  assign n349 = n343 & n467 ;
  assign n345 = n344 ^ x111 ;
  assign n346 = n345 ^ x109 ;
  assign n347 = n344 & n346 ;
  assign n350 = n349 ^ n347 ;
  assign n351 = n350 ^ n345 ;
  assign n352 = ~x114 & ~x115 ;
  assign n392 = ~x112 & ~x113 ;
  assign n393 = n352 & n392 ;
  assign n357 = n351 & n393 ;
  assign n353 = n352 ^ x115 ;
  assign n354 = n353 ^ x113 ;
  assign n355 = n352 & n354 ;
  assign n358 = n357 ^ n355 ;
  assign n359 = n358 ^ n353 ;
  assign n360 = ~x118 & ~x119 ;
  assign n388 = ~x116 & ~x117 ;
  assign n389 = n360 & n388 ;
  assign n365 = n359 & n389 ;
  assign n361 = n360 ^ x119 ;
  assign n362 = n361 ^ x117 ;
  assign n363 = n360 & n362 ;
  assign n366 = n365 ^ n363 ;
  assign n367 = n366 ^ n361 ;
  assign n368 = ~x122 & ~x123 ;
  assign n386 = ~x120 & ~x121 ;
  assign n387 = n368 & n386 ;
  assign n373 = n367 & n387 ;
  assign n369 = n368 ^ x123 ;
  assign n370 = n369 ^ x121 ;
  assign n371 = n368 & n370 ;
  assign n374 = n373 ^ n371 ;
  assign n375 = n374 ^ n369 ;
  assign n376 = ~x126 & ~x127 ;
  assign n384 = ~x124 & ~x125 ;
  assign n385 = n376 & n384 ;
  assign n381 = n375 & n385 ;
  assign n377 = n376 ^ x127 ;
  assign n378 = n377 ^ x125 ;
  assign n379 = n376 & n378 ;
  assign n382 = n381 ^ n379 ;
  assign n383 = n382 ^ n377 ;
  assign n593 = n385 ^ n376 ;
  assign n390 = n387 & n389 ;
  assign n391 = n385 & n390 ;
  assign n397 = n396 ^ n336 ;
  assign n399 = n398 ^ n320 ;
  assign n401 = n400 ^ n304 ;
  assign n404 = n402 & n403 ;
  assign n462 = n402 & n461 ;
  assign n465 = n462 & n464 ;
  assign n466 = n460 & n465 ;
  assign n556 = ~n288 & n296 ;
  assign n557 = n459 & n556 ;
  assign n406 = n405 ^ n272 ;
  assign n408 = n407 ^ n256 ;
  assign n480 = n477 & n479 ;
  assign n484 = n481 & n483 ;
  assign n485 = n480 & n484 ;
  assign n411 = n409 ^ n240 ;
  assign n413 = ~n224 & n232 ;
  assign n414 = n412 & n413 ;
  assign n415 = n414 ^ n232 ;
  assign n534 = n415 ^ n411 ;
  assign n418 = n410 & n417 ;
  assign n422 = n419 & n421 ;
  assign n423 = n418 & n422 ;
  assign n428 = n426 ^ n208 ;
  assign n522 = n208 ^ n200 ;
  assign n523 = n522 ^ n426 ;
  assign n488 = n427 & n487 ;
  assign n493 = n490 & n492 ;
  assign n494 = n488 & n493 ;
  assign n495 = n423 & n494 ;
  assign n433 = n430 & n432 ;
  assign n436 = n433 & n435 ;
  assign n450 = n436 & n449 ;
  assign n454 = n451 ^ n144 ;
  assign n455 = n452 & ~n454 ;
  assign n458 = n452 & n457 ;
  assign n470 = n467 & n469 ;
  assign n474 = n471 & n473 ;
  assign n475 = n470 & n474 ;
  assign n476 = n466 & n475 ;
  assign n500 = ~n450 & n495 ;
  assign n501 = n500 ^ n423 ;
  assign n502 = n485 & ~n501 ;
  assign n503 = n476 & ~n502 ;
  assign n504 = n503 ^ n475 ;
  assign n505 = ~n458 & ~n504 ;
  assign n506 = n136 & ~n505 ;
  assign n510 = n506 ^ n505 ;
  assign n507 = ~x4 & ~x5 ;
  assign n508 = ~n131 & n507 ;
  assign n509 = n506 & n508 ;
  assign n511 = n510 ^ n509 ;
  assign n512 = n455 & n511 ;
  assign n453 = n452 ^ n152 ;
  assign n513 = n512 ^ n453 ;
  assign n514 = n450 & ~n513 ;
  assign n437 = ~n160 & n436 ;
  assign n438 = n437 ^ n184 ;
  assign n439 = n430 & n438 ;
  assign n444 = ~n168 & n432 ;
  assign n445 = n444 ^ n176 ;
  assign n446 = n439 & ~n445 ;
  assign n447 = n446 ^ n438 ;
  assign n516 = n514 ^ n447 ;
  assign n518 = n495 & ~n516 ;
  assign n519 = n518 ^ n192 ;
  assign n521 = n490 & ~n519 ;
  assign n524 = n523 ^ n521 ;
  assign n525 = ~n428 & ~n524 ;
  assign n526 = n487 ^ n216 ;
  assign n527 = n526 ^ n426 ;
  assign n528 = n525 & n527 ;
  assign n529 = n528 ^ n428 ;
  assign n530 = n427 & n529 ;
  assign n424 = n232 ^ n216 ;
  assign n425 = n424 ^ n423 ;
  assign n531 = n530 ^ n425 ;
  assign n532 = n423 & ~n531 ;
  assign n535 = n534 ^ n532 ;
  assign n536 = ~n411 & ~n535 ;
  assign n537 = n417 ^ n248 ;
  assign n538 = n537 ^ n409 ;
  assign n539 = n536 & n538 ;
  assign n540 = n539 ^ n411 ;
  assign n541 = n410 & n540 ;
  assign n542 = n541 ^ n248 ;
  assign n544 = n485 & ~n542 ;
  assign n545 = n544 ^ n481 ;
  assign n546 = ~n408 & n545 ;
  assign n547 = n546 ^ n481 ;
  assign n548 = n547 ^ n264 ;
  assign n549 = n477 & n478 ;
  assign n550 = ~n548 & n549 ;
  assign n551 = n550 ^ n477 ;
  assign n552 = ~n406 & n551 ;
  assign n553 = n552 ^ n477 ;
  assign n554 = n553 ^ n280 ;
  assign n555 = n554 ^ n466 ;
  assign n558 = n557 ^ n555 ;
  assign n561 = n466 & n558 ;
  assign n559 = n557 ^ n296 ;
  assign n562 = n561 ^ n559 ;
  assign n563 = n404 & ~n562 ;
  assign n564 = n563 ^ n402 ;
  assign n565 = ~n401 & n564 ;
  assign n566 = n565 ^ n402 ;
  assign n567 = n566 ^ n312 ;
  assign n568 = n471 & n472 ;
  assign n569 = ~n567 & n568 ;
  assign n570 = n569 ^ n471 ;
  assign n571 = ~n399 & n570 ;
  assign n572 = n571 ^ n471 ;
  assign n573 = n572 ^ n328 ;
  assign n574 = n467 & n468 ;
  assign n575 = ~n573 & n574 ;
  assign n576 = n575 ^ n467 ;
  assign n577 = ~n397 & n576 ;
  assign n578 = n577 ^ n467 ;
  assign n579 = n578 ^ n344 ;
  assign n580 = n352 & ~n579 ;
  assign n394 = n390 & n393 ;
  assign n595 = n385 & n387 ;
  assign n654 = n394 & n595 ;
  assign n581 = n580 & n654 ;
  assign n582 = n581 ^ n352 ;
  assign n583 = n391 & ~n582 ;
  assign n584 = n583 ^ n385 ;
  assign n590 = ~n360 & n387 ;
  assign n585 = n384 ^ n368 ;
  assign n591 = n590 ^ n585 ;
  assign n592 = n584 & ~n591 ;
  assign n594 = n593 ^ n592 ;
  assign n625 = n462 ^ n402 ;
  assign n596 = n449 & n452 ;
  assign n600 = n506 & n507 ;
  assign n601 = n600 ^ n505 ;
  assign n602 = n596 & n601 ;
  assign n603 = n602 ^ n449 ;
  assign n609 = n436 & ~n603 ;
  assign n604 = n433 ^ n430 ;
  assign n610 = n609 ^ n604 ;
  assign n611 = n493 & ~n610 ;
  assign n612 = n611 ^ n490 ;
  assign n613 = n488 & ~n612 ;
  assign n614 = n613 ^ n427 ;
  assign n615 = n422 & ~n614 ;
  assign n616 = n615 ^ n419 ;
  assign n617 = n418 & ~n616 ;
  assign n618 = n617 ^ n410 ;
  assign n619 = n484 & ~n618 ;
  assign n620 = n619 ^ n481 ;
  assign n621 = n480 & ~n620 ;
  assign n622 = n621 ^ n477 ;
  assign n623 = n465 & ~n622 ;
  assign n624 = n623 ^ n460 ;
  assign n626 = n625 ^ n624 ;
  assign n627 = n462 ^ n460 ;
  assign n628 = n627 ^ n625 ;
  assign n629 = n626 & ~n628 ;
  assign n630 = n629 ^ n625 ;
  assign n631 = n474 & ~n630 ;
  assign n632 = n631 ^ n471 ;
  assign n633 = n470 & ~n632 ;
  assign n634 = n633 ^ n467 ;
  assign n636 = n394 & ~n634 ;
  assign n637 = n636 ^ n389 ;
  assign n638 = n595 & ~n637 ;
  assign n639 = n638 ^ n385 ;
  assign n640 = n466 & n485 ;
  assign n642 = n433 & n495 ;
  assign n643 = ~n505 & n642 ;
  assign n644 = n643 ^ n495 ;
  assign n645 = n644 ^ n418 ;
  assign n641 = n423 & ~n488 ;
  assign n646 = n645 ^ n641 ;
  assign n647 = n466 & ~n480 ;
  assign n648 = n647 ^ n462 ;
  assign n649 = ~n646 & n648 ;
  assign n650 = n640 & n649 ;
  assign n651 = n650 ^ n648 ;
  assign n652 = n475 & ~n651 ;
  assign n653 = n652 ^ n470 ;
  assign n655 = ~n653 & n654 ;
  assign n656 = n655 ^ n595 ;
  assign n657 = ~n504 & n654 ;
  assign n658 = n475 & n654 ;
  assign n659 = n640 & n658 ;
  assign n660 = ~n495 & n659 ;
  assign n661 = n660 ^ n658 ;
  assign n662 = ~x0 & ~x1 ;
  assign n663 = n495 & n662 ;
  assign n664 = n659 & n663 ;
  assign n665 = ~n502 & n664 ;
  assign n666 = n511 & n665 ;
  assign n667 = ~n644 & n666 ;
  assign n668 = ~n603 & n667 ;
  assign y0 = n383 ;
  assign y1 = ~n594 ;
  assign y2 = ~n639 ;
  assign y3 = ~n656 ;
  assign y4 = ~n657 ;
  assign y5 = ~n661 ;
  assign y6 = ~n659 ;
  assign y7 = ~n668 ;
endmodule
