module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n212 , n213 , n214 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n255 , n256 , n257 , n258 , n262 , n263 , n264 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n303 , n304 , n305 , n306 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n396 , n397 , n398 , n399 , n400 , n401 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n471 , n472 , n475 , n476 , n477 , n478 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n497 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n520 , n521 , n522 , n523 , n524 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n541 , n542 , n543 , n544 , n545 , n546 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n653 , n654 , n655 , n656 , n657 , n658 , n663 , n664 , n665 , n666 , n668 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n689 , n692 , n693 , n694 , n695 , n696 , n697 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n810 , n811 , n812 , n813 , n814 , n815 , n818 , n819 , n820 , n821 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n847 , n848 , n849 , n850 , n853 , n854 , n855 , n856 , n859 , n860 , n861 , n862 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n874 , n875 , n876 , n877 , n880 , n881 , n882 , n883 , n886 , n887 , n888 , n889 , n892 , n893 , n894 , n895 , n898 , n899 , n900 , n901 , n904 , n905 , n906 , n907 , n910 , n911 , n912 , n913 , n916 , n917 , n918 , n919 , n922 , n923 , n924 , n925 , n928 , n929 , n930 , n931 , n934 , n935 , n936 , n937 , n940 , n941 , n942 , n943 , n944 , n947 , n948 , n949 , n950 , n953 , n954 , n955 , n956 , n959 , n960 , n961 , n962 , n965 , n966 , n967 , n968 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n1000 , n1001 , n1002 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1013 , n1014 , n1015 , n1016 , n1019 , n1020 , n1021 , n1022 , n1023 , n1026 , n1027 , n1028 , n1029 , n1032 , n1033 , n1034 , n1035 , n1038 , n1039 , n1040 , n1041 , n1044 , n1045 , n1046 , n1047 , n1050 , n1051 , n1052 , n1053 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1065 , n1066 , n1067 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1079 , n1080 , n1081 , n1082 , n1083 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1094 , n1095 , n1096 , n1097 , n1100 , n1101 , n1102 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1167 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1210 , n1211 , n1212 , n1213 , n1214 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1263 , n1264 , n1265 , n1266 , n1267 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1295 , n1296 , n1297 , n1298 , n1301 , n1302 , n1303 , n1304 , n1307 , n1308 , n1309 , n1310 , n1313 , n1314 , n1315 , n1316 , n1317 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 ;
  assign n148 = ~x3 & ~x129 ;
  assign n149 = x54 & ~x56 ;
  assign n155 = ~x9 & ~x11 ;
  assign n150 = ~x5 & ~x22 ;
  assign n156 = n155 ^ n150 ;
  assign n157 = n149 & n156 ;
  assign n183 = ~x11 & n150 ;
  assign n158 = ~x17 & x54 ;
  assign n164 = ~x4 & ~x9 ;
  assign n165 = ~x12 & n164 ;
  assign n192 = ~x6 & n165 ;
  assign n184 = ~x18 & ~x19 ;
  assign n185 = x16 & n184 ;
  assign n186 = n185 ^ n184 ;
  assign n198 = x10 ^ x8 ;
  assign n160 = ~x8 & ~x10 ;
  assign n193 = x21 ^ x14 ;
  assign n194 = x14 ^ x13 ;
  assign n195 = n193 & n194 ;
  assign n196 = n195 ^ x14 ;
  assign n197 = n160 & ~n196 ;
  assign n199 = n198 ^ n197 ;
  assign n161 = ~x14 & ~x21 ;
  assign n200 = ~x13 & n161 ;
  assign n201 = n199 & n200 ;
  assign n162 = n160 & n161 ;
  assign n163 = ~x13 & n162 ;
  assign n203 = n201 ^ n163 ;
  assign n204 = n203 ^ n197 ;
  assign n205 = x7 & n204 ;
  assign n202 = n201 ^ n197 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n186 & n206 ;
  assign n208 = n192 & n207 ;
  assign n212 = n158 & n208 ;
  assign n213 = n183 & n212 ;
  assign n166 = ~x7 & n165 ;
  assign n167 = n163 & n166 ;
  assign n168 = x7 ^ x6 ;
  assign n169 = n168 ^ x9 ;
  assign n170 = n169 ^ x12 ;
  assign n171 = n170 ^ x13 ;
  assign n172 = x13 ^ x12 ;
  assign n173 = x9 ^ x7 ;
  assign n174 = n173 ^ x12 ;
  assign n175 = n172 & n174 ;
  assign n176 = n175 ^ x12 ;
  assign n177 = n171 & n176 ;
  assign n178 = n177 ^ n171 ;
  assign n179 = x7 & x9 ;
  assign n180 = n178 & n179 ;
  assign n181 = n180 ^ n178 ;
  assign n182 = n167 & ~n181 ;
  assign n187 = n183 & n186 ;
  assign n188 = n182 & n187 ;
  assign n189 = n158 & ~n188 ;
  assign n159 = n158 ^ x54 ;
  assign n190 = n189 ^ n159 ;
  assign n191 = ~x0 & ~n190 ;
  assign n214 = n213 ^ n191 ;
  assign n216 = ~n157 & ~n214 ;
  assign n217 = n148 & ~n216 ;
  assign n218 = ~x1 & n148 ;
  assign n234 = ~n189 & n218 ;
  assign n219 = ~x4 & n162 ;
  assign n220 = x54 & n148 ;
  assign n221 = x17 & n220 ;
  assign n222 = n221 ^ n220 ;
  assign n223 = n186 & n222 ;
  assign n224 = ~x11 & ~x22 ;
  assign n225 = n223 & n224 ;
  assign n226 = n219 & n225 ;
  assign n227 = ~x5 & n226 ;
  assign n228 = ~n181 & n227 ;
  assign n229 = n228 ^ n226 ;
  assign n231 = ~x5 & n229 ;
  assign n230 = n182 & n229 ;
  assign n232 = n231 ^ n230 ;
  assign n235 = n234 ^ n232 ;
  assign n243 = ~x15 & ~x20 ;
  assign n241 = ~x24 & ~x45 ;
  assign n242 = ~x49 & n241 ;
  assign n237 = ~x43 & ~x47 ;
  assign n238 = ~x41 & ~x46 ;
  assign n239 = ~x48 & n238 ;
  assign n240 = n237 & n239 ;
  assign n248 = ~x38 & ~x50 ;
  assign n251 = ~x42 & ~x44 ;
  assign n252 = ~x40 & n251 ;
  assign n262 = n248 & n252 ;
  assign n263 = n240 & n262 ;
  assign n264 = n242 & n263 ;
  assign n267 = n243 & n264 ;
  assign n268 = x82 & n267 ;
  assign n269 = n268 ^ x82 ;
  assign n236 = x122 & x127 ;
  assign n257 = ~x82 & ~n236 ;
  assign n258 = n257 ^ x82 ;
  assign n270 = n269 ^ n258 ;
  assign n271 = x2 & ~n270 ;
  assign n272 = ~x129 & ~n271 ;
  assign n275 = n272 ^ x129 ;
  assign n418 = x82 & n263 ;
  assign n419 = ~x45 & n418 ;
  assign n704 = n419 ^ x82 ;
  assign n244 = ~x2 & n243 ;
  assign n245 = n242 & n244 ;
  assign n705 = x82 & ~n245 ;
  assign n706 = ~n704 & ~n705 ;
  assign n255 = n236 & n706 ;
  assign n256 = n706 ^ n255 ;
  assign n273 = ~x65 & n272 ;
  assign n274 = n256 & n273 ;
  assign n276 = n275 ^ n274 ;
  assign n277 = x0 & ~x113 ;
  assign n278 = x123 & ~x129 ;
  assign n279 = n278 ^ x129 ;
  assign n280 = ~x61 & ~x118 ;
  assign n281 = ~x17 & n188 ;
  assign n282 = ~x129 & ~n281 ;
  assign n283 = n280 & n282 ;
  assign n284 = ~n279 & ~n283 ;
  assign n285 = n277 & n284 ;
  assign n286 = n285 ^ n283 ;
  assign n290 = n220 ^ n148 ;
  assign n291 = x4 & n290 ;
  assign n287 = n183 & n222 ;
  assign n288 = n208 & n287 ;
  assign n289 = x10 & n288 ;
  assign n292 = n291 ^ n289 ;
  assign n301 = x5 & n290 ;
  assign n293 = ~x29 & ~x59 ;
  assign n294 = n182 & n287 ;
  assign n295 = ~x16 & n294 ;
  assign n296 = n184 & n295 ;
  assign n297 = n293 & n296 ;
  assign n298 = ~x25 & ~x28 ;
  assign n299 = n298 ^ x25 ;
  assign n300 = n297 & ~n299 ;
  assign n303 = n301 ^ n300 ;
  assign n306 = x6 & n290 ;
  assign n304 = n298 ^ x28 ;
  assign n305 = n297 & ~n304 ;
  assign n308 = n306 ^ n305 ;
  assign n310 = x7 & n290 ;
  assign n309 = x8 & n288 ;
  assign n311 = n310 ^ n309 ;
  assign n313 = x8 & n290 ;
  assign n312 = x21 & n288 ;
  assign n314 = n313 ^ n312 ;
  assign n319 = x9 & n290 ;
  assign n315 = ~x5 & n182 ;
  assign n316 = n223 & n315 ;
  assign n317 = x11 & ~x22 ;
  assign n318 = n316 & n317 ;
  assign n320 = n319 ^ n318 ;
  assign n322 = x10 & n290 ;
  assign n321 = x14 & n288 ;
  assign n323 = n322 ^ n321 ;
  assign n328 = x22 & n316 ;
  assign n329 = n328 ^ n290 ;
  assign n330 = ~x11 & n329 ;
  assign n331 = n330 ^ n290 ;
  assign n333 = ~x18 & n295 ;
  assign n334 = n333 ^ n295 ;
  assign n335 = ~x19 & n334 ;
  assign n332 = x12 & n290 ;
  assign n336 = n335 ^ n332 ;
  assign n343 = x13 & n290 ;
  assign n338 = x29 & x54 ;
  assign n339 = ~x59 & n298 ;
  assign n340 = n338 & n339 ;
  assign n341 = n281 & n340 ;
  assign n342 = n148 & n341 ;
  assign n344 = n343 ^ n342 ;
  assign n346 = x14 & n290 ;
  assign n345 = x13 & n288 ;
  assign n347 = n346 ^ n345 ;
  assign n348 = n264 ^ x15 ;
  assign n349 = n348 ^ x70 ;
  assign n350 = n349 ^ n264 ;
  assign n353 = ~n236 & ~n350 ;
  assign n354 = n353 ^ n264 ;
  assign n355 = ~x82 & n354 ;
  assign n356 = n355 ^ n348 ;
  assign n357 = ~x129 & n244 ;
  assign n365 = ~x70 & n357 ;
  assign n366 = ~n236 & n365 ;
  assign n367 = n366 ^ n236 ;
  assign n358 = n357 ^ x129 ;
  assign n359 = n358 ^ n236 ;
  assign n368 = n367 ^ n359 ;
  assign n369 = n356 & ~n368 ;
  assign n371 = x16 & n290 ;
  assign n370 = x6 & n232 ;
  assign n372 = n371 ^ n370 ;
  assign n374 = ~x29 & n298 ;
  assign n375 = n188 & n374 ;
  assign n376 = x59 & n222 ;
  assign n377 = n375 & n376 ;
  assign n373 = x17 & n290 ;
  assign n378 = n377 ^ n373 ;
  assign n380 = n185 & n294 ;
  assign n379 = x18 & n290 ;
  assign n381 = n380 ^ n379 ;
  assign n383 = x19 & n290 ;
  assign n382 = n188 & n221 ;
  assign n384 = n383 ^ n382 ;
  assign n385 = x71 ^ x20 ;
  assign n386 = ~n236 & ~n385 ;
  assign n387 = n386 ^ x20 ;
  assign n388 = x82 & ~n387 ;
  assign n396 = ~n386 & n388 ;
  assign n397 = ~x2 & n396 ;
  assign n398 = n397 ^ x2 ;
  assign n389 = n388 ^ n387 ;
  assign n390 = n389 ^ x2 ;
  assign n399 = n398 ^ n390 ;
  assign n400 = ~x129 & n399 ;
  assign n401 = x82 & n400 ;
  assign n406 = ~x15 & n264 ;
  assign n407 = n406 ^ x20 ;
  assign n408 = n401 & ~n407 ;
  assign n409 = n408 ^ n400 ;
  assign n411 = x19 & n333 ;
  assign n410 = x21 & n290 ;
  assign n412 = n411 ^ n410 ;
  assign n413 = x22 & n290 ;
  assign n414 = n413 ^ n230 ;
  assign n415 = ~x23 & x55 ;
  assign n416 = x61 & ~x129 ;
  assign n417 = ~n415 & n416 ;
  assign n420 = n419 ^ n255 ;
  assign n421 = n420 ^ x82 ;
  assign n422 = n421 ^ n419 ;
  assign n425 = ~x24 & n422 ;
  assign n426 = n425 ^ n419 ;
  assign n427 = ~x129 & ~n426 ;
  assign n428 = x63 & n256 ;
  assign n429 = n427 & n428 ;
  assign n430 = n429 ^ n427 ;
  assign n431 = ~x26 & x27 ;
  assign n432 = n431 ^ x26 ;
  assign n449 = x58 ^ x53 ;
  assign n439 = ~x53 & ~x58 ;
  assign n450 = n449 ^ n439 ;
  assign n451 = ~x85 & n450 ;
  assign n452 = n451 ^ n439 ;
  assign n453 = ~n432 & n452 ;
  assign n443 = ~x85 & n439 ;
  assign n447 = ~n432 & n443 ;
  assign n444 = n432 ^ x27 ;
  assign n445 = n444 ^ x26 ;
  assign n446 = n443 & ~n445 ;
  assign n448 = n447 ^ n446 ;
  assign n454 = n453 ^ n448 ;
  assign n455 = ~x116 & n454 ;
  assign n456 = x27 & x116 ;
  assign n457 = ~x39 & ~x51 ;
  assign n458 = ~x52 & n457 ;
  assign n459 = n148 & ~n458 ;
  assign n460 = n456 & n459 ;
  assign n461 = n460 ^ n148 ;
  assign n462 = ~n455 & n461 ;
  assign n471 = x26 & x116 ;
  assign n472 = n458 & n471 ;
  assign n475 = n446 & ~n472 ;
  assign n463 = ~x95 & ~x100 ;
  assign n464 = ~x97 & ~x110 ;
  assign n465 = n463 & n464 ;
  assign n466 = n465 ^ x110 ;
  assign n467 = n447 & n466 ;
  assign n468 = n467 ^ n447 ;
  assign n476 = n475 ^ n468 ;
  assign n477 = n462 & ~n476 ;
  assign n478 = n477 ^ n461 ;
  assign n434 = ~x96 & ~x110 ;
  assign n435 = n434 ^ x116 ;
  assign n436 = ~x85 & n435 ;
  assign n437 = n436 ^ x116 ;
  assign n438 = x100 & n437 ;
  assign n440 = n148 & ~n432 ;
  assign n441 = n439 & n440 ;
  assign n442 = n438 & n441 ;
  assign n482 = n478 ^ n442 ;
  assign n433 = x116 & n432 ;
  assign n480 = ~x25 & n478 ;
  assign n481 = ~n433 & n480 ;
  assign n483 = n482 ^ n481 ;
  assign n484 = n148 & n444 ;
  assign n485 = x116 & n458 ;
  assign n486 = n443 & n485 ;
  assign n487 = n486 ^ n443 ;
  assign n488 = n484 & n487 ;
  assign n489 = n488 ^ n442 ;
  assign n490 = ~x100 & n437 ;
  assign n491 = ~n432 & n439 ;
  assign n492 = n490 & n491 ;
  assign n497 = x85 & x116 ;
  assign n500 = ~x95 & ~n497 ;
  assign n493 = n492 ^ n431 ;
  assign n494 = n493 ^ n487 ;
  assign n501 = n500 ^ n494 ;
  assign n502 = n492 & n501 ;
  assign n503 = n502 ^ n494 ;
  assign n505 = n503 ^ n431 ;
  assign n506 = n503 ^ n492 ;
  assign n507 = ~n505 & ~n506 ;
  assign n504 = n503 ^ n487 ;
  assign n509 = n507 ^ n504 ;
  assign n510 = n509 ^ n487 ;
  assign n511 = n148 & ~n510 ;
  assign n512 = ~x27 & n443 ;
  assign n513 = ~x26 & x28 ;
  assign n514 = n466 & n513 ;
  assign n515 = n514 ^ n472 ;
  assign n516 = n512 & n515 ;
  assign n517 = n511 ^ x28 ;
  assign n520 = ~n455 & n517 ;
  assign n521 = n520 ^ x28 ;
  assign n522 = ~n516 & ~n521 ;
  assign n523 = n148 & ~n522 ;
  assign n524 = n440 & n451 ;
  assign n528 = n434 & n463 ;
  assign n529 = n528 ^ x116 ;
  assign n530 = ~x58 & n529 ;
  assign n531 = n530 ^ x116 ;
  assign n532 = x97 & n531 ;
  assign n533 = n532 ^ x116 ;
  assign n534 = ~x53 & ~n533 ;
  assign n535 = n534 ^ x116 ;
  assign n536 = n524 & ~n535 ;
  assign n537 = n536 ^ x29 ;
  assign n538 = n467 ^ n455 ;
  assign n541 = n537 & ~n538 ;
  assign n542 = n541 ^ x29 ;
  assign n543 = n148 & n542 ;
  assign n545 = x88 ^ x60 ;
  assign n544 = x88 ^ x30 ;
  assign n546 = n545 ^ n544 ;
  assign n549 = ~x109 & n546 ;
  assign n550 = n549 ^ n545 ;
  assign n551 = ~x106 & n550 ;
  assign n552 = n551 ^ x88 ;
  assign n553 = ~x129 & n552 ;
  assign n555 = x89 ^ x31 ;
  assign n554 = x89 ^ x30 ;
  assign n556 = n555 ^ n554 ;
  assign n559 = x109 & n556 ;
  assign n560 = n559 ^ n555 ;
  assign n561 = ~x106 & n560 ;
  assign n562 = n561 ^ x89 ;
  assign n563 = ~x129 & n562 ;
  assign n565 = x99 ^ x32 ;
  assign n564 = x99 ^ x31 ;
  assign n566 = n565 ^ n564 ;
  assign n569 = x109 & n566 ;
  assign n570 = n569 ^ n565 ;
  assign n571 = ~x106 & n570 ;
  assign n572 = n571 ^ x99 ;
  assign n573 = ~x129 & n572 ;
  assign n575 = x90 ^ x33 ;
  assign n574 = x90 ^ x32 ;
  assign n576 = n575 ^ n574 ;
  assign n579 = x109 & n576 ;
  assign n580 = n579 ^ n575 ;
  assign n581 = ~x106 & n580 ;
  assign n582 = n581 ^ x90 ;
  assign n583 = ~x129 & n582 ;
  assign n585 = x91 ^ x34 ;
  assign n584 = x91 ^ x33 ;
  assign n586 = n585 ^ n584 ;
  assign n589 = x109 & n586 ;
  assign n590 = n589 ^ n585 ;
  assign n591 = ~x106 & n590 ;
  assign n592 = n591 ^ x91 ;
  assign n593 = ~x129 & n592 ;
  assign n595 = x92 ^ x35 ;
  assign n594 = x92 ^ x34 ;
  assign n596 = n595 ^ n594 ;
  assign n599 = x109 & n596 ;
  assign n600 = n599 ^ n595 ;
  assign n601 = ~x106 & n600 ;
  assign n602 = n601 ^ x92 ;
  assign n603 = ~x129 & n602 ;
  assign n605 = x98 ^ x36 ;
  assign n604 = x98 ^ x35 ;
  assign n606 = n605 ^ n604 ;
  assign n609 = x109 & n606 ;
  assign n610 = n609 ^ n605 ;
  assign n611 = ~x106 & n610 ;
  assign n612 = n611 ^ x98 ;
  assign n613 = ~x129 & n612 ;
  assign n615 = x93 ^ x37 ;
  assign n614 = x93 ^ x36 ;
  assign n616 = n615 ^ n614 ;
  assign n619 = x109 & n616 ;
  assign n620 = n619 ^ n615 ;
  assign n621 = ~x106 & n620 ;
  assign n622 = n621 ^ x93 ;
  assign n623 = ~x129 & n622 ;
  assign n624 = n252 ^ x38 ;
  assign n246 = n240 & n245 ;
  assign n247 = x82 & ~n246 ;
  assign n249 = x82 & ~n248 ;
  assign n250 = ~n247 & ~n249 ;
  assign n625 = ~x129 & n250 ;
  assign n626 = x74 ^ x38 ;
  assign n629 = ~n236 & ~n626 ;
  assign n630 = n629 ^ x38 ;
  assign n631 = n625 & ~n630 ;
  assign n632 = n631 ^ x129 ;
  assign n633 = x82 & ~n632 ;
  assign n634 = ~n624 & n633 ;
  assign n635 = n634 ^ n632 ;
  assign n636 = ~x106 & ~x129 ;
  assign n637 = ~x51 & x109 ;
  assign n642 = ~x52 & n637 ;
  assign n643 = n642 ^ x39 ;
  assign n644 = n636 & ~n643 ;
  assign n645 = n644 ^ x129 ;
  assign n253 = x82 & ~n252 ;
  assign n648 = n706 ^ n253 ;
  assign n646 = ~x73 & ~n236 ;
  assign n647 = n646 & n706 ;
  assign n649 = n648 ^ n647 ;
  assign n650 = x40 & n649 ;
  assign n653 = x82 & ~n251 ;
  assign n654 = n653 ^ n258 ;
  assign n655 = n650 & ~n654 ;
  assign n656 = n655 ^ n649 ;
  assign n657 = ~x129 & ~n656 ;
  assign n668 = x76 ^ x41 ;
  assign n671 = ~n236 & ~n668 ;
  assign n672 = n671 ^ x41 ;
  assign n658 = x82 & ~x129 ;
  assign n717 = n262 ^ x46 ;
  assign n718 = n658 & ~n717 ;
  assign n719 = n718 ^ x129 ;
  assign n720 = n706 & ~n719 ;
  assign n673 = ~n672 & n720 ;
  assign n663 = ~x46 & n262 ;
  assign n664 = n663 ^ x41 ;
  assign n665 = n658 & ~n664 ;
  assign n666 = n665 ^ x129 ;
  assign n674 = n673 ^ n666 ;
  assign n681 = x42 & ~n257 ;
  assign n675 = ~x72 & ~n236 ;
  assign n679 = n675 & n706 ;
  assign n676 = x44 & x82 ;
  assign n677 = n706 ^ n676 ;
  assign n680 = n679 ^ n677 ;
  assign n682 = n681 ^ n680 ;
  assign n683 = ~x129 & ~n682 ;
  assign n689 = x77 ^ x43 ;
  assign n692 = ~n236 & ~n689 ;
  assign n693 = n692 ^ x43 ;
  assign n694 = ~n693 & n720 ;
  assign n684 = n238 & n262 ;
  assign n685 = n684 ^ x43 ;
  assign n686 = n658 & ~n685 ;
  assign n687 = n686 ^ x129 ;
  assign n695 = n694 ^ n687 ;
  assign n696 = ~x129 & ~n676 ;
  assign n697 = x67 ^ x44 ;
  assign n700 = n236 & ~n697 ;
  assign n701 = n700 ^ x67 ;
  assign n702 = n701 & n706 ;
  assign n703 = n696 & ~n702 ;
  assign n707 = ~x68 & n706 ;
  assign n708 = ~n236 & n707 ;
  assign n709 = n708 ^ n706 ;
  assign n710 = n709 ^ n704 ;
  assign n711 = ~n257 & ~n418 ;
  assign n712 = x45 & n711 ;
  assign n713 = n712 ^ x129 ;
  assign n714 = ~x129 & ~n713 ;
  assign n715 = n710 & n714 ;
  assign n716 = n715 ^ x129 ;
  assign n721 = x75 ^ x46 ;
  assign n724 = ~n236 & ~n721 ;
  assign n725 = n724 ^ x46 ;
  assign n726 = n720 & ~n725 ;
  assign n727 = n726 ^ n719 ;
  assign n728 = ~x43 & n684 ;
  assign n729 = n728 ^ x47 ;
  assign n730 = ~x129 & ~n247 ;
  assign n731 = x64 ^ x47 ;
  assign n734 = ~n236 & ~n731 ;
  assign n735 = n734 ^ x47 ;
  assign n736 = n730 & ~n735 ;
  assign n737 = n736 ^ x129 ;
  assign n738 = x82 & ~n737 ;
  assign n739 = ~n729 & n738 ;
  assign n740 = n739 ^ n737 ;
  assign n741 = ~x47 & n728 ;
  assign n742 = n741 ^ x48 ;
  assign n743 = x62 ^ x48 ;
  assign n744 = ~n236 & ~n743 ;
  assign n745 = n744 ^ x48 ;
  assign n746 = ~x129 & ~n705 ;
  assign n747 = ~n745 & n746 ;
  assign n752 = ~n744 & n747 ;
  assign n753 = n752 ^ x129 ;
  assign n754 = n742 & ~n753 ;
  assign n748 = n747 ^ x129 ;
  assign n755 = n754 ^ n748 ;
  assign n756 = x82 & ~n755 ;
  assign n757 = n756 ^ n748 ;
  assign n764 = x49 & ~n257 ;
  assign n759 = n706 ^ x24 ;
  assign n762 = n419 & ~n759 ;
  assign n758 = ~x69 & ~n236 ;
  assign n761 = n706 & n758 ;
  assign n763 = n762 ^ n761 ;
  assign n765 = n764 ^ n763 ;
  assign n766 = ~x129 & n765 ;
  assign n767 = n258 ^ n249 ;
  assign n768 = ~n253 & n767 ;
  assign n769 = n246 & n768 ;
  assign n777 = ~x66 & n769 ;
  assign n778 = ~n236 & n777 ;
  assign n779 = n778 ^ n236 ;
  assign n770 = n769 ^ n768 ;
  assign n771 = n770 ^ n236 ;
  assign n780 = n779 ^ n771 ;
  assign n781 = ~x50 & ~n780 ;
  assign n782 = n249 & n252 ;
  assign n783 = ~x38 & n782 ;
  assign n784 = n783 ^ x129 ;
  assign n785 = ~x129 & ~n784 ;
  assign n786 = ~n781 & n785 ;
  assign n787 = x66 & n257 ;
  assign n788 = n786 & n787 ;
  assign n789 = n788 ^ n786 ;
  assign n790 = x109 ^ x51 ;
  assign n791 = n636 & ~n790 ;
  assign n792 = n791 ^ x129 ;
  assign n793 = n637 ^ x52 ;
  assign n794 = n636 & ~n793 ;
  assign n795 = n794 ^ x129 ;
  assign n796 = ~x129 & ~n256 ;
  assign n797 = ~x114 & ~x122 ;
  assign n798 = n797 ^ x122 ;
  assign n799 = ~n279 & ~n798 ;
  assign n800 = n453 ^ n446 ;
  assign n801 = n148 & n800 ;
  assign n803 = x58 & x116 ;
  assign n802 = n471 ^ x58 ;
  assign n804 = n803 ^ n802 ;
  assign n805 = n471 ^ x94 ;
  assign n806 = n805 ^ n803 ;
  assign n807 = n806 ^ x94 ;
  assign n810 = ~x37 & ~n807 ;
  assign n811 = n810 ^ x94 ;
  assign n812 = ~n804 & ~n811 ;
  assign n813 = n812 ^ x94 ;
  assign n814 = n801 & n813 ;
  assign n815 = x60 ^ x57 ;
  assign n818 = ~n803 & n815 ;
  assign n819 = n818 ^ x60 ;
  assign n820 = n801 & n819 ;
  assign n826 = n433 & n458 ;
  assign n821 = n803 ^ x58 ;
  assign n827 = n826 ^ n821 ;
  assign n828 = n801 & n827 ;
  assign n830 = x96 & n468 ;
  assign n829 = x59 & n538 ;
  assign n831 = n830 ^ n829 ;
  assign n832 = n148 & n831 ;
  assign n833 = ~x117 & ~x122 ;
  assign n834 = x123 ^ x60 ;
  assign n835 = n833 & n834 ;
  assign n836 = n835 ^ x60 ;
  assign n837 = n278 & n797 ;
  assign n838 = x140 ^ x62 ;
  assign n839 = x132 & x133 ;
  assign n840 = x131 & n839 ;
  assign n841 = ~x138 & n840 ;
  assign n842 = x136 & x137 ;
  assign n843 = n842 ^ x136 ;
  assign n844 = n841 & n843 ;
  assign n847 = ~n838 & n844 ;
  assign n848 = n847 ^ x62 ;
  assign n849 = ~x129 & n848 ;
  assign n850 = x142 ^ x63 ;
  assign n853 = n844 & ~n850 ;
  assign n854 = n853 ^ x63 ;
  assign n855 = ~x129 & n854 ;
  assign n856 = x139 ^ x64 ;
  assign n859 = n844 & ~n856 ;
  assign n860 = n859 ^ x64 ;
  assign n861 = ~x129 & n860 ;
  assign n862 = x146 ^ x65 ;
  assign n865 = n844 & ~n862 ;
  assign n866 = n865 ^ x65 ;
  assign n867 = ~x129 & n866 ;
  assign n868 = x143 ^ x66 ;
  assign n869 = n842 ^ x137 ;
  assign n870 = n869 ^ x136 ;
  assign n871 = n841 & ~n870 ;
  assign n874 = ~n868 & n871 ;
  assign n875 = n874 ^ x66 ;
  assign n876 = ~x129 & n875 ;
  assign n877 = x139 ^ x67 ;
  assign n880 = n871 & ~n877 ;
  assign n881 = n880 ^ x67 ;
  assign n882 = ~x129 & n881 ;
  assign n883 = x141 ^ x68 ;
  assign n886 = n844 & ~n883 ;
  assign n887 = n886 ^ x68 ;
  assign n888 = ~x129 & n887 ;
  assign n889 = x143 ^ x69 ;
  assign n892 = n844 & ~n889 ;
  assign n893 = n892 ^ x69 ;
  assign n894 = ~x129 & n893 ;
  assign n895 = x144 ^ x70 ;
  assign n898 = n844 & ~n895 ;
  assign n899 = n898 ^ x70 ;
  assign n900 = ~x129 & n899 ;
  assign n901 = x145 ^ x71 ;
  assign n904 = n844 & ~n901 ;
  assign n905 = n904 ^ x71 ;
  assign n906 = ~x129 & n905 ;
  assign n907 = x140 ^ x72 ;
  assign n910 = n871 & ~n907 ;
  assign n911 = n910 ^ x72 ;
  assign n912 = ~x129 & n911 ;
  assign n913 = x141 ^ x73 ;
  assign n916 = n871 & ~n913 ;
  assign n917 = n916 ^ x73 ;
  assign n918 = ~x129 & n917 ;
  assign n919 = x142 ^ x74 ;
  assign n922 = n871 & ~n919 ;
  assign n923 = n922 ^ x74 ;
  assign n924 = ~x129 & n923 ;
  assign n925 = x144 ^ x75 ;
  assign n928 = n871 & ~n925 ;
  assign n929 = n928 ^ x75 ;
  assign n930 = ~x129 & n929 ;
  assign n931 = x145 ^ x76 ;
  assign n934 = n871 & ~n931 ;
  assign n935 = n934 ^ x76 ;
  assign n936 = ~x129 & n935 ;
  assign n937 = x146 ^ x77 ;
  assign n940 = n871 & ~n937 ;
  assign n941 = n940 ^ x77 ;
  assign n942 = ~x129 & n941 ;
  assign n943 = x142 ^ x78 ;
  assign n944 = n841 & n869 ;
  assign n947 = n943 & n944 ;
  assign n948 = n947 ^ x78 ;
  assign n949 = ~x129 & n948 ;
  assign n950 = x143 ^ x79 ;
  assign n953 = n944 & n950 ;
  assign n954 = n953 ^ x79 ;
  assign n955 = ~x129 & n954 ;
  assign n956 = x144 ^ x80 ;
  assign n959 = n944 & n956 ;
  assign n960 = n959 ^ x80 ;
  assign n961 = ~x129 & n960 ;
  assign n962 = x145 ^ x81 ;
  assign n965 = n944 & n962 ;
  assign n966 = n965 ^ x81 ;
  assign n967 = ~x129 & n966 ;
  assign n968 = x146 ^ x82 ;
  assign n971 = n944 & n968 ;
  assign n972 = n971 ^ x82 ;
  assign n973 = ~x129 & n972 ;
  assign n991 = x89 & ~x137 ;
  assign n983 = x138 ^ x136 ;
  assign n984 = x89 ^ x62 ;
  assign n985 = n984 ^ x31 ;
  assign n988 = ~x137 & ~n985 ;
  assign n989 = n988 ^ x31 ;
  assign n990 = n983 & n989 ;
  assign n992 = n991 ^ n990 ;
  assign n974 = x115 ^ x87 ;
  assign n975 = x138 & ~n974 ;
  assign n976 = n975 ^ x87 ;
  assign n993 = n992 ^ n976 ;
  assign n977 = n976 ^ x72 ;
  assign n978 = n977 ^ x119 ;
  assign n979 = n978 ^ n976 ;
  assign n980 = x138 & ~n979 ;
  assign n981 = n980 ^ n977 ;
  assign n982 = ~x137 & ~n981 ;
  assign n994 = n993 ^ n982 ;
  assign n995 = ~x136 & n994 ;
  assign n996 = n995 ^ n992 ;
  assign n997 = x141 ^ x84 ;
  assign n1000 = n944 & n997 ;
  assign n1001 = n1000 ^ x84 ;
  assign n1002 = ~x129 & n1001 ;
  assign n1005 = x96 & ~n466 ;
  assign n1006 = n1005 ^ x116 ;
  assign n1007 = ~x85 & ~n1006 ;
  assign n1008 = n1007 ^ x116 ;
  assign n1009 = n441 & ~n1008 ;
  assign n1010 = x139 ^ x86 ;
  assign n1013 = n944 & n1010 ;
  assign n1014 = n1013 ^ x86 ;
  assign n1015 = ~x129 & n1014 ;
  assign n1016 = x140 ^ x87 ;
  assign n1019 = n944 & n1016 ;
  assign n1020 = n1019 ^ x87 ;
  assign n1021 = ~x129 & n1020 ;
  assign n1022 = x139 ^ x88 ;
  assign n1023 = n841 & n842 ;
  assign n1026 = n1022 & n1023 ;
  assign n1027 = n1026 ^ x88 ;
  assign n1028 = ~x129 & n1027 ;
  assign n1029 = x140 ^ x89 ;
  assign n1032 = n1023 & n1029 ;
  assign n1033 = n1032 ^ x89 ;
  assign n1034 = ~x129 & n1033 ;
  assign n1035 = x142 ^ x90 ;
  assign n1038 = n1023 & n1035 ;
  assign n1039 = n1038 ^ x90 ;
  assign n1040 = ~x129 & n1039 ;
  assign n1041 = x143 ^ x91 ;
  assign n1044 = n1023 & n1041 ;
  assign n1045 = n1044 ^ x91 ;
  assign n1046 = ~x129 & n1045 ;
  assign n1047 = x144 ^ x92 ;
  assign n1050 = n1023 & n1047 ;
  assign n1051 = n1050 ^ x92 ;
  assign n1052 = ~x129 & n1051 ;
  assign n1053 = x146 ^ x93 ;
  assign n1056 = n1023 & n1053 ;
  assign n1057 = n1056 ^ x93 ;
  assign n1058 = ~x129 & n1057 ;
  assign n1059 = x142 ^ x94 ;
  assign n1060 = x82 & x138 ;
  assign n1061 = ~n870 & n1060 ;
  assign n1062 = n840 & n1061 ;
  assign n1065 = n1059 & n1062 ;
  assign n1066 = n1065 ^ x94 ;
  assign n1067 = ~x129 & n1066 ;
  assign n1070 = ~x3 & ~x110 ;
  assign n1071 = ~n840 & ~n1070 ;
  assign n1072 = x95 & ~n1071 ;
  assign n1073 = n1072 ^ x143 ;
  assign n1074 = ~n1062 & n1073 ;
  assign n1075 = n1074 ^ x143 ;
  assign n1076 = ~x129 & n1075 ;
  assign n1079 = x96 & ~n1071 ;
  assign n1080 = n1079 ^ x146 ;
  assign n1081 = ~n1062 & n1080 ;
  assign n1082 = n1081 ^ x146 ;
  assign n1083 = ~x129 & n1082 ;
  assign n1086 = x97 & ~n1071 ;
  assign n1087 = n1086 ^ x145 ;
  assign n1088 = ~n1062 & n1087 ;
  assign n1089 = n1088 ^ x145 ;
  assign n1090 = ~x129 & n1089 ;
  assign n1091 = x145 ^ x98 ;
  assign n1094 = n1023 & n1091 ;
  assign n1095 = n1094 ^ x98 ;
  assign n1096 = ~x129 & n1095 ;
  assign n1097 = x141 ^ x99 ;
  assign n1100 = n1023 & n1097 ;
  assign n1101 = n1100 ^ x99 ;
  assign n1102 = ~x129 & n1101 ;
  assign n1105 = x100 & ~n1071 ;
  assign n1106 = n1105 ^ x144 ;
  assign n1107 = ~n1062 & n1106 ;
  assign n1108 = n1107 ^ x144 ;
  assign n1109 = ~x129 & n1108 ;
  assign n1110 = x124 ^ x77 ;
  assign n1111 = x138 & ~n1110 ;
  assign n1112 = n1111 ^ x77 ;
  assign n1113 = ~n870 & ~n1112 ;
  assign n1122 = x138 ^ x137 ;
  assign n1123 = x82 ^ x65 ;
  assign n1124 = n1123 ^ x37 ;
  assign n1125 = x136 & ~n1124 ;
  assign n1126 = n1125 ^ x82 ;
  assign n1127 = n1122 & n1126 ;
  assign n1121 = ~x65 & x136 ;
  assign n1128 = n1127 ^ n1121 ;
  assign n1114 = x137 ^ x136 ;
  assign n1115 = x96 ^ x93 ;
  assign n1118 = ~x137 & n1115 ;
  assign n1119 = n1118 ^ x96 ;
  assign n1120 = n1114 & n1119 ;
  assign n1129 = n1128 ^ n1120 ;
  assign n1130 = x138 & n1129 ;
  assign n1131 = n1130 ^ n1128 ;
  assign n1132 = ~n1113 & ~n1131 ;
  assign n1139 = x69 ^ x66 ;
  assign n1140 = x136 & n1139 ;
  assign n1141 = n1140 ^ x66 ;
  assign n1143 = n1141 ^ x34 ;
  assign n1142 = n1141 ^ x79 ;
  assign n1144 = n1143 ^ n1142 ;
  assign n1147 = x136 & n1144 ;
  assign n1148 = n1147 ^ n1142 ;
  assign n1149 = x137 & ~n1148 ;
  assign n1150 = n1149 ^ n1141 ;
  assign n1133 = x95 ^ x91 ;
  assign n1136 = ~x137 & n1133 ;
  assign n1137 = n1136 ^ x95 ;
  assign n1138 = n1114 & n1137 ;
  assign n1151 = n1150 ^ n1138 ;
  assign n1152 = x138 & ~n1151 ;
  assign n1153 = n1152 ^ n1150 ;
  assign n1159 = ~x74 & ~x137 ;
  assign n1154 = x63 ^ x33 ;
  assign n1155 = ~x137 & ~n1154 ;
  assign n1156 = n1155 ^ x33 ;
  assign n1160 = n1159 ^ n1156 ;
  assign n1161 = ~x136 & n1160 ;
  assign n1162 = n1161 ^ n1156 ;
  assign n1163 = ~x138 & n1162 ;
  assign n1164 = n1163 ^ x138 ;
  assign n1175 = x78 & n869 ;
  assign n1176 = ~n1164 & n1175 ;
  assign n1167 = x94 ^ x90 ;
  assign n1170 = x137 & n1167 ;
  assign n1171 = n1170 ^ x90 ;
  assign n1172 = n1114 & n1171 ;
  assign n1173 = x138 & n1172 ;
  assign n1174 = n1173 ^ n1163 ;
  assign n1177 = n1176 ^ n1174 ;
  assign n1185 = x73 ^ x68 ;
  assign n1186 = ~x136 & n1185 ;
  assign n1187 = n1186 ^ x68 ;
  assign n1189 = n1187 ^ x32 ;
  assign n1188 = n1187 ^ x84 ;
  assign n1190 = n1189 ^ n1188 ;
  assign n1193 = x136 & n1190 ;
  assign n1194 = n1193 ^ n1188 ;
  assign n1195 = x137 & ~n1194 ;
  assign n1196 = n1195 ^ n1187 ;
  assign n1178 = x138 ^ x112 ;
  assign n1179 = n1178 ^ x99 ;
  assign n1182 = x137 & n1179 ;
  assign n1183 = n1182 ^ x99 ;
  assign n1184 = n1114 & n1183 ;
  assign n1197 = n1196 ^ n1184 ;
  assign n1198 = x138 & ~n1197 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1218 = x125 ^ x92 ;
  assign n1219 = n1218 ^ x100 ;
  assign n1220 = ~x137 & n1219 ;
  assign n1221 = n1220 ^ x100 ;
  assign n1222 = x136 & n1221 ;
  assign n1202 = x80 ^ x75 ;
  assign n1203 = x137 & ~n1202 ;
  assign n1204 = n1203 ^ x75 ;
  assign n1206 = n1204 ^ x35 ;
  assign n1205 = n1204 ^ x70 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1210 = x137 & ~n1207 ;
  assign n1211 = n1210 ^ n1205 ;
  assign n1212 = x136 & n1211 ;
  assign n1213 = n1212 ^ n1204 ;
  assign n1214 = n1213 ^ x100 ;
  assign n1223 = n1222 ^ n1214 ;
  assign n1200 = x125 ^ x100 ;
  assign n1201 = ~x137 & n1200 ;
  assign n1224 = n1223 ^ n1201 ;
  assign n1225 = x138 & ~n1224 ;
  assign n1226 = n1225 ^ n1213 ;
  assign n1227 = n497 ^ n468 ;
  assign n1228 = n148 & n1227 ;
  assign n1247 = x98 & ~x137 ;
  assign n1240 = x71 ^ x36 ;
  assign n1241 = ~x137 & ~n1240 ;
  assign n1242 = n1241 ^ x36 ;
  assign n1248 = n1247 ^ n1242 ;
  assign n1249 = x138 & n1248 ;
  assign n1250 = n1249 ^ n1242 ;
  assign n1229 = x76 ^ x23 ;
  assign n1230 = ~x138 & ~n1229 ;
  assign n1231 = n1230 ^ x23 ;
  assign n1251 = n1250 ^ n1231 ;
  assign n1233 = n1231 ^ x81 ;
  assign n1232 = n1231 ^ x97 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1237 = ~x138 & n1234 ;
  assign n1238 = n1237 ^ n1232 ;
  assign n1239 = x137 & n1238 ;
  assign n1252 = n1251 ^ n1239 ;
  assign n1253 = ~x136 & n1252 ;
  assign n1254 = n1253 ^ n1250 ;
  assign n1273 = x88 & ~x137 ;
  assign n1266 = x88 ^ x64 ;
  assign n1267 = n1266 ^ x30 ;
  assign n1270 = ~x137 & ~n1267 ;
  assign n1271 = n1270 ^ x30 ;
  assign n1272 = n983 & n1271 ;
  assign n1274 = n1273 ^ n1272 ;
  assign n1255 = x120 ^ x67 ;
  assign n1256 = x138 & ~n1255 ;
  assign n1257 = n1256 ^ x67 ;
  assign n1275 = n1274 ^ n1257 ;
  assign n1259 = n1257 ^ x86 ;
  assign n1258 = n1257 ^ x111 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n1263 = ~x138 & n1260 ;
  assign n1264 = n1263 ^ n1258 ;
  assign n1265 = x137 & ~n1264 ;
  assign n1276 = n1275 ^ n1265 ;
  assign n1277 = ~x136 & ~n1276 ;
  assign n1278 = n1277 ^ n1274 ;
  assign n1279 = x116 & n148 ;
  assign n1284 = n431 & ~n458 ;
  assign n1285 = n1284 ^ n444 ;
  assign n1286 = n1279 & n1285 ;
  assign n1287 = n449 & n1279 ;
  assign n1288 = ~x53 & x97 ;
  assign n1289 = n1287 & n1288 ;
  assign n1290 = n1289 ^ n1287 ;
  assign n1291 = ~x129 & n840 ;
  assign n1292 = x139 ^ x111 ;
  assign n1295 = ~n1061 & n1292 ;
  assign n1296 = n1295 ^ x139 ;
  assign n1297 = n1291 & n1296 ;
  assign n1298 = x141 ^ x112 ;
  assign n1301 = ~n1061 & ~n1298 ;
  assign n1302 = n1301 ^ x141 ;
  assign n1303 = n1291 & n1302 ;
  assign n1304 = n224 ^ x113 ;
  assign n1307 = x54 & n1304 ;
  assign n1308 = n1307 ^ x113 ;
  assign n1309 = n148 & ~n1308 ;
  assign n1310 = x140 ^ x115 ;
  assign n1313 = ~n1061 & ~n1310 ;
  assign n1314 = n1313 ^ x140 ;
  assign n1315 = n1291 & n1314 ;
  assign n1316 = ~n166 & n220 ;
  assign n1317 = x122 & ~x129 ;
  assign n1322 = ~x54 & x118 ;
  assign n1323 = n1322 ^ n340 ;
  assign n1324 = ~x129 & n1323 ;
  assign n1325 = ~x129 & ~n463 ;
  assign n1326 = ~x111 & ~x129 ;
  assign n1327 = ~x120 & n1070 ;
  assign n1328 = n1326 & n1327 ;
  assign n1329 = n1328 ^ n1326 ;
  assign n1330 = x81 & x120 ;
  assign n1331 = ~x129 & n1330 ;
  assign n1332 = ~x129 & ~x134 ;
  assign n1333 = ~x129 & ~x135 ;
  assign n1334 = x57 & ~x129 ;
  assign n1337 = n148 ^ x129 ;
  assign n1335 = ~x96 & x125 ;
  assign n1336 = n148 & n1335 ;
  assign n1338 = n1337 ^ n1336 ;
  assign n1339 = ~x126 & n839 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n217 ;
  assign y16 = ~n235 ;
  assign y17 = ~n276 ;
  assign y18 = n286 ;
  assign y19 = n292 ;
  assign y20 = n303 ;
  assign y21 = n308 ;
  assign y22 = n311 ;
  assign y23 = n314 ;
  assign y24 = n320 ;
  assign y25 = n323 ;
  assign y26 = n331 ;
  assign y27 = n336 ;
  assign y28 = n344 ;
  assign y29 = n347 ;
  assign y30 = n369 ;
  assign y31 = n372 ;
  assign y32 = n378 ;
  assign y33 = n381 ;
  assign y34 = n384 ;
  assign y35 = n409 ;
  assign y36 = n412 ;
  assign y37 = n414 ;
  assign y38 = n417 ;
  assign y39 = n430 ;
  assign y40 = n483 ;
  assign y41 = n489 ;
  assign y42 = n511 ;
  assign y43 = n523 ;
  assign y44 = n543 ;
  assign y45 = n553 ;
  assign y46 = n563 ;
  assign y47 = n573 ;
  assign y48 = n583 ;
  assign y49 = n593 ;
  assign y50 = n603 ;
  assign y51 = n613 ;
  assign y52 = n623 ;
  assign y53 = ~n635 ;
  assign y54 = ~n645 ;
  assign y55 = n657 ;
  assign y56 = ~n674 ;
  assign y57 = n683 ;
  assign y58 = ~n695 ;
  assign y59 = n703 ;
  assign y60 = ~n716 ;
  assign y61 = ~n727 ;
  assign y62 = ~n740 ;
  assign y63 = ~n757 ;
  assign y64 = n766 ;
  assign y65 = n789 ;
  assign y66 = ~n792 ;
  assign y67 = ~n795 ;
  assign y68 = n536 ;
  assign y69 = ~n796 ;
  assign y70 = n799 ;
  assign y71 = n814 ;
  assign y72 = n820 ;
  assign y73 = n828 ;
  assign y74 = n832 ;
  assign y75 = n836 ;
  assign y76 = n837 ;
  assign y77 = ~n849 ;
  assign y78 = ~n855 ;
  assign y79 = ~n861 ;
  assign y80 = ~n867 ;
  assign y81 = ~n876 ;
  assign y82 = ~n882 ;
  assign y83 = ~n888 ;
  assign y84 = ~n894 ;
  assign y85 = ~n900 ;
  assign y86 = ~n906 ;
  assign y87 = ~n912 ;
  assign y88 = ~n918 ;
  assign y89 = ~n924 ;
  assign y90 = ~n930 ;
  assign y91 = ~n936 ;
  assign y92 = ~n942 ;
  assign y93 = n949 ;
  assign y94 = n955 ;
  assign y95 = n961 ;
  assign y96 = n967 ;
  assign y97 = n973 ;
  assign y98 = n996 ;
  assign y99 = n1002 ;
  assign y100 = n1009 ;
  assign y101 = n1015 ;
  assign y102 = n1021 ;
  assign y103 = n1028 ;
  assign y104 = n1034 ;
  assign y105 = n1040 ;
  assign y106 = n1046 ;
  assign y107 = n1052 ;
  assign y108 = n1058 ;
  assign y109 = n1067 ;
  assign y110 = n1076 ;
  assign y111 = n1083 ;
  assign y112 = n1090 ;
  assign y113 = n1096 ;
  assign y114 = n1102 ;
  assign y115 = n1109 ;
  assign y116 = ~n1132 ;
  assign y117 = ~n1153 ;
  assign y118 = n1177 ;
  assign y119 = ~n1199 ;
  assign y120 = ~n1226 ;
  assign y121 = n1228 ;
  assign y122 = n1254 ;
  assign y123 = n1278 ;
  assign y124 = n1286 ;
  assign y125 = n1290 ;
  assign y126 = n1297 ;
  assign y127 = n1303 ;
  assign y128 = n1309 ;
  assign y129 = n279 ;
  assign y130 = n1315 ;
  assign y131 = n1316 ;
  assign y132 = ~n1317 ;
  assign y133 = n1324 ;
  assign y134 = n1325 ;
  assign y135 = n1329 ;
  assign y136 = n1331 ;
  assign y137 = ~n1332 ;
  assign y138 = ~n1333 ;
  assign y139 = n1334 ;
  assign y140 = ~n1338 ;
  assign y141 = n1339 ;
endmodule
