module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, y0, y64, y16, y80, y32, y96, y48, y112, y4, y68, y20, y84, y36, y100, y52, y116, y8, y72, y24, y88, y40, y104, y56, y120, y12, y76, y28, y92, y44, y108, y60, y124, y3, y67, y19, y83, y35, y99, y51, y115, y15, y79, y63, y127, y31, y95, y47, y111, y7, y71, y23, y87, y39, y103, y55, y119, y11, y75, y27, y91, y43, y107, y59, y123, y1, y65, y17, y81, y33, y97, y49, y113, y5, y69, y21, y85, y37, y101, y53, y117, y9, y73, y25, y89, y41, y105, y57, y121, y13, y77, y29, y93, y45, y109, y61, y125, y2, y66, y18, y82, y34, y98, y50, y114, y6, y70, y22, y86, y38, y102, y54, y118, y10, y74, y26, y90, y42, y106, y58, y122, y14, y78, y30, y94, y46, y110, y62, y126;
assign n_0 = x2 ^ x0;
assign n_1 = x3 ^ x1;
assign n_2 = x4 ^ x2;
assign n_3 = x5 ^ x3;
assign n_4 = x6 ^ x4;
assign n_5 = x7 ^ x5;
assign n_6 = x8 ^ x6;
assign n_7 = x9 ^ x7;
assign n_8 = x10 ^ x8;
assign n_9 = x11 ^ x9;
assign n_10 = x12 ^ x10;
assign n_11 = x13 ^ x11;
assign n_12 = x14 ^ x12;
assign n_13 = x15 ^ x13;
assign n_14 = x16 ^ x14;
assign n_15 = x17 ^ x15;
assign n_16 = x18 ^ x16;
assign n_17 = x19 ^ x17;
assign n_18 = x20 ^ x18;
assign n_19 = x21 ^ x19;
assign n_20 = x22 ^ x20;
assign n_21 = x23 ^ x21;
assign n_22 = x24 ^ x22;
assign n_23 = x25 ^ x23;
assign n_24 = x26 ^ x24;
assign n_25 = x27 ^ x25;
assign n_26 = x28 ^ x26;
assign n_27 = x29 ^ x27;
assign n_28 = x30 ^ x28;
assign n_29 = x31 ^ x29;
assign n_30 = x32 ^ x30;
assign n_31 = x33 ^ x31;
assign n_32 = x34 ^ x32;
assign n_33 = x35 ^ x33;
assign n_34 = x36 ^ x34;
assign n_35 = x37 ^ x35;
assign n_36 = x38 ^ x36;
assign n_37 = x39 ^ x37;
assign n_38 = x40 ^ x38;
assign n_39 = x41 ^ x39;
assign n_40 = x42 ^ x40;
assign n_41 = x43 ^ x41;
assign n_42 = x44 ^ x42;
assign n_43 = x45 ^ x43;
assign n_44 = x46 ^ x44;
assign n_45 = x47 ^ x45;
assign n_46 = x48 ^ x46;
assign n_47 = x49 ^ x47;
assign n_48 = x50 ^ x48;
assign n_49 = x51 ^ x49;
assign n_50 = x52 ^ x50;
assign n_51 = x53 ^ x51;
assign n_52 = x54 ^ x52;
assign n_53 = x55 ^ x53;
assign n_54 = x56 ^ x54;
assign n_55 = x57 ^ x55;
assign n_56 = x58 ^ x56;
assign n_57 = x59 ^ x57;
assign n_58 = x60 ^ x58;
assign n_59 = x61 ^ x59;
assign n_60 = x62 ^ x60;
assign n_61 = x63 ^ x61;
assign n_62 = x64 ^ x62;
assign n_63 = x65 ^ x63;
assign n_64 = x66 ^ x64;
assign n_65 = x67 ^ x65;
assign n_66 = x68 ^ x66;
assign n_67 = x69 ^ x67;
assign n_68 = x70 ^ x68;
assign n_69 = x71 ^ x69;
assign n_70 = x72 ^ x70;
assign n_71 = x73 ^ x71;
assign n_72 = x74 ^ x72;
assign n_73 = x75 ^ x73;
assign n_74 = x76 ^ x74;
assign n_75 = x77 ^ x75;
assign n_76 = x78 ^ x76;
assign n_77 = x79 ^ x77;
assign n_78 = x80 ^ x78;
assign n_79 = x81 ^ x79;
assign n_80 = x82 ^ x80;
assign n_81 = x83 ^ x81;
assign n_82 = x84 ^ x82;
assign n_83 = x85 ^ x83;
assign n_84 = x86 ^ x84;
assign n_85 = x87 ^ x85;
assign n_86 = x88 ^ x86;
assign n_87 = x89 ^ x87;
assign n_88 = x90 ^ x88;
assign n_89 = x91 ^ x89;
assign n_90 = x92 ^ x90;
assign n_91 = x93 ^ x91;
assign n_92 = x94 ^ x92;
assign n_93 = x95 ^ x93;
assign n_94 = x96 ^ x94;
assign n_95 = x97 ^ x95;
assign n_96 = x98 ^ x96;
assign n_97 = x99 ^ x97;
assign n_98 = x100 ^ x98;
assign n_99 = x101 ^ x99;
assign n_100 = x102 ^ x100;
assign n_101 = x103 ^ x101;
assign n_102 = x104 ^ x102;
assign n_103 = x105 ^ x103;
assign n_104 = x106 ^ x104;
assign n_105 = x107 ^ x105;
assign n_106 = x108 ^ x106;
assign n_107 = x109 ^ x107;
assign n_108 = x110 ^ x108;
assign n_109 = x111 ^ x109;
assign n_110 = x112 ^ x110;
assign n_111 = x113 ^ x111;
assign n_112 = x114 ^ x112;
assign n_113 = x115 ^ x113;
assign n_114 = x116 ^ x114;
assign n_115 = x117 ^ x115;
assign n_116 = x118 ^ x116;
assign n_117 = x119 ^ x117;
assign n_118 = x120 ^ x118;
assign n_119 = x121 ^ x119;
assign n_120 = x122 ^ x120;
assign n_121 = x123 ^ x121;
assign n_122 = x124 ^ x122;
assign n_123 = x125 ^ x123;
assign n_124 = x126 ^ x0;
assign n_125 = x126 ^ x124;
assign n_126 = x127 ^ x125;
assign n_127 = x127 ^ x1;
assign n_128 = ~x129 & n_0;
assign n_129 = ~x129 & n_1;
assign n_130 = ~x129 & n_2;
assign n_131 = ~x129 & n_3;
assign n_132 = ~x129 & n_4;
assign n_133 = ~x129 & n_5;
assign n_134 = ~x129 & n_6;
assign n_135 = ~x129 & n_7;
assign n_136 = ~x129 & n_8;
assign n_137 = ~x129 & n_9;
assign n_138 = ~x129 & n_10;
assign n_139 = ~x129 & n_11;
assign n_140 = ~x129 & n_12;
assign n_141 = ~x129 & n_13;
assign n_142 = ~x129 & n_14;
assign n_143 = ~x129 & n_15;
assign n_144 = ~x129 & n_16;
assign n_145 = ~x129 & n_17;
assign n_146 = ~x129 & n_18;
assign n_147 = ~x129 & n_19;
assign n_148 = ~x129 & n_20;
assign n_149 = ~x129 & n_21;
assign n_150 = ~x129 & n_22;
assign n_151 = ~x129 & n_23;
assign n_152 = ~x129 & n_24;
assign n_153 = ~x129 & n_25;
assign n_154 = ~x129 & n_26;
assign n_155 = ~x129 & n_27;
assign n_156 = ~x129 & n_28;
assign n_157 = ~x129 & n_29;
assign n_158 = ~x129 & n_30;
assign n_159 = ~x129 & n_31;
assign n_160 = ~x129 & n_32;
assign n_161 = ~x129 & n_33;
assign n_162 = ~x129 & n_34;
assign n_163 = ~x129 & n_35;
assign n_164 = ~x129 & n_36;
assign n_165 = ~x129 & n_37;
assign n_166 = ~x129 & n_38;
assign n_167 = ~x129 & n_39;
assign n_168 = ~x129 & n_40;
assign n_169 = ~x129 & n_41;
assign n_170 = ~x129 & n_42;
assign n_171 = ~x129 & n_43;
assign n_172 = ~x129 & n_44;
assign n_173 = ~x129 & n_45;
assign n_174 = ~x129 & n_46;
assign n_175 = ~x129 & n_47;
assign n_176 = ~x129 & n_48;
assign n_177 = ~x129 & n_49;
assign n_178 = ~x129 & n_50;
assign n_179 = ~x129 & n_51;
assign n_180 = ~x129 & n_52;
assign n_181 = ~x129 & n_53;
assign n_182 = ~x129 & n_54;
assign n_183 = ~x129 & n_55;
assign n_184 = ~x129 & n_56;
assign n_185 = ~x129 & n_57;
assign n_186 = ~x129 & n_58;
assign n_187 = ~x129 & n_59;
assign n_188 = ~x129 & n_60;
assign n_189 = ~x129 & n_61;
assign n_190 = ~x129 & n_62;
assign n_191 = ~x129 & n_63;
assign n_192 = ~x129 & n_64;
assign n_193 = ~x129 & n_65;
assign n_194 = ~x129 & n_66;
assign n_195 = ~x129 & n_67;
assign n_196 = ~x129 & n_68;
assign n_197 = ~x129 & n_69;
assign n_198 = ~x129 & n_70;
assign n_199 = ~x129 & n_71;
assign n_200 = ~x129 & n_72;
assign n_201 = ~x129 & n_73;
assign n_202 = ~x129 & n_74;
assign n_203 = ~x129 & n_75;
assign n_204 = ~x129 & n_76;
assign n_205 = ~x129 & n_77;
assign n_206 = ~x129 & n_78;
assign n_207 = ~x129 & n_79;
assign n_208 = ~x129 & n_80;
assign n_209 = ~x129 & n_81;
assign n_210 = ~x129 & n_82;
assign n_211 = ~x129 & n_83;
assign n_212 = ~x129 & n_84;
assign n_213 = ~x129 & n_85;
assign n_214 = ~x129 & n_86;
assign n_215 = ~x129 & n_87;
assign n_216 = ~x129 & n_88;
assign n_217 = ~x129 & n_89;
assign n_218 = ~x129 & n_90;
assign n_219 = ~x129 & n_91;
assign n_220 = ~x129 & n_92;
assign n_221 = ~x129 & n_93;
assign n_222 = ~x129 & n_94;
assign n_223 = ~x129 & n_95;
assign n_224 = ~x129 & n_96;
assign n_225 = ~x129 & n_97;
assign n_226 = ~x129 & n_98;
assign n_227 = ~x129 & n_99;
assign n_228 = ~x129 & n_100;
assign n_229 = ~x129 & n_101;
assign n_230 = ~x129 & n_102;
assign n_231 = ~x129 & n_103;
assign n_232 = ~x129 & n_104;
assign n_233 = ~x129 & n_105;
assign n_234 = ~x129 & n_106;
assign n_235 = ~x129 & n_107;
assign n_236 = ~x129 & n_108;
assign n_237 = ~x129 & n_109;
assign n_238 = ~x129 & n_110;
assign n_239 = ~x129 & n_111;
assign n_240 = ~x129 & n_112;
assign n_241 = ~x129 & n_113;
assign n_242 = ~x129 & n_114;
assign n_243 = ~x129 & n_115;
assign n_244 = ~x129 & n_116;
assign n_245 = ~x129 & n_117;
assign n_246 = ~x129 & n_118;
assign n_247 = ~x129 & n_119;
assign n_248 = ~x129 & n_120;
assign n_249 = ~x129 & n_121;
assign n_250 = ~x129 & n_122;
assign n_251 = ~x129 & n_123;
assign n_252 = x129 & n_124;
assign n_253 = ~x129 & n_125;
assign n_254 = ~x129 & n_126;
assign n_255 = x129 & n_127;
assign n_256 = n_128 ^ x0;
assign n_257 = n_129 ^ x1;
assign n_258 = n_130 ^ x2;
assign n_259 = n_131 ^ x3;
assign n_260 = n_132 ^ x4;
assign n_261 = n_133 ^ x5;
assign n_262 = n_134 ^ x6;
assign n_263 = n_135 ^ x7;
assign n_264 = n_136 ^ x8;
assign n_265 = n_137 ^ x9;
assign n_266 = n_138 ^ x10;
assign n_267 = n_139 ^ x11;
assign n_268 = n_140 ^ x12;
assign n_269 = n_141 ^ x13;
assign n_270 = n_142 ^ x14;
assign n_271 = n_143 ^ x15;
assign n_272 = n_144 ^ x16;
assign n_273 = n_145 ^ x17;
assign n_274 = n_146 ^ x18;
assign n_275 = n_147 ^ x19;
assign n_276 = n_148 ^ x20;
assign n_277 = n_149 ^ x21;
assign n_278 = n_150 ^ x22;
assign n_279 = n_151 ^ x23;
assign n_280 = n_152 ^ x24;
assign n_281 = n_153 ^ x25;
assign n_282 = n_154 ^ x26;
assign n_283 = n_155 ^ x27;
assign n_284 = n_156 ^ x28;
assign n_285 = n_157 ^ x29;
assign n_286 = n_158 ^ x30;
assign n_287 = n_159 ^ x31;
assign n_288 = n_160 ^ x32;
assign n_289 = n_161 ^ x33;
assign n_290 = n_162 ^ x34;
assign n_291 = n_163 ^ x35;
assign n_292 = n_164 ^ x36;
assign n_293 = n_165 ^ x37;
assign n_294 = n_166 ^ x38;
assign n_295 = n_167 ^ x39;
assign n_296 = n_168 ^ x40;
assign n_297 = n_169 ^ x41;
assign n_298 = n_170 ^ x42;
assign n_299 = n_171 ^ x43;
assign n_300 = n_172 ^ x44;
assign n_301 = n_173 ^ x45;
assign n_302 = n_174 ^ x46;
assign n_303 = n_175 ^ x47;
assign n_304 = n_176 ^ x48;
assign n_305 = n_177 ^ x49;
assign n_306 = n_178 ^ x50;
assign n_307 = n_179 ^ x51;
assign n_308 = n_180 ^ x52;
assign n_309 = n_181 ^ x53;
assign n_310 = n_182 ^ x54;
assign n_311 = n_183 ^ x55;
assign n_312 = n_184 ^ x56;
assign n_313 = n_185 ^ x57;
assign n_314 = n_186 ^ x58;
assign n_315 = n_187 ^ x59;
assign n_316 = n_188 ^ x60;
assign n_317 = n_189 ^ x61;
assign n_318 = n_190 ^ x62;
assign n_319 = n_191 ^ x63;
assign n_320 = n_192 ^ x64;
assign n_321 = n_193 ^ x65;
assign n_322 = n_194 ^ x66;
assign n_323 = n_195 ^ x67;
assign n_324 = n_196 ^ x68;
assign n_325 = n_197 ^ x69;
assign n_326 = n_198 ^ x70;
assign n_327 = n_199 ^ x71;
assign n_328 = n_200 ^ x72;
assign n_329 = n_201 ^ x73;
assign n_330 = n_202 ^ x74;
assign n_331 = n_203 ^ x75;
assign n_332 = n_204 ^ x76;
assign n_333 = n_205 ^ x77;
assign n_334 = n_206 ^ x78;
assign n_335 = n_207 ^ x79;
assign n_336 = n_208 ^ x80;
assign n_337 = n_209 ^ x81;
assign n_338 = n_210 ^ x82;
assign n_339 = n_211 ^ x83;
assign n_340 = n_212 ^ x84;
assign n_341 = n_213 ^ x85;
assign n_342 = n_214 ^ x86;
assign n_343 = n_215 ^ x87;
assign n_344 = n_216 ^ x88;
assign n_345 = n_217 ^ x89;
assign n_346 = n_218 ^ x90;
assign n_347 = n_219 ^ x91;
assign n_348 = n_220 ^ x92;
assign n_349 = n_221 ^ x93;
assign n_350 = n_222 ^ x94;
assign n_351 = n_223 ^ x95;
assign n_352 = n_224 ^ x96;
assign n_353 = n_225 ^ x97;
assign n_354 = n_226 ^ x98;
assign n_355 = n_227 ^ x99;
assign n_356 = n_228 ^ x100;
assign n_357 = n_229 ^ x101;
assign n_358 = n_230 ^ x102;
assign n_359 = n_231 ^ x103;
assign n_360 = n_232 ^ x104;
assign n_361 = n_233 ^ x105;
assign n_362 = n_234 ^ x106;
assign n_363 = n_235 ^ x107;
assign n_364 = n_236 ^ x108;
assign n_365 = n_237 ^ x109;
assign n_366 = n_238 ^ x110;
assign n_367 = n_239 ^ x111;
assign n_368 = n_240 ^ x112;
assign n_369 = n_241 ^ x113;
assign n_370 = n_242 ^ x114;
assign n_371 = n_243 ^ x115;
assign n_372 = n_244 ^ x116;
assign n_373 = n_245 ^ x117;
assign n_374 = n_246 ^ x118;
assign n_375 = n_247 ^ x119;
assign n_376 = n_248 ^ x120;
assign n_377 = n_249 ^ x121;
assign n_378 = n_250 ^ x122;
assign n_379 = n_251 ^ x123;
assign n_380 = n_252 ^ x0;
assign n_381 = n_253 ^ x124;
assign n_382 = n_254 ^ x125;
assign n_383 = n_255 ^ x1;
assign n_384 = n_256 ^ n_257;
assign n_385 = n_258 ^ n_257;
assign n_386 = n_259 ^ n_258;
assign n_387 = n_260 ^ n_259;
assign n_388 = n_260 ^ n_261;
assign n_389 = n_262 ^ n_261;
assign n_390 = n_263 ^ n_262;
assign n_391 = n_264 ^ n_263;
assign n_392 = n_264 ^ n_265;
assign n_393 = n_266 ^ n_265;
assign n_394 = n_267 ^ n_266;
assign n_395 = n_268 ^ n_267;
assign n_396 = n_268 ^ n_269;
assign n_397 = n_270 ^ n_269;
assign n_398 = n_271 ^ n_270;
assign n_399 = n_272 ^ n_271;
assign n_400 = n_272 ^ n_273;
assign n_401 = n_274 ^ n_273;
assign n_402 = n_275 ^ n_274;
assign n_403 = n_276 ^ n_275;
assign n_404 = n_276 ^ n_277;
assign n_405 = n_278 ^ n_277;
assign n_406 = n_279 ^ n_278;
assign n_407 = n_280 ^ n_279;
assign n_408 = n_280 ^ n_281;
assign n_409 = n_282 ^ n_281;
assign n_410 = n_283 ^ n_282;
assign n_411 = n_284 ^ n_283;
assign n_412 = n_284 ^ n_285;
assign n_413 = n_286 ^ n_285;
assign n_414 = n_287 ^ n_286;
assign n_415 = n_288 ^ n_287;
assign n_416 = n_288 ^ n_289;
assign n_417 = n_290 ^ n_289;
assign n_418 = n_291 ^ n_290;
assign n_419 = n_292 ^ n_291;
assign n_420 = n_292 ^ n_293;
assign n_421 = n_294 ^ n_293;
assign n_422 = n_295 ^ n_294;
assign n_423 = n_296 ^ n_295;
assign n_424 = n_296 ^ n_297;
assign n_425 = n_298 ^ n_297;
assign n_426 = n_299 ^ n_298;
assign n_427 = n_300 ^ n_299;
assign n_428 = n_300 ^ n_301;
assign n_429 = n_302 ^ n_301;
assign n_430 = n_303 ^ n_302;
assign n_431 = n_304 ^ n_303;
assign n_432 = n_304 ^ n_305;
assign n_433 = n_306 ^ n_305;
assign n_434 = n_307 ^ n_306;
assign n_435 = n_308 ^ n_307;
assign n_436 = n_308 ^ n_309;
assign n_437 = n_310 ^ n_309;
assign n_438 = n_311 ^ n_310;
assign n_439 = n_312 ^ n_311;
assign n_440 = n_312 ^ n_313;
assign n_441 = n_314 ^ n_313;
assign n_442 = n_315 ^ n_314;
assign n_443 = n_316 ^ n_315;
assign n_444 = n_316 ^ n_317;
assign n_445 = n_318 ^ n_317;
assign n_446 = n_319 ^ n_318;
assign n_447 = n_320 ^ n_319;
assign n_448 = n_320 ^ n_321;
assign n_449 = n_322 ^ n_321;
assign n_450 = n_323 ^ n_322;
assign n_451 = n_324 ^ n_323;
assign n_452 = n_324 ^ n_325;
assign n_453 = n_326 ^ n_325;
assign n_454 = n_327 ^ n_326;
assign n_455 = n_328 ^ n_327;
assign n_456 = n_328 ^ n_329;
assign n_457 = n_330 ^ n_329;
assign n_458 = n_331 ^ n_330;
assign n_459 = n_332 ^ n_331;
assign n_460 = n_332 ^ n_333;
assign n_461 = n_334 ^ n_333;
assign n_462 = n_335 ^ n_334;
assign n_463 = n_336 ^ n_335;
assign n_464 = n_336 ^ n_337;
assign n_465 = n_338 ^ n_337;
assign n_466 = n_339 ^ n_338;
assign n_467 = n_340 ^ n_339;
assign n_468 = n_340 ^ n_341;
assign n_469 = n_342 ^ n_341;
assign n_470 = n_343 ^ n_342;
assign n_471 = n_344 ^ n_343;
assign n_472 = n_344 ^ n_345;
assign n_473 = n_346 ^ n_345;
assign n_474 = n_347 ^ n_346;
assign n_475 = n_348 ^ n_347;
assign n_476 = n_348 ^ n_349;
assign n_477 = n_350 ^ n_349;
assign n_478 = n_351 ^ n_350;
assign n_479 = n_352 ^ n_351;
assign n_480 = n_352 ^ n_353;
assign n_481 = n_354 ^ n_353;
assign n_482 = n_355 ^ n_354;
assign n_483 = n_356 ^ n_355;
assign n_484 = n_356 ^ n_357;
assign n_485 = n_358 ^ n_357;
assign n_486 = n_359 ^ n_358;
assign n_487 = n_360 ^ n_359;
assign n_488 = n_360 ^ n_361;
assign n_489 = n_362 ^ n_361;
assign n_490 = n_363 ^ n_362;
assign n_491 = n_364 ^ n_363;
assign n_492 = n_364 ^ n_365;
assign n_493 = n_366 ^ n_365;
assign n_494 = n_367 ^ n_366;
assign n_495 = n_368 ^ n_367;
assign n_496 = n_368 ^ n_369;
assign n_497 = n_370 ^ n_369;
assign n_498 = n_371 ^ n_370;
assign n_499 = n_372 ^ n_371;
assign n_500 = n_372 ^ n_373;
assign n_501 = n_374 ^ n_373;
assign n_502 = n_375 ^ n_374;
assign n_503 = n_376 ^ n_375;
assign n_504 = n_376 ^ n_377;
assign n_505 = n_378 ^ n_377;
assign n_506 = n_379 ^ n_378;
assign n_507 = n_381 ^ n_379;
assign n_508 = n_382 ^ n_380;
assign n_509 = n_381 ^ n_382;
assign n_510 = n_383 ^ n_380;
assign n_511 = n_256 ^ n_383;
assign n_512 = x128 & n_384;
assign n_513 = x128 & n_385;
assign n_514 = ~x128 & n_386;
assign n_515 = ~x128 & n_387;
assign n_516 = x128 & n_388;
assign n_517 = x128 & n_389;
assign n_518 = ~x128 & n_390;
assign n_519 = ~x128 & n_391;
assign n_520 = x128 & n_392;
assign n_521 = x128 & n_393;
assign n_522 = ~x128 & n_394;
assign n_523 = ~x128 & n_395;
assign n_524 = x128 & n_396;
assign n_525 = x128 & n_397;
assign n_526 = ~x128 & n_398;
assign n_527 = ~x128 & n_399;
assign n_528 = x128 & n_400;
assign n_529 = x128 & n_401;
assign n_530 = ~x128 & n_402;
assign n_531 = ~x128 & n_403;
assign n_532 = x128 & n_404;
assign n_533 = x128 & n_405;
assign n_534 = ~x128 & n_406;
assign n_535 = ~x128 & n_407;
assign n_536 = x128 & n_408;
assign n_537 = x128 & n_409;
assign n_538 = ~x128 & n_410;
assign n_539 = ~x128 & n_411;
assign n_540 = x128 & n_412;
assign n_541 = x128 & n_413;
assign n_542 = ~x128 & n_414;
assign n_543 = ~x128 & n_415;
assign n_544 = x128 & n_416;
assign n_545 = x128 & n_417;
assign n_546 = ~x128 & n_418;
assign n_547 = ~x128 & n_419;
assign n_548 = x128 & n_420;
assign n_549 = x128 & n_421;
assign n_550 = ~x128 & n_422;
assign n_551 = ~x128 & n_423;
assign n_552 = x128 & n_424;
assign n_553 = x128 & n_425;
assign n_554 = ~x128 & n_426;
assign n_555 = ~x128 & n_427;
assign n_556 = x128 & n_428;
assign n_557 = x128 & n_429;
assign n_558 = ~x128 & n_430;
assign n_559 = ~x128 & n_431;
assign n_560 = x128 & n_432;
assign n_561 = x128 & n_433;
assign n_562 = ~x128 & n_434;
assign n_563 = ~x128 & n_435;
assign n_564 = x128 & n_436;
assign n_565 = x128 & n_437;
assign n_566 = ~x128 & n_438;
assign n_567 = ~x128 & n_439;
assign n_568 = x128 & n_440;
assign n_569 = x128 & n_441;
assign n_570 = ~x128 & n_442;
assign n_571 = ~x128 & n_443;
assign n_572 = x128 & n_444;
assign n_573 = x128 & n_445;
assign n_574 = ~x128 & n_446;
assign n_575 = ~x128 & n_447;
assign n_576 = x128 & n_448;
assign n_577 = x128 & n_449;
assign n_578 = ~x128 & n_450;
assign n_579 = ~x128 & n_451;
assign n_580 = x128 & n_452;
assign n_581 = x128 & n_453;
assign n_582 = ~x128 & n_454;
assign n_583 = ~x128 & n_455;
assign n_584 = x128 & n_456;
assign n_585 = x128 & n_457;
assign n_586 = ~x128 & n_458;
assign n_587 = ~x128 & n_459;
assign n_588 = x128 & n_460;
assign n_589 = x128 & n_461;
assign n_590 = ~x128 & n_462;
assign n_591 = ~x128 & n_463;
assign n_592 = x128 & n_464;
assign n_593 = x128 & n_465;
assign n_594 = ~x128 & n_466;
assign n_595 = ~x128 & n_467;
assign n_596 = x128 & n_468;
assign n_597 = x128 & n_469;
assign n_598 = ~x128 & n_470;
assign n_599 = ~x128 & n_471;
assign n_600 = x128 & n_472;
assign n_601 = x128 & n_473;
assign n_602 = ~x128 & n_474;
assign n_603 = ~x128 & n_475;
assign n_604 = x128 & n_476;
assign n_605 = x128 & n_477;
assign n_606 = ~x128 & n_478;
assign n_607 = ~x128 & n_479;
assign n_608 = x128 & n_480;
assign n_609 = x128 & n_481;
assign n_610 = ~x128 & n_482;
assign n_611 = ~x128 & n_483;
assign n_612 = x128 & n_484;
assign n_613 = x128 & n_485;
assign n_614 = ~x128 & n_486;
assign n_615 = ~x128 & n_487;
assign n_616 = x128 & n_488;
assign n_617 = x128 & n_489;
assign n_618 = ~x128 & n_490;
assign n_619 = ~x128 & n_491;
assign n_620 = x128 & n_492;
assign n_621 = x128 & n_493;
assign n_622 = ~x128 & n_494;
assign n_623 = ~x128 & n_495;
assign n_624 = x128 & n_496;
assign n_625 = x128 & n_497;
assign n_626 = ~x128 & n_498;
assign n_627 = ~x128 & n_499;
assign n_628 = x128 & n_500;
assign n_629 = x128 & n_501;
assign n_630 = ~x128 & n_502;
assign n_631 = ~x128 & n_503;
assign n_632 = x128 & n_504;
assign n_633 = x128 & n_505;
assign n_634 = ~x128 & n_506;
assign n_635 = ~x128 & n_507;
assign n_636 = x128 & n_508;
assign n_637 = x128 & n_509;
assign n_638 = ~x128 & n_510;
assign n_639 = ~x128 & n_511;
assign n_640 = n_512 ^ n_257;
assign n_641 = n_513 ^ n_258;
assign n_642 = n_514 ^ n_258;
assign n_643 = n_515 ^ n_259;
assign n_644 = n_516 ^ n_261;
assign n_645 = n_517 ^ n_262;
assign n_646 = n_518 ^ n_262;
assign n_647 = n_519 ^ n_263;
assign n_648 = n_520 ^ n_265;
assign n_649 = n_521 ^ n_266;
assign n_650 = n_522 ^ n_266;
assign n_651 = n_523 ^ n_267;
assign n_652 = n_524 ^ n_269;
assign n_653 = n_525 ^ n_270;
assign n_654 = n_526 ^ n_270;
assign n_655 = n_527 ^ n_271;
assign n_656 = n_528 ^ n_273;
assign n_657 = n_529 ^ n_274;
assign n_658 = n_530 ^ n_274;
assign n_659 = n_531 ^ n_275;
assign n_660 = n_532 ^ n_277;
assign n_661 = n_533 ^ n_278;
assign n_662 = n_534 ^ n_278;
assign n_663 = n_535 ^ n_279;
assign n_664 = n_536 ^ n_281;
assign n_665 = n_537 ^ n_282;
assign n_666 = n_538 ^ n_282;
assign n_667 = n_539 ^ n_283;
assign n_668 = n_540 ^ n_285;
assign n_669 = n_541 ^ n_286;
assign n_670 = n_542 ^ n_286;
assign n_671 = n_543 ^ n_287;
assign n_672 = n_544 ^ n_289;
assign n_673 = n_545 ^ n_290;
assign n_674 = n_546 ^ n_290;
assign n_675 = n_547 ^ n_291;
assign n_676 = n_548 ^ n_293;
assign n_677 = n_549 ^ n_294;
assign n_678 = n_550 ^ n_294;
assign n_679 = n_551 ^ n_295;
assign n_680 = n_552 ^ n_297;
assign n_681 = n_553 ^ n_298;
assign n_682 = n_554 ^ n_298;
assign n_683 = n_555 ^ n_299;
assign n_684 = n_556 ^ n_301;
assign n_685 = n_557 ^ n_302;
assign n_686 = n_558 ^ n_302;
assign n_687 = n_559 ^ n_303;
assign n_688 = n_560 ^ n_305;
assign n_689 = n_561 ^ n_306;
assign n_690 = n_562 ^ n_306;
assign n_691 = n_563 ^ n_307;
assign n_692 = n_564 ^ n_309;
assign n_693 = n_565 ^ n_310;
assign n_694 = n_566 ^ n_310;
assign n_695 = n_567 ^ n_311;
assign n_696 = n_568 ^ n_313;
assign n_697 = n_569 ^ n_314;
assign n_698 = n_570 ^ n_314;
assign n_699 = n_571 ^ n_315;
assign n_700 = n_572 ^ n_317;
assign n_701 = n_573 ^ n_318;
assign n_702 = n_574 ^ n_318;
assign n_703 = n_575 ^ n_319;
assign n_704 = n_576 ^ n_321;
assign n_705 = n_577 ^ n_322;
assign n_706 = n_578 ^ n_322;
assign n_707 = n_579 ^ n_323;
assign n_708 = n_580 ^ n_325;
assign n_709 = n_581 ^ n_326;
assign n_710 = n_582 ^ n_326;
assign n_711 = n_583 ^ n_327;
assign n_712 = n_584 ^ n_329;
assign n_713 = n_585 ^ n_330;
assign n_714 = n_586 ^ n_330;
assign n_715 = n_587 ^ n_331;
assign n_716 = n_588 ^ n_333;
assign n_717 = n_589 ^ n_334;
assign n_718 = n_590 ^ n_334;
assign n_719 = n_591 ^ n_335;
assign n_720 = n_592 ^ n_337;
assign n_721 = n_593 ^ n_338;
assign n_722 = n_594 ^ n_338;
assign n_723 = n_595 ^ n_339;
assign n_724 = n_596 ^ n_341;
assign n_725 = n_597 ^ n_342;
assign n_726 = n_598 ^ n_342;
assign n_727 = n_599 ^ n_343;
assign n_728 = n_600 ^ n_345;
assign n_729 = n_601 ^ n_346;
assign n_730 = n_602 ^ n_346;
assign n_731 = n_603 ^ n_347;
assign n_732 = n_604 ^ n_349;
assign n_733 = n_605 ^ n_350;
assign n_734 = n_606 ^ n_350;
assign n_735 = n_607 ^ n_351;
assign n_736 = n_608 ^ n_353;
assign n_737 = n_609 ^ n_354;
assign n_738 = n_610 ^ n_354;
assign n_739 = n_611 ^ n_355;
assign n_740 = n_612 ^ n_357;
assign n_741 = n_613 ^ n_358;
assign n_742 = n_614 ^ n_358;
assign n_743 = n_615 ^ n_359;
assign n_744 = n_616 ^ n_361;
assign n_745 = n_617 ^ n_362;
assign n_746 = n_618 ^ n_362;
assign n_747 = n_619 ^ n_363;
assign n_748 = n_620 ^ n_365;
assign n_749 = n_621 ^ n_366;
assign n_750 = n_622 ^ n_366;
assign n_751 = n_623 ^ n_367;
assign n_752 = n_624 ^ n_369;
assign n_753 = n_625 ^ n_370;
assign n_754 = n_626 ^ n_370;
assign n_755 = n_627 ^ n_371;
assign n_756 = n_628 ^ n_373;
assign n_757 = n_629 ^ n_374;
assign n_758 = n_630 ^ n_374;
assign n_759 = n_631 ^ n_375;
assign n_760 = n_632 ^ n_377;
assign n_761 = n_633 ^ n_378;
assign n_762 = n_634 ^ n_378;
assign n_763 = n_635 ^ n_379;
assign n_764 = n_636 ^ n_380;
assign n_765 = n_637 ^ n_382;
assign n_766 = n_638 ^ n_380;
assign n_767 = n_639 ^ n_383;
assign n_768 = n_640 ^ n_648;
assign n_769 = n_649 ^ n_641;
assign n_770 = n_650 ^ n_642;
assign n_771 = n_651 ^ n_643;
assign n_772 = n_652 ^ n_644;
assign n_773 = n_653 ^ n_645;
assign n_774 = n_654 ^ n_646;
assign n_775 = n_655 ^ n_647;
assign n_776 = n_656 ^ n_648;
assign n_777 = n_657 ^ n_649;
assign n_778 = n_658 ^ n_650;
assign n_779 = n_659 ^ n_651;
assign n_780 = n_660 ^ n_652;
assign n_781 = n_661 ^ n_653;
assign n_782 = n_662 ^ n_654;
assign n_783 = n_663 ^ n_655;
assign n_784 = n_664 ^ n_656;
assign n_785 = n_665 ^ n_657;
assign n_786 = n_666 ^ n_658;
assign n_787 = n_667 ^ n_659;
assign n_788 = n_668 ^ n_660;
assign n_789 = n_669 ^ n_661;
assign n_790 = n_670 ^ n_662;
assign n_791 = n_671 ^ n_663;
assign n_792 = n_672 ^ n_664;
assign n_793 = n_665 ^ n_673;
assign n_794 = n_666 ^ n_674;
assign n_795 = n_667 ^ n_675;
assign n_796 = n_668 ^ n_676;
assign n_797 = n_669 ^ n_677;
assign n_798 = n_670 ^ n_678;
assign n_799 = n_671 ^ n_679;
assign n_800 = n_672 ^ n_680;
assign n_801 = n_681 ^ n_673;
assign n_802 = n_682 ^ n_674;
assign n_803 = n_683 ^ n_675;
assign n_804 = n_684 ^ n_676;
assign n_805 = n_685 ^ n_677;
assign n_806 = n_686 ^ n_678;
assign n_807 = n_687 ^ n_679;
assign n_808 = n_688 ^ n_680;
assign n_809 = n_689 ^ n_681;
assign n_810 = n_690 ^ n_682;
assign n_811 = n_691 ^ n_683;
assign n_812 = n_692 ^ n_684;
assign n_813 = n_693 ^ n_685;
assign n_814 = n_694 ^ n_686;
assign n_815 = n_695 ^ n_687;
assign n_816 = n_696 ^ n_688;
assign n_817 = n_697 ^ n_689;
assign n_818 = n_698 ^ n_690;
assign n_819 = n_699 ^ n_691;
assign n_820 = n_700 ^ n_692;
assign n_821 = n_701 ^ n_693;
assign n_822 = n_702 ^ n_694;
assign n_823 = n_703 ^ n_695;
assign n_824 = n_704 ^ n_696;
assign n_825 = n_705 ^ n_697;
assign n_826 = n_706 ^ n_698;
assign n_827 = n_707 ^ n_699;
assign n_828 = n_708 ^ n_700;
assign n_829 = n_709 ^ n_701;
assign n_830 = n_710 ^ n_702;
assign n_831 = n_711 ^ n_703;
assign n_832 = n_712 ^ n_704;
assign n_833 = n_713 ^ n_705;
assign n_834 = n_714 ^ n_706;
assign n_835 = n_715 ^ n_707;
assign n_836 = n_716 ^ n_708;
assign n_837 = n_717 ^ n_709;
assign n_838 = n_718 ^ n_710;
assign n_839 = n_719 ^ n_711;
assign n_840 = n_720 ^ n_712;
assign n_841 = n_721 ^ n_713;
assign n_842 = n_722 ^ n_714;
assign n_843 = n_723 ^ n_715;
assign n_844 = n_724 ^ n_716;
assign n_845 = n_725 ^ n_717;
assign n_846 = n_726 ^ n_718;
assign n_847 = n_727 ^ n_719;
assign n_848 = n_728 ^ n_720;
assign n_849 = n_729 ^ n_721;
assign n_850 = n_730 ^ n_722;
assign n_851 = n_731 ^ n_723;
assign n_852 = n_732 ^ n_724;
assign n_853 = n_733 ^ n_725;
assign n_854 = n_734 ^ n_726;
assign n_855 = n_735 ^ n_727;
assign n_856 = n_736 ^ n_728;
assign n_857 = n_729 ^ n_737;
assign n_858 = n_730 ^ n_738;
assign n_859 = n_731 ^ n_739;
assign n_860 = n_732 ^ n_740;
assign n_861 = n_733 ^ n_741;
assign n_862 = n_734 ^ n_742;
assign n_863 = n_735 ^ n_743;
assign n_864 = n_736 ^ n_744;
assign n_865 = n_745 ^ n_737;
assign n_866 = n_746 ^ n_738;
assign n_867 = n_747 ^ n_739;
assign n_868 = n_748 ^ n_740;
assign n_869 = n_749 ^ n_741;
assign n_870 = n_750 ^ n_742;
assign n_871 = n_751 ^ n_743;
assign n_872 = n_752 ^ n_744;
assign n_873 = n_753 ^ n_745;
assign n_874 = n_754 ^ n_746;
assign n_875 = n_755 ^ n_747;
assign n_876 = n_756 ^ n_748;
assign n_877 = n_757 ^ n_749;
assign n_878 = n_758 ^ n_750;
assign n_879 = n_759 ^ n_751;
assign n_880 = n_760 ^ n_640;
assign n_881 = n_760 ^ n_752;
assign n_882 = n_761 ^ n_753;
assign n_883 = n_761 ^ n_641;
assign n_884 = n_762 ^ n_754;
assign n_885 = n_762 ^ n_642;
assign n_886 = n_763 ^ n_755;
assign n_887 = n_763 ^ n_643;
assign n_888 = n_764 ^ n_757;
assign n_889 = n_764 ^ n_645;
assign n_890 = n_765 ^ n_756;
assign n_891 = n_765 ^ n_644;
assign n_892 = n_766 ^ n_758;
assign n_893 = n_766 ^ n_646;
assign n_894 = n_767 ^ n_759;
assign n_895 = n_767 ^ n_647;
assign n_896 = x131 & n_768;
assign n_897 = x131 & n_769;
assign n_898 = x131 & n_770;
assign n_899 = x131 & n_771;
assign n_900 = x131 & n_772;
assign n_901 = x131 & n_773;
assign n_902 = x131 & n_774;
assign n_903 = x131 & n_775;
assign n_904 = x131 & n_776;
assign n_905 = x131 & n_777;
assign n_906 = x131 & n_778;
assign n_907 = x131 & n_779;
assign n_908 = x131 & n_780;
assign n_909 = x131 & n_781;
assign n_910 = x131 & n_782;
assign n_911 = x131 & n_783;
assign n_912 = x131 & n_784;
assign n_913 = x131 & n_785;
assign n_914 = x131 & n_786;
assign n_915 = x131 & n_787;
assign n_916 = x131 & n_788;
assign n_917 = x131 & n_789;
assign n_918 = x131 & n_790;
assign n_919 = x131 & n_791;
assign n_920 = x131 & n_792;
assign n_921 = ~x131 & n_793;
assign n_922 = ~x131 & n_794;
assign n_923 = ~x131 & n_795;
assign n_924 = ~x131 & n_796;
assign n_925 = ~x131 & n_797;
assign n_926 = ~x131 & n_798;
assign n_927 = ~x131 & n_799;
assign n_928 = ~x131 & n_800;
assign n_929 = x131 & n_801;
assign n_930 = x131 & n_802;
assign n_931 = x131 & n_803;
assign n_932 = x131 & n_804;
assign n_933 = x131 & n_805;
assign n_934 = x131 & n_806;
assign n_935 = x131 & n_807;
assign n_936 = x131 & n_808;
assign n_937 = x131 & n_809;
assign n_938 = x131 & n_810;
assign n_939 = x131 & n_811;
assign n_940 = x131 & n_812;
assign n_941 = x131 & n_813;
assign n_942 = x131 & n_814;
assign n_943 = x131 & n_815;
assign n_944 = x131 & n_816;
assign n_945 = x131 & n_817;
assign n_946 = x131 & n_818;
assign n_947 = x131 & n_819;
assign n_948 = x131 & n_820;
assign n_949 = x131 & n_821;
assign n_950 = x131 & n_822;
assign n_951 = x131 & n_823;
assign n_952 = x131 & n_824;
assign n_953 = ~x131 & n_825;
assign n_954 = ~x131 & n_826;
assign n_955 = ~x131 & n_827;
assign n_956 = ~x131 & n_828;
assign n_957 = ~x131 & n_829;
assign n_958 = ~x131 & n_830;
assign n_959 = ~x131 & n_831;
assign n_960 = ~x131 & n_832;
assign n_961 = x131 & n_833;
assign n_962 = x131 & n_834;
assign n_963 = x131 & n_835;
assign n_964 = x131 & n_836;
assign n_965 = x131 & n_837;
assign n_966 = x131 & n_838;
assign n_967 = x131 & n_839;
assign n_968 = x131 & n_840;
assign n_969 = x131 & n_841;
assign n_970 = x131 & n_842;
assign n_971 = x131 & n_843;
assign n_972 = x131 & n_844;
assign n_973 = x131 & n_845;
assign n_974 = x131 & n_846;
assign n_975 = x131 & n_847;
assign n_976 = x131 & n_848;
assign n_977 = x131 & n_849;
assign n_978 = x131 & n_850;
assign n_979 = x131 & n_851;
assign n_980 = x131 & n_852;
assign n_981 = x131 & n_853;
assign n_982 = x131 & n_854;
assign n_983 = x131 & n_855;
assign n_984 = x131 & n_856;
assign n_985 = ~x131 & n_857;
assign n_986 = ~x131 & n_858;
assign n_987 = ~x131 & n_859;
assign n_988 = ~x131 & n_860;
assign n_989 = ~x131 & n_861;
assign n_990 = ~x131 & n_862;
assign n_991 = ~x131 & n_863;
assign n_992 = ~x131 & n_864;
assign n_993 = x131 & n_865;
assign n_994 = x131 & n_866;
assign n_995 = x131 & n_867;
assign n_996 = x131 & n_868;
assign n_997 = x131 & n_869;
assign n_998 = x131 & n_870;
assign n_999 = x131 & n_871;
assign n_1000 = x131 & n_872;
assign n_1001 = x131 & n_873;
assign n_1002 = x131 & n_874;
assign n_1003 = x131 & n_875;
assign n_1004 = x131 & n_876;
assign n_1005 = x131 & n_877;
assign n_1006 = x131 & n_878;
assign n_1007 = x131 & n_879;
assign n_1008 = x131 & n_880;
assign n_1009 = x131 & n_881;
assign n_1010 = x131 & n_882;
assign n_1011 = x131 & n_883;
assign n_1012 = x131 & n_884;
assign n_1013 = x131 & n_885;
assign n_1014 = x131 & n_886;
assign n_1015 = x131 & n_887;
assign n_1016 = x131 & n_888;
assign n_1017 = x131 & n_889;
assign n_1018 = x131 & n_890;
assign n_1019 = x131 & n_891;
assign n_1020 = x131 & n_892;
assign n_1021 = x131 & n_893;
assign n_1022 = x131 & n_894;
assign n_1023 = x131 & n_895;
assign n_1024 = n_896 ^ n_648;
assign n_1025 = n_897 ^ n_649;
assign n_1026 = n_898 ^ n_650;
assign n_1027 = n_899 ^ n_651;
assign n_1028 = n_900 ^ n_652;
assign n_1029 = n_901 ^ n_653;
assign n_1030 = n_902 ^ n_654;
assign n_1031 = n_903 ^ n_655;
assign n_1032 = n_904 ^ n_656;
assign n_1033 = n_905 ^ n_657;
assign n_1034 = n_906 ^ n_658;
assign n_1035 = n_907 ^ n_659;
assign n_1036 = n_908 ^ n_660;
assign n_1037 = n_909 ^ n_661;
assign n_1038 = n_910 ^ n_662;
assign n_1039 = n_911 ^ n_663;
assign n_1040 = n_912 ^ n_664;
assign n_1041 = n_913 ^ n_665;
assign n_1042 = n_914 ^ n_666;
assign n_1043 = n_915 ^ n_667;
assign n_1044 = n_916 ^ n_668;
assign n_1045 = n_917 ^ n_669;
assign n_1046 = n_918 ^ n_670;
assign n_1047 = n_919 ^ n_671;
assign n_1048 = n_920 ^ n_672;
assign n_1049 = n_921 ^ n_665;
assign n_1050 = n_922 ^ n_666;
assign n_1051 = n_923 ^ n_667;
assign n_1052 = n_924 ^ n_668;
assign n_1053 = n_925 ^ n_669;
assign n_1054 = n_926 ^ n_670;
assign n_1055 = n_927 ^ n_671;
assign n_1056 = n_928 ^ n_672;
assign n_1057 = n_929 ^ n_681;
assign n_1058 = n_930 ^ n_682;
assign n_1059 = n_931 ^ n_683;
assign n_1060 = n_932 ^ n_684;
assign n_1061 = n_933 ^ n_685;
assign n_1062 = n_934 ^ n_686;
assign n_1063 = n_935 ^ n_687;
assign n_1064 = n_936 ^ n_688;
assign n_1065 = n_937 ^ n_689;
assign n_1066 = n_938 ^ n_690;
assign n_1067 = n_939 ^ n_691;
assign n_1068 = n_940 ^ n_692;
assign n_1069 = n_941 ^ n_693;
assign n_1070 = n_942 ^ n_694;
assign n_1071 = n_943 ^ n_695;
assign n_1072 = n_944 ^ n_696;
assign n_1073 = n_945 ^ n_697;
assign n_1074 = n_946 ^ n_698;
assign n_1075 = n_947 ^ n_699;
assign n_1076 = n_948 ^ n_700;
assign n_1077 = n_949 ^ n_701;
assign n_1078 = n_950 ^ n_702;
assign n_1079 = n_951 ^ n_703;
assign n_1080 = n_952 ^ n_704;
assign n_1081 = n_953 ^ n_697;
assign n_1082 = n_954 ^ n_698;
assign n_1083 = n_955 ^ n_699;
assign n_1084 = n_956 ^ n_700;
assign n_1085 = n_957 ^ n_701;
assign n_1086 = n_958 ^ n_702;
assign n_1087 = n_959 ^ n_703;
assign n_1088 = n_960 ^ n_704;
assign n_1089 = n_961 ^ n_713;
assign n_1090 = n_962 ^ n_714;
assign n_1091 = n_963 ^ n_715;
assign n_1092 = n_964 ^ n_716;
assign n_1093 = n_965 ^ n_717;
assign n_1094 = n_966 ^ n_718;
assign n_1095 = n_967 ^ n_719;
assign n_1096 = n_968 ^ n_720;
assign n_1097 = n_969 ^ n_721;
assign n_1098 = n_970 ^ n_722;
assign n_1099 = n_971 ^ n_723;
assign n_1100 = n_972 ^ n_724;
assign n_1101 = n_973 ^ n_725;
assign n_1102 = n_974 ^ n_726;
assign n_1103 = n_975 ^ n_727;
assign n_1104 = n_976 ^ n_728;
assign n_1105 = n_977 ^ n_729;
assign n_1106 = n_978 ^ n_730;
assign n_1107 = n_979 ^ n_731;
assign n_1108 = n_980 ^ n_732;
assign n_1109 = n_981 ^ n_733;
assign n_1110 = n_982 ^ n_734;
assign n_1111 = n_983 ^ n_735;
assign n_1112 = n_984 ^ n_736;
assign n_1113 = n_985 ^ n_729;
assign n_1114 = n_986 ^ n_730;
assign n_1115 = n_987 ^ n_731;
assign n_1116 = n_988 ^ n_732;
assign n_1117 = n_989 ^ n_733;
assign n_1118 = n_990 ^ n_734;
assign n_1119 = n_991 ^ n_735;
assign n_1120 = n_992 ^ n_736;
assign n_1121 = n_993 ^ n_745;
assign n_1122 = n_994 ^ n_746;
assign n_1123 = n_995 ^ n_747;
assign n_1124 = n_996 ^ n_748;
assign n_1125 = n_997 ^ n_749;
assign n_1126 = n_998 ^ n_750;
assign n_1127 = n_999 ^ n_751;
assign n_1128 = n_1000 ^ n_752;
assign n_1129 = n_1001 ^ n_753;
assign n_1130 = n_1002 ^ n_754;
assign n_1131 = n_1003 ^ n_755;
assign n_1132 = n_1004 ^ n_756;
assign n_1133 = n_1005 ^ n_757;
assign n_1134 = n_1006 ^ n_758;
assign n_1135 = n_1007 ^ n_759;
assign n_1136 = n_1008 ^ n_640;
assign n_1137 = n_1009 ^ n_760;
assign n_1138 = n_1010 ^ n_761;
assign n_1139 = n_1011 ^ n_641;
assign n_1140 = n_1012 ^ n_762;
assign n_1141 = n_1013 ^ n_642;
assign n_1142 = n_1014 ^ n_763;
assign n_1143 = n_1015 ^ n_643;
assign n_1144 = n_1016 ^ n_764;
assign n_1145 = n_1017 ^ n_645;
assign n_1146 = n_1018 ^ n_765;
assign n_1147 = n_1019 ^ n_644;
assign n_1148 = n_1020 ^ n_766;
assign n_1149 = n_1021 ^ n_646;
assign n_1150 = n_1022 ^ n_767;
assign n_1151 = n_1023 ^ n_647;
assign n_1152 = n_1024 ^ n_1028;
assign n_1153 = n_1029 ^ n_1025;
assign n_1154 = n_1030 ^ n_1026;
assign n_1155 = n_1031 ^ n_1027;
assign n_1156 = n_1032 ^ n_1028;
assign n_1157 = n_1033 ^ n_1029;
assign n_1158 = n_1034 ^ n_1030;
assign n_1159 = n_1035 ^ n_1031;
assign n_1160 = n_1036 ^ n_1032;
assign n_1161 = n_1037 ^ n_1033;
assign n_1162 = n_1038 ^ n_1034;
assign n_1163 = n_1039 ^ n_1035;
assign n_1164 = n_1040 ^ n_1036;
assign n_1165 = n_1037 ^ n_1041;
assign n_1166 = n_1038 ^ n_1042;
assign n_1167 = n_1039 ^ n_1043;
assign n_1168 = n_1040 ^ n_1044;
assign n_1169 = n_1045 ^ n_1041;
assign n_1170 = n_1046 ^ n_1042;
assign n_1171 = n_1047 ^ n_1043;
assign n_1172 = n_1048 ^ n_1044;
assign n_1173 = n_1049 ^ n_1045;
assign n_1174 = n_1050 ^ n_1046;
assign n_1175 = n_1051 ^ n_1047;
assign n_1176 = n_1052 ^ n_1048;
assign n_1177 = n_1053 ^ n_1049;
assign n_1178 = n_1054 ^ n_1050;
assign n_1179 = n_1055 ^ n_1051;
assign n_1180 = n_1056 ^ n_1052;
assign n_1181 = n_1053 ^ n_1057;
assign n_1182 = n_1054 ^ n_1058;
assign n_1183 = n_1055 ^ n_1059;
assign n_1184 = n_1056 ^ n_1060;
assign n_1185 = n_1061 ^ n_1057;
assign n_1186 = n_1062 ^ n_1058;
assign n_1187 = n_1063 ^ n_1059;
assign n_1188 = n_1064 ^ n_1060;
assign n_1189 = n_1065 ^ n_1061;
assign n_1190 = n_1066 ^ n_1062;
assign n_1191 = n_1067 ^ n_1063;
assign n_1192 = n_1068 ^ n_1064;
assign n_1193 = n_1069 ^ n_1065;
assign n_1194 = n_1070 ^ n_1066;
assign n_1195 = n_1071 ^ n_1067;
assign n_1196 = n_1072 ^ n_1068;
assign n_1197 = n_1069 ^ n_1073;
assign n_1198 = n_1070 ^ n_1074;
assign n_1199 = n_1071 ^ n_1075;
assign n_1200 = n_1072 ^ n_1076;
assign n_1201 = n_1077 ^ n_1073;
assign n_1202 = n_1078 ^ n_1074;
assign n_1203 = n_1079 ^ n_1075;
assign n_1204 = n_1080 ^ n_1076;
assign n_1205 = n_1081 ^ n_1077;
assign n_1206 = n_1082 ^ n_1078;
assign n_1207 = n_1083 ^ n_1079;
assign n_1208 = n_1084 ^ n_1080;
assign n_1209 = n_1085 ^ n_1081;
assign n_1210 = n_1086 ^ n_1082;
assign n_1211 = n_1087 ^ n_1083;
assign n_1212 = n_1088 ^ n_1084;
assign n_1213 = n_1085 ^ n_1089;
assign n_1214 = n_1086 ^ n_1090;
assign n_1215 = n_1087 ^ n_1091;
assign n_1216 = n_1088 ^ n_1092;
assign n_1217 = n_1093 ^ n_1089;
assign n_1218 = n_1094 ^ n_1090;
assign n_1219 = n_1095 ^ n_1091;
assign n_1220 = n_1096 ^ n_1092;
assign n_1221 = n_1097 ^ n_1093;
assign n_1222 = n_1098 ^ n_1094;
assign n_1223 = n_1099 ^ n_1095;
assign n_1224 = n_1100 ^ n_1096;
assign n_1225 = n_1101 ^ n_1097;
assign n_1226 = n_1102 ^ n_1098;
assign n_1227 = n_1103 ^ n_1099;
assign n_1228 = n_1104 ^ n_1100;
assign n_1229 = n_1101 ^ n_1105;
assign n_1230 = n_1102 ^ n_1106;
assign n_1231 = n_1103 ^ n_1107;
assign n_1232 = n_1104 ^ n_1108;
assign n_1233 = n_1109 ^ n_1105;
assign n_1234 = n_1110 ^ n_1106;
assign n_1235 = n_1111 ^ n_1107;
assign n_1236 = n_1112 ^ n_1108;
assign n_1237 = n_1113 ^ n_1109;
assign n_1238 = n_1114 ^ n_1110;
assign n_1239 = n_1115 ^ n_1111;
assign n_1240 = n_1116 ^ n_1112;
assign n_1241 = n_1117 ^ n_1113;
assign n_1242 = n_1118 ^ n_1114;
assign n_1243 = n_1119 ^ n_1115;
assign n_1244 = n_1120 ^ n_1116;
assign n_1245 = n_1117 ^ n_1121;
assign n_1246 = n_1118 ^ n_1122;
assign n_1247 = n_1119 ^ n_1123;
assign n_1248 = n_1120 ^ n_1124;
assign n_1249 = n_1125 ^ n_1121;
assign n_1250 = n_1126 ^ n_1122;
assign n_1251 = n_1127 ^ n_1123;
assign n_1252 = n_1128 ^ n_1124;
assign n_1253 = n_1129 ^ n_1125;
assign n_1254 = n_1130 ^ n_1126;
assign n_1255 = n_1131 ^ n_1127;
assign n_1256 = n_1132 ^ n_1128;
assign n_1257 = n_1133 ^ n_1129;
assign n_1258 = n_1134 ^ n_1130;
assign n_1259 = n_1135 ^ n_1131;
assign n_1260 = n_1137 ^ n_1132;
assign n_1261 = n_1133 ^ n_1138;
assign n_1262 = n_1134 ^ n_1140;
assign n_1263 = n_1135 ^ n_1142;
assign n_1264 = n_1144 ^ n_1138;
assign n_1265 = n_1139 ^ n_1144;
assign n_1266 = n_1145 ^ n_1139;
assign n_1267 = n_1145 ^ n_1025;
assign n_1268 = n_1146 ^ n_1136;
assign n_1269 = n_1137 ^ n_1146;
assign n_1270 = n_1147 ^ n_1136;
assign n_1271 = n_1024 ^ n_1147;
assign n_1272 = n_1148 ^ n_1140;
assign n_1273 = n_1141 ^ n_1148;
assign n_1274 = n_1149 ^ n_1141;
assign n_1275 = n_1149 ^ n_1026;
assign n_1276 = n_1150 ^ n_1142;
assign n_1277 = n_1143 ^ n_1150;
assign n_1278 = n_1151 ^ n_1143;
assign n_1279 = n_1151 ^ n_1027;
assign n_1280 = x130 & n_1152;
assign n_1281 = x130 & n_1153;
assign n_1282 = x130 & n_1154;
assign n_1283 = x130 & n_1155;
assign n_1284 = x130 & n_1156;
assign n_1285 = ~x130 & n_1157;
assign n_1286 = ~x130 & n_1158;
assign n_1287 = ~x130 & n_1159;
assign n_1288 = ~x130 & n_1160;
assign n_1289 = ~x130 & n_1161;
assign n_1290 = ~x130 & n_1162;
assign n_1291 = ~x130 & n_1163;
assign n_1292 = ~x130 & n_1164;
assign n_1293 = x130 & n_1165;
assign n_1294 = x130 & n_1166;
assign n_1295 = x130 & n_1167;
assign n_1296 = x130 & n_1168;
assign n_1297 = x130 & n_1169;
assign n_1298 = x130 & n_1170;
assign n_1299 = x130 & n_1171;
assign n_1300 = x130 & n_1172;
assign n_1301 = ~x130 & n_1173;
assign n_1302 = ~x130 & n_1174;
assign n_1303 = ~x130 & n_1175;
assign n_1304 = ~x130 & n_1176;
assign n_1305 = ~x130 & n_1177;
assign n_1306 = ~x130 & n_1178;
assign n_1307 = ~x130 & n_1179;
assign n_1308 = ~x130 & n_1180;
assign n_1309 = x130 & n_1181;
assign n_1310 = x130 & n_1182;
assign n_1311 = x130 & n_1183;
assign n_1312 = x130 & n_1184;
assign n_1313 = x130 & n_1185;
assign n_1314 = x130 & n_1186;
assign n_1315 = x130 & n_1187;
assign n_1316 = x130 & n_1188;
assign n_1317 = ~x130 & n_1189;
assign n_1318 = ~x130 & n_1190;
assign n_1319 = ~x130 & n_1191;
assign n_1320 = ~x130 & n_1192;
assign n_1321 = ~x130 & n_1193;
assign n_1322 = ~x130 & n_1194;
assign n_1323 = ~x130 & n_1195;
assign n_1324 = ~x130 & n_1196;
assign n_1325 = x130 & n_1197;
assign n_1326 = x130 & n_1198;
assign n_1327 = x130 & n_1199;
assign n_1328 = x130 & n_1200;
assign n_1329 = x130 & n_1201;
assign n_1330 = x130 & n_1202;
assign n_1331 = x130 & n_1203;
assign n_1332 = x130 & n_1204;
assign n_1333 = ~x130 & n_1205;
assign n_1334 = ~x130 & n_1206;
assign n_1335 = ~x130 & n_1207;
assign n_1336 = ~x130 & n_1208;
assign n_1337 = ~x130 & n_1209;
assign n_1338 = ~x130 & n_1210;
assign n_1339 = ~x130 & n_1211;
assign n_1340 = ~x130 & n_1212;
assign n_1341 = x130 & n_1213;
assign n_1342 = x130 & n_1214;
assign n_1343 = x130 & n_1215;
assign n_1344 = x130 & n_1216;
assign n_1345 = x130 & n_1217;
assign n_1346 = x130 & n_1218;
assign n_1347 = x130 & n_1219;
assign n_1348 = x130 & n_1220;
assign n_1349 = ~x130 & n_1221;
assign n_1350 = ~x130 & n_1222;
assign n_1351 = ~x130 & n_1223;
assign n_1352 = ~x130 & n_1224;
assign n_1353 = ~x130 & n_1225;
assign n_1354 = ~x130 & n_1226;
assign n_1355 = ~x130 & n_1227;
assign n_1356 = ~x130 & n_1228;
assign n_1357 = x130 & n_1229;
assign n_1358 = x130 & n_1230;
assign n_1359 = x130 & n_1231;
assign n_1360 = x130 & n_1232;
assign n_1361 = x130 & n_1233;
assign n_1362 = x130 & n_1234;
assign n_1363 = x130 & n_1235;
assign n_1364 = x130 & n_1236;
assign n_1365 = ~x130 & n_1237;
assign n_1366 = ~x130 & n_1238;
assign n_1367 = ~x130 & n_1239;
assign n_1368 = ~x130 & n_1240;
assign n_1369 = ~x130 & n_1241;
assign n_1370 = ~x130 & n_1242;
assign n_1371 = ~x130 & n_1243;
assign n_1372 = ~x130 & n_1244;
assign n_1373 = x130 & n_1245;
assign n_1374 = x130 & n_1246;
assign n_1375 = x130 & n_1247;
assign n_1376 = x130 & n_1248;
assign n_1377 = x130 & n_1249;
assign n_1378 = x130 & n_1250;
assign n_1379 = x130 & n_1251;
assign n_1380 = x130 & n_1252;
assign n_1381 = ~x130 & n_1253;
assign n_1382 = ~x130 & n_1254;
assign n_1383 = ~x130 & n_1255;
assign n_1384 = ~x130 & n_1256;
assign n_1385 = ~x130 & n_1257;
assign n_1386 = ~x130 & n_1258;
assign n_1387 = ~x130 & n_1259;
assign n_1388 = ~x130 & n_1260;
assign n_1389 = x130 & n_1261;
assign n_1390 = x130 & n_1262;
assign n_1391 = x130 & n_1263;
assign n_1392 = x130 & n_1264;
assign n_1393 = ~x130 & n_1265;
assign n_1394 = ~x130 & n_1266;
assign n_1395 = x130 & n_1267;
assign n_1396 = x130 & n_1268;
assign n_1397 = x130 & n_1269;
assign n_1398 = ~x130 & n_1270;
assign n_1399 = ~x130 & n_1271;
assign n_1400 = x130 & n_1272;
assign n_1401 = ~x130 & n_1273;
assign n_1402 = ~x130 & n_1274;
assign n_1403 = x130 & n_1275;
assign n_1404 = x130 & n_1276;
assign n_1405 = ~x130 & n_1277;
assign n_1406 = ~x130 & n_1278;
assign n_1407 = x130 & n_1279;
assign n_1408 = n_1280 ^ n_1028;
assign n_1409 = n_1281 ^ n_1029;
assign n_1410 = n_1282 ^ n_1030;
assign n_1411 = n_1283 ^ n_1031;
assign n_1412 = n_1284 ^ n_1032;
assign n_1413 = n_1285 ^ n_1029;
assign n_1414 = n_1286 ^ n_1030;
assign n_1415 = n_1287 ^ n_1031;
assign n_1416 = n_1288 ^ n_1032;
assign n_1417 = n_1289 ^ n_1033;
assign n_1418 = n_1290 ^ n_1034;
assign n_1419 = n_1291 ^ n_1035;
assign n_1420 = n_1292 ^ n_1036;
assign n_1421 = n_1293 ^ n_1041;
assign n_1422 = n_1294 ^ n_1042;
assign n_1423 = n_1295 ^ n_1043;
assign n_1424 = n_1296 ^ n_1044;
assign n_1425 = n_1297 ^ n_1045;
assign n_1426 = n_1298 ^ n_1046;
assign n_1427 = n_1299 ^ n_1047;
assign n_1428 = n_1300 ^ n_1048;
assign n_1429 = n_1301 ^ n_1045;
assign n_1430 = n_1302 ^ n_1046;
assign n_1431 = n_1303 ^ n_1047;
assign n_1432 = n_1304 ^ n_1048;
assign n_1433 = n_1305 ^ n_1049;
assign n_1434 = n_1306 ^ n_1050;
assign n_1435 = n_1307 ^ n_1051;
assign n_1436 = n_1308 ^ n_1052;
assign n_1437 = n_1309 ^ n_1057;
assign n_1438 = n_1310 ^ n_1058;
assign n_1439 = n_1311 ^ n_1059;
assign n_1440 = n_1312 ^ n_1060;
assign n_1441 = n_1313 ^ n_1061;
assign n_1442 = n_1314 ^ n_1062;
assign n_1443 = n_1315 ^ n_1063;
assign n_1444 = n_1316 ^ n_1064;
assign n_1445 = n_1317 ^ n_1061;
assign n_1446 = n_1318 ^ n_1062;
assign n_1447 = n_1319 ^ n_1063;
assign n_1448 = n_1320 ^ n_1064;
assign n_1449 = n_1321 ^ n_1065;
assign n_1450 = n_1322 ^ n_1066;
assign n_1451 = n_1323 ^ n_1067;
assign n_1452 = n_1324 ^ n_1068;
assign n_1453 = n_1325 ^ n_1073;
assign n_1454 = n_1326 ^ n_1074;
assign n_1455 = n_1327 ^ n_1075;
assign n_1456 = n_1328 ^ n_1076;
assign n_1457 = n_1329 ^ n_1077;
assign n_1458 = n_1330 ^ n_1078;
assign n_1459 = n_1331 ^ n_1079;
assign n_1460 = n_1332 ^ n_1080;
assign n_1461 = n_1333 ^ n_1077;
assign n_1462 = n_1334 ^ n_1078;
assign n_1463 = n_1335 ^ n_1079;
assign n_1464 = n_1336 ^ n_1080;
assign n_1465 = n_1337 ^ n_1081;
assign n_1466 = n_1338 ^ n_1082;
assign n_1467 = n_1339 ^ n_1083;
assign n_1468 = n_1340 ^ n_1084;
assign n_1469 = n_1341 ^ n_1089;
assign n_1470 = n_1342 ^ n_1090;
assign n_1471 = n_1343 ^ n_1091;
assign n_1472 = n_1344 ^ n_1092;
assign n_1473 = n_1345 ^ n_1093;
assign n_1474 = n_1346 ^ n_1094;
assign n_1475 = n_1347 ^ n_1095;
assign n_1476 = n_1348 ^ n_1096;
assign n_1477 = n_1349 ^ n_1093;
assign n_1478 = n_1350 ^ n_1094;
assign n_1479 = n_1351 ^ n_1095;
assign n_1480 = n_1352 ^ n_1096;
assign n_1481 = n_1353 ^ n_1097;
assign n_1482 = n_1354 ^ n_1098;
assign n_1483 = n_1355 ^ n_1099;
assign n_1484 = n_1356 ^ n_1100;
assign n_1485 = n_1357 ^ n_1105;
assign n_1486 = n_1358 ^ n_1106;
assign n_1487 = n_1359 ^ n_1107;
assign n_1488 = n_1360 ^ n_1108;
assign n_1489 = n_1361 ^ n_1109;
assign n_1490 = n_1362 ^ n_1110;
assign n_1491 = n_1363 ^ n_1111;
assign n_1492 = n_1364 ^ n_1112;
assign n_1493 = n_1365 ^ n_1109;
assign n_1494 = n_1366 ^ n_1110;
assign n_1495 = n_1367 ^ n_1111;
assign n_1496 = n_1368 ^ n_1112;
assign n_1497 = n_1369 ^ n_1113;
assign n_1498 = n_1370 ^ n_1114;
assign n_1499 = n_1371 ^ n_1115;
assign n_1500 = n_1372 ^ n_1116;
assign n_1501 = n_1373 ^ n_1121;
assign n_1502 = n_1374 ^ n_1122;
assign n_1503 = n_1375 ^ n_1123;
assign n_1504 = n_1376 ^ n_1124;
assign n_1505 = n_1377 ^ n_1125;
assign n_1506 = n_1378 ^ n_1126;
assign n_1507 = n_1379 ^ n_1127;
assign n_1508 = n_1380 ^ n_1128;
assign n_1509 = n_1381 ^ n_1125;
assign n_1510 = n_1382 ^ n_1126;
assign n_1511 = n_1383 ^ n_1127;
assign n_1512 = n_1384 ^ n_1128;
assign n_1513 = n_1385 ^ n_1129;
assign n_1514 = n_1386 ^ n_1130;
assign n_1515 = n_1387 ^ n_1131;
assign n_1516 = n_1388 ^ n_1132;
assign n_1517 = n_1389 ^ n_1138;
assign n_1518 = n_1390 ^ n_1140;
assign n_1519 = n_1391 ^ n_1142;
assign n_1520 = n_1392 ^ n_1144;
assign n_1521 = n_1393 ^ n_1144;
assign n_1522 = n_1394 ^ n_1139;
assign n_1523 = n_1395 ^ n_1025;
assign n_1524 = n_1396 ^ n_1136;
assign n_1525 = n_1397 ^ n_1146;
assign n_1526 = n_1398 ^ n_1136;
assign n_1527 = n_1399 ^ n_1147;
assign n_1528 = n_1400 ^ n_1148;
assign n_1529 = n_1401 ^ n_1148;
assign n_1530 = n_1402 ^ n_1141;
assign n_1531 = n_1403 ^ n_1026;
assign n_1532 = n_1404 ^ n_1150;
assign n_1533 = n_1405 ^ n_1150;
assign n_1534 = n_1406 ^ n_1143;
assign n_1535 = n_1407 ^ n_1027;
assign n_1536 = n_1408 ^ n_1440;
assign n_1537 = n_1441 ^ n_1409;
assign n_1538 = n_1442 ^ n_1410;
assign n_1539 = n_1443 ^ n_1411;
assign n_1540 = n_1444 ^ n_1412;
assign n_1541 = n_1445 ^ n_1413;
assign n_1542 = n_1446 ^ n_1414;
assign n_1543 = n_1447 ^ n_1415;
assign n_1544 = n_1448 ^ n_1416;
assign n_1545 = n_1449 ^ n_1417;
assign n_1546 = n_1450 ^ n_1418;
assign n_1547 = n_1451 ^ n_1419;
assign n_1548 = n_1452 ^ n_1420;
assign n_1549 = n_1453 ^ n_1421;
assign n_1550 = n_1454 ^ n_1422;
assign n_1551 = n_1455 ^ n_1423;
assign n_1552 = n_1456 ^ n_1424;
assign n_1553 = n_1457 ^ n_1425;
assign n_1554 = n_1458 ^ n_1426;
assign n_1555 = n_1459 ^ n_1427;
assign n_1556 = n_1460 ^ n_1428;
assign n_1557 = n_1461 ^ n_1429;
assign n_1558 = n_1462 ^ n_1430;
assign n_1559 = n_1463 ^ n_1431;
assign n_1560 = n_1464 ^ n_1432;
assign n_1561 = n_1465 ^ n_1433;
assign n_1562 = n_1466 ^ n_1434;
assign n_1563 = n_1467 ^ n_1435;
assign n_1564 = n_1468 ^ n_1436;
assign n_1565 = n_1469 ^ n_1437;
assign n_1566 = n_1470 ^ n_1438;
assign n_1567 = n_1471 ^ n_1439;
assign n_1568 = n_1472 ^ n_1440;
assign n_1569 = n_1473 ^ n_1441;
assign n_1570 = n_1474 ^ n_1442;
assign n_1571 = n_1475 ^ n_1443;
assign n_1572 = n_1476 ^ n_1444;
assign n_1573 = n_1477 ^ n_1445;
assign n_1574 = n_1478 ^ n_1446;
assign n_1575 = n_1479 ^ n_1447;
assign n_1576 = n_1480 ^ n_1448;
assign n_1577 = n_1481 ^ n_1449;
assign n_1578 = n_1482 ^ n_1450;
assign n_1579 = n_1483 ^ n_1451;
assign n_1580 = n_1484 ^ n_1452;
assign n_1581 = n_1485 ^ n_1453;
assign n_1582 = n_1486 ^ n_1454;
assign n_1583 = n_1487 ^ n_1455;
assign n_1584 = n_1488 ^ n_1456;
assign n_1585 = n_1489 ^ n_1457;
assign n_1586 = n_1490 ^ n_1458;
assign n_1587 = n_1491 ^ n_1459;
assign n_1588 = n_1492 ^ n_1460;
assign n_1589 = n_1493 ^ n_1461;
assign n_1590 = n_1494 ^ n_1462;
assign n_1591 = n_1495 ^ n_1463;
assign n_1592 = n_1496 ^ n_1464;
assign n_1593 = n_1497 ^ n_1465;
assign n_1594 = n_1498 ^ n_1466;
assign n_1595 = n_1499 ^ n_1467;
assign n_1596 = n_1500 ^ n_1468;
assign n_1597 = n_1501 ^ n_1469;
assign n_1598 = n_1502 ^ n_1470;
assign n_1599 = n_1503 ^ n_1471;
assign n_1600 = n_1504 ^ n_1408;
assign n_1601 = n_1504 ^ n_1472;
assign n_1602 = n_1505 ^ n_1473;
assign n_1603 = n_1505 ^ n_1409;
assign n_1604 = n_1506 ^ n_1474;
assign n_1605 = n_1506 ^ n_1410;
assign n_1606 = n_1507 ^ n_1475;
assign n_1607 = n_1507 ^ n_1411;
assign n_1608 = n_1508 ^ n_1476;
assign n_1609 = n_1508 ^ n_1412;
assign n_1610 = n_1509 ^ n_1477;
assign n_1611 = n_1509 ^ n_1413;
assign n_1612 = n_1510 ^ n_1478;
assign n_1613 = n_1510 ^ n_1414;
assign n_1614 = n_1511 ^ n_1479;
assign n_1615 = n_1511 ^ n_1415;
assign n_1616 = n_1512 ^ n_1480;
assign n_1617 = n_1512 ^ n_1416;
assign n_1618 = n_1513 ^ n_1481;
assign n_1619 = n_1513 ^ n_1417;
assign n_1620 = n_1514 ^ n_1482;
assign n_1621 = n_1514 ^ n_1418;
assign n_1622 = n_1515 ^ n_1483;
assign n_1623 = n_1515 ^ n_1419;
assign n_1624 = n_1516 ^ n_1484;
assign n_1625 = n_1516 ^ n_1420;
assign n_1626 = n_1517 ^ n_1485;
assign n_1627 = n_1517 ^ n_1421;
assign n_1628 = n_1518 ^ n_1486;
assign n_1629 = n_1518 ^ n_1422;
assign n_1630 = n_1519 ^ n_1487;
assign n_1631 = n_1519 ^ n_1423;
assign n_1632 = n_1520 ^ n_1489;
assign n_1633 = n_1520 ^ n_1425;
assign n_1634 = n_1521 ^ n_1493;
assign n_1635 = n_1521 ^ n_1429;
assign n_1636 = n_1522 ^ n_1497;
assign n_1637 = n_1522 ^ n_1433;
assign n_1638 = n_1523 ^ n_1501;
assign n_1639 = n_1523 ^ n_1437;
assign n_1640 = n_1524 ^ n_1492;
assign n_1641 = n_1524 ^ n_1428;
assign n_1642 = n_1525 ^ n_1488;
assign n_1643 = n_1525 ^ n_1424;
assign n_1644 = n_1526 ^ n_1496;
assign n_1645 = n_1526 ^ n_1432;
assign n_1646 = n_1527 ^ n_1500;
assign n_1647 = n_1527 ^ n_1436;
assign n_1648 = n_1528 ^ n_1490;
assign n_1649 = n_1528 ^ n_1426;
assign n_1650 = n_1529 ^ n_1494;
assign n_1651 = n_1529 ^ n_1430;
assign n_1652 = n_1530 ^ n_1498;
assign n_1653 = n_1530 ^ n_1434;
assign n_1654 = n_1531 ^ n_1502;
assign n_1655 = n_1531 ^ n_1438;
assign n_1656 = n_1532 ^ n_1491;
assign n_1657 = n_1532 ^ n_1427;
assign n_1658 = n_1533 ^ n_1495;
assign n_1659 = n_1533 ^ n_1431;
assign n_1660 = n_1534 ^ n_1499;
assign n_1661 = n_1534 ^ n_1435;
assign n_1662 = n_1535 ^ n_1503;
assign n_1663 = n_1535 ^ n_1439;
assign n_1664 = x133 & n_1536;
assign n_1665 = x133 & n_1537;
assign n_1666 = x133 & n_1538;
assign n_1667 = x133 & n_1539;
assign n_1668 = x133 & n_1540;
assign n_1669 = x133 & n_1541;
assign n_1670 = x133 & n_1542;
assign n_1671 = x133 & n_1543;
assign n_1672 = x133 & n_1544;
assign n_1673 = x133 & n_1545;
assign n_1674 = x133 & n_1546;
assign n_1675 = x133 & n_1547;
assign n_1676 = x133 & n_1548;
assign n_1677 = x133 & n_1549;
assign n_1678 = x133 & n_1550;
assign n_1679 = x133 & n_1551;
assign n_1680 = x133 & n_1552;
assign n_1681 = x133 & n_1553;
assign n_1682 = x133 & n_1554;
assign n_1683 = x133 & n_1555;
assign n_1684 = x133 & n_1556;
assign n_1685 = x133 & n_1557;
assign n_1686 = x133 & n_1558;
assign n_1687 = x133 & n_1559;
assign n_1688 = x133 & n_1560;
assign n_1689 = x133 & n_1561;
assign n_1690 = x133 & n_1562;
assign n_1691 = x133 & n_1563;
assign n_1692 = x133 & n_1564;
assign n_1693 = x133 & n_1565;
assign n_1694 = x133 & n_1566;
assign n_1695 = x133 & n_1567;
assign n_1696 = x133 & n_1568;
assign n_1697 = ~x133 & n_1569;
assign n_1698 = ~x133 & n_1570;
assign n_1699 = ~x133 & n_1571;
assign n_1700 = ~x133 & n_1572;
assign n_1701 = ~x133 & n_1573;
assign n_1702 = ~x133 & n_1574;
assign n_1703 = ~x133 & n_1575;
assign n_1704 = ~x133 & n_1576;
assign n_1705 = ~x133 & n_1577;
assign n_1706 = ~x133 & n_1578;
assign n_1707 = ~x133 & n_1579;
assign n_1708 = ~x133 & n_1580;
assign n_1709 = ~x133 & n_1581;
assign n_1710 = ~x133 & n_1582;
assign n_1711 = ~x133 & n_1583;
assign n_1712 = ~x133 & n_1584;
assign n_1713 = ~x133 & n_1585;
assign n_1714 = ~x133 & n_1586;
assign n_1715 = ~x133 & n_1587;
assign n_1716 = ~x133 & n_1588;
assign n_1717 = ~x133 & n_1589;
assign n_1718 = ~x133 & n_1590;
assign n_1719 = ~x133 & n_1591;
assign n_1720 = ~x133 & n_1592;
assign n_1721 = ~x133 & n_1593;
assign n_1722 = ~x133 & n_1594;
assign n_1723 = ~x133 & n_1595;
assign n_1724 = ~x133 & n_1596;
assign n_1725 = ~x133 & n_1597;
assign n_1726 = ~x133 & n_1598;
assign n_1727 = ~x133 & n_1599;
assign n_1728 = x133 & n_1600;
assign n_1729 = ~x133 & n_1601;
assign n_1730 = x133 & n_1602;
assign n_1731 = x133 & n_1603;
assign n_1732 = x133 & n_1604;
assign n_1733 = x133 & n_1605;
assign n_1734 = x133 & n_1606;
assign n_1735 = x133 & n_1607;
assign n_1736 = x133 & n_1608;
assign n_1737 = x133 & n_1609;
assign n_1738 = x133 & n_1610;
assign n_1739 = x133 & n_1611;
assign n_1740 = x133 & n_1612;
assign n_1741 = x133 & n_1613;
assign n_1742 = x133 & n_1614;
assign n_1743 = x133 & n_1615;
assign n_1744 = x133 & n_1616;
assign n_1745 = x133 & n_1617;
assign n_1746 = x133 & n_1618;
assign n_1747 = x133 & n_1619;
assign n_1748 = x133 & n_1620;
assign n_1749 = x133 & n_1621;
assign n_1750 = x133 & n_1622;
assign n_1751 = x133 & n_1623;
assign n_1752 = x133 & n_1624;
assign n_1753 = x133 & n_1625;
assign n_1754 = x133 & n_1626;
assign n_1755 = x133 & n_1627;
assign n_1756 = x133 & n_1628;
assign n_1757 = x133 & n_1629;
assign n_1758 = x133 & n_1630;
assign n_1759 = x133 & n_1631;
assign n_1760 = x133 & n_1632;
assign n_1761 = x133 & n_1633;
assign n_1762 = x133 & n_1634;
assign n_1763 = x133 & n_1635;
assign n_1764 = x133 & n_1636;
assign n_1765 = x133 & n_1637;
assign n_1766 = x133 & n_1638;
assign n_1767 = x133 & n_1639;
assign n_1768 = x133 & n_1640;
assign n_1769 = x133 & n_1641;
assign n_1770 = x133 & n_1642;
assign n_1771 = x133 & n_1643;
assign n_1772 = x133 & n_1644;
assign n_1773 = x133 & n_1645;
assign n_1774 = x133 & n_1646;
assign n_1775 = x133 & n_1647;
assign n_1776 = x133 & n_1648;
assign n_1777 = x133 & n_1649;
assign n_1778 = x133 & n_1650;
assign n_1779 = x133 & n_1651;
assign n_1780 = x133 & n_1652;
assign n_1781 = x133 & n_1653;
assign n_1782 = x133 & n_1654;
assign n_1783 = x133 & n_1655;
assign n_1784 = x133 & n_1656;
assign n_1785 = x133 & n_1657;
assign n_1786 = x133 & n_1658;
assign n_1787 = x133 & n_1659;
assign n_1788 = x133 & n_1660;
assign n_1789 = x133 & n_1661;
assign n_1790 = x133 & n_1662;
assign n_1791 = x133 & n_1663;
assign n_1792 = n_1664 ^ n_1440;
assign n_1793 = n_1665 ^ n_1441;
assign n_1794 = n_1666 ^ n_1442;
assign n_1795 = n_1667 ^ n_1443;
assign n_1796 = n_1668 ^ n_1444;
assign n_1797 = n_1669 ^ n_1445;
assign n_1798 = n_1670 ^ n_1446;
assign n_1799 = n_1671 ^ n_1447;
assign n_1800 = n_1672 ^ n_1448;
assign n_1801 = n_1673 ^ n_1449;
assign n_1802 = n_1674 ^ n_1450;
assign n_1803 = n_1675 ^ n_1451;
assign n_1804 = n_1676 ^ n_1452;
assign n_1805 = n_1677 ^ n_1453;
assign n_1806 = n_1678 ^ n_1454;
assign n_1807 = n_1679 ^ n_1455;
assign n_1808 = n_1680 ^ n_1456;
assign n_1809 = n_1681 ^ n_1457;
assign n_1810 = n_1682 ^ n_1458;
assign n_1811 = n_1683 ^ n_1459;
assign n_1812 = n_1684 ^ n_1460;
assign n_1813 = n_1685 ^ n_1461;
assign n_1814 = n_1686 ^ n_1462;
assign n_1815 = n_1687 ^ n_1463;
assign n_1816 = n_1688 ^ n_1464;
assign n_1817 = n_1689 ^ n_1465;
assign n_1818 = n_1690 ^ n_1466;
assign n_1819 = n_1691 ^ n_1467;
assign n_1820 = n_1692 ^ n_1468;
assign n_1821 = n_1693 ^ n_1469;
assign n_1822 = n_1694 ^ n_1470;
assign n_1823 = n_1695 ^ n_1471;
assign n_1824 = n_1696 ^ n_1472;
assign n_1825 = n_1697 ^ n_1441;
assign n_1826 = n_1698 ^ n_1442;
assign n_1827 = n_1699 ^ n_1443;
assign n_1828 = n_1700 ^ n_1444;
assign n_1829 = n_1701 ^ n_1445;
assign n_1830 = n_1702 ^ n_1446;
assign n_1831 = n_1703 ^ n_1447;
assign n_1832 = n_1704 ^ n_1448;
assign n_1833 = n_1705 ^ n_1449;
assign n_1834 = n_1706 ^ n_1450;
assign n_1835 = n_1707 ^ n_1451;
assign n_1836 = n_1708 ^ n_1452;
assign n_1837 = n_1709 ^ n_1453;
assign n_1838 = n_1710 ^ n_1454;
assign n_1839 = n_1711 ^ n_1455;
assign n_1840 = n_1712 ^ n_1456;
assign n_1841 = n_1713 ^ n_1457;
assign n_1842 = n_1714 ^ n_1458;
assign n_1843 = n_1715 ^ n_1459;
assign n_1844 = n_1716 ^ n_1460;
assign n_1845 = n_1717 ^ n_1461;
assign n_1846 = n_1718 ^ n_1462;
assign n_1847 = n_1719 ^ n_1463;
assign n_1848 = n_1720 ^ n_1464;
assign n_1849 = n_1721 ^ n_1465;
assign n_1850 = n_1722 ^ n_1466;
assign n_1851 = n_1723 ^ n_1467;
assign n_1852 = n_1724 ^ n_1468;
assign n_1853 = n_1725 ^ n_1469;
assign n_1854 = n_1726 ^ n_1470;
assign n_1855 = n_1727 ^ n_1471;
assign n_1856 = n_1728 ^ n_1408;
assign n_1857 = n_1729 ^ n_1472;
assign n_1858 = n_1730 ^ n_1505;
assign n_1859 = n_1731 ^ n_1409;
assign n_1860 = n_1732 ^ n_1506;
assign n_1861 = n_1733 ^ n_1410;
assign n_1862 = n_1734 ^ n_1507;
assign n_1863 = n_1735 ^ n_1411;
assign n_1864 = n_1736 ^ n_1508;
assign n_1865 = n_1737 ^ n_1412;
assign n_1866 = n_1738 ^ n_1509;
assign n_1867 = n_1739 ^ n_1413;
assign n_1868 = n_1740 ^ n_1510;
assign n_1869 = n_1741 ^ n_1414;
assign n_1870 = n_1742 ^ n_1511;
assign n_1871 = n_1743 ^ n_1415;
assign n_1872 = n_1744 ^ n_1512;
assign n_1873 = n_1745 ^ n_1416;
assign n_1874 = n_1746 ^ n_1513;
assign n_1875 = n_1747 ^ n_1417;
assign n_1876 = n_1748 ^ n_1514;
assign n_1877 = n_1749 ^ n_1418;
assign n_1878 = n_1750 ^ n_1515;
assign n_1879 = n_1751 ^ n_1419;
assign n_1880 = n_1752 ^ n_1516;
assign n_1881 = n_1753 ^ n_1420;
assign n_1882 = n_1754 ^ n_1517;
assign n_1883 = n_1755 ^ n_1421;
assign n_1884 = n_1756 ^ n_1518;
assign n_1885 = n_1757 ^ n_1422;
assign n_1886 = n_1758 ^ n_1519;
assign n_1887 = n_1759 ^ n_1423;
assign n_1888 = n_1760 ^ n_1520;
assign n_1889 = n_1761 ^ n_1425;
assign n_1890 = n_1762 ^ n_1521;
assign n_1891 = n_1763 ^ n_1429;
assign n_1892 = n_1764 ^ n_1522;
assign n_1893 = n_1765 ^ n_1433;
assign n_1894 = n_1766 ^ n_1523;
assign n_1895 = n_1767 ^ n_1437;
assign n_1896 = n_1768 ^ n_1524;
assign n_1897 = n_1769 ^ n_1428;
assign n_1898 = n_1770 ^ n_1525;
assign n_1899 = n_1771 ^ n_1424;
assign n_1900 = n_1772 ^ n_1526;
assign n_1901 = n_1773 ^ n_1432;
assign n_1902 = n_1774 ^ n_1527;
assign n_1903 = n_1775 ^ n_1436;
assign n_1904 = n_1776 ^ n_1528;
assign n_1905 = n_1777 ^ n_1426;
assign n_1906 = n_1778 ^ n_1529;
assign n_1907 = n_1779 ^ n_1430;
assign n_1908 = n_1780 ^ n_1530;
assign n_1909 = n_1781 ^ n_1434;
assign n_1910 = n_1782 ^ n_1531;
assign n_1911 = n_1783 ^ n_1438;
assign n_1912 = n_1784 ^ n_1532;
assign n_1913 = n_1785 ^ n_1427;
assign n_1914 = n_1786 ^ n_1533;
assign n_1915 = n_1787 ^ n_1431;
assign n_1916 = n_1788 ^ n_1534;
assign n_1917 = n_1789 ^ n_1435;
assign n_1918 = n_1790 ^ n_1535;
assign n_1919 = n_1791 ^ n_1439;
assign n_1920 = n_1792 ^ n_1808;
assign n_1921 = n_1809 ^ n_1793;
assign n_1922 = n_1810 ^ n_1794;
assign n_1923 = n_1811 ^ n_1795;
assign n_1924 = n_1812 ^ n_1796;
assign n_1925 = n_1813 ^ n_1797;
assign n_1926 = n_1814 ^ n_1798;
assign n_1927 = n_1815 ^ n_1799;
assign n_1928 = n_1816 ^ n_1800;
assign n_1929 = n_1817 ^ n_1801;
assign n_1930 = n_1818 ^ n_1802;
assign n_1931 = n_1819 ^ n_1803;
assign n_1932 = n_1820 ^ n_1804;
assign n_1933 = n_1821 ^ n_1805;
assign n_1934 = n_1822 ^ n_1806;
assign n_1935 = n_1823 ^ n_1807;
assign n_1936 = n_1824 ^ n_1808;
assign n_1937 = n_1825 ^ n_1809;
assign n_1938 = n_1826 ^ n_1810;
assign n_1939 = n_1827 ^ n_1811;
assign n_1940 = n_1828 ^ n_1812;
assign n_1941 = n_1829 ^ n_1813;
assign n_1942 = n_1830 ^ n_1814;
assign n_1943 = n_1831 ^ n_1815;
assign n_1944 = n_1832 ^ n_1816;
assign n_1945 = n_1833 ^ n_1817;
assign n_1946 = n_1834 ^ n_1818;
assign n_1947 = n_1835 ^ n_1819;
assign n_1948 = n_1836 ^ n_1820;
assign n_1949 = n_1837 ^ n_1821;
assign n_1950 = n_1838 ^ n_1822;
assign n_1951 = n_1839 ^ n_1823;
assign n_1952 = n_1840 ^ n_1824;
assign n_1953 = n_1841 ^ n_1825;
assign n_1954 = n_1842 ^ n_1826;
assign n_1955 = n_1843 ^ n_1827;
assign n_1956 = n_1844 ^ n_1828;
assign n_1957 = n_1845 ^ n_1829;
assign n_1958 = n_1846 ^ n_1830;
assign n_1959 = n_1847 ^ n_1831;
assign n_1960 = n_1848 ^ n_1832;
assign n_1961 = n_1849 ^ n_1833;
assign n_1962 = n_1850 ^ n_1834;
assign n_1963 = n_1851 ^ n_1835;
assign n_1964 = n_1852 ^ n_1836;
assign n_1965 = n_1853 ^ n_1837;
assign n_1966 = n_1854 ^ n_1838;
assign n_1967 = n_1855 ^ n_1839;
assign n_1968 = n_1857 ^ n_1840;
assign n_1969 = n_1841 ^ n_1858;
assign n_1970 = n_1842 ^ n_1860;
assign n_1971 = n_1843 ^ n_1862;
assign n_1972 = n_1844 ^ n_1864;
assign n_1973 = n_1845 ^ n_1866;
assign n_1974 = n_1846 ^ n_1868;
assign n_1975 = n_1847 ^ n_1870;
assign n_1976 = n_1848 ^ n_1872;
assign n_1977 = n_1849 ^ n_1874;
assign n_1978 = n_1850 ^ n_1876;
assign n_1979 = n_1851 ^ n_1878;
assign n_1980 = n_1852 ^ n_1880;
assign n_1981 = n_1853 ^ n_1882;
assign n_1982 = n_1854 ^ n_1884;
assign n_1983 = n_1855 ^ n_1886;
assign n_1984 = n_1888 ^ n_1858;
assign n_1985 = n_1859 ^ n_1888;
assign n_1986 = n_1889 ^ n_1859;
assign n_1987 = n_1889 ^ n_1793;
assign n_1988 = n_1890 ^ n_1866;
assign n_1989 = n_1867 ^ n_1890;
assign n_1990 = n_1891 ^ n_1867;
assign n_1991 = n_1891 ^ n_1797;
assign n_1992 = n_1892 ^ n_1874;
assign n_1993 = n_1875 ^ n_1892;
assign n_1994 = n_1893 ^ n_1875;
assign n_1995 = n_1893 ^ n_1801;
assign n_1996 = n_1894 ^ n_1882;
assign n_1997 = n_1883 ^ n_1894;
assign n_1998 = n_1895 ^ n_1883;
assign n_1999 = n_1895 ^ n_1805;
assign n_2000 = n_1896 ^ n_1864;
assign n_2001 = n_1865 ^ n_1896;
assign n_2002 = n_1897 ^ n_1865;
assign n_2003 = n_1897 ^ n_1796;
assign n_2004 = n_1898 ^ n_1856;
assign n_2005 = n_1857 ^ n_1898;
assign n_2006 = n_1899 ^ n_1856;
assign n_2007 = n_1792 ^ n_1899;
assign n_2008 = n_1900 ^ n_1872;
assign n_2009 = n_1873 ^ n_1900;
assign n_2010 = n_1901 ^ n_1873;
assign n_2011 = n_1901 ^ n_1800;
assign n_2012 = n_1902 ^ n_1880;
assign n_2013 = n_1881 ^ n_1902;
assign n_2014 = n_1903 ^ n_1881;
assign n_2015 = n_1903 ^ n_1804;
assign n_2016 = n_1904 ^ n_1860;
assign n_2017 = n_1861 ^ n_1904;
assign n_2018 = n_1905 ^ n_1861;
assign n_2019 = n_1905 ^ n_1794;
assign n_2020 = n_1906 ^ n_1868;
assign n_2021 = n_1869 ^ n_1906;
assign n_2022 = n_1907 ^ n_1869;
assign n_2023 = n_1907 ^ n_1798;
assign n_2024 = n_1908 ^ n_1876;
assign n_2025 = n_1877 ^ n_1908;
assign n_2026 = n_1909 ^ n_1877;
assign n_2027 = n_1909 ^ n_1802;
assign n_2028 = n_1910 ^ n_1884;
assign n_2029 = n_1885 ^ n_1910;
assign n_2030 = n_1911 ^ n_1885;
assign n_2031 = n_1911 ^ n_1806;
assign n_2032 = n_1912 ^ n_1862;
assign n_2033 = n_1863 ^ n_1912;
assign n_2034 = n_1913 ^ n_1863;
assign n_2035 = n_1913 ^ n_1795;
assign n_2036 = n_1914 ^ n_1870;
assign n_2037 = n_1871 ^ n_1914;
assign n_2038 = n_1915 ^ n_1871;
assign n_2039 = n_1915 ^ n_1799;
assign n_2040 = n_1916 ^ n_1878;
assign n_2041 = n_1879 ^ n_1916;
assign n_2042 = n_1917 ^ n_1879;
assign n_2043 = n_1917 ^ n_1803;
assign n_2044 = n_1918 ^ n_1886;
assign n_2045 = n_1887 ^ n_1918;
assign n_2046 = n_1919 ^ n_1887;
assign n_2047 = n_1919 ^ n_1807;
assign n_2048 = x132 & n_1920;
assign n_2049 = x132 & n_1921;
assign n_2050 = x132 & n_1922;
assign n_2051 = x132 & n_1923;
assign n_2052 = x132 & n_1924;
assign n_2053 = x132 & n_1925;
assign n_2054 = x132 & n_1926;
assign n_2055 = x132 & n_1927;
assign n_2056 = x132 & n_1928;
assign n_2057 = x132 & n_1929;
assign n_2058 = x132 & n_1930;
assign n_2059 = x132 & n_1931;
assign n_2060 = x132 & n_1932;
assign n_2061 = x132 & n_1933;
assign n_2062 = x132 & n_1934;
assign n_2063 = x132 & n_1935;
assign n_2064 = x132 & n_1936;
assign n_2065 = ~x132 & n_1937;
assign n_2066 = ~x132 & n_1938;
assign n_2067 = ~x132 & n_1939;
assign n_2068 = ~x132 & n_1940;
assign n_2069 = ~x132 & n_1941;
assign n_2070 = ~x132 & n_1942;
assign n_2071 = ~x132 & n_1943;
assign n_2072 = ~x132 & n_1944;
assign n_2073 = ~x132 & n_1945;
assign n_2074 = ~x132 & n_1946;
assign n_2075 = ~x132 & n_1947;
assign n_2076 = ~x132 & n_1948;
assign n_2077 = ~x132 & n_1949;
assign n_2078 = ~x132 & n_1950;
assign n_2079 = ~x132 & n_1951;
assign n_2080 = ~x132 & n_1952;
assign n_2081 = ~x132 & n_1953;
assign n_2082 = ~x132 & n_1954;
assign n_2083 = ~x132 & n_1955;
assign n_2084 = ~x132 & n_1956;
assign n_2085 = ~x132 & n_1957;
assign n_2086 = ~x132 & n_1958;
assign n_2087 = ~x132 & n_1959;
assign n_2088 = ~x132 & n_1960;
assign n_2089 = ~x132 & n_1961;
assign n_2090 = ~x132 & n_1962;
assign n_2091 = ~x132 & n_1963;
assign n_2092 = ~x132 & n_1964;
assign n_2093 = ~x132 & n_1965;
assign n_2094 = ~x132 & n_1966;
assign n_2095 = ~x132 & n_1967;
assign n_2096 = ~x132 & n_1968;
assign n_2097 = x132 & n_1969;
assign n_2098 = x132 & n_1970;
assign n_2099 = x132 & n_1971;
assign n_2100 = x132 & n_1972;
assign n_2101 = x132 & n_1973;
assign n_2102 = x132 & n_1974;
assign n_2103 = x132 & n_1975;
assign n_2104 = x132 & n_1976;
assign n_2105 = x132 & n_1977;
assign n_2106 = x132 & n_1978;
assign n_2107 = x132 & n_1979;
assign n_2108 = x132 & n_1980;
assign n_2109 = x132 & n_1981;
assign n_2110 = x132 & n_1982;
assign n_2111 = x132 & n_1983;
assign n_2112 = x132 & n_1984;
assign n_2113 = ~x132 & n_1985;
assign n_2114 = ~x132 & n_1986;
assign n_2115 = x132 & n_1987;
assign n_2116 = x132 & n_1988;
assign n_2117 = ~x132 & n_1989;
assign n_2118 = ~x132 & n_1990;
assign n_2119 = x132 & n_1991;
assign n_2120 = x132 & n_1992;
assign n_2121 = ~x132 & n_1993;
assign n_2122 = ~x132 & n_1994;
assign n_2123 = x132 & n_1995;
assign n_2124 = x132 & n_1996;
assign n_2125 = ~x132 & n_1997;
assign n_2126 = ~x132 & n_1998;
assign n_2127 = x132 & n_1999;
assign n_2128 = x132 & n_2000;
assign n_2129 = ~x132 & n_2001;
assign n_2130 = ~x132 & n_2002;
assign n_2131 = x132 & n_2003;
assign n_2132 = x132 & n_2004;
assign n_2133 = x132 & n_2005;
assign n_2134 = ~x132 & n_2006;
assign n_2135 = ~x132 & n_2007;
assign n_2136 = x132 & n_2008;
assign n_2137 = ~x132 & n_2009;
assign n_2138 = ~x132 & n_2010;
assign n_2139 = x132 & n_2011;
assign n_2140 = x132 & n_2012;
assign n_2141 = ~x132 & n_2013;
assign n_2142 = ~x132 & n_2014;
assign n_2143 = x132 & n_2015;
assign n_2144 = x132 & n_2016;
assign n_2145 = ~x132 & n_2017;
assign n_2146 = ~x132 & n_2018;
assign n_2147 = x132 & n_2019;
assign n_2148 = x132 & n_2020;
assign n_2149 = ~x132 & n_2021;
assign n_2150 = ~x132 & n_2022;
assign n_2151 = x132 & n_2023;
assign n_2152 = x132 & n_2024;
assign n_2153 = ~x132 & n_2025;
assign n_2154 = ~x132 & n_2026;
assign n_2155 = x132 & n_2027;
assign n_2156 = x132 & n_2028;
assign n_2157 = ~x132 & n_2029;
assign n_2158 = ~x132 & n_2030;
assign n_2159 = x132 & n_2031;
assign n_2160 = x132 & n_2032;
assign n_2161 = ~x132 & n_2033;
assign n_2162 = ~x132 & n_2034;
assign n_2163 = x132 & n_2035;
assign n_2164 = x132 & n_2036;
assign n_2165 = ~x132 & n_2037;
assign n_2166 = ~x132 & n_2038;
assign n_2167 = x132 & n_2039;
assign n_2168 = x132 & n_2040;
assign n_2169 = ~x132 & n_2041;
assign n_2170 = ~x132 & n_2042;
assign n_2171 = x132 & n_2043;
assign n_2172 = x132 & n_2044;
assign n_2173 = ~x132 & n_2045;
assign n_2174 = ~x132 & n_2046;
assign n_2175 = x132 & n_2047;
assign n_2176 = n_2048 ^ n_1808;
assign n_2177 = n_2049 ^ n_1809;
assign n_2178 = n_2050 ^ n_1810;
assign n_2179 = n_2051 ^ n_1811;
assign n_2180 = n_2052 ^ n_1812;
assign n_2181 = n_2053 ^ n_1813;
assign n_2182 = n_2054 ^ n_1814;
assign n_2183 = n_2055 ^ n_1815;
assign n_2184 = n_2056 ^ n_1816;
assign n_2185 = n_2057 ^ n_1817;
assign n_2186 = n_2058 ^ n_1818;
assign n_2187 = n_2059 ^ n_1819;
assign n_2188 = n_2060 ^ n_1820;
assign n_2189 = n_2061 ^ n_1821;
assign n_2190 = n_2062 ^ n_1822;
assign n_2191 = n_2063 ^ n_1823;
assign n_2192 = n_2064 ^ n_1824;
assign n_2193 = n_2065 ^ n_1809;
assign n_2194 = n_2066 ^ n_1810;
assign n_2195 = n_2067 ^ n_1811;
assign n_2196 = n_2068 ^ n_1812;
assign n_2197 = n_2069 ^ n_1813;
assign n_2198 = n_2070 ^ n_1814;
assign n_2199 = n_2071 ^ n_1815;
assign n_2200 = n_2072 ^ n_1816;
assign n_2201 = n_2073 ^ n_1817;
assign n_2202 = n_2074 ^ n_1818;
assign n_2203 = n_2075 ^ n_1819;
assign n_2204 = n_2076 ^ n_1820;
assign n_2205 = n_2077 ^ n_1821;
assign n_2206 = n_2078 ^ n_1822;
assign n_2207 = n_2079 ^ n_1823;
assign n_2208 = n_2080 ^ n_1824;
assign n_2209 = n_2081 ^ n_1825;
assign n_2210 = n_2082 ^ n_1826;
assign n_2211 = n_2083 ^ n_1827;
assign n_2212 = n_2084 ^ n_1828;
assign n_2213 = n_2085 ^ n_1829;
assign n_2214 = n_2086 ^ n_1830;
assign n_2215 = n_2087 ^ n_1831;
assign n_2216 = n_2088 ^ n_1832;
assign n_2217 = n_2089 ^ n_1833;
assign n_2218 = n_2090 ^ n_1834;
assign n_2219 = n_2091 ^ n_1835;
assign n_2220 = n_2092 ^ n_1836;
assign n_2221 = n_2093 ^ n_1837;
assign n_2222 = n_2094 ^ n_1838;
assign n_2223 = n_2095 ^ n_1839;
assign n_2224 = n_2096 ^ n_1840;
assign n_2225 = n_2097 ^ n_1858;
assign n_2226 = n_2098 ^ n_1860;
assign n_2227 = n_2099 ^ n_1862;
assign n_2228 = n_2100 ^ n_1864;
assign n_2229 = n_2101 ^ n_1866;
assign n_2230 = n_2102 ^ n_1868;
assign n_2231 = n_2103 ^ n_1870;
assign n_2232 = n_2104 ^ n_1872;
assign n_2233 = n_2105 ^ n_1874;
assign n_2234 = n_2106 ^ n_1876;
assign n_2235 = n_2107 ^ n_1878;
assign n_2236 = n_2108 ^ n_1880;
assign n_2237 = n_2109 ^ n_1882;
assign n_2238 = n_2110 ^ n_1884;
assign n_2239 = n_2111 ^ n_1886;
assign n_2240 = n_2112 ^ n_1888;
assign n_2241 = n_2113 ^ n_1888;
assign n_2242 = n_2114 ^ n_1859;
assign n_2243 = n_2115 ^ n_1793;
assign n_2244 = n_2116 ^ n_1890;
assign n_2245 = n_2117 ^ n_1890;
assign n_2246 = n_2118 ^ n_1867;
assign n_2247 = n_2119 ^ n_1797;
assign n_2248 = n_2120 ^ n_1892;
assign n_2249 = n_2121 ^ n_1892;
assign n_2250 = n_2122 ^ n_1875;
assign n_2251 = n_2123 ^ n_1801;
assign n_2252 = n_2124 ^ n_1894;
assign n_2253 = n_2125 ^ n_1894;
assign n_2254 = n_2126 ^ n_1883;
assign n_2255 = n_2127 ^ n_1805;
assign n_2256 = n_2128 ^ n_1896;
assign n_2257 = n_2129 ^ n_1896;
assign n_2258 = n_2130 ^ n_1865;
assign n_2259 = n_2131 ^ n_1796;
assign n_2260 = n_2132 ^ n_1856;
assign n_2261 = n_2133 ^ n_1898;
assign n_2262 = n_2134 ^ n_1856;
assign n_2263 = n_2135 ^ n_1899;
assign n_2264 = n_2136 ^ n_1900;
assign n_2265 = n_2137 ^ n_1900;
assign n_2266 = n_2138 ^ n_1873;
assign n_2267 = n_2139 ^ n_1800;
assign n_2268 = n_2140 ^ n_1902;
assign n_2269 = n_2141 ^ n_1902;
assign n_2270 = n_2142 ^ n_1881;
assign n_2271 = n_2143 ^ n_1804;
assign n_2272 = n_2144 ^ n_1904;
assign n_2273 = n_2145 ^ n_1904;
assign n_2274 = n_2146 ^ n_1861;
assign n_2275 = n_2147 ^ n_1794;
assign n_2276 = n_2148 ^ n_1906;
assign n_2277 = n_2149 ^ n_1906;
assign n_2278 = n_2150 ^ n_1869;
assign n_2279 = n_2151 ^ n_1798;
assign n_2280 = n_2152 ^ n_1908;
assign n_2281 = n_2153 ^ n_1908;
assign n_2282 = n_2154 ^ n_1877;
assign n_2283 = n_2155 ^ n_1802;
assign n_2284 = n_2156 ^ n_1910;
assign n_2285 = n_2157 ^ n_1910;
assign n_2286 = n_2158 ^ n_1885;
assign n_2287 = n_2159 ^ n_1806;
assign n_2288 = n_2160 ^ n_1912;
assign n_2289 = n_2161 ^ n_1912;
assign n_2290 = n_2162 ^ n_1863;
assign n_2291 = n_2163 ^ n_1795;
assign n_2292 = n_2164 ^ n_1914;
assign n_2293 = n_2165 ^ n_1914;
assign n_2294 = n_2166 ^ n_1871;
assign n_2295 = n_2167 ^ n_1799;
assign n_2296 = n_2168 ^ n_1916;
assign n_2297 = n_2169 ^ n_1916;
assign n_2298 = n_2170 ^ n_1879;
assign n_2299 = n_2171 ^ n_1803;
assign n_2300 = n_2172 ^ n_1918;
assign n_2301 = n_2173 ^ n_1918;
assign n_2302 = n_2174 ^ n_1887;
assign n_2303 = n_2175 ^ n_1807;
assign n_2304 = n_2240 ^ n_2177;
assign n_2305 = n_2241 ^ n_2193;
assign n_2306 = n_2242 ^ n_2209;
assign n_2307 = n_2243 ^ n_2225;
assign n_2308 = n_2244 ^ n_2181;
assign n_2309 = n_2245 ^ n_2197;
assign n_2310 = n_2246 ^ n_2213;
assign n_2311 = n_2247 ^ n_2229;
assign n_2312 = n_2248 ^ n_2185;
assign n_2313 = n_2249 ^ n_2201;
assign n_2314 = n_2250 ^ n_2217;
assign n_2315 = n_2251 ^ n_2233;
assign n_2316 = n_2252 ^ n_2189;
assign n_2317 = n_2253 ^ n_2205;
assign n_2318 = n_2254 ^ n_2221;
assign n_2319 = n_2255 ^ n_2237;
assign n_2320 = n_2256 ^ n_2180;
assign n_2321 = n_2257 ^ n_2196;
assign n_2322 = n_2258 ^ n_2212;
assign n_2323 = n_2259 ^ n_2228;
assign n_2324 = n_2260 ^ n_2192;
assign n_2325 = n_2261 ^ n_2176;
assign n_2326 = n_2262 ^ n_2208;
assign n_2327 = n_2263 ^ n_2224;
assign n_2328 = n_2264 ^ n_2184;
assign n_2329 = n_2265 ^ n_2200;
assign n_2330 = n_2266 ^ n_2216;
assign n_2331 = n_2267 ^ n_2232;
assign n_2332 = n_2268 ^ n_2188;
assign n_2333 = n_2269 ^ n_2204;
assign n_2334 = n_2270 ^ n_2220;
assign n_2335 = n_2271 ^ n_2236;
assign n_2336 = n_2272 ^ n_2178;
assign n_2337 = n_2273 ^ n_2194;
assign n_2338 = n_2274 ^ n_2210;
assign n_2339 = n_2275 ^ n_2226;
assign n_2340 = n_2276 ^ n_2182;
assign n_2341 = n_2277 ^ n_2198;
assign n_2342 = n_2278 ^ n_2214;
assign n_2343 = n_2279 ^ n_2230;
assign n_2344 = n_2280 ^ n_2186;
assign n_2345 = n_2281 ^ n_2202;
assign n_2346 = n_2282 ^ n_2218;
assign n_2347 = n_2283 ^ n_2234;
assign n_2348 = n_2284 ^ n_2190;
assign n_2349 = n_2285 ^ n_2206;
assign n_2350 = n_2286 ^ n_2222;
assign n_2351 = n_2287 ^ n_2238;
assign n_2352 = n_2288 ^ n_2179;
assign n_2353 = n_2289 ^ n_2195;
assign n_2354 = n_2290 ^ n_2211;
assign n_2355 = n_2291 ^ n_2227;
assign n_2356 = n_2292 ^ n_2183;
assign n_2357 = n_2293 ^ n_2199;
assign n_2358 = n_2294 ^ n_2215;
assign n_2359 = n_2295 ^ n_2231;
assign n_2360 = n_2296 ^ n_2187;
assign n_2361 = n_2297 ^ n_2203;
assign n_2362 = n_2298 ^ n_2219;
assign n_2363 = n_2299 ^ n_2235;
assign n_2364 = n_2300 ^ n_2191;
assign n_2365 = n_2301 ^ n_2207;
assign n_2366 = n_2302 ^ n_2223;
assign n_2367 = n_2303 ^ n_2239;
assign n_2368 = x134 & n_2304;
assign n_2369 = x134 & n_2305;
assign n_2370 = x134 & n_2306;
assign n_2371 = x134 & n_2307;
assign n_2372 = x134 & n_2308;
assign n_2373 = x134 & n_2309;
assign n_2374 = x134 & n_2310;
assign n_2375 = x134 & n_2311;
assign n_2376 = x134 & n_2312;
assign n_2377 = x134 & n_2313;
assign n_2378 = x134 & n_2314;
assign n_2379 = x134 & n_2315;
assign n_2380 = x134 & n_2316;
assign n_2381 = x134 & n_2317;
assign n_2382 = x134 & n_2318;
assign n_2383 = x134 & n_2319;
assign n_2384 = x134 & n_2320;
assign n_2385 = x134 & n_2321;
assign n_2386 = x134 & n_2322;
assign n_2387 = x134 & n_2323;
assign n_2388 = x134 & n_2324;
assign n_2389 = x134 & n_2325;
assign n_2390 = x134 & n_2326;
assign n_2391 = x134 & n_2327;
assign n_2392 = x134 & n_2328;
assign n_2393 = x134 & n_2329;
assign n_2394 = x134 & n_2330;
assign n_2395 = x134 & n_2331;
assign n_2396 = x134 & n_2332;
assign n_2397 = x134 & n_2333;
assign n_2398 = x134 & n_2334;
assign n_2399 = x134 & n_2335;
assign n_2400 = x134 & n_2336;
assign n_2401 = x134 & n_2337;
assign n_2402 = x134 & n_2338;
assign n_2403 = x134 & n_2339;
assign n_2404 = x134 & n_2340;
assign n_2405 = x134 & n_2341;
assign n_2406 = x134 & n_2342;
assign n_2407 = x134 & n_2343;
assign n_2408 = x134 & n_2344;
assign n_2409 = x134 & n_2345;
assign n_2410 = x134 & n_2346;
assign n_2411 = x134 & n_2347;
assign n_2412 = x134 & n_2348;
assign n_2413 = x134 & n_2349;
assign n_2414 = x134 & n_2350;
assign n_2415 = x134 & n_2351;
assign n_2416 = x134 & n_2352;
assign n_2417 = x134 & n_2353;
assign n_2418 = x134 & n_2354;
assign n_2419 = x134 & n_2355;
assign n_2420 = x134 & n_2356;
assign n_2421 = x134 & n_2357;
assign n_2422 = x134 & n_2358;
assign n_2423 = x134 & n_2359;
assign n_2424 = x134 & n_2360;
assign n_2425 = x134 & n_2361;
assign n_2426 = x134 & n_2362;
assign n_2427 = x134 & n_2363;
assign n_2428 = x134 & n_2364;
assign n_2429 = x134 & n_2365;
assign n_2430 = x134 & n_2366;
assign n_2431 = x134 & n_2367;
assign n_2432 = n_2368 ^ n_2240;
assign n_2433 = n_2368 ^ n_2177;
assign n_2434 = n_2369 ^ n_2241;
assign n_2435 = n_2369 ^ n_2193;
assign n_2436 = n_2370 ^ n_2242;
assign n_2437 = n_2370 ^ n_2209;
assign n_2438 = n_2371 ^ n_2243;
assign n_2439 = n_2371 ^ n_2225;
assign n_2440 = n_2372 ^ n_2244;
assign n_2441 = n_2372 ^ n_2181;
assign n_2442 = n_2373 ^ n_2245;
assign n_2443 = n_2373 ^ n_2197;
assign n_2444 = n_2374 ^ n_2246;
assign n_2445 = n_2374 ^ n_2213;
assign n_2446 = n_2375 ^ n_2247;
assign n_2447 = n_2375 ^ n_2229;
assign n_2448 = n_2376 ^ n_2248;
assign n_2449 = n_2376 ^ n_2185;
assign n_2450 = n_2377 ^ n_2249;
assign n_2451 = n_2377 ^ n_2201;
assign n_2452 = n_2378 ^ n_2250;
assign n_2453 = n_2378 ^ n_2217;
assign n_2454 = n_2379 ^ n_2251;
assign n_2455 = n_2379 ^ n_2233;
assign n_2456 = n_2380 ^ n_2252;
assign n_2457 = n_2380 ^ n_2189;
assign n_2458 = n_2381 ^ n_2253;
assign n_2459 = n_2381 ^ n_2205;
assign n_2460 = n_2382 ^ n_2254;
assign n_2461 = n_2382 ^ n_2221;
assign n_2462 = n_2383 ^ n_2255;
assign n_2463 = n_2383 ^ n_2237;
assign n_2464 = n_2384 ^ n_2256;
assign n_2465 = n_2384 ^ n_2180;
assign n_2466 = n_2385 ^ n_2257;
assign n_2467 = n_2385 ^ n_2196;
assign n_2468 = n_2386 ^ n_2258;
assign n_2469 = n_2386 ^ n_2212;
assign n_2470 = n_2387 ^ n_2259;
assign n_2471 = n_2387 ^ n_2228;
assign n_2472 = n_2388 ^ n_2260;
assign n_2473 = n_2388 ^ n_2192;
assign n_2474 = n_2389 ^ n_2176;
assign n_2475 = n_2389 ^ n_2261;
assign n_2476 = n_2390 ^ n_2262;
assign n_2477 = n_2390 ^ n_2208;
assign n_2478 = n_2391 ^ n_2263;
assign n_2479 = n_2391 ^ n_2224;
assign n_2480 = n_2392 ^ n_2264;
assign n_2481 = n_2392 ^ n_2184;
assign n_2482 = n_2393 ^ n_2265;
assign n_2483 = n_2393 ^ n_2200;
assign n_2484 = n_2394 ^ n_2266;
assign n_2485 = n_2394 ^ n_2216;
assign n_2486 = n_2395 ^ n_2267;
assign n_2487 = n_2395 ^ n_2232;
assign n_2488 = n_2396 ^ n_2268;
assign n_2489 = n_2396 ^ n_2188;
assign n_2490 = n_2397 ^ n_2269;
assign n_2491 = n_2397 ^ n_2204;
assign n_2492 = n_2398 ^ n_2270;
assign n_2493 = n_2398 ^ n_2220;
assign n_2494 = n_2399 ^ n_2271;
assign n_2495 = n_2399 ^ n_2236;
assign n_2496 = n_2400 ^ n_2272;
assign n_2497 = n_2400 ^ n_2178;
assign n_2498 = n_2401 ^ n_2273;
assign n_2499 = n_2401 ^ n_2194;
assign n_2500 = n_2402 ^ n_2274;
assign n_2501 = n_2402 ^ n_2210;
assign n_2502 = n_2403 ^ n_2275;
assign n_2503 = n_2403 ^ n_2226;
assign n_2504 = n_2404 ^ n_2276;
assign n_2505 = n_2404 ^ n_2182;
assign n_2506 = n_2405 ^ n_2277;
assign n_2507 = n_2405 ^ n_2198;
assign n_2508 = n_2406 ^ n_2278;
assign n_2509 = n_2406 ^ n_2214;
assign n_2510 = n_2407 ^ n_2279;
assign n_2511 = n_2407 ^ n_2230;
assign n_2512 = n_2408 ^ n_2280;
assign n_2513 = n_2408 ^ n_2186;
assign n_2514 = n_2409 ^ n_2281;
assign n_2515 = n_2409 ^ n_2202;
assign n_2516 = n_2410 ^ n_2282;
assign n_2517 = n_2410 ^ n_2218;
assign n_2518 = n_2411 ^ n_2283;
assign n_2519 = n_2411 ^ n_2234;
assign n_2520 = n_2412 ^ n_2284;
assign n_2521 = n_2412 ^ n_2190;
assign n_2522 = n_2413 ^ n_2285;
assign n_2523 = n_2413 ^ n_2206;
assign n_2524 = n_2414 ^ n_2286;
assign n_2525 = n_2414 ^ n_2222;
assign n_2526 = n_2415 ^ n_2287;
assign n_2527 = n_2415 ^ n_2238;
assign n_2528 = n_2416 ^ n_2288;
assign n_2529 = n_2416 ^ n_2179;
assign n_2530 = n_2417 ^ n_2289;
assign n_2531 = n_2417 ^ n_2195;
assign n_2532 = n_2418 ^ n_2290;
assign n_2533 = n_2418 ^ n_2211;
assign n_2534 = n_2419 ^ n_2291;
assign n_2535 = n_2419 ^ n_2227;
assign n_2536 = n_2420 ^ n_2292;
assign n_2537 = n_2420 ^ n_2183;
assign n_2538 = n_2421 ^ n_2293;
assign n_2539 = n_2421 ^ n_2199;
assign n_2540 = n_2422 ^ n_2294;
assign n_2541 = n_2422 ^ n_2215;
assign n_2542 = n_2423 ^ n_2295;
assign n_2543 = n_2423 ^ n_2231;
assign n_2544 = n_2424 ^ n_2296;
assign n_2545 = n_2424 ^ n_2187;
assign n_2546 = n_2425 ^ n_2297;
assign n_2547 = n_2425 ^ n_2203;
assign n_2548 = n_2426 ^ n_2298;
assign n_2549 = n_2426 ^ n_2219;
assign n_2550 = n_2427 ^ n_2299;
assign n_2551 = n_2427 ^ n_2235;
assign n_2552 = n_2428 ^ n_2300;
assign n_2553 = n_2428 ^ n_2191;
assign n_2554 = n_2429 ^ n_2301;
assign n_2555 = n_2429 ^ n_2207;
assign n_2556 = n_2430 ^ n_2302;
assign n_2557 = n_2430 ^ n_2223;
assign n_2558 = n_2431 ^ n_2303;
assign n_2559 = n_2431 ^ n_2239;
assign y0 = n_2432;
assign y64 = n_2433;
assign y16 = n_2434;
assign y80 = n_2435;
assign y32 = n_2436;
assign y96 = n_2437;
assign y48 = n_2438;
assign y112 = n_2439;
assign y4 = n_2440;
assign y68 = n_2441;
assign y20 = n_2442;
assign y84 = n_2443;
assign y36 = n_2444;
assign y100 = n_2445;
assign y52 = n_2446;
assign y116 = n_2447;
assign y8 = n_2448;
assign y72 = n_2449;
assign y24 = n_2450;
assign y88 = n_2451;
assign y40 = n_2452;
assign y104 = n_2453;
assign y56 = n_2454;
assign y120 = n_2455;
assign y12 = n_2456;
assign y76 = n_2457;
assign y28 = n_2458;
assign y92 = n_2459;
assign y44 = n_2460;
assign y108 = n_2461;
assign y60 = n_2462;
assign y124 = n_2463;
assign y3 = n_2464;
assign y67 = n_2465;
assign y19 = n_2466;
assign y83 = n_2467;
assign y35 = n_2468;
assign y99 = n_2469;
assign y51 = n_2470;
assign y115 = n_2471;
assign y15 = n_2472;
assign y79 = n_2473;
assign y63 = n_2474;
assign y127 = n_2475;
assign y31 = n_2476;
assign y95 = n_2477;
assign y47 = n_2478;
assign y111 = n_2479;
assign y7 = n_2480;
assign y71 = n_2481;
assign y23 = n_2482;
assign y87 = n_2483;
assign y39 = n_2484;
assign y103 = n_2485;
assign y55 = n_2486;
assign y119 = n_2487;
assign y11 = n_2488;
assign y75 = n_2489;
assign y27 = n_2490;
assign y91 = n_2491;
assign y43 = n_2492;
assign y107 = n_2493;
assign y59 = n_2494;
assign y123 = n_2495;
assign y1 = n_2496;
assign y65 = n_2497;
assign y17 = n_2498;
assign y81 = n_2499;
assign y33 = n_2500;
assign y97 = n_2501;
assign y49 = n_2502;
assign y113 = n_2503;
assign y5 = n_2504;
assign y69 = n_2505;
assign y21 = n_2506;
assign y85 = n_2507;
assign y37 = n_2508;
assign y101 = n_2509;
assign y53 = n_2510;
assign y117 = n_2511;
assign y9 = n_2512;
assign y73 = n_2513;
assign y25 = n_2514;
assign y89 = n_2515;
assign y41 = n_2516;
assign y105 = n_2517;
assign y57 = n_2518;
assign y121 = n_2519;
assign y13 = n_2520;
assign y77 = n_2521;
assign y29 = n_2522;
assign y93 = n_2523;
assign y45 = n_2524;
assign y109 = n_2525;
assign y61 = n_2526;
assign y125 = n_2527;
assign y2 = n_2528;
assign y66 = n_2529;
assign y18 = n_2530;
assign y82 = n_2531;
assign y34 = n_2532;
assign y98 = n_2533;
assign y50 = n_2534;
assign y114 = n_2535;
assign y6 = n_2536;
assign y70 = n_2537;
assign y22 = n_2538;
assign y86 = n_2539;
assign y38 = n_2540;
assign y102 = n_2541;
assign y54 = n_2542;
assign y118 = n_2543;
assign y10 = n_2544;
assign y74 = n_2545;
assign y26 = n_2546;
assign y90 = n_2547;
assign y42 = n_2548;
assign y106 = n_2549;
assign y58 = n_2550;
assign y122 = n_2551;
assign y14 = n_2552;
assign y78 = n_2553;
assign y30 = n_2554;
assign y94 = n_2555;
assign y46 = n_2556;
assign y110 = n_2557;
assign y62 = n_2558;
assign y126 = n_2559;
endmodule