module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n245 , n246 , n247 , n249 , n250 , n251 , n252 , n253 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n293 , n294 , n295 , n296 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n464 , n465 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n523 , n524 , n525 , n526 , n527 , n528 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n611 , n614 , n615 , n616 , n617 , n618 , n619 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n636 , n637 , n638 , n639 , n640 , n645 , n646 , n647 , n648 , n650 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n671 , n674 , n675 , n676 , n677 , n678 , n679 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n706 , n707 , n708 , n709 , n710 , n711 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n743 , n744 , n745 , n746 , n747 , n748 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n795 , n796 , n797 , n798 , n799 , n800 , n803 , n804 , n805 , n806 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n832 , n833 , n834 , n835 , n838 , n839 , n840 , n841 , n844 , n845 , n846 , n847 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n859 , n860 , n861 , n862 , n865 , n866 , n867 , n868 , n871 , n872 , n873 , n874 , n877 , n878 , n879 , n880 , n883 , n884 , n885 , n886 , n889 , n890 , n891 , n892 , n895 , n896 , n897 , n898 , n901 , n902 , n903 , n904 , n907 , n908 , n909 , n910 , n913 , n914 , n915 , n916 , n919 , n920 , n921 , n922 , n925 , n926 , n927 , n928 , n929 , n932 , n933 , n934 , n935 , n938 , n939 , n940 , n941 , n944 , n945 , n946 , n947 , n950 , n951 , n952 , n953 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n985 , n986 , n987 , n990 , n991 , n992 , n993 , n994 , n995 , n998 , n999 , n1000 , n1001 , n1004 , n1005 , n1006 , n1007 , n1008 , n1011 , n1012 , n1013 , n1014 , n1017 , n1018 , n1019 , n1020 , n1023 , n1024 , n1025 , n1026 , n1029 , n1030 , n1031 , n1032 , n1035 , n1036 , n1037 , n1038 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1050 , n1051 , n1052 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1064 , n1065 , n1066 , n1067 , n1068 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1079 , n1080 , n1081 , n1082 , n1085 , n1086 , n1087 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1117 , n1118 , n1119 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1153 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1196 , n1197 , n1198 , n1199 , n1200 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1249 , n1250 , n1251 , n1252 , n1253 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1281 , n1282 , n1283 , n1284 , n1287 , n1288 , n1289 , n1290 , n1293 , n1294 , n1295 , n1296 , n1299 , n1300 , n1301 , n1302 , n1303 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 ;
  assign n148 = ~x17 & x54 ;
  assign n150 = ~x8 & ~x10 ;
  assign n151 = ~x14 & ~x21 ;
  assign n152 = n150 & n151 ;
  assign n153 = ~x13 & n152 ;
  assign n154 = ~x4 & ~x9 ;
  assign n155 = ~x12 & n154 ;
  assign n156 = ~x7 & n155 ;
  assign n157 = n153 & n156 ;
  assign n158 = x7 ^ x6 ;
  assign n159 = n158 ^ x9 ;
  assign n160 = n159 ^ x12 ;
  assign n161 = n160 ^ x13 ;
  assign n162 = x13 ^ x12 ;
  assign n163 = x9 ^ x7 ;
  assign n164 = n163 ^ x12 ;
  assign n165 = n162 & n164 ;
  assign n166 = n165 ^ x12 ;
  assign n167 = n161 & n166 ;
  assign n168 = n167 ^ n161 ;
  assign n169 = x7 & x9 ;
  assign n170 = n168 & n169 ;
  assign n171 = n170 ^ n168 ;
  assign n172 = n157 & ~n171 ;
  assign n173 = ~x5 & ~x22 ;
  assign n174 = ~x11 & n173 ;
  assign n175 = ~x18 & ~x19 ;
  assign n176 = x16 & n175 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n174 & n177 ;
  assign n179 = n172 & n178 ;
  assign n180 = n148 & ~n179 ;
  assign n149 = n148 ^ x54 ;
  assign n181 = n180 ^ n149 ;
  assign n182 = ~x0 & ~n181 ;
  assign n183 = ~x6 & n177 ;
  assign n184 = n155 & n183 ;
  assign n190 = x10 ^ x8 ;
  assign n185 = x21 ^ x14 ;
  assign n186 = x14 ^ x13 ;
  assign n187 = n185 & n186 ;
  assign n188 = n187 ^ x14 ;
  assign n189 = n150 & ~n188 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = ~x13 & n151 ;
  assign n193 = n191 & n192 ;
  assign n194 = n193 ^ n153 ;
  assign n195 = n194 ^ n189 ;
  assign n196 = x7 & n195 ;
  assign n197 = n196 ^ n193 ;
  assign n198 = n197 ^ n189 ;
  assign n202 = n184 & n198 ;
  assign n203 = n148 & n174 ;
  assign n204 = n202 & n203 ;
  assign n205 = ~x9 & ~x11 ;
  assign n206 = n205 ^ n173 ;
  assign n207 = x54 & ~x56 ;
  assign n208 = n206 & n207 ;
  assign n209 = ~n204 & ~n208 ;
  assign n210 = ~n182 & n209 ;
  assign n211 = ~x3 & ~x129 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = ~x1 & ~n180 ;
  assign n214 = ~x5 & ~n171 ;
  assign n215 = x54 & n211 ;
  assign n216 = x17 & n215 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = n177 & n217 ;
  assign n219 = ~x11 & ~x22 ;
  assign n220 = ~x4 & n219 ;
  assign n221 = n152 & n220 ;
  assign n222 = n218 & n221 ;
  assign n223 = ~n214 & n222 ;
  assign n225 = ~x5 & n223 ;
  assign n224 = n172 & n223 ;
  assign n226 = n225 ^ n224 ;
  assign n227 = n211 & ~n226 ;
  assign n228 = n213 & n227 ;
  assign n229 = n228 ^ n226 ;
  assign n231 = ~x41 & ~x46 ;
  assign n232 = ~x47 & ~x48 ;
  assign n233 = n231 & n232 ;
  assign n234 = ~x43 & n233 ;
  assign n242 = ~x38 & ~x50 ;
  assign n245 = ~x42 & ~x44 ;
  assign n246 = ~x40 & n245 ;
  assign n256 = n242 & n246 ;
  assign n257 = n234 & n256 ;
  assign n408 = x82 & n257 ;
  assign n409 = ~x45 & n408 ;
  assign n686 = n409 ^ x82 ;
  assign n235 = ~x24 & ~x49 ;
  assign n236 = ~x45 & n235 ;
  assign n237 = ~x15 & ~x20 ;
  assign n238 = ~x2 & n237 ;
  assign n239 = n236 & n238 ;
  assign n687 = x82 & ~n239 ;
  assign n688 = ~n686 & ~n687 ;
  assign n230 = x122 & x127 ;
  assign n249 = n230 & n688 ;
  assign n250 = n688 ^ n249 ;
  assign n251 = x2 & ~x129 ;
  assign n258 = n236 & n257 ;
  assign n259 = n237 & n258 ;
  assign n260 = x82 & n259 ;
  assign n252 = ~x82 & ~n230 ;
  assign n261 = n260 ^ n252 ;
  assign n262 = n251 & ~n261 ;
  assign n263 = n262 ^ x129 ;
  assign n264 = ~x65 & ~n263 ;
  assign n265 = n250 & n264 ;
  assign n267 = n265 ^ n262 ;
  assign n268 = ~x17 & n179 ;
  assign n269 = ~x61 & ~x118 ;
  assign n270 = ~x129 & n269 ;
  assign n271 = ~n268 & n270 ;
  assign n272 = x0 & ~x113 ;
  assign n273 = x123 & ~x129 ;
  assign n274 = n273 ^ x129 ;
  assign n275 = n272 & ~n274 ;
  assign n276 = ~n271 & ~n275 ;
  assign n280 = n215 ^ n211 ;
  assign n281 = x4 & n280 ;
  assign n277 = n174 & n217 ;
  assign n278 = n202 & n277 ;
  assign n279 = x10 & n278 ;
  assign n282 = n281 ^ n279 ;
  assign n291 = x5 & n280 ;
  assign n283 = ~x25 & ~x28 ;
  assign n284 = n283 ^ x25 ;
  assign n285 = ~x29 & ~x59 ;
  assign n286 = n172 & n277 ;
  assign n287 = ~x16 & n286 ;
  assign n288 = n175 & n287 ;
  assign n289 = n285 & n288 ;
  assign n290 = ~n284 & n289 ;
  assign n293 = n291 ^ n290 ;
  assign n296 = x6 & n280 ;
  assign n294 = n283 ^ x28 ;
  assign n295 = n289 & ~n294 ;
  assign n298 = n296 ^ n295 ;
  assign n300 = x7 & n280 ;
  assign n299 = x8 & n278 ;
  assign n301 = n300 ^ n299 ;
  assign n303 = x8 & n280 ;
  assign n302 = x21 & n278 ;
  assign n304 = n303 ^ n302 ;
  assign n309 = x9 & n280 ;
  assign n305 = ~x5 & n218 ;
  assign n306 = n172 & n305 ;
  assign n307 = x11 & ~x22 ;
  assign n308 = n306 & n307 ;
  assign n310 = n309 ^ n308 ;
  assign n312 = x10 & n280 ;
  assign n311 = x14 & n278 ;
  assign n313 = n312 ^ n311 ;
  assign n318 = x22 & n306 ;
  assign n319 = n318 ^ n280 ;
  assign n320 = ~x11 & n319 ;
  assign n321 = n320 ^ n280 ;
  assign n323 = ~x18 & n287 ;
  assign n324 = n323 ^ n287 ;
  assign n325 = ~x19 & n324 ;
  assign n322 = x12 & n280 ;
  assign n326 = n325 ^ n322 ;
  assign n333 = x13 & n280 ;
  assign n327 = x29 & x54 ;
  assign n328 = ~x59 & n327 ;
  assign n329 = n283 & n328 ;
  assign n330 = n268 & n329 ;
  assign n332 = n211 & n330 ;
  assign n334 = n333 ^ n332 ;
  assign n336 = x14 & n280 ;
  assign n335 = x13 & n278 ;
  assign n337 = n336 ^ n335 ;
  assign n338 = n258 ^ x15 ;
  assign n339 = n338 ^ x70 ;
  assign n340 = n339 ^ n258 ;
  assign n343 = ~n230 & ~n340 ;
  assign n344 = n343 ^ n258 ;
  assign n345 = ~x82 & n344 ;
  assign n346 = n345 ^ n338 ;
  assign n347 = ~x129 & n238 ;
  assign n355 = ~x70 & n347 ;
  assign n356 = ~n230 & n355 ;
  assign n357 = n356 ^ n230 ;
  assign n348 = n347 ^ x129 ;
  assign n349 = n348 ^ n230 ;
  assign n358 = n357 ^ n349 ;
  assign n359 = n346 & ~n358 ;
  assign n361 = x16 & n280 ;
  assign n360 = x6 & n226 ;
  assign n362 = n361 ^ n360 ;
  assign n364 = ~x29 & n283 ;
  assign n365 = n179 & n364 ;
  assign n366 = x59 & n217 ;
  assign n367 = n365 & n366 ;
  assign n363 = x17 & n280 ;
  assign n368 = n367 ^ n363 ;
  assign n370 = n176 & n286 ;
  assign n369 = x18 & n280 ;
  assign n371 = n370 ^ n369 ;
  assign n373 = x19 & n280 ;
  assign n372 = n179 & n216 ;
  assign n374 = n373 ^ n372 ;
  assign n379 = ~x15 & n258 ;
  assign n380 = n379 ^ x20 ;
  assign n381 = x82 & ~n380 ;
  assign n382 = x71 ^ x20 ;
  assign n383 = ~n230 & ~n382 ;
  assign n384 = n383 ^ x20 ;
  assign n385 = x82 & ~n384 ;
  assign n393 = ~n383 & n385 ;
  assign n394 = ~x2 & n393 ;
  assign n395 = n394 ^ x2 ;
  assign n386 = n385 ^ n384 ;
  assign n387 = n386 ^ x2 ;
  assign n396 = n395 ^ n387 ;
  assign n397 = ~x129 & n396 ;
  assign n398 = ~n381 & n397 ;
  assign n400 = x19 & n323 ;
  assign n399 = x21 & n280 ;
  assign n401 = n400 ^ n399 ;
  assign n402 = x22 & n280 ;
  assign n403 = n402 ^ n224 ;
  assign n404 = ~x23 & x55 ;
  assign n405 = x61 & ~x129 ;
  assign n406 = ~n404 & n405 ;
  assign n407 = x63 & n250 ;
  assign n410 = n409 ^ n249 ;
  assign n411 = n410 ^ x82 ;
  assign n412 = n411 ^ n409 ;
  assign n415 = ~x24 & n412 ;
  assign n416 = n415 ^ n409 ;
  assign n417 = ~x129 & ~n416 ;
  assign n418 = ~n407 & n417 ;
  assign n419 = ~x26 & x27 ;
  assign n420 = n419 ^ x26 ;
  assign n448 = x58 ^ x53 ;
  assign n427 = ~x53 & ~x58 ;
  assign n449 = n448 ^ n427 ;
  assign n450 = ~x85 & n449 ;
  assign n451 = n450 ^ n427 ;
  assign n452 = ~n420 & n451 ;
  assign n442 = ~x85 & n427 ;
  assign n446 = ~n420 & n442 ;
  assign n443 = n420 ^ x27 ;
  assign n444 = n443 ^ x26 ;
  assign n445 = n442 & ~n444 ;
  assign n447 = n446 ^ n445 ;
  assign n453 = n452 ^ n447 ;
  assign n454 = ~x116 & n453 ;
  assign n431 = x27 & x116 ;
  assign n432 = ~x39 & ~x52 ;
  assign n433 = ~x51 & n432 ;
  assign n434 = n211 & ~n433 ;
  assign n435 = n431 & n434 ;
  assign n436 = n435 ^ n211 ;
  assign n455 = n454 ^ n436 ;
  assign n421 = x116 & n420 ;
  assign n422 = ~x96 & ~x110 ;
  assign n423 = n422 ^ x116 ;
  assign n424 = ~x85 & n423 ;
  assign n425 = n424 ^ x116 ;
  assign n426 = x100 & n425 ;
  assign n428 = n211 & ~n420 ;
  assign n429 = n427 & n428 ;
  assign n430 = n426 & n429 ;
  assign n437 = ~n430 & n436 ;
  assign n438 = ~n421 & n437 ;
  assign n439 = ~x25 & n438 ;
  assign n440 = n439 ^ n437 ;
  assign n464 = x26 & x116 ;
  assign n465 = n433 & n464 ;
  assign n468 = n445 & ~n465 ;
  assign n456 = ~x95 & ~x100 ;
  assign n457 = ~x97 & ~x110 ;
  assign n458 = n456 & n457 ;
  assign n459 = n458 ^ x110 ;
  assign n460 = n446 & n459 ;
  assign n461 = n460 ^ n446 ;
  assign n469 = n468 ^ n461 ;
  assign n470 = n440 & ~n469 ;
  assign n471 = n455 & n470 ;
  assign n441 = n440 ^ n430 ;
  assign n472 = n471 ^ n441 ;
  assign n473 = n211 & n443 ;
  assign n474 = x116 & n433 ;
  assign n475 = n442 & n474 ;
  assign n476 = n475 ^ n442 ;
  assign n477 = n473 & n476 ;
  assign n478 = n477 ^ n430 ;
  assign n479 = n419 & n476 ;
  assign n480 = x85 & x116 ;
  assign n481 = ~x95 & ~n480 ;
  assign n482 = ~n420 & n427 ;
  assign n483 = ~n481 & n482 ;
  assign n484 = ~x100 & n483 ;
  assign n485 = n425 & n484 ;
  assign n486 = ~n479 & ~n485 ;
  assign n487 = n211 & ~n486 ;
  assign n488 = ~x27 & n442 ;
  assign n489 = n487 ^ x28 ;
  assign n490 = ~n454 & n489 ;
  assign n491 = n490 ^ x28 ;
  assign n498 = ~x26 & x28 ;
  assign n499 = n459 & n498 ;
  assign n500 = n499 ^ n459 ;
  assign n492 = n465 ^ n459 ;
  assign n501 = n500 ^ n492 ;
  assign n502 = ~n491 & n501 ;
  assign n503 = n488 & n502 ;
  assign n504 = n503 ^ n491 ;
  assign n505 = n211 & n504 ;
  assign n506 = n428 & n450 ;
  assign n510 = n422 & n456 ;
  assign n511 = n510 ^ x116 ;
  assign n512 = ~x58 & n511 ;
  assign n513 = n512 ^ x116 ;
  assign n514 = x97 & n513 ;
  assign n515 = n514 ^ x116 ;
  assign n516 = ~x53 & ~n515 ;
  assign n517 = n516 ^ x116 ;
  assign n518 = n506 & ~n517 ;
  assign n519 = n518 ^ x29 ;
  assign n520 = n460 ^ n454 ;
  assign n523 = n519 & ~n520 ;
  assign n524 = n523 ^ x29 ;
  assign n525 = n211 & n524 ;
  assign n527 = x88 ^ x60 ;
  assign n526 = x88 ^ x30 ;
  assign n528 = n527 ^ n526 ;
  assign n531 = ~x109 & n528 ;
  assign n532 = n531 ^ n527 ;
  assign n533 = ~x106 & n532 ;
  assign n534 = n533 ^ x88 ;
  assign n535 = ~x129 & n534 ;
  assign n537 = x89 ^ x31 ;
  assign n536 = x89 ^ x30 ;
  assign n538 = n537 ^ n536 ;
  assign n541 = x109 & n538 ;
  assign n542 = n541 ^ n537 ;
  assign n543 = ~x106 & n542 ;
  assign n544 = n543 ^ x89 ;
  assign n545 = ~x129 & n544 ;
  assign n547 = x99 ^ x32 ;
  assign n546 = x99 ^ x31 ;
  assign n548 = n547 ^ n546 ;
  assign n551 = x109 & n548 ;
  assign n552 = n551 ^ n547 ;
  assign n553 = ~x106 & n552 ;
  assign n554 = n553 ^ x99 ;
  assign n555 = ~x129 & n554 ;
  assign n557 = x90 ^ x33 ;
  assign n556 = x90 ^ x32 ;
  assign n558 = n557 ^ n556 ;
  assign n561 = x109 & n558 ;
  assign n562 = n561 ^ n557 ;
  assign n563 = ~x106 & n562 ;
  assign n564 = n563 ^ x90 ;
  assign n565 = ~x129 & n564 ;
  assign n567 = x91 ^ x34 ;
  assign n566 = x91 ^ x33 ;
  assign n568 = n567 ^ n566 ;
  assign n571 = x109 & n568 ;
  assign n572 = n571 ^ n567 ;
  assign n573 = ~x106 & n572 ;
  assign n574 = n573 ^ x91 ;
  assign n575 = ~x129 & n574 ;
  assign n577 = x92 ^ x35 ;
  assign n576 = x92 ^ x34 ;
  assign n578 = n577 ^ n576 ;
  assign n581 = x109 & n578 ;
  assign n582 = n581 ^ n577 ;
  assign n583 = ~x106 & n582 ;
  assign n584 = n583 ^ x92 ;
  assign n585 = ~x129 & n584 ;
  assign n587 = x98 ^ x36 ;
  assign n586 = x98 ^ x35 ;
  assign n588 = n587 ^ n586 ;
  assign n591 = x109 & n588 ;
  assign n592 = n591 ^ n587 ;
  assign n593 = ~x106 & n592 ;
  assign n594 = n593 ^ x98 ;
  assign n595 = ~x129 & n594 ;
  assign n597 = x93 ^ x37 ;
  assign n596 = x93 ^ x36 ;
  assign n598 = n597 ^ n596 ;
  assign n601 = x109 & n598 ;
  assign n602 = n601 ^ n597 ;
  assign n603 = ~x106 & n602 ;
  assign n604 = n603 ^ x93 ;
  assign n605 = ~x129 & n604 ;
  assign n611 = x74 ^ x38 ;
  assign n614 = ~n230 & ~n611 ;
  assign n615 = n614 ^ x38 ;
  assign n607 = x82 & ~x129 ;
  assign n699 = n256 ^ x46 ;
  assign n700 = n607 & ~n699 ;
  assign n701 = n700 ^ x129 ;
  assign n702 = n688 & ~n701 ;
  assign n616 = ~n615 & n702 ;
  assign n606 = n246 ^ x38 ;
  assign n608 = ~n606 & n607 ;
  assign n609 = n608 ^ x129 ;
  assign n617 = n616 ^ n609 ;
  assign n618 = ~x106 & ~x129 ;
  assign n619 = ~x51 & x109 ;
  assign n624 = ~x52 & n619 ;
  assign n625 = n624 ^ x39 ;
  assign n626 = n618 & ~n625 ;
  assign n627 = n626 ^ x129 ;
  assign n247 = x82 & ~n246 ;
  assign n630 = n688 ^ n247 ;
  assign n628 = ~x73 & ~n230 ;
  assign n629 = n628 & n688 ;
  assign n631 = n630 ^ n629 ;
  assign n632 = x40 & n631 ;
  assign n636 = x82 & n245 ;
  assign n637 = n636 ^ n252 ;
  assign n638 = n632 & ~n637 ;
  assign n639 = n638 ^ n631 ;
  assign n640 = ~x129 & ~n639 ;
  assign n650 = x76 ^ x41 ;
  assign n653 = ~n230 & ~n650 ;
  assign n654 = n653 ^ x41 ;
  assign n655 = ~n654 & n702 ;
  assign n645 = ~x46 & n256 ;
  assign n646 = n645 ^ x41 ;
  assign n647 = n607 & ~n646 ;
  assign n648 = n647 ^ x129 ;
  assign n656 = n655 ^ n648 ;
  assign n663 = x42 & ~n252 ;
  assign n657 = x72 & n688 ;
  assign n661 = ~n249 & n657 ;
  assign n658 = x44 & x82 ;
  assign n659 = n658 ^ n249 ;
  assign n662 = n661 ^ n659 ;
  assign n664 = n663 ^ n662 ;
  assign n665 = ~x129 & ~n664 ;
  assign n671 = x77 ^ x43 ;
  assign n674 = ~n230 & ~n671 ;
  assign n675 = n674 ^ x43 ;
  assign n676 = ~n675 & n702 ;
  assign n666 = n231 & n256 ;
  assign n667 = n666 ^ x43 ;
  assign n668 = n607 & ~n667 ;
  assign n669 = n668 ^ x129 ;
  assign n677 = n676 ^ n669 ;
  assign n678 = ~x129 & ~n658 ;
  assign n679 = x67 ^ x44 ;
  assign n682 = n230 & ~n679 ;
  assign n683 = n682 ^ x67 ;
  assign n684 = n683 & n688 ;
  assign n685 = n678 & ~n684 ;
  assign n689 = ~x68 & n688 ;
  assign n690 = ~n230 & n689 ;
  assign n691 = n690 ^ n688 ;
  assign n692 = n691 ^ n686 ;
  assign n693 = ~n252 & ~n408 ;
  assign n694 = x45 & n693 ;
  assign n695 = n694 ^ x129 ;
  assign n696 = ~x129 & ~n695 ;
  assign n697 = n692 & n696 ;
  assign n698 = n697 ^ x129 ;
  assign n703 = x75 ^ x46 ;
  assign n706 = ~n230 & ~n703 ;
  assign n707 = n706 ^ x46 ;
  assign n708 = n702 & ~n707 ;
  assign n709 = n708 ^ n701 ;
  assign n718 = ~x43 & n666 ;
  assign n719 = n718 ^ x47 ;
  assign n240 = n234 & n239 ;
  assign n241 = x82 & ~n240 ;
  assign n710 = ~x129 & ~n241 ;
  assign n711 = x64 ^ x47 ;
  assign n714 = ~n230 & ~n711 ;
  assign n715 = n714 ^ x47 ;
  assign n716 = n710 & ~n715 ;
  assign n717 = n716 ^ x129 ;
  assign n720 = x82 & ~n717 ;
  assign n721 = ~n719 & n720 ;
  assign n722 = n721 ^ n717 ;
  assign n723 = ~x47 & n718 ;
  assign n724 = n723 ^ x48 ;
  assign n725 = x62 ^ x48 ;
  assign n726 = ~n230 & ~n725 ;
  assign n727 = n726 ^ x48 ;
  assign n728 = ~n687 & ~n727 ;
  assign n729 = ~x129 & n728 ;
  assign n734 = ~n726 & n729 ;
  assign n735 = n734 ^ x129 ;
  assign n736 = n724 & ~n735 ;
  assign n730 = n729 ^ x129 ;
  assign n737 = n736 ^ n730 ;
  assign n738 = x82 & ~n737 ;
  assign n739 = n738 ^ n730 ;
  assign n746 = x49 & ~n252 ;
  assign n743 = ~x69 & ~n230 ;
  assign n744 = n688 & n743 ;
  assign n740 = n688 ^ x24 ;
  assign n741 = n409 & ~n740 ;
  assign n745 = n744 ^ n741 ;
  assign n747 = n746 ^ n745 ;
  assign n748 = ~x129 & n747 ;
  assign n253 = n252 ^ x82 ;
  assign n243 = x82 & ~n242 ;
  assign n751 = n253 ^ n243 ;
  assign n752 = n240 & n751 ;
  assign n753 = ~x66 & n752 ;
  assign n754 = ~n230 & n753 ;
  assign n755 = n754 ^ n752 ;
  assign n756 = n755 ^ n751 ;
  assign n757 = n756 ^ x50 ;
  assign n758 = n757 ^ n246 ;
  assign n759 = n758 ^ n756 ;
  assign n760 = ~x82 & ~n759 ;
  assign n761 = n760 ^ n246 ;
  assign n762 = n756 ^ x38 ;
  assign n763 = n760 ^ n759 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = n764 ^ x38 ;
  assign n766 = n765 ^ n762 ;
  assign n767 = ~n761 & n766 ;
  assign n768 = n767 ^ n764 ;
  assign n769 = n768 ^ x50 ;
  assign n770 = n769 ^ n756 ;
  assign n771 = ~x129 & n770 ;
  assign n772 = x66 & n252 ;
  assign n773 = n771 & n772 ;
  assign n774 = n773 ^ n771 ;
  assign n775 = x109 ^ x51 ;
  assign n776 = n618 & ~n775 ;
  assign n777 = n776 ^ x129 ;
  assign n778 = n619 ^ x52 ;
  assign n779 = n618 & ~n778 ;
  assign n780 = n779 ^ x129 ;
  assign n781 = ~x129 & ~n250 ;
  assign n782 = ~x114 & ~x122 ;
  assign n783 = n782 ^ x122 ;
  assign n784 = ~n274 & ~n783 ;
  assign n785 = n452 ^ n445 ;
  assign n786 = n211 & n785 ;
  assign n788 = x58 & x116 ;
  assign n787 = n464 ^ x58 ;
  assign n789 = n788 ^ n787 ;
  assign n790 = n464 ^ x94 ;
  assign n791 = n790 ^ n788 ;
  assign n792 = n791 ^ x94 ;
  assign n795 = ~x37 & ~n792 ;
  assign n796 = n795 ^ x94 ;
  assign n797 = ~n789 & ~n796 ;
  assign n798 = n797 ^ x94 ;
  assign n799 = n786 & n798 ;
  assign n800 = x60 ^ x57 ;
  assign n803 = ~n788 & n800 ;
  assign n804 = n803 ^ x60 ;
  assign n805 = n786 & n804 ;
  assign n811 = n421 & n433 ;
  assign n806 = n788 ^ x58 ;
  assign n812 = n811 ^ n806 ;
  assign n813 = n786 & n812 ;
  assign n815 = x96 & n461 ;
  assign n814 = x59 & n520 ;
  assign n816 = n815 ^ n814 ;
  assign n817 = n211 & n816 ;
  assign n818 = ~x117 & ~x122 ;
  assign n819 = x123 ^ x60 ;
  assign n820 = n818 & n819 ;
  assign n821 = n820 ^ x60 ;
  assign n822 = n273 & n782 ;
  assign n823 = x140 ^ x62 ;
  assign n824 = x132 & x133 ;
  assign n825 = x131 & n824 ;
  assign n826 = ~x138 & n825 ;
  assign n827 = x136 & x137 ;
  assign n828 = n827 ^ x136 ;
  assign n829 = n826 & n828 ;
  assign n832 = ~n823 & n829 ;
  assign n833 = n832 ^ x62 ;
  assign n834 = ~x129 & n833 ;
  assign n835 = x142 ^ x63 ;
  assign n838 = n829 & ~n835 ;
  assign n839 = n838 ^ x63 ;
  assign n840 = ~x129 & n839 ;
  assign n841 = x139 ^ x64 ;
  assign n844 = n829 & ~n841 ;
  assign n845 = n844 ^ x64 ;
  assign n846 = ~x129 & n845 ;
  assign n847 = x146 ^ x65 ;
  assign n850 = n829 & ~n847 ;
  assign n851 = n850 ^ x65 ;
  assign n852 = ~x129 & n851 ;
  assign n853 = x143 ^ x66 ;
  assign n854 = n827 ^ x137 ;
  assign n855 = n854 ^ x136 ;
  assign n856 = n826 & ~n855 ;
  assign n859 = ~n853 & n856 ;
  assign n860 = n859 ^ x66 ;
  assign n861 = ~x129 & n860 ;
  assign n862 = x139 ^ x67 ;
  assign n865 = n856 & ~n862 ;
  assign n866 = n865 ^ x67 ;
  assign n867 = ~x129 & n866 ;
  assign n868 = x141 ^ x68 ;
  assign n871 = n829 & ~n868 ;
  assign n872 = n871 ^ x68 ;
  assign n873 = ~x129 & n872 ;
  assign n874 = x143 ^ x69 ;
  assign n877 = n829 & ~n874 ;
  assign n878 = n877 ^ x69 ;
  assign n879 = ~x129 & n878 ;
  assign n880 = x144 ^ x70 ;
  assign n883 = n829 & ~n880 ;
  assign n884 = n883 ^ x70 ;
  assign n885 = ~x129 & n884 ;
  assign n886 = x145 ^ x71 ;
  assign n889 = n829 & ~n886 ;
  assign n890 = n889 ^ x71 ;
  assign n891 = ~x129 & n890 ;
  assign n892 = x140 ^ x72 ;
  assign n895 = n856 & ~n892 ;
  assign n896 = n895 ^ x72 ;
  assign n897 = ~x129 & n896 ;
  assign n898 = x141 ^ x73 ;
  assign n901 = n856 & ~n898 ;
  assign n902 = n901 ^ x73 ;
  assign n903 = ~x129 & n902 ;
  assign n904 = x142 ^ x74 ;
  assign n907 = n856 & ~n904 ;
  assign n908 = n907 ^ x74 ;
  assign n909 = ~x129 & n908 ;
  assign n910 = x144 ^ x75 ;
  assign n913 = n856 & ~n910 ;
  assign n914 = n913 ^ x75 ;
  assign n915 = ~x129 & n914 ;
  assign n916 = x145 ^ x76 ;
  assign n919 = n856 & ~n916 ;
  assign n920 = n919 ^ x76 ;
  assign n921 = ~x129 & n920 ;
  assign n922 = x146 ^ x77 ;
  assign n925 = n856 & ~n922 ;
  assign n926 = n925 ^ x77 ;
  assign n927 = ~x129 & n926 ;
  assign n928 = x142 ^ x78 ;
  assign n929 = n826 & n854 ;
  assign n932 = n928 & n929 ;
  assign n933 = n932 ^ x78 ;
  assign n934 = ~x129 & n933 ;
  assign n935 = x143 ^ x79 ;
  assign n938 = n929 & n935 ;
  assign n939 = n938 ^ x79 ;
  assign n940 = ~x129 & n939 ;
  assign n941 = x144 ^ x80 ;
  assign n944 = n929 & n941 ;
  assign n945 = n944 ^ x80 ;
  assign n946 = ~x129 & n945 ;
  assign n947 = x145 ^ x81 ;
  assign n950 = n929 & n947 ;
  assign n951 = n950 ^ x81 ;
  assign n952 = ~x129 & n951 ;
  assign n953 = x146 ^ x82 ;
  assign n956 = n929 & n953 ;
  assign n957 = n956 ^ x82 ;
  assign n958 = ~x129 & n957 ;
  assign n976 = x89 & ~x137 ;
  assign n968 = x138 ^ x136 ;
  assign n969 = x89 ^ x62 ;
  assign n970 = n969 ^ x31 ;
  assign n973 = ~x137 & ~n970 ;
  assign n974 = n973 ^ x31 ;
  assign n975 = n968 & n974 ;
  assign n977 = n976 ^ n975 ;
  assign n959 = x115 ^ x87 ;
  assign n960 = x138 & ~n959 ;
  assign n961 = n960 ^ x87 ;
  assign n978 = n977 ^ n961 ;
  assign n962 = n961 ^ x72 ;
  assign n963 = n962 ^ x119 ;
  assign n964 = n963 ^ n961 ;
  assign n965 = x138 & ~n964 ;
  assign n966 = n965 ^ n962 ;
  assign n967 = ~x137 & ~n966 ;
  assign n979 = n978 ^ n967 ;
  assign n980 = ~x136 & n979 ;
  assign n981 = n980 ^ n977 ;
  assign n982 = x141 ^ x84 ;
  assign n985 = n929 & n982 ;
  assign n986 = n985 ^ x84 ;
  assign n987 = ~x129 & n986 ;
  assign n990 = x96 & ~n459 ;
  assign n991 = n990 ^ x116 ;
  assign n992 = ~x85 & ~n991 ;
  assign n993 = n992 ^ x116 ;
  assign n994 = n429 & ~n993 ;
  assign n995 = x139 ^ x86 ;
  assign n998 = n929 & n995 ;
  assign n999 = n998 ^ x86 ;
  assign n1000 = ~x129 & n999 ;
  assign n1001 = x140 ^ x87 ;
  assign n1004 = n929 & n1001 ;
  assign n1005 = n1004 ^ x87 ;
  assign n1006 = ~x129 & n1005 ;
  assign n1007 = x139 ^ x88 ;
  assign n1008 = n826 & n827 ;
  assign n1011 = n1007 & n1008 ;
  assign n1012 = n1011 ^ x88 ;
  assign n1013 = ~x129 & n1012 ;
  assign n1014 = x140 ^ x89 ;
  assign n1017 = n1008 & n1014 ;
  assign n1018 = n1017 ^ x89 ;
  assign n1019 = ~x129 & n1018 ;
  assign n1020 = x142 ^ x90 ;
  assign n1023 = n1008 & n1020 ;
  assign n1024 = n1023 ^ x90 ;
  assign n1025 = ~x129 & n1024 ;
  assign n1026 = x143 ^ x91 ;
  assign n1029 = n1008 & n1026 ;
  assign n1030 = n1029 ^ x91 ;
  assign n1031 = ~x129 & n1030 ;
  assign n1032 = x144 ^ x92 ;
  assign n1035 = n1008 & n1032 ;
  assign n1036 = n1035 ^ x92 ;
  assign n1037 = ~x129 & n1036 ;
  assign n1038 = x146 ^ x93 ;
  assign n1041 = n1008 & n1038 ;
  assign n1042 = n1041 ^ x93 ;
  assign n1043 = ~x129 & n1042 ;
  assign n1044 = x142 ^ x94 ;
  assign n1045 = x82 & x138 ;
  assign n1046 = ~n855 & n1045 ;
  assign n1047 = n825 & n1046 ;
  assign n1050 = n1044 & n1047 ;
  assign n1051 = n1050 ^ x94 ;
  assign n1052 = ~x129 & n1051 ;
  assign n1055 = ~x3 & ~x110 ;
  assign n1056 = ~n825 & ~n1055 ;
  assign n1057 = x95 & ~n1056 ;
  assign n1058 = n1057 ^ x143 ;
  assign n1059 = ~n1047 & n1058 ;
  assign n1060 = n1059 ^ x143 ;
  assign n1061 = ~x129 & n1060 ;
  assign n1064 = x96 & ~n1056 ;
  assign n1065 = n1064 ^ x146 ;
  assign n1066 = ~n1047 & n1065 ;
  assign n1067 = n1066 ^ x146 ;
  assign n1068 = ~x129 & n1067 ;
  assign n1071 = x97 & ~n1056 ;
  assign n1072 = n1071 ^ x145 ;
  assign n1073 = ~n1047 & n1072 ;
  assign n1074 = n1073 ^ x145 ;
  assign n1075 = ~x129 & n1074 ;
  assign n1076 = x145 ^ x98 ;
  assign n1079 = n1008 & n1076 ;
  assign n1080 = n1079 ^ x98 ;
  assign n1081 = ~x129 & n1080 ;
  assign n1082 = x141 ^ x99 ;
  assign n1085 = n1008 & n1082 ;
  assign n1086 = n1085 ^ x99 ;
  assign n1087 = ~x129 & n1086 ;
  assign n1090 = x100 & ~n1056 ;
  assign n1091 = n1090 ^ x144 ;
  assign n1092 = ~n1047 & n1091 ;
  assign n1093 = n1092 ^ x144 ;
  assign n1094 = ~x129 & n1093 ;
  assign n1095 = x124 ^ x77 ;
  assign n1096 = x138 & ~n1095 ;
  assign n1097 = n1096 ^ x77 ;
  assign n1117 = ~n855 & ~n1097 ;
  assign n1106 = x138 ^ x137 ;
  assign n1107 = x82 ^ x65 ;
  assign n1108 = n1107 ^ x37 ;
  assign n1109 = x136 & ~n1108 ;
  assign n1110 = n1109 ^ x82 ;
  assign n1111 = n1106 & n1110 ;
  assign n1105 = ~x65 & x136 ;
  assign n1112 = n1111 ^ n1105 ;
  assign n1098 = x137 ^ x136 ;
  assign n1099 = x96 ^ x93 ;
  assign n1102 = ~x137 & n1099 ;
  assign n1103 = n1102 ^ x96 ;
  assign n1104 = n1098 & n1103 ;
  assign n1113 = n1112 ^ n1104 ;
  assign n1114 = x138 & n1113 ;
  assign n1115 = n1114 ^ n1112 ;
  assign n1118 = n1117 ^ n1115 ;
  assign n1125 = x69 ^ x66 ;
  assign n1126 = x136 & n1125 ;
  assign n1127 = n1126 ^ x66 ;
  assign n1129 = n1127 ^ x34 ;
  assign n1128 = n1127 ^ x79 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1133 = x136 & n1130 ;
  assign n1134 = n1133 ^ n1128 ;
  assign n1135 = x137 & ~n1134 ;
  assign n1136 = n1135 ^ n1127 ;
  assign n1119 = x95 ^ x91 ;
  assign n1122 = ~x137 & n1119 ;
  assign n1123 = n1122 ^ x95 ;
  assign n1124 = n1098 & n1123 ;
  assign n1137 = n1136 ^ n1124 ;
  assign n1138 = x138 & ~n1137 ;
  assign n1139 = n1138 ^ n1136 ;
  assign n1145 = ~x74 & ~x137 ;
  assign n1140 = x63 ^ x33 ;
  assign n1141 = ~x137 & ~n1140 ;
  assign n1142 = n1141 ^ x33 ;
  assign n1146 = n1145 ^ n1142 ;
  assign n1147 = ~x136 & n1146 ;
  assign n1148 = n1147 ^ n1142 ;
  assign n1149 = ~x138 & n1148 ;
  assign n1150 = n1149 ^ x138 ;
  assign n1161 = x78 & n854 ;
  assign n1162 = ~n1150 & n1161 ;
  assign n1153 = x94 ^ x90 ;
  assign n1156 = x137 & n1153 ;
  assign n1157 = n1156 ^ x90 ;
  assign n1158 = n1098 & n1157 ;
  assign n1159 = x138 & n1158 ;
  assign n1160 = n1159 ^ n1149 ;
  assign n1163 = n1162 ^ n1160 ;
  assign n1171 = x73 ^ x68 ;
  assign n1172 = ~x136 & n1171 ;
  assign n1173 = n1172 ^ x68 ;
  assign n1175 = n1173 ^ x32 ;
  assign n1174 = n1173 ^ x84 ;
  assign n1176 = n1175 ^ n1174 ;
  assign n1179 = x136 & n1176 ;
  assign n1180 = n1179 ^ n1174 ;
  assign n1181 = x137 & ~n1180 ;
  assign n1182 = n1181 ^ n1173 ;
  assign n1164 = x138 ^ x112 ;
  assign n1165 = n1164 ^ x99 ;
  assign n1168 = x137 & n1165 ;
  assign n1169 = n1168 ^ x99 ;
  assign n1170 = n1098 & n1169 ;
  assign n1183 = n1182 ^ n1170 ;
  assign n1184 = x138 & ~n1183 ;
  assign n1185 = n1184 ^ n1182 ;
  assign n1204 = x125 ^ x92 ;
  assign n1205 = n1204 ^ x100 ;
  assign n1206 = ~x137 & n1205 ;
  assign n1207 = n1206 ^ x100 ;
  assign n1208 = x136 & n1207 ;
  assign n1188 = x80 ^ x75 ;
  assign n1189 = x137 & ~n1188 ;
  assign n1190 = n1189 ^ x75 ;
  assign n1192 = n1190 ^ x35 ;
  assign n1191 = n1190 ^ x70 ;
  assign n1193 = n1192 ^ n1191 ;
  assign n1196 = x137 & ~n1193 ;
  assign n1197 = n1196 ^ n1191 ;
  assign n1198 = x136 & n1197 ;
  assign n1199 = n1198 ^ n1190 ;
  assign n1200 = n1199 ^ x100 ;
  assign n1209 = n1208 ^ n1200 ;
  assign n1186 = x125 ^ x100 ;
  assign n1187 = ~x137 & n1186 ;
  assign n1210 = n1209 ^ n1187 ;
  assign n1211 = x138 & ~n1210 ;
  assign n1212 = n1211 ^ n1199 ;
  assign n1213 = n480 ^ n461 ;
  assign n1214 = n211 & n1213 ;
  assign n1233 = x98 & ~x137 ;
  assign n1226 = x71 ^ x36 ;
  assign n1227 = ~x137 & ~n1226 ;
  assign n1228 = n1227 ^ x36 ;
  assign n1234 = n1233 ^ n1228 ;
  assign n1235 = x138 & n1234 ;
  assign n1236 = n1235 ^ n1228 ;
  assign n1215 = x76 ^ x23 ;
  assign n1216 = ~x138 & ~n1215 ;
  assign n1217 = n1216 ^ x23 ;
  assign n1237 = n1236 ^ n1217 ;
  assign n1219 = n1217 ^ x81 ;
  assign n1218 = n1217 ^ x97 ;
  assign n1220 = n1219 ^ n1218 ;
  assign n1223 = ~x138 & n1220 ;
  assign n1224 = n1223 ^ n1218 ;
  assign n1225 = x137 & n1224 ;
  assign n1238 = n1237 ^ n1225 ;
  assign n1239 = ~x136 & n1238 ;
  assign n1240 = n1239 ^ n1236 ;
  assign n1259 = x88 & ~x137 ;
  assign n1252 = x88 ^ x64 ;
  assign n1253 = n1252 ^ x30 ;
  assign n1256 = ~x137 & ~n1253 ;
  assign n1257 = n1256 ^ x30 ;
  assign n1258 = n968 & n1257 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n1241 = x120 ^ x67 ;
  assign n1242 = x138 & ~n1241 ;
  assign n1243 = n1242 ^ x67 ;
  assign n1261 = n1260 ^ n1243 ;
  assign n1245 = n1243 ^ x86 ;
  assign n1244 = n1243 ^ x111 ;
  assign n1246 = n1245 ^ n1244 ;
  assign n1249 = ~x138 & n1246 ;
  assign n1250 = n1249 ^ n1244 ;
  assign n1251 = x137 & ~n1250 ;
  assign n1262 = n1261 ^ n1251 ;
  assign n1263 = ~x136 & ~n1262 ;
  assign n1264 = n1263 ^ n1260 ;
  assign n1265 = x116 & n211 ;
  assign n1270 = n419 & ~n433 ;
  assign n1271 = n1270 ^ n443 ;
  assign n1272 = n1265 & n1271 ;
  assign n1273 = n448 & n1265 ;
  assign n1274 = ~x53 & x97 ;
  assign n1275 = n1273 & n1274 ;
  assign n1276 = n1275 ^ n1273 ;
  assign n1277 = ~x129 & n825 ;
  assign n1278 = x139 ^ x111 ;
  assign n1281 = ~n1046 & n1278 ;
  assign n1282 = n1281 ^ x139 ;
  assign n1283 = n1277 & n1282 ;
  assign n1284 = x141 ^ x112 ;
  assign n1287 = ~n1046 & ~n1284 ;
  assign n1288 = n1287 ^ x141 ;
  assign n1289 = n1277 & n1288 ;
  assign n1290 = n219 ^ x113 ;
  assign n1293 = x54 & n1290 ;
  assign n1294 = n1293 ^ x113 ;
  assign n1295 = n211 & ~n1294 ;
  assign n1296 = x140 ^ x115 ;
  assign n1299 = ~n1046 & ~n1296 ;
  assign n1300 = n1299 ^ x140 ;
  assign n1301 = n1277 & n1300 ;
  assign n1302 = ~n156 & n215 ;
  assign n1303 = x122 & ~x129 ;
  assign n1308 = ~x54 & x118 ;
  assign n1309 = n1308 ^ n329 ;
  assign n1310 = ~x129 & n1309 ;
  assign n1311 = ~x129 & ~n456 ;
  assign n1312 = ~x120 & n1055 ;
  assign n1313 = ~x111 & ~x129 ;
  assign n1314 = ~n1312 & n1313 ;
  assign n1315 = x81 & x120 ;
  assign n1316 = ~x129 & n1315 ;
  assign n1317 = ~x129 & ~x134 ;
  assign n1318 = ~x129 & ~x135 ;
  assign n1319 = x57 & ~x129 ;
  assign n1322 = n211 ^ x129 ;
  assign n1320 = ~x96 & x125 ;
  assign n1321 = n211 & n1320 ;
  assign n1323 = n1322 ^ n1321 ;
  assign n1324 = ~x126 & n824 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = ~n212 ;
  assign y16 = ~n229 ;
  assign y17 = n267 ;
  assign y18 = ~n276 ;
  assign y19 = n282 ;
  assign y20 = n293 ;
  assign y21 = n298 ;
  assign y22 = n301 ;
  assign y23 = n304 ;
  assign y24 = n310 ;
  assign y25 = n313 ;
  assign y26 = n321 ;
  assign y27 = n326 ;
  assign y28 = n334 ;
  assign y29 = n337 ;
  assign y30 = n359 ;
  assign y31 = n362 ;
  assign y32 = n368 ;
  assign y33 = n371 ;
  assign y34 = n374 ;
  assign y35 = n398 ;
  assign y36 = n401 ;
  assign y37 = n403 ;
  assign y38 = n406 ;
  assign y39 = n418 ;
  assign y40 = n472 ;
  assign y41 = n478 ;
  assign y42 = n487 ;
  assign y43 = n505 ;
  assign y44 = n525 ;
  assign y45 = n535 ;
  assign y46 = n545 ;
  assign y47 = n555 ;
  assign y48 = n565 ;
  assign y49 = n575 ;
  assign y50 = n585 ;
  assign y51 = n595 ;
  assign y52 = n605 ;
  assign y53 = ~n617 ;
  assign y54 = ~n627 ;
  assign y55 = n640 ;
  assign y56 = ~n656 ;
  assign y57 = n665 ;
  assign y58 = ~n677 ;
  assign y59 = n685 ;
  assign y60 = ~n698 ;
  assign y61 = ~n709 ;
  assign y62 = ~n722 ;
  assign y63 = ~n739 ;
  assign y64 = n748 ;
  assign y65 = n774 ;
  assign y66 = ~n777 ;
  assign y67 = ~n780 ;
  assign y68 = n518 ;
  assign y69 = ~n781 ;
  assign y70 = n784 ;
  assign y71 = n799 ;
  assign y72 = n805 ;
  assign y73 = n813 ;
  assign y74 = n817 ;
  assign y75 = n821 ;
  assign y76 = n822 ;
  assign y77 = ~n834 ;
  assign y78 = ~n840 ;
  assign y79 = ~n846 ;
  assign y80 = ~n852 ;
  assign y81 = ~n861 ;
  assign y82 = ~n867 ;
  assign y83 = ~n873 ;
  assign y84 = ~n879 ;
  assign y85 = ~n885 ;
  assign y86 = ~n891 ;
  assign y87 = ~n897 ;
  assign y88 = ~n903 ;
  assign y89 = ~n909 ;
  assign y90 = ~n915 ;
  assign y91 = ~n921 ;
  assign y92 = ~n927 ;
  assign y93 = n934 ;
  assign y94 = n940 ;
  assign y95 = n946 ;
  assign y96 = n952 ;
  assign y97 = n958 ;
  assign y98 = n981 ;
  assign y99 = n987 ;
  assign y100 = n994 ;
  assign y101 = n1000 ;
  assign y102 = n1006 ;
  assign y103 = n1013 ;
  assign y104 = n1019 ;
  assign y105 = n1025 ;
  assign y106 = n1031 ;
  assign y107 = n1037 ;
  assign y108 = n1043 ;
  assign y109 = n1052 ;
  assign y110 = n1061 ;
  assign y111 = n1068 ;
  assign y112 = n1075 ;
  assign y113 = n1081 ;
  assign y114 = n1087 ;
  assign y115 = n1094 ;
  assign y116 = n1118 ;
  assign y117 = ~n1139 ;
  assign y118 = n1163 ;
  assign y119 = ~n1185 ;
  assign y120 = ~n1212 ;
  assign y121 = n1214 ;
  assign y122 = n1240 ;
  assign y123 = n1264 ;
  assign y124 = n1272 ;
  assign y125 = n1276 ;
  assign y126 = n1283 ;
  assign y127 = n1289 ;
  assign y128 = n1295 ;
  assign y129 = n274 ;
  assign y130 = n1301 ;
  assign y131 = n1302 ;
  assign y132 = ~n1303 ;
  assign y133 = n1310 ;
  assign y134 = n1311 ;
  assign y135 = n1314 ;
  assign y136 = n1316 ;
  assign y137 = ~n1317 ;
  assign y138 = ~n1318 ;
  assign y139 = n1319 ;
  assign y140 = ~n1323 ;
  assign y141 = n1324 ;
endmodule
