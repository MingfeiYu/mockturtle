module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 ;
  output y0 ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1056 , n1057 , n1058 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1072 , n1073 , n1074 , n1075 , n1076 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1287 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1373 , n1374 , n1375 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1417 , n1424 , n1425 , n1426 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1442 , n1443 , n1446 , n1447 , n1448 , n1450 , n1451 , n1452 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1578 , n1579 , n1580 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1633 , n1634 , n1635 , n1636 , n1637 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1681 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1721 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1761 , n1762 , n1763 , n1764 , n1767 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1793 , n1794 , n1795 , n1796 , n1799 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1834 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1875 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2195 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2240 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2282 , n2283 , n2284 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2313 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2431 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2474 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2562 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2702 , n2703 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2768 , n2769 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2917 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3114 , n3115 , n3116 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3144 , n3146 , n3148 , n3149 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3166 , n3167 , n3168 , n3171 , n3172 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3317 , n3318 , n3319 , n3320 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3364 , n3365 , n3366 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3478 , n3479 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3509 , n3510 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3572 , n3573 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3623 , n3630 , n3631 , n3632 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3648 , n3649 , n3652 , n3653 , n3654 , n3656 , n3657 , n3658 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3683 , n3684 , n3685 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3697 , n3698 , n3699 , n3700 , n3702 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3896 , n3897 , n3898 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4194 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4212 , n4217 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4346 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4371 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4415 , n4416 , n4417 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4490 , n4491 , n4492 , n4493 , n4494 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4621 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4663 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4693 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4706 , n4707 , n4708 , n4709 , n4710 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4746 , n4750 , n4751 , n4758 , n4760 , n4761 , n4762 , n4763 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4911 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4936 , n4939 , n4940 , n4941 , n4942 , n4943 , n4945 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4970 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5078 , n5079 , n5080 , n5081 , n5082 , n5087 , n5094 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5124 , n5125 , n5128 , n5129 , n5130 , n5132 , n5133 , n5134 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5192 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5216 , n5217 , n5218 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5263 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5288 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5454 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5491 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5554 , n5555 , n5556 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5639 , n5640 , n5641 , n5642 , n5643 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5803 , n5804 , n5805 , n5806 , n5807 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5837 , n5838 , n5839 , n5840 , n5841 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5916 , n5917 , n5920 , n5921 , n5922 , n5924 , n5925 , n5926 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5972 , n5973 , n5976 , n5977 , n5978 , n5980 , n5981 , n5982 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5998 , n5999 , n6001 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6031 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6265 , n6266 , n6267 , n6268 , n6269 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6363 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6406 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6712 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6750 , n6751 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6770 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6795 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6922 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7144 , n7148 , n7160 , n7161 , n7162 , n7179 , n7180 , n7181 , n7182 , n7185 , n7186 , n7187 , n7189 , n7190 , n7191 , n7192 , n7193 , n7198 , n7203 , n7206 , n7207 , n7214 , n7215 , n7218 , n7219 , n7220 , n7221 , n7222 , n7227 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7449 , n7450 , n7451 , n7452 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7523 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7577 , n7579 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7714 , n7715 , n7716 , n7717 , n7718 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7771 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7796 , n7799 , n7800 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7814 , n7815 , n7818 , n7819 , n7820 , n7822 , n7823 , n7824 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7915 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7940 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7961 , n7963 , n7966 , n7967 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8033 , n8034 , n8035 , n8036 , n8038 , n8039 , n8040 , n8041 , n8042 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8139 , n8140 , n8143 , n8144 , n8145 , n8147 , n8151 , n8152 , n8153 , n8154 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8169 , n8170 , n8171 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8188 , n8189 , n8190 , n8191 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8232 , n8233 , n8234 , n8237 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8331 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8374 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8443 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8491 , n8494 , n8495 , n8496 , n8498 , n8502 , n8503 , n8504 , n8505 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8520 , n8521 , n8522 , n8523 , n8524 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8558 , n8559 , n8560 , n8561 , n8562 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8807 , n8808 , n8809 , n8810 , n8813 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8834 , n8835 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8865 , n8866 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8899 , n8900 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8927 , n8928 , n8931 , n8932 , n8933 , n8935 , n8936 , n8937 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8950 , n8951 , n8954 , n8955 , n8956 , n8958 , n8959 , n8960 , n8963 , n8964 , n8965 , n8966 , n8967 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9075 , n9076 , n9077 , n9078 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9162 , n9163 , n9164 , n9165 , n9166 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9285 , n9286 , n9289 , n9290 , n9291 , n9292 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9303 , n9304 , n9305 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9401 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9444 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9538 , n9539 , n9540 , n9541 , n9542 , n9548 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9560 , n9561 , n9562 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9573 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9598 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9616 , n9617 , n9618 , n9619 , n9622 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9680 , n9681 , n9682 , n9683 , n9684 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9712 , n9713 , n9719 , n9720 , n9723 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9749 , n9750 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9769 , n9770 , n9771 , n9772 , n9773 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9845 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9856 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10016 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10041 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10084 , n10085 , n10088 , n10089 , n10090 , n10092 , n10093 , n10094 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10154 , n10155 , n10156 , n10157 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10169 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10255 , n10256 , n10257 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10334 , n10335 , n10336 , n10337 , n10340 , n10341 , n10342 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10365 , n10366 , n10367 , n10369 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10424 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10449 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10608 , n10611 , n10612 , n10613 , n10614 , n10615 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10677 , n10678 , n10679 , n10680 , n10681 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10744 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10963 , n10964 , n10965 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11157 , n11158 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11197 , n11200 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11235 , n11236 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11273 , n11274 , n11275 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11456 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11496 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11626 , n11627 , n11628 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11689 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11714 , n11717 , n11718 , n11719 , n11720 , n11721 , n11723 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11748 , n11751 , n11752 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11768 , n11769 , n11770 , n11771 , n11773 , n11774 , n11775 , n11776 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11792 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11999 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12097 , n12098 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12123 , n12124 , n12125 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12164 , n12165 , n12166 , n12167 , n12168 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12190 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12424 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12480 , n12481 , n12483 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12493 , n12494 , n12495 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12543 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12557 , n12558 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12573 , n12574 , n12575 , n12576 , n12579 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12629 , n12630 , n12631 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12663 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12678 , n12679 , n12680 , n12681 , n12684 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12705 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12718 , n12719 , n12720 , n12721 , n12722 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12741 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12900 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12925 , n12928 , n12929 , n12930 , n12931 , n12932 , n12934 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12959 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n13003 , n13004 , n13005 , n13008 , n13009 , n13014 , n13015 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13050 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13140 , n13141 , n13145 , n13146 , n13147 , n13148 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13215 , n13216 , n13217 , n13219 , n13221 , n13223 , n13224 , n13227 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13518 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 ;
  assign n5361 = x197 & x198 ;
  assign n5362 = x195 & x196 ;
  assign n5363 = n5361 & n5362 ;
  assign n5371 = n5362 ^ n5361 ;
  assign n5372 = n5371 ^ n5363 ;
  assign n5366 = x198 ^ x197 ;
  assign n5367 = n5366 ^ n5361 ;
  assign n5364 = x196 ^ x195 ;
  assign n5365 = n5364 ^ n5362 ;
  assign n5369 = n5367 ^ n5365 ;
  assign n5368 = ~n5365 & ~n5367 ;
  assign n5370 = n5369 ^ n5368 ;
  assign n5373 = n5372 ^ n5370 ;
  assign n5374 = x194 ^ x193 ;
  assign n5375 = n5374 ^ n5372 ;
  assign n5376 = n5373 & ~n5375 ;
  assign n5377 = x193 & x194 ;
  assign n5378 = ~n5363 & n5377 ;
  assign n5379 = n5378 ^ n5374 ;
  assign n5380 = n5376 & n5379 ;
  assign n5381 = n5380 ^ n5378 ;
  assign n5382 = ~n5363 & ~n5381 ;
  assign n5394 = n5382 ^ n5381 ;
  assign n5390 = n5374 ^ n5365 ;
  assign n5391 = n5390 ^ n5367 ;
  assign n5392 = ~n5368 & ~n5391 ;
  assign n5393 = n5373 & ~n5392 ;
  assign n5395 = n5394 ^ n5393 ;
  assign n5396 = n5395 ^ n5377 ;
  assign n5322 = x190 ^ x189 ;
  assign n5319 = x192 ^ x191 ;
  assign n5385 = n5322 ^ n5319 ;
  assign n5384 = x188 ^ x187 ;
  assign n5386 = n5385 ^ n5384 ;
  assign n5387 = n5374 ^ n5366 ;
  assign n5388 = n5387 ^ n5364 ;
  assign n5389 = n5386 & n5388 ;
  assign n5397 = n5396 ^ n5389 ;
  assign n5318 = ~x191 & ~x192 ;
  assign n5325 = n5318 ^ x188 ;
  assign n5321 = ~x189 & ~x190 ;
  assign n5326 = n5325 ^ n5321 ;
  assign n5328 = n5321 ^ n5318 ;
  assign n5327 = n5318 & n5321 ;
  assign n5329 = n5328 ^ n5327 ;
  assign n5330 = n5326 & n5329 ;
  assign n5412 = n5327 ^ x187 ;
  assign n5413 = ~n5330 & ~n5412 ;
  assign n5337 = x191 ^ x188 ;
  assign n5338 = n5337 ^ x190 ;
  assign n5339 = n5338 ^ x192 ;
  assign n5335 = x191 ^ x189 ;
  assign n5340 = n5339 ^ n5335 ;
  assign n5341 = n5340 ^ x192 ;
  assign n5342 = n5341 ^ x191 ;
  assign n5343 = n5342 ^ n5335 ;
  assign n5349 = n5385 ^ n5335 ;
  assign n5350 = ~n5343 & ~n5349 ;
  assign n5351 = ~x191 & n5350 ;
  assign n5354 = n5351 ^ n5350 ;
  assign n5352 = n5351 ^ n5335 ;
  assign n5353 = n5340 & n5352 ;
  assign n5355 = n5354 ^ n5353 ;
  assign n5356 = n5355 ^ x191 ;
  assign n5358 = ~x187 & ~n5356 ;
  assign n5409 = n5396 ^ n5358 ;
  assign n5357 = n5356 ^ x187 ;
  assign n5323 = n5322 ^ n5321 ;
  assign n5320 = n5319 ^ n5318 ;
  assign n5324 = n5323 ^ n5320 ;
  assign n5331 = n5326 ^ n5320 ;
  assign n5332 = n5331 ^ n5330 ;
  assign n5333 = n5324 & n5332 ;
  assign n5334 = n5333 ^ n5323 ;
  assign n5400 = n5357 ^ n5334 ;
  assign n5401 = n5400 ^ n5356 ;
  assign n5405 = n5334 & ~n5355 ;
  assign n5406 = n5405 ^ x191 ;
  assign n5407 = n5401 & ~n5406 ;
  assign n5408 = n5407 ^ n5357 ;
  assign n5410 = n5409 ^ n5408 ;
  assign n5398 = n5320 & n5323 ;
  assign n5399 = n5358 & n5398 ;
  assign n5411 = n5410 ^ n5399 ;
  assign n5414 = n5413 ^ n5411 ;
  assign n5415 = n5397 & n5414 ;
  assign n5416 = n5415 ^ n5396 ;
  assign n5359 = n5358 ^ n5357 ;
  assign n5360 = n5334 & n5359 ;
  assign n5383 = n5382 ^ n5360 ;
  assign n5458 = n5416 ^ n5383 ;
  assign n5421 = x179 & x180 ;
  assign n5420 = x180 ^ x179 ;
  assign n5422 = n5421 ^ n5420 ;
  assign n5424 = x177 & x178 ;
  assign n5423 = x178 ^ x177 ;
  assign n5425 = n5424 ^ n5423 ;
  assign n5426 = n5422 & n5425 ;
  assign n5427 = n5426 ^ x176 ;
  assign n5431 = n5424 ^ x176 ;
  assign n5429 = n5424 ^ n5421 ;
  assign n5428 = n5424 ^ x175 ;
  assign n5430 = n5429 ^ n5428 ;
  assign n5432 = n5431 ^ n5430 ;
  assign n5442 = n5427 & n5432 ;
  assign n5448 = n5442 ^ x175 ;
  assign n5444 = n5426 ^ n5421 ;
  assign n5445 = n5444 ^ n5442 ;
  assign n5446 = ~n5429 & n5445 ;
  assign n5449 = n5426 & n5446 ;
  assign n5450 = n5448 & n5449 ;
  assign n5443 = n5442 ^ n5427 ;
  assign n5447 = n5446 ^ n5443 ;
  assign n5451 = n5450 ^ n5447 ;
  assign n5454 = n5451 ^ n5424 ;
  assign n5457 = n5454 ^ n5431 ;
  assign n5459 = n5458 ^ n5457 ;
  assign n5503 = x176 ^ x175 ;
  assign n5504 = n5503 ^ n5423 ;
  assign n5505 = n5504 ^ n5420 ;
  assign n5479 = x182 ^ x181 ;
  assign n5469 = x184 ^ x183 ;
  assign n5506 = n5479 ^ n5469 ;
  assign n5465 = x186 ^ x185 ;
  assign n5507 = n5506 ^ n5465 ;
  assign n5508 = n5505 & n5507 ;
  assign n5461 = x185 ^ x184 ;
  assign n5466 = ~n5461 & ~n5465 ;
  assign n5460 = x183 ^ x182 ;
  assign n5462 = n5461 ^ x183 ;
  assign n5463 = n5462 ^ x186 ;
  assign n5464 = ~n5460 & n5463 ;
  assign n5467 = n5466 ^ n5464 ;
  assign n5468 = ~x181 & n5467 ;
  assign n5470 = x184 ^ x182 ;
  assign n5471 = x186 ^ x181 ;
  assign n5474 = ~x184 & ~n5471 ;
  assign n5475 = n5474 ^ x181 ;
  assign n5476 = ~n5470 & n5475 ;
  assign n5477 = ~n5469 & n5476 ;
  assign n5478 = ~x185 & n5477 ;
  assign n5480 = ~x183 & ~x184 ;
  assign n5486 = ~x185 & ~x186 ;
  assign n5487 = ~n5480 & ~n5486 ;
  assign n5481 = n5480 ^ n5469 ;
  assign n5482 = x181 & x182 ;
  assign n5483 = x186 & n5482 ;
  assign n5484 = ~n5481 & n5483 ;
  assign n5485 = n5484 ^ n5482 ;
  assign n5488 = n5487 ^ n5485 ;
  assign n5491 = n5486 ^ n5465 ;
  assign n5494 = n5481 & n5491 ;
  assign n5495 = n5494 ^ n5485 ;
  assign n5496 = n5488 & ~n5495 ;
  assign n5497 = n5496 ^ n5485 ;
  assign n5498 = ~n5479 & n5497 ;
  assign n5499 = n5496 & n5498 ;
  assign n5500 = n5499 ^ n5497 ;
  assign n5501 = ~n5478 & ~n5500 ;
  assign n5502 = ~n5468 & n5501 ;
  assign n5509 = n5508 ^ n5502 ;
  assign n5515 = n5503 ^ n5424 ;
  assign n5516 = n5515 ^ n5426 ;
  assign n5517 = ~n5429 & ~n5516 ;
  assign n5514 = n5502 ^ x175 ;
  assign n5518 = n5517 ^ n5514 ;
  assign n5519 = n5518 ^ n5426 ;
  assign n5520 = n5519 ^ n5502 ;
  assign n5521 = n5520 ^ n5517 ;
  assign n5522 = ~n5427 & n5521 ;
  assign n5523 = n5522 ^ n5518 ;
  assign n5511 = n5429 ^ n5426 ;
  assign n5510 = n5423 ^ n5420 ;
  assign n5512 = n5511 ^ n5510 ;
  assign n5513 = n5503 & ~n5512 ;
  assign n5526 = n5523 ^ n5513 ;
  assign n5527 = n5509 & n5526 ;
  assign n5528 = n5527 ^ n5508 ;
  assign n5529 = n5528 ^ n5457 ;
  assign n5530 = n5459 & ~n5529 ;
  assign n5531 = n5530 ^ n5458 ;
  assign n5541 = n5491 ^ n5481 ;
  assign n5542 = x182 & n5487 ;
  assign n5543 = n5542 ^ n5481 ;
  assign n5544 = n5541 & ~n5543 ;
  assign n5545 = n5544 ^ n5481 ;
  assign n5546 = ~n5500 & ~n5545 ;
  assign n5547 = n5546 ^ n5500 ;
  assign n5548 = n5547 ^ n5457 ;
  assign n5549 = n5548 ^ n5528 ;
  assign n5550 = n5549 ^ n5458 ;
  assign n5533 = n5414 ^ n5389 ;
  assign n5532 = n5526 ^ n5508 ;
  assign n5534 = n5533 ^ n5532 ;
  assign n5535 = n5388 ^ n5386 ;
  assign n5536 = n5507 ^ n5505 ;
  assign n5537 = n5535 & n5536 ;
  assign n5538 = n5537 ^ n5532 ;
  assign n5539 = ~n5534 & n5538 ;
  assign n5540 = n5539 ^ n5533 ;
  assign n5551 = n5550 ^ n5540 ;
  assign n5552 = n5551 ^ n5547 ;
  assign n5554 = n5550 & ~n5552 ;
  assign n5555 = n5554 ^ n5547 ;
  assign n5588 = ~n5531 & ~n5555 ;
  assign n5417 = n5416 ^ n5360 ;
  assign n5418 = n5383 & n5417 ;
  assign n5419 = n5418 ^ n5382 ;
  assign n5556 = n5555 ^ n5531 ;
  assign n5587 = n5419 & n5556 ;
  assign n5589 = n5588 ^ n5587 ;
  assign n5043 = x209 & x210 ;
  assign n5042 = x210 ^ x209 ;
  assign n5044 = n5043 ^ n5042 ;
  assign n5047 = x207 & x208 ;
  assign n5048 = ~n5044 & ~n5047 ;
  assign n5049 = x205 & x206 ;
  assign n5050 = ~n5048 & n5049 ;
  assign n5051 = x208 ^ x207 ;
  assign n5052 = n5043 ^ x208 ;
  assign n5053 = ~n5051 & ~n5052 ;
  assign n5054 = n5050 & ~n5053 ;
  assign n5045 = x206 ^ x205 ;
  assign n5046 = n5044 & n5045 ;
  assign n5055 = n5053 ^ n5052 ;
  assign n5056 = n5055 ^ x207 ;
  assign n5057 = n5046 & ~n5056 ;
  assign n5058 = ~n5054 & ~n5057 ;
  assign n5299 = n5043 & n5047 ;
  assign n5300 = n5058 & n5299 ;
  assign n5301 = n5300 ^ n5058 ;
  assign n5149 = x222 ^ x221 ;
  assign n5174 = x221 ^ x220 ;
  assign n5178 = ~n5149 & ~n5174 ;
  assign n5173 = x219 ^ x218 ;
  assign n5175 = n5174 ^ x219 ;
  assign n5176 = n5175 ^ x222 ;
  assign n5177 = ~n5173 & n5176 ;
  assign n5179 = n5178 ^ n5177 ;
  assign n5180 = ~x217 & n5179 ;
  assign n5181 = ~x219 & ~x220 ;
  assign n5187 = ~x221 & ~x222 ;
  assign n5188 = ~n5181 & ~n5187 ;
  assign n5152 = x220 ^ x219 ;
  assign n5182 = n5181 ^ n5152 ;
  assign n5183 = x217 & x218 ;
  assign n5184 = x222 & n5183 ;
  assign n5185 = ~n5182 & n5184 ;
  assign n5186 = n5185 ^ n5183 ;
  assign n5189 = n5188 ^ n5186 ;
  assign n5192 = n5187 ^ n5149 ;
  assign n5195 = n5182 & n5192 ;
  assign n5196 = n5195 ^ n5186 ;
  assign n5197 = n5189 & ~n5196 ;
  assign n5150 = x218 ^ x217 ;
  assign n5198 = n5197 ^ n5186 ;
  assign n5199 = ~n5150 & n5198 ;
  assign n5200 = n5197 & n5199 ;
  assign n5201 = n5200 ^ n5198 ;
  assign n5202 = x220 ^ x218 ;
  assign n5203 = x222 ^ x217 ;
  assign n5206 = ~x220 & ~n5203 ;
  assign n5207 = n5206 ^ x217 ;
  assign n5208 = ~n5202 & n5207 ;
  assign n5209 = ~n5152 & n5208 ;
  assign n5210 = ~x221 & n5209 ;
  assign n5211 = ~n5201 & ~n5210 ;
  assign n5212 = ~n5180 & n5211 ;
  assign n5165 = x215 & x216 ;
  assign n5164 = x213 & x214 ;
  assign n5166 = n5165 ^ n5164 ;
  assign n5157 = x214 ^ x213 ;
  assign n5167 = n5164 ^ n5157 ;
  assign n5155 = x216 ^ x215 ;
  assign n5168 = n5165 ^ n5155 ;
  assign n5169 = n5167 & n5168 ;
  assign n5170 = n5169 ^ n5165 ;
  assign n5171 = ~n5166 & ~n5170 ;
  assign n5154 = x212 ^ x211 ;
  assign n5160 = n5157 ^ x212 ;
  assign n5161 = n5160 ^ n5155 ;
  assign n5162 = n5154 & ~n5161 ;
  assign n5163 = n5162 ^ x211 ;
  assign n5172 = n5171 ^ n5163 ;
  assign n5213 = n5212 ^ n5172 ;
  assign n5151 = n5150 ^ n5149 ;
  assign n5153 = n5152 ^ n5151 ;
  assign n5156 = n5155 ^ n5154 ;
  assign n5158 = n5157 ^ n5156 ;
  assign n5159 = n5153 & n5158 ;
  assign n5293 = n5172 ^ n5159 ;
  assign n5294 = ~n5213 & ~n5293 ;
  assign n5295 = n5294 ^ n5172 ;
  assign n5260 = n5164 ^ x211 ;
  assign n5263 = n5260 ^ n5166 ;
  assign n5258 = n5164 ^ x212 ;
  assign n5268 = n5263 ^ n5258 ;
  assign n5259 = n5170 ^ n5166 ;
  assign n5261 = n5260 ^ n5259 ;
  assign n5269 = n5268 ^ n5261 ;
  assign n5270 = n5269 ^ n5166 ;
  assign n5272 = n5268 & n5270 ;
  assign n5265 = n5261 ^ n5166 ;
  assign n5266 = n5265 ^ n5165 ;
  assign n5267 = ~n5169 & n5266 ;
  assign n5273 = n5272 ^ n5267 ;
  assign n5274 = n5273 ^ n5265 ;
  assign n5275 = n5272 ^ n5263 ;
  assign n5276 = n5275 ^ n5265 ;
  assign n5277 = n5274 & n5276 ;
  assign n5278 = ~n5166 & n5277 ;
  assign n5279 = n5278 ^ n5272 ;
  assign n5280 = n5279 ^ n5270 ;
  assign n5288 = n5280 ^ n5164 ;
  assign n5291 = n5288 ^ n5258 ;
  assign n5252 = n5192 ^ n5182 ;
  assign n5253 = x218 & n5188 ;
  assign n5254 = n5253 ^ n5182 ;
  assign n5255 = n5252 & ~n5254 ;
  assign n5256 = n5255 ^ n5182 ;
  assign n5257 = ~n5201 & n5256 ;
  assign n5292 = n5291 ^ n5257 ;
  assign n5296 = n5295 ^ n5292 ;
  assign n5103 = x201 & x202 ;
  assign n5075 = x202 ^ x201 ;
  assign n5104 = n5103 ^ n5075 ;
  assign n5105 = ~x203 & ~x204 ;
  assign n5076 = x204 ^ x203 ;
  assign n5106 = n5105 ^ n5076 ;
  assign n5107 = n5106 ^ n5103 ;
  assign n5108 = x200 & ~n5105 ;
  assign n5109 = n5108 ^ n5103 ;
  assign n5110 = ~n5107 & n5109 ;
  assign n5111 = n5110 ^ n5103 ;
  assign n5112 = n5104 & n5111 ;
  assign n5082 = n5075 ^ x203 ;
  assign n5081 = x204 ^ x200 ;
  assign n5128 = x204 ^ x202 ;
  assign n5096 = ~n5081 & ~n5128 ;
  assign n5097 = ~n5082 & n5096 ;
  assign n5100 = n5097 ^ n5096 ;
  assign n5087 = x203 ^ x201 ;
  assign n5098 = n5097 ^ n5087 ;
  assign n5132 = n5081 ^ n5075 ;
  assign n5099 = n5098 & n5132 ;
  assign n5101 = n5100 ^ n5099 ;
  assign n5102 = n5101 ^ x203 ;
  assign n5146 = x199 & n5102 ;
  assign n5147 = ~n5112 & n5146 ;
  assign n5072 = n5051 ^ n5045 ;
  assign n5073 = n5072 ^ n5042 ;
  assign n5094 = n5082 ^ x204 ;
  assign n5074 = x200 ^ x199 ;
  assign n5078 = n5094 ^ n5074 ;
  assign n5079 = n5073 & n5078 ;
  assign n5059 = ~n5046 & n5058 ;
  assign n5060 = n5051 ^ x205 ;
  assign n5066 = ~x206 & n5048 ;
  assign n5061 = ~x205 & ~n5052 ;
  assign n5067 = n5066 ^ n5061 ;
  assign n5068 = n5060 & n5067 ;
  assign n5069 = n5068 ^ n5061 ;
  assign n5070 = n5059 & n5069 ;
  assign n5071 = n5070 ^ n5058 ;
  assign n5080 = n5079 ^ n5071 ;
  assign n5113 = ~n5104 & n5106 ;
  assign n5114 = ~n5108 & n5113 ;
  assign n5115 = n5114 ^ n5112 ;
  assign n5116 = n5115 ^ n5102 ;
  assign n5117 = x199 & n5116 ;
  assign n5118 = n5117 ^ n5115 ;
  assign n5140 = n5118 ^ n5071 ;
  assign n5119 = ~x203 & ~n5118 ;
  assign n5120 = x204 ^ x201 ;
  assign n5121 = n5120 ^ n5081 ;
  assign n5122 = n5121 ^ x204 ;
  assign n5124 = x200 & n5122 ;
  assign n5125 = n5124 ^ x204 ;
  assign n5129 = n5128 ^ n5081 ;
  assign n5130 = n5129 ^ n5074 ;
  assign n5133 = n5132 ^ x204 ;
  assign n5134 = ~n5130 & n5133 ;
  assign n5137 = n5134 ^ x201 ;
  assign n5138 = ~n5125 & ~n5137 ;
  assign n5139 = n5119 & n5138 ;
  assign n5141 = n5140 ^ n5139 ;
  assign n5142 = n5080 & n5141 ;
  assign n5143 = n5142 ^ n5079 ;
  assign n5144 = n5143 ^ n5112 ;
  assign n5148 = n5147 ^ n5144 ;
  assign n5297 = n5296 ^ n5148 ;
  assign n5216 = n5158 ^ n5153 ;
  assign n5217 = n5078 ^ n5073 ;
  assign n5218 = n5216 & n5217 ;
  assign n5563 = n5218 ^ n5159 ;
  assign n5564 = n5563 ^ n5079 ;
  assign n5565 = n5564 ^ n5141 ;
  assign n5566 = n5565 ^ n5213 ;
  assign n5221 = n5218 ^ n5079 ;
  assign n5225 = n5566 ^ n5221 ;
  assign n5230 = n5225 ^ n5079 ;
  assign n5234 = n5141 & n5230 ;
  assign n5222 = n5141 ^ n5079 ;
  assign n5223 = n5222 ^ n5221 ;
  assign n5224 = n5223 ^ n5159 ;
  assign n5227 = n5566 ^ n5223 ;
  assign n5226 = n5225 ^ n5159 ;
  assign n5228 = n5227 ^ n5226 ;
  assign n5229 = ~n5224 & n5228 ;
  assign n5235 = n5234 ^ n5229 ;
  assign n5236 = n5235 ^ n5227 ;
  assign n5237 = n5234 ^ n5225 ;
  assign n5238 = n5237 ^ n5227 ;
  assign n5239 = n5236 & ~n5238 ;
  assign n5240 = n5239 & n5566 ;
  assign n5241 = n5240 ^ n5234 ;
  assign n5242 = n5241 ^ n5141 ;
  assign n5214 = n5213 ^ n5159 ;
  assign n5243 = n5242 ^ n5214 ;
  assign n5244 = n5243 ^ n5079 ;
  assign n5248 = n5244 ^ n5214 ;
  assign n5298 = n5297 ^ n5248 ;
  assign n5302 = n5301 ^ n5298 ;
  assign n5249 = n5248 ^ n5143 ;
  assign n5250 = ~n5148 & ~n5249 ;
  assign n5251 = n5250 ^ n5248 ;
  assign n5591 = ~n5251 & n5296 ;
  assign n5592 = ~n5302 & n5591 ;
  assign n5307 = n5251 & ~n5301 ;
  assign n5308 = n5307 ^ n5302 ;
  assign n5309 = n5296 ^ n5251 ;
  assign n5310 = n5309 ^ n5302 ;
  assign n5311 = n5310 ^ n5251 ;
  assign n5312 = n5308 & ~n5311 ;
  assign n5313 = n5312 ^ n5309 ;
  assign n5314 = n5295 ^ n5291 ;
  assign n5315 = ~n5292 & ~n5314 ;
  assign n5316 = n5315 ^ n5291 ;
  assign n5590 = ~n5313 & n5316 ;
  assign n5593 = n5592 ^ n5590 ;
  assign n5594 = ~n5589 & n5593 ;
  assign n5596 = n5594 ^ n5589 ;
  assign n5597 = n5596 ^ n5593 ;
  assign n5560 = n5556 ^ n5419 ;
  assign n5317 = n5316 ^ n5313 ;
  assign n5561 = n5560 ^ n5317 ;
  assign n5562 = n5551 ^ n5302 ;
  assign n5573 = n5566 ^ n5537 ;
  assign n5576 = n5573 ^ n5302 ;
  assign n5567 = n5566 ^ n5534 ;
  assign n5568 = n5536 ^ n5535 ;
  assign n5569 = n5217 ^ n5216 ;
  assign n5570 = n5569 ^ n5536 ;
  assign n5571 = n5568 & ~n5570 ;
  assign n5572 = n5571 ^ n5535 ;
  assign n5574 = n5573 ^ n5572 ;
  assign n5575 = ~n5567 & n5574 ;
  assign n5577 = n5576 ^ n5575 ;
  assign n5578 = n5577 ^ n5302 ;
  assign n5579 = n5537 & ~n5575 ;
  assign n5580 = n5578 & n5579 ;
  assign n5581 = n5580 ^ n5577 ;
  assign n5582 = n5562 & ~n5581 ;
  assign n5583 = n5582 ^ n5551 ;
  assign n5584 = n5583 ^ n5317 ;
  assign n5585 = n5561 & n5584 ;
  assign n5586 = n5585 ^ n5560 ;
  assign n5598 = n5586 & ~n5594 ;
  assign n5599 = ~n5597 & ~n5598 ;
  assign n5601 = n5598 ^ n5597 ;
  assign n5602 = n5601 ^ n5599 ;
  assign n4865 = x233 & x234 ;
  assign n4864 = x231 & x232 ;
  assign n4866 = n4865 ^ n4864 ;
  assign n4942 = n4864 ^ x229 ;
  assign n4945 = n4942 ^ n4866 ;
  assign n4940 = n4864 ^ x230 ;
  assign n4950 = n4945 ^ n4940 ;
  assign n4854 = x232 ^ x231 ;
  assign n4867 = n4864 ^ n4854 ;
  assign n4851 = x234 ^ x233 ;
  assign n4868 = n4865 ^ n4851 ;
  assign n4869 = n4867 & n4868 ;
  assign n4870 = n4869 ^ n4865 ;
  assign n4941 = n4870 ^ n4866 ;
  assign n4943 = n4942 ^ n4941 ;
  assign n4951 = n4950 ^ n4943 ;
  assign n4952 = n4951 ^ n4866 ;
  assign n4954 = n4950 & n4952 ;
  assign n4947 = n4943 ^ n4866 ;
  assign n4948 = n4947 ^ n4865 ;
  assign n4949 = ~n4869 & n4948 ;
  assign n4955 = n4954 ^ n4949 ;
  assign n4956 = n4955 ^ n4947 ;
  assign n4957 = n4954 ^ n4945 ;
  assign n4958 = n4957 ^ n4947 ;
  assign n4959 = n4956 & n4958 ;
  assign n4960 = ~n4866 & n4959 ;
  assign n4961 = n4960 ^ n4954 ;
  assign n4962 = n4961 ^ n4952 ;
  assign n4970 = n4962 ^ n4864 ;
  assign n4973 = n4970 ^ n4940 ;
  assign n4884 = x227 & x228 ;
  assign n4883 = x225 & x226 ;
  assign n4885 = n4884 ^ n4883 ;
  assign n4908 = n4883 ^ x223 ;
  assign n4911 = n4908 ^ n4885 ;
  assign n4906 = n4883 ^ x224 ;
  assign n4916 = n4911 ^ n4906 ;
  assign n4859 = x226 ^ x225 ;
  assign n4886 = n4883 ^ n4859 ;
  assign n4857 = x228 ^ x227 ;
  assign n4887 = n4884 ^ n4857 ;
  assign n4888 = n4886 & n4887 ;
  assign n4889 = n4888 ^ n4884 ;
  assign n4907 = n4889 ^ n4885 ;
  assign n4909 = n4908 ^ n4907 ;
  assign n4917 = n4916 ^ n4909 ;
  assign n4918 = n4917 ^ n4885 ;
  assign n4920 = n4916 & n4918 ;
  assign n4913 = n4909 ^ n4885 ;
  assign n4914 = n4913 ^ n4884 ;
  assign n4915 = ~n4888 & n4914 ;
  assign n4921 = n4920 ^ n4915 ;
  assign n4922 = n4921 ^ n4913 ;
  assign n4923 = n4920 ^ n4911 ;
  assign n4924 = n4923 ^ n4913 ;
  assign n4925 = n4922 & n4924 ;
  assign n4926 = ~n4885 & n4925 ;
  assign n4927 = n4926 ^ n4920 ;
  assign n4928 = n4927 ^ n4918 ;
  assign n4936 = n4928 ^ n4883 ;
  assign n4939 = n4936 ^ n4906 ;
  assign n4974 = n4973 ^ n4939 ;
  assign n4890 = ~n4885 & ~n4889 ;
  assign n4862 = n4857 ^ x224 ;
  assign n4863 = n4862 ^ n4859 ;
  assign n4852 = x230 ^ x229 ;
  assign n4872 = n4851 ^ x230 ;
  assign n4873 = n4872 ^ n4854 ;
  assign n4874 = n4852 & ~n4873 ;
  assign n4875 = n4874 ^ x229 ;
  assign n4871 = ~n4866 & ~n4870 ;
  assign n4876 = n4875 ^ n4871 ;
  assign n4877 = n4876 ^ x223 ;
  assign n4878 = n4877 ^ n4857 ;
  assign n4879 = n4878 ^ n4859 ;
  assign n4880 = n4879 ^ n4876 ;
  assign n4881 = ~n4863 & n4880 ;
  assign n4882 = n4881 ^ n4877 ;
  assign n4891 = n4890 ^ n4882 ;
  assign n4853 = n4852 ^ n4851 ;
  assign n4855 = n4854 ^ n4853 ;
  assign n4856 = x224 ^ x223 ;
  assign n4858 = n4857 ^ n4856 ;
  assign n4860 = n4859 ^ n4858 ;
  assign n4861 = n4855 & n4860 ;
  assign n4975 = n4876 ^ n4861 ;
  assign n4976 = n4891 & ~n4975 ;
  assign n4977 = n4976 ^ n4876 ;
  assign n5024 = n4977 ^ n4973 ;
  assign n5025 = ~n4974 & ~n5024 ;
  assign n5026 = n5025 ^ n4977 ;
  assign n4978 = n4977 ^ n4974 ;
  assign n4781 = x245 & x246 ;
  assign n4782 = x243 & x244 ;
  assign n4783 = ~n4781 & ~n4782 ;
  assign n4786 = x244 ^ x243 ;
  assign n4787 = n4786 ^ n4782 ;
  assign n4784 = x246 ^ x245 ;
  assign n4785 = n4784 ^ n4781 ;
  assign n4789 = n4787 ^ n4785 ;
  assign n4788 = ~n4785 & ~n4787 ;
  assign n4790 = n4789 ^ n4788 ;
  assign n4791 = n4790 ^ n4783 ;
  assign n4793 = n4782 ^ n4781 ;
  assign n4794 = n4793 ^ n4783 ;
  assign n4795 = x241 & x242 ;
  assign n4796 = n4794 & n4795 ;
  assign n4792 = x242 ^ x241 ;
  assign n4797 = n4796 ^ n4792 ;
  assign n4798 = ~n4791 & ~n4797 ;
  assign n4799 = n4783 & n4798 ;
  assign n4828 = n4796 ^ n4790 ;
  assign n4829 = n4796 ^ n4783 ;
  assign n4830 = n4829 ^ n4798 ;
  assign n4831 = ~n4828 & n4830 ;
  assign n4832 = n4831 ^ n4790 ;
  assign n4833 = n4788 ^ x241 ;
  assign n4834 = n4833 ^ n4832 ;
  assign n4835 = n4794 ^ x242 ;
  assign n4836 = ~n4788 & ~n4835 ;
  assign n4837 = n4836 ^ x242 ;
  assign n4838 = n4834 & n4837 ;
  assign n4839 = n4838 ^ n4788 ;
  assign n4840 = n4832 & ~n4839 ;
  assign n4843 = n4799 & n4840 ;
  assign n4806 = x237 & x238 ;
  assign n4802 = x239 & x240 ;
  assign n4815 = n4806 ^ n4802 ;
  assign n4810 = ~n4802 & ~n4806 ;
  assign n4816 = n4815 ^ n4810 ;
  assign n4801 = x240 ^ x239 ;
  assign n4803 = n4802 ^ n4801 ;
  assign n4805 = x238 ^ x237 ;
  assign n4807 = n4806 ^ n4805 ;
  assign n4811 = n4803 & n4807 ;
  assign n4814 = n4811 ^ n4810 ;
  assign n4800 = x236 ^ x235 ;
  assign n4812 = n4811 ^ n4800 ;
  assign n4817 = x235 & x236 ;
  assign n4818 = n4816 & n4817 ;
  assign n4819 = n4818 ^ n4811 ;
  assign n4820 = ~n4812 & n4819 ;
  assign n4821 = n4814 & n4820 ;
  assign n4822 = n4821 ^ n4818 ;
  assign n4823 = n4816 & ~n4822 ;
  assign n4824 = n4823 ^ x235 ;
  assign n4825 = n4824 ^ n4822 ;
  assign n4813 = n4810 & ~n4812 ;
  assign n4826 = n4825 ^ n4813 ;
  assign n4804 = n4803 ^ x236 ;
  assign n4808 = n4807 ^ n4804 ;
  assign n4809 = n4800 & n4808 ;
  assign n4827 = n4826 ^ n4809 ;
  assign n4841 = n4840 ^ n4827 ;
  assign n4844 = n4843 ^ n4841 ;
  assign n4845 = n4792 ^ n4784 ;
  assign n4846 = n4845 ^ n4786 ;
  assign n4847 = n4801 ^ n4800 ;
  assign n4848 = n4847 ^ n4805 ;
  assign n4849 = n4846 & n4848 ;
  assign n4902 = n4849 ^ n4827 ;
  assign n4903 = ~n4844 & n4902 ;
  assign n4904 = n4903 ^ n4849 ;
  assign n4900 = n4794 & n4832 ;
  assign n4901 = n4900 ^ n4823 ;
  assign n4905 = n4904 ^ n4901 ;
  assign n4979 = n4978 ^ n4905 ;
  assign n4892 = n4891 ^ n4861 ;
  assign n4850 = n4849 ^ n4844 ;
  assign n4893 = n4892 ^ n4850 ;
  assign n4894 = n4860 ^ n4855 ;
  assign n4895 = n4848 ^ n4846 ;
  assign n4896 = n4894 & n4895 ;
  assign n4897 = n4896 ^ n4850 ;
  assign n4898 = n4893 & n4897 ;
  assign n4899 = n4898 ^ n4850 ;
  assign n4980 = n4979 ^ n4899 ;
  assign n5014 = ~n4904 & n4978 ;
  assign n5015 = n4980 & n5014 ;
  assign n5016 = n5015 ^ n4980 ;
  assign n5012 = ~n4823 & ~n4900 ;
  assign n5017 = ~n5012 & ~n5016 ;
  assign n5013 = n5012 ^ n4901 ;
  assign n5018 = n5017 ^ n5013 ;
  assign n5019 = n5017 ^ n4978 ;
  assign n5020 = ~n5018 & ~n5019 ;
  assign n5021 = n5020 ^ n4978 ;
  assign n5027 = n5021 ^ n5017 ;
  assign n5028 = n5027 ^ n5026 ;
  assign n5022 = ~n4899 & ~n4904 ;
  assign n5023 = ~n5021 & n5022 ;
  assign n5029 = n5028 ^ n5023 ;
  assign n5036 = ~n5012 & ~n5029 ;
  assign n5037 = ~n5016 & ~n5036 ;
  assign n5038 = n5026 & n5037 ;
  assign n5039 = n5038 ^ n5036 ;
  assign n4654 = x255 & x256 ;
  assign n4651 = x257 & x258 ;
  assign n4657 = n4654 ^ n4651 ;
  assign n4650 = x258 ^ x257 ;
  assign n4652 = n4651 ^ n4650 ;
  assign n4653 = x256 ^ x255 ;
  assign n4655 = n4654 ^ n4653 ;
  assign n4656 = n4652 & n4655 ;
  assign n4668 = x254 & n4656 ;
  assign n4669 = n4668 ^ n4654 ;
  assign n4670 = n4657 & ~n4669 ;
  assign n4671 = n4670 ^ n4651 ;
  assign n4672 = n4656 ^ x254 ;
  assign n4673 = n4672 ^ n4657 ;
  assign n4676 = ~n4656 & ~n4657 ;
  assign n4677 = ~n4673 & n4676 ;
  assign n4674 = n4673 ^ n4671 ;
  assign n4678 = n4677 ^ n4674 ;
  assign n4733 = x253 & ~n4678 ;
  assign n4734 = ~n4671 & n4733 ;
  assign n4687 = x249 & x250 ;
  assign n4684 = x251 & x252 ;
  assign n4690 = n4687 ^ n4684 ;
  assign n4683 = x252 ^ x251 ;
  assign n4685 = n4684 ^ n4683 ;
  assign n4686 = x250 ^ x249 ;
  assign n4688 = n4687 ^ n4686 ;
  assign n4689 = n4685 & n4688 ;
  assign n4698 = x248 & n4689 ;
  assign n4699 = n4698 ^ n4687 ;
  assign n4700 = n4690 & ~n4699 ;
  assign n4701 = n4700 ^ n4684 ;
  assign n4702 = n4689 ^ x248 ;
  assign n4703 = n4702 ^ n4690 ;
  assign n4706 = ~n4689 & ~n4690 ;
  assign n4707 = ~n4703 & n4706 ;
  assign n4704 = n4703 ^ n4701 ;
  assign n4708 = n4707 ^ n4704 ;
  assign n4728 = x247 & ~n4708 ;
  assign n4729 = ~n4701 & n4728 ;
  assign n4730 = n4729 ^ n4701 ;
  assign n4731 = n4730 ^ n4671 ;
  assign n4735 = n4734 ^ n4731 ;
  assign n4591 = x269 ^ x268 ;
  assign n4595 = x270 ^ x269 ;
  assign n4596 = ~n4591 & ~n4595 ;
  assign n4590 = x267 ^ x266 ;
  assign n4592 = n4591 ^ x267 ;
  assign n4593 = n4592 ^ x270 ;
  assign n4594 = ~n4590 & n4593 ;
  assign n4597 = n4596 ^ n4594 ;
  assign n4598 = ~x265 & n4597 ;
  assign n4599 = x268 ^ x267 ;
  assign n4600 = x268 ^ x266 ;
  assign n4601 = x270 ^ x265 ;
  assign n4604 = ~x268 & ~n4601 ;
  assign n4605 = n4604 ^ x265 ;
  assign n4606 = ~n4600 & n4605 ;
  assign n4607 = ~n4599 & n4606 ;
  assign n4608 = ~x269 & n4607 ;
  assign n4610 = ~x267 & ~x268 ;
  assign n4616 = ~x269 & ~x270 ;
  assign n4617 = ~n4610 & ~n4616 ;
  assign n4611 = n4610 ^ n4599 ;
  assign n4612 = x265 & x266 ;
  assign n4613 = x270 & n4612 ;
  assign n4614 = ~n4611 & n4613 ;
  assign n4615 = n4614 ^ n4612 ;
  assign n4618 = n4617 ^ n4615 ;
  assign n4621 = n4616 ^ n4595 ;
  assign n4624 = n4611 & n4621 ;
  assign n4625 = n4624 ^ n4615 ;
  assign n4626 = n4618 & ~n4625 ;
  assign n4609 = x266 ^ x265 ;
  assign n4627 = n4626 ^ n4615 ;
  assign n4628 = ~n4609 & n4627 ;
  assign n4629 = n4626 & n4628 ;
  assign n4630 = n4629 ^ n4627 ;
  assign n4631 = ~n4608 & ~n4630 ;
  assign n4632 = ~n4598 & n4631 ;
  assign n4544 = ~x263 & ~x264 ;
  assign n4546 = x259 & x260 ;
  assign n4545 = x260 ^ x259 ;
  assign n4547 = n4546 ^ n4545 ;
  assign n4548 = n4547 ^ x262 ;
  assign n4549 = n4547 ^ x261 ;
  assign n4550 = ~n4548 & ~n4549 ;
  assign n4551 = n4550 ^ n4547 ;
  assign n4552 = x264 ^ x263 ;
  assign n4553 = n4552 ^ n4544 ;
  assign n4554 = n4553 ^ n4548 ;
  assign n4555 = n4554 ^ n4549 ;
  assign n4557 = n4548 ^ n4546 ;
  assign n4558 = n4557 ^ n4549 ;
  assign n4559 = n4555 & n4558 ;
  assign n4560 = n4559 ^ n4547 ;
  assign n4561 = n4551 & n4560 ;
  assign n4562 = n4561 ^ n4547 ;
  assign n4563 = n4562 ^ n4546 ;
  assign n4564 = ~n4544 & n4563 ;
  assign n4565 = x262 ^ x261 ;
  assign n4566 = ~x259 & ~n4565 ;
  assign n4567 = x261 & x262 ;
  assign n4573 = ~n4546 & n4553 ;
  assign n4574 = n4567 & n4573 ;
  assign n4575 = n4574 ^ n4567 ;
  assign n4569 = ~x260 & n4544 ;
  assign n4570 = n4565 ^ n4545 ;
  assign n4571 = ~n4567 & n4570 ;
  assign n4572 = n4569 & n4571 ;
  assign n4576 = n4575 ^ n4572 ;
  assign n4568 = ~n4553 & n4567 ;
  assign n4577 = n4576 ^ n4568 ;
  assign n4578 = x263 ^ x262 ;
  assign n4581 = n4578 ^ x264 ;
  assign n4582 = ~x260 & n4581 ;
  assign n4583 = n4582 ^ n4578 ;
  assign n4584 = n4552 & ~n4583 ;
  assign n4585 = n4584 ^ n4578 ;
  assign n4586 = ~n4577 & ~n4585 ;
  assign n4587 = n4566 & n4586 ;
  assign n4588 = n4587 ^ n4577 ;
  assign n4589 = ~n4564 & ~n4588 ;
  assign n4633 = n4632 ^ n4589 ;
  assign n4635 = n4609 ^ n4599 ;
  assign n4636 = n4635 ^ n4595 ;
  assign n4634 = n4570 ^ n4552 ;
  assign n4738 = n4636 ^ n4634 ;
  assign n4712 = x248 ^ x247 ;
  assign n4722 = n4712 ^ n4686 ;
  assign n4723 = n4722 ^ n4683 ;
  assign n4661 = x254 ^ x253 ;
  assign n4720 = n4661 ^ n4653 ;
  assign n4721 = n4720 ^ n4650 ;
  assign n4739 = n4723 ^ n4721 ;
  assign n4740 = n4739 ^ n4636 ;
  assign n4741 = n4738 & ~n4740 ;
  assign n4742 = n4741 ^ n4634 ;
  assign n4724 = n4721 & n4723 ;
  assign n4982 = n4742 ^ n4724 ;
  assign n4693 = ~x247 & ~n4703 ;
  assign n4709 = n4708 ^ n4693 ;
  assign n4713 = n4686 ^ n4683 ;
  assign n4691 = n4690 ^ n4689 ;
  assign n4714 = n4713 ^ n4691 ;
  assign n4715 = n4714 ^ n4708 ;
  assign n4716 = n4715 ^ n4693 ;
  assign n4717 = n4712 & n4716 ;
  assign n4718 = n4709 & n4717 ;
  assign n4658 = n4657 ^ n4656 ;
  assign n4659 = n4658 ^ n4653 ;
  assign n4660 = n4659 ^ n4650 ;
  assign n4663 = ~x253 & ~n4673 ;
  assign n4679 = n4678 ^ n4663 ;
  assign n4680 = n4661 & n4679 ;
  assign n4681 = ~n4660 & n4680 ;
  assign n4682 = n4681 ^ n4679 ;
  assign n4710 = n4709 ^ n4682 ;
  assign n4719 = n4718 ^ n4710 ;
  assign n4983 = n4982 ^ n4719 ;
  assign n4637 = n4634 & n4636 ;
  assign n4750 = n4637 ^ n4633 ;
  assign n4751 = n4750 ^ n4742 ;
  assign n4767 = n4983 ^ n4751 ;
  assign n4768 = ~n4633 & n4767 ;
  assign n4758 = n4751 ^ n4724 ;
  assign n4984 = n4983 ^ n4633 ;
  assign n4761 = n4984 ^ n4751 ;
  assign n4746 = n4984 ^ n4742 ;
  assign n4760 = n4746 ^ n4724 ;
  assign n4762 = n4761 ^ n4760 ;
  assign n4763 = n4758 & ~n4762 ;
  assign n4769 = n4768 ^ n4763 ;
  assign n4770 = n4769 ^ n4761 ;
  assign n4771 = n4768 ^ n4746 ;
  assign n4772 = n4771 ^ n4761 ;
  assign n4773 = ~n4770 & n4772 ;
  assign n4774 = n4773 & n4984 ;
  assign n4775 = n4774 ^ n4768 ;
  assign n4776 = n4775 ^ n4633 ;
  assign n4777 = n4776 ^ n4637 ;
  assign n4725 = n4724 ^ n4682 ;
  assign n4726 = ~n4719 & n4725 ;
  assign n4727 = n4726 ^ n4724 ;
  assign n4736 = n4735 ^ n4727 ;
  assign n4998 = n4777 ^ n4736 ;
  assign n4638 = n4637 ^ n4589 ;
  assign n4639 = n4633 & ~n4638 ;
  assign n4640 = n4639 ^ n4632 ;
  assign n4999 = n4736 ^ n4640 ;
  assign n5000 = n4998 & ~n4999 ;
  assign n5001 = n5000 ^ n4777 ;
  assign n5002 = n5001 ^ n4730 ;
  assign n5003 = n5002 ^ n4727 ;
  assign n5004 = n5003 ^ n5001 ;
  assign n5005 = n4735 & n5004 ;
  assign n5006 = n5005 ^ n5002 ;
  assign n4647 = ~n4564 & ~n4575 ;
  assign n4641 = n4621 ^ n4611 ;
  assign n4642 = x266 & n4617 ;
  assign n4643 = n4642 ^ n4611 ;
  assign n4644 = n4641 & ~n4643 ;
  assign n4645 = n4644 ^ n4611 ;
  assign n4646 = ~n4630 & n4645 ;
  assign n4648 = n4647 ^ n4646 ;
  assign n4649 = n4648 ^ n4640 ;
  assign n4737 = n4736 ^ n4649 ;
  assign n4780 = n4777 ^ n4737 ;
  assign n5007 = n4780 ^ n4647 ;
  assign n5008 = n4648 & n5007 ;
  assign n5009 = n5008 ^ n4647 ;
  assign n5033 = n5009 ^ n5001 ;
  assign n5034 = ~n5006 & ~n5033 ;
  assign n5035 = n5034 ^ n5009 ;
  assign n5040 = n5039 ^ n5035 ;
  assign n5010 = n5009 ^ n5006 ;
  assign n4981 = n4980 ^ n4780 ;
  assign n4991 = n4984 ^ n4896 ;
  assign n4985 = n4895 ^ n4894 ;
  assign n4986 = n4739 ^ n4738 ;
  assign n4987 = n4986 ^ n4895 ;
  assign n4988 = n4985 & ~n4987 ;
  assign n4989 = n4988 ^ n4894 ;
  assign n4992 = n4991 ^ n4989 ;
  assign n4993 = n4893 & n4992 ;
  assign n4990 = n4984 & n4989 ;
  assign n4994 = n4993 ^ n4990 ;
  assign n4995 = n4994 ^ n4780 ;
  assign n4996 = ~n4981 & ~n4995 ;
  assign n4997 = n4996 ^ n4980 ;
  assign n5011 = n5010 ^ n4997 ;
  assign n5030 = n5029 ^ n4997 ;
  assign n5031 = ~n5011 & n5030 ;
  assign n5032 = n5031 ^ n5029 ;
  assign n5041 = n5040 ^ n5032 ;
  assign n5667 = n5602 ^ n5041 ;
  assign n5668 = ~n5599 & ~n5667 ;
  assign n5609 = n5583 ^ n5561 ;
  assign n5608 = n5029 ^ n5011 ;
  assign n5610 = n5609 ^ n5608 ;
  assign n5612 = n5581 ^ n5551 ;
  assign n5611 = n4994 ^ n4981 ;
  assign n5613 = n5612 ^ n5611 ;
  assign n5616 = n5572 ^ n5534 ;
  assign n5617 = n5616 ^ n5566 ;
  assign n5614 = n4984 ^ n4893 ;
  assign n5615 = n5614 ^ n4989 ;
  assign n5618 = n5617 ^ n5615 ;
  assign n5619 = n4986 ^ n4985 ;
  assign n5620 = n5569 ^ n5568 ;
  assign n5621 = n5619 & n5620 ;
  assign n5622 = n5621 ^ n5615 ;
  assign n5623 = ~n5618 & ~n5622 ;
  assign n5624 = n5623 ^ n5617 ;
  assign n5625 = n5624 ^ n5612 ;
  assign n5626 = ~n5613 & ~n5625 ;
  assign n5627 = n5626 ^ n5612 ;
  assign n5628 = n5627 ^ n5608 ;
  assign n5629 = ~n5610 & n5628 ;
  assign n5630 = n5629 ^ n5609 ;
  assign n5669 = n5630 ^ n5602 ;
  assign n5670 = n5668 & n5669 ;
  assign n5671 = n5670 ^ n5602 ;
  assign n5604 = n5035 ^ n5032 ;
  assign n5605 = n5040 & ~n5604 ;
  assign n5606 = n5605 ^ n5039 ;
  assign n5595 = n5594 ^ n5586 ;
  assign n5600 = n5599 ^ n5595 ;
  assign n5603 = n5602 ^ n5600 ;
  assign n5607 = ~n5603 & n5606 ;
  assign n5631 = n5607 & n5630 ;
  assign n5632 = ~n5041 & n5631 ;
  assign n5633 = n5632 ^ n5607 ;
  assign n5634 = n5633 ^ n5603 ;
  assign n5635 = n5634 ^ n5586 ;
  assign n5657 = n5593 ^ n5589 ;
  assign n5658 = n5657 ^ n5586 ;
  assign n5659 = n5658 ^ n5041 ;
  assign n5660 = n5659 ^ n5630 ;
  assign n5661 = ~n5594 & ~n5660 ;
  assign n5636 = ~n5039 & n5594 ;
  assign n5637 = n5636 ^ n5589 ;
  assign n5649 = ~n5035 & ~n5039 ;
  assign n5650 = n5637 & n5649 ;
  assign n5651 = n5650 ^ n5637 ;
  assign n5639 = ~n5035 & n5592 ;
  assign n5640 = ~n5637 & n5639 ;
  assign n5641 = n5640 ^ n5636 ;
  assign n5642 = n5641 ^ n5594 ;
  assign n5643 = n5642 ^ n5637 ;
  assign n5652 = n5651 ^ n5643 ;
  assign n5653 = ~n5032 & n5652 ;
  assign n5654 = n5653 ^ n5641 ;
  assign n5662 = n5661 ^ n5654 ;
  assign n5663 = ~n5634 & n5662 ;
  assign n5664 = n5663 ^ n5654 ;
  assign n5665 = n5635 & n5664 ;
  assign n5666 = n5665 ^ n5634 ;
  assign n5719 = n5606 & n5666 ;
  assign n5720 = n5671 & n5719 ;
  assign n5721 = n5720 ^ n5671 ;
  assign n5672 = n5671 ^ n5606 ;
  assign n5673 = n5672 ^ n5671 ;
  assign n5674 = n5602 & n5630 ;
  assign n5675 = n5674 ^ n5671 ;
  assign n5676 = ~n5673 & ~n5675 ;
  assign n5677 = n5676 ^ n5671 ;
  assign n5678 = n5666 & ~n5677 ;
  assign n5679 = n5678 ^ n5666 ;
  assign n4026 = ~x83 & ~x84 ;
  assign n3920 = x82 ^ x81 ;
  assign n3919 = x84 ^ x83 ;
  assign n4027 = n4026 ^ n3919 ;
  assign n4028 = n4027 ^ x82 ;
  assign n4029 = n3920 & n4028 ;
  assign n4030 = n4029 ^ x81 ;
  assign n4032 = ~n4026 & n4030 ;
  assign n4031 = n4030 ^ n4026 ;
  assign n4033 = n4032 ^ n4031 ;
  assign n4045 = n4029 ^ n4028 ;
  assign n4053 = ~n4033 & ~n4045 ;
  assign n4054 = n4053 ^ n4032 ;
  assign n4055 = x80 & n4054 ;
  assign n4056 = n4055 ^ n4032 ;
  assign n4035 = x81 & x82 ;
  assign n4039 = ~n4027 & n4035 ;
  assign n4040 = x80 & ~n4026 ;
  assign n4041 = n4030 & ~n4040 ;
  assign n4042 = ~n4039 & n4041 ;
  assign n4043 = n4042 ^ n4030 ;
  assign n4101 = x79 & ~n4043 ;
  assign n4102 = n4056 & n4101 ;
  assign n4103 = n4102 ^ n4043 ;
  assign n4062 = ~x87 & ~x88 ;
  assign n3924 = x88 ^ x87 ;
  assign n4068 = n4062 ^ n3924 ;
  assign n4061 = ~x89 & ~x90 ;
  assign n4066 = ~n4061 & ~n4062 ;
  assign n4063 = x85 & x86 ;
  assign n4067 = n4066 ^ n4063 ;
  assign n4069 = n4068 ^ n4067 ;
  assign n3926 = x90 ^ x89 ;
  assign n4070 = n4061 ^ n3926 ;
  assign n4071 = n4070 ^ n4068 ;
  assign n4072 = n4071 ^ n4063 ;
  assign n3923 = x86 ^ x85 ;
  assign n4073 = n4072 ^ n3923 ;
  assign n4074 = ~n4066 & n4073 ;
  assign n4075 = n4074 ^ n4073 ;
  assign n4076 = ~n4069 & n4075 ;
  assign n4077 = n4076 ^ n4067 ;
  assign n4078 = n4074 ^ n3923 ;
  assign n4079 = n4078 ^ n4076 ;
  assign n4080 = n4077 & n4079 ;
  assign n4081 = n4080 ^ n4063 ;
  assign n4064 = n4062 & ~n4063 ;
  assign n4065 = n4061 & n4064 ;
  assign n4082 = n4081 ^ n4065 ;
  assign n4085 = ~n4068 & ~n4070 ;
  assign n4086 = n4085 ^ n4071 ;
  assign n4087 = ~x86 & ~n4066 ;
  assign n4088 = ~n4086 & n4087 ;
  assign n4089 = n4088 ^ n4085 ;
  assign n4090 = ~x85 & n4089 ;
  assign n4091 = ~n4082 & n4090 ;
  assign n4034 = ~x80 & n4033 ;
  assign n4036 = n4035 ^ n3920 ;
  assign n4037 = n4034 & ~n4036 ;
  assign n4046 = n4045 ^ n4039 ;
  assign n4047 = ~n4040 & n4046 ;
  assign n4038 = n4037 ^ n4034 ;
  assign n4044 = n4043 ^ n4038 ;
  assign n4048 = n4047 ^ n4044 ;
  assign n4057 = n4056 ^ n4048 ;
  assign n4058 = x79 & n4057 ;
  assign n4059 = n4058 ^ n4048 ;
  assign n4060 = ~n4037 & ~n4059 ;
  assign n4083 = n4082 ^ n4060 ;
  assign n4092 = n4091 ^ n4083 ;
  assign n3921 = n3920 ^ n3919 ;
  assign n3918 = x80 ^ x79 ;
  assign n3922 = n3921 ^ n3918 ;
  assign n3925 = n3924 ^ n3923 ;
  assign n3927 = n3926 ^ n3925 ;
  assign n4022 = n3922 & n3927 ;
  assign n4106 = n4060 ^ n4022 ;
  assign n4107 = n4092 & n4106 ;
  assign n4108 = n4107 ^ n4022 ;
  assign n4384 = ~n4103 & ~n4108 ;
  assign n3910 = x102 ^ x101 ;
  assign n3908 = x98 ^ x97 ;
  assign n3907 = x100 ^ x99 ;
  assign n3909 = n3908 ^ n3907 ;
  assign n3911 = n3910 ^ n3909 ;
  assign n3915 = x96 ^ x95 ;
  assign n3913 = x92 ^ x91 ;
  assign n3912 = x94 ^ x93 ;
  assign n3914 = n3913 ^ n3912 ;
  assign n3916 = n3915 ^ n3914 ;
  assign n4021 = n3911 & n3916 ;
  assign n4023 = n4021 & n4022 ;
  assign n3977 = x95 & x96 ;
  assign n3978 = n3977 ^ n3915 ;
  assign n3979 = x91 & x92 ;
  assign n3980 = n3979 ^ n3913 ;
  assign n3981 = n3980 ^ x94 ;
  assign n3982 = n3980 ^ x93 ;
  assign n3983 = ~n3981 & ~n3982 ;
  assign n3984 = n3983 ^ n3980 ;
  assign n3985 = n3981 ^ n3977 ;
  assign n3986 = n3985 ^ n3982 ;
  assign n3988 = n3981 ^ n3979 ;
  assign n3989 = n3988 ^ n3982 ;
  assign n3990 = ~n3986 & n3989 ;
  assign n3991 = n3990 ^ n3980 ;
  assign n3992 = n3984 & n3991 ;
  assign n3993 = n3992 ^ n3980 ;
  assign n3994 = n3993 ^ n3979 ;
  assign n3995 = n3978 & n3994 ;
  assign n3996 = ~x91 & ~n3912 ;
  assign n3998 = x93 & x94 ;
  assign n4005 = n3977 & n3998 ;
  assign n4001 = ~n3977 & ~n3979 ;
  assign n4002 = n3998 & n4001 ;
  assign n4003 = n4002 ^ n3998 ;
  assign n3997 = ~x92 & ~n3978 ;
  assign n3999 = n3914 & ~n3998 ;
  assign n4000 = n3997 & n3999 ;
  assign n4004 = n4003 ^ n4000 ;
  assign n4006 = n4005 ^ n4004 ;
  assign n4007 = x95 ^ x94 ;
  assign n4010 = n4007 ^ x96 ;
  assign n4011 = ~x92 & n4010 ;
  assign n4012 = n4011 ^ n4007 ;
  assign n4013 = n3915 & ~n4012 ;
  assign n4014 = n4013 ^ n4007 ;
  assign n4015 = ~n4006 & ~n4014 ;
  assign n4016 = n3996 & n4015 ;
  assign n4017 = n4016 ^ n4006 ;
  assign n4018 = ~n3995 & ~n4017 ;
  assign n3935 = x101 & x102 ;
  assign n3936 = n3935 ^ n3910 ;
  assign n3937 = x97 & x98 ;
  assign n3938 = n3937 ^ n3908 ;
  assign n3939 = n3938 ^ x100 ;
  assign n3940 = n3938 ^ x99 ;
  assign n3941 = ~n3939 & ~n3940 ;
  assign n3942 = n3941 ^ n3938 ;
  assign n3943 = n3939 ^ n3935 ;
  assign n3944 = n3943 ^ n3940 ;
  assign n3946 = n3939 ^ n3937 ;
  assign n3947 = n3946 ^ n3940 ;
  assign n3948 = ~n3944 & n3947 ;
  assign n3949 = n3948 ^ n3938 ;
  assign n3950 = n3942 & n3949 ;
  assign n3951 = n3950 ^ n3938 ;
  assign n3952 = n3951 ^ n3937 ;
  assign n3953 = n3936 & n3952 ;
  assign n3954 = ~x97 & ~n3907 ;
  assign n3956 = x99 & x100 ;
  assign n3963 = n3935 & n3956 ;
  assign n3959 = ~n3935 & ~n3937 ;
  assign n3960 = n3956 & n3959 ;
  assign n3961 = n3960 ^ n3956 ;
  assign n3955 = ~x98 & ~n3936 ;
  assign n3957 = n3909 & ~n3956 ;
  assign n3958 = n3955 & n3957 ;
  assign n3962 = n3961 ^ n3958 ;
  assign n3964 = n3963 ^ n3962 ;
  assign n3965 = x101 ^ x100 ;
  assign n3968 = n3965 ^ x102 ;
  assign n3969 = ~x98 & n3968 ;
  assign n3970 = n3969 ^ n3965 ;
  assign n3971 = n3910 & ~n3970 ;
  assign n3972 = n3971 ^ n3965 ;
  assign n3973 = ~n3964 & ~n3972 ;
  assign n3974 = n3954 & n3973 ;
  assign n3975 = n3974 ^ n3964 ;
  assign n3976 = ~n3953 & ~n3975 ;
  assign n4019 = n4018 ^ n3976 ;
  assign n3917 = n3916 ^ n3911 ;
  assign n3928 = n3927 ^ n3922 ;
  assign n3929 = n3928 ^ n3911 ;
  assign n3930 = ~n3917 & n3929 ;
  assign n3931 = n3930 ^ n3928 ;
  assign n3932 = n3922 & ~n3931 ;
  assign n3933 = ~n3930 & n3932 ;
  assign n3934 = n3933 ^ n3931 ;
  assign n4020 = n4019 ^ n3934 ;
  assign n4024 = n4023 ^ n4020 ;
  assign n4025 = n4024 ^ n4022 ;
  assign n4093 = n4025 & n4092 ;
  assign n4094 = n4093 ^ n4022 ;
  assign n4095 = n4021 ^ n3934 ;
  assign n4098 = ~n4019 & ~n4095 ;
  assign n4099 = n4098 ^ n4021 ;
  assign n4100 = ~n4094 & ~n4099 ;
  assign n4104 = ~n4081 & ~n4085 ;
  assign n4383 = ~n4100 & n4104 ;
  assign n4385 = n4384 ^ n4383 ;
  assign n4105 = n4104 ^ n4103 ;
  assign n4109 = n4108 ^ n4105 ;
  assign n4110 = n4109 ^ n4100 ;
  assign n4115 = ~n3995 & ~n4003 ;
  assign n4114 = ~n3953 & ~n3961 ;
  assign n4116 = n4115 ^ n4114 ;
  assign n4111 = n4021 ^ n4018 ;
  assign n4112 = n4019 & n4111 ;
  assign n4113 = n4112 ^ n4018 ;
  assign n4117 = n4116 ^ n4113 ;
  assign n4386 = ~n4110 & ~n4117 ;
  assign n4387 = n4386 ^ n4383 ;
  assign n4388 = n4385 & ~n4387 ;
  assign n4389 = n4388 ^ n4384 ;
  assign n4380 = n4115 ^ n4113 ;
  assign n4381 = n4116 & ~n4380 ;
  assign n4382 = n4381 ^ n4115 ;
  assign n4390 = ~n4383 & ~n4384 ;
  assign n4391 = n4386 ^ n4110 ;
  assign n4392 = n4390 & ~n4391 ;
  assign n4467 = n4382 & ~n4392 ;
  assign n4473 = ~n4389 & n4467 ;
  assign n4300 = x119 & x120 ;
  assign n4299 = x117 & x118 ;
  assign n4301 = n4300 ^ n4299 ;
  assign n4343 = n4299 ^ x115 ;
  assign n4346 = n4343 ^ n4301 ;
  assign n4341 = n4299 ^ x116 ;
  assign n4351 = n4346 ^ n4341 ;
  assign n4137 = x118 ^ x117 ;
  assign n4302 = n4299 ^ n4137 ;
  assign n4135 = x120 ^ x119 ;
  assign n4303 = n4300 ^ n4135 ;
  assign n4304 = n4302 & n4303 ;
  assign n4305 = n4304 ^ n4300 ;
  assign n4342 = n4305 ^ n4301 ;
  assign n4344 = n4343 ^ n4342 ;
  assign n4352 = n4351 ^ n4344 ;
  assign n4353 = n4352 ^ n4301 ;
  assign n4355 = n4351 & n4353 ;
  assign n4348 = n4344 ^ n4301 ;
  assign n4349 = n4348 ^ n4300 ;
  assign n4350 = ~n4304 & n4349 ;
  assign n4356 = n4355 ^ n4350 ;
  assign n4357 = n4356 ^ n4348 ;
  assign n4358 = n4355 ^ n4346 ;
  assign n4359 = n4358 ^ n4348 ;
  assign n4360 = n4357 & n4359 ;
  assign n4361 = ~n4301 & n4360 ;
  assign n4362 = n4361 ^ n4355 ;
  assign n4363 = n4362 ^ n4353 ;
  assign n4371 = n4363 ^ n4299 ;
  assign n4374 = n4371 ^ n4341 ;
  assign n4266 = x121 & x122 ;
  assign n4258 = x123 & x124 ;
  assign n4259 = x125 & x126 ;
  assign n4267 = n4258 & ~n4259 ;
  assign n4268 = ~n4266 & n4267 ;
  assign n4269 = n4268 ^ n4258 ;
  assign n4130 = x126 ^ x125 ;
  assign n4260 = n4259 ^ n4130 ;
  assign n4131 = x122 ^ x121 ;
  assign n4271 = n4266 ^ n4131 ;
  assign n4272 = n4271 ^ x124 ;
  assign n4273 = n4271 ^ x123 ;
  assign n4274 = ~n4272 & ~n4273 ;
  assign n4275 = n4274 ^ n4271 ;
  assign n4276 = n4266 ^ n4259 ;
  assign n4277 = n4272 ^ n4266 ;
  assign n4278 = n4277 ^ n4273 ;
  assign n4279 = n4276 & n4278 ;
  assign n4280 = n4279 ^ n4271 ;
  assign n4281 = n4275 & n4280 ;
  assign n4282 = n4281 ^ n4271 ;
  assign n4283 = n4282 ^ n4266 ;
  assign n4284 = n4260 & n4283 ;
  assign n4340 = ~n4269 & ~n4284 ;
  assign n4375 = n4374 ^ n4340 ;
  assign n4136 = x116 ^ x115 ;
  assign n4307 = n4137 ^ x116 ;
  assign n4308 = n4307 ^ n4135 ;
  assign n4309 = n4136 & ~n4308 ;
  assign n4310 = n4309 ^ x115 ;
  assign n4306 = ~n4301 & ~n4305 ;
  assign n4311 = n4310 ^ n4306 ;
  assign n4286 = n4284 ^ x121 ;
  assign n4297 = n4286 ^ n4259 ;
  assign n4133 = x124 ^ x123 ;
  assign n4132 = n4131 ^ n4130 ;
  assign n4134 = n4133 ^ n4132 ;
  assign n4285 = n4284 ^ n4134 ;
  assign n4287 = n4286 ^ n4285 ;
  assign n4294 = ~n4284 & n4286 ;
  assign n4288 = n4258 ^ n4133 ;
  assign n4289 = ~n4259 & ~n4288 ;
  assign n4295 = n4294 ^ n4289 ;
  assign n4296 = n4287 & ~n4295 ;
  assign n4298 = n4297 ^ n4296 ;
  assign n4312 = n4311 ^ n4298 ;
  assign n4270 = n4134 & ~n4269 ;
  assign n4313 = n4312 ^ n4270 ;
  assign n4263 = x122 & ~n4260 ;
  assign n4264 = n4263 ^ n4130 ;
  assign n4265 = ~n4258 & ~n4264 ;
  assign n4314 = n4313 ^ n4265 ;
  assign n4138 = n4137 ^ n4136 ;
  assign n4139 = n4138 ^ n4135 ;
  assign n4140 = n4134 & n4139 ;
  assign n4337 = n4311 ^ n4140 ;
  assign n4338 = ~n4314 & ~n4337 ;
  assign n4339 = n4338 ^ n4140 ;
  assign n4376 = n4375 ^ n4339 ;
  assign n4120 = x112 ^ x111 ;
  assign n4119 = x114 ^ x113 ;
  assign n4121 = n4120 ^ n4119 ;
  assign n4145 = ~x111 & ~x112 ;
  assign n4146 = n4145 ^ n4120 ;
  assign n4147 = ~x113 & ~x114 ;
  assign n4148 = n4147 ^ n4119 ;
  assign n4149 = n4146 & n4148 ;
  assign n4150 = n4149 ^ x110 ;
  assign n4151 = ~n4121 & ~n4150 ;
  assign n4152 = n4151 ^ x110 ;
  assign n4153 = ~n4145 & ~n4147 ;
  assign n4156 = n4153 ^ n4149 ;
  assign n4157 = x109 & x110 ;
  assign n4158 = x114 & ~n4146 ;
  assign n4159 = n4157 & n4158 ;
  assign n4160 = n4159 ^ n4157 ;
  assign n4161 = n4160 ^ n4149 ;
  assign n4162 = n4156 & ~n4161 ;
  assign n4122 = x110 ^ x109 ;
  assign n4163 = n4162 ^ n4160 ;
  assign n4164 = ~n4122 & n4163 ;
  assign n4165 = n4162 & n4164 ;
  assign n4166 = n4165 ^ n4163 ;
  assign n4333 = n4153 & ~n4166 ;
  assign n4334 = n4152 & n4333 ;
  assign n4335 = n4334 ^ n4166 ;
  assign n4411 = n4376 ^ n4335 ;
  assign n4126 = x106 ^ x105 ;
  assign n4125 = x108 ^ x107 ;
  assign n4127 = n4126 ^ n4125 ;
  assign n4124 = x104 ^ x103 ;
  assign n4128 = n4127 ^ n4124 ;
  assign n4123 = n4122 ^ n4121 ;
  assign n4129 = n4128 ^ n4123 ;
  assign n4142 = n4139 ^ n4134 ;
  assign n4141 = n4140 ^ n4123 ;
  assign n4143 = n4142 ^ n4141 ;
  assign n4144 = n4143 ^ n4123 ;
  assign n4178 = x106 ^ x104 ;
  assign n4179 = x108 ^ x103 ;
  assign n4182 = ~x106 & ~n4179 ;
  assign n4183 = n4182 ^ x103 ;
  assign n4184 = ~n4178 & n4183 ;
  assign n4185 = ~n4126 & n4184 ;
  assign n4186 = ~x107 & n4185 ;
  assign n4187 = ~x105 & ~x106 ;
  assign n4188 = n4187 ^ n4126 ;
  assign n4189 = n4188 ^ n4125 ;
  assign n4230 = n4126 ^ x108 ;
  assign n4235 = n4125 & n4230 ;
  assign n4236 = ~n4189 & n4235 ;
  assign n4231 = n4230 ^ n4187 ;
  assign n4190 = ~x107 & ~x108 ;
  assign n4225 = n4190 ^ n4188 ;
  assign n4226 = n4225 ^ x103 ;
  assign n4204 = n4187 ^ n4125 ;
  assign n4201 = n4190 ^ n4125 ;
  assign n4202 = n4187 & n4201 ;
  assign n4203 = n4202 ^ n4190 ;
  assign n4205 = n4204 ^ n4203 ;
  assign n4217 = n4190 ^ x104 ;
  assign n4227 = n4205 & ~n4217 ;
  assign n4228 = ~n4226 & n4227 ;
  assign n4229 = n4228 ^ n4190 ;
  assign n4232 = n4231 ^ n4229 ;
  assign n4237 = n4236 ^ n4232 ;
  assign n4238 = x104 & n4237 ;
  assign n4239 = n4238 ^ n4229 ;
  assign n4199 = x104 & n4190 ;
  assign n4191 = n4190 ^ n4189 ;
  assign n4192 = n4191 ^ x104 ;
  assign n4194 = n4201 ^ n4192 ;
  assign n4200 = n4199 ^ n4194 ;
  assign n4206 = n4205 ^ n4191 ;
  assign n4207 = n4199 ^ x104 ;
  assign n4208 = ~n4206 & n4207 ;
  assign n4209 = n4208 ^ n4191 ;
  assign n4210 = ~n4200 & n4209 ;
  assign n4212 = n4210 ^ n4188 ;
  assign n4220 = n4188 & n4217 ;
  assign n4221 = n4203 & n4220 ;
  assign n4222 = n4221 ^ n4203 ;
  assign n4223 = n4222 ^ n4190 ;
  assign n4224 = n4212 & ~n4223 ;
  assign n4240 = n4239 ^ n4224 ;
  assign n4241 = ~x103 & n4240 ;
  assign n4242 = n4241 ^ n4239 ;
  assign n4243 = ~n4186 & n4242 ;
  assign n4154 = n4153 ^ n4152 ;
  assign n4155 = ~x109 & ~n4154 ;
  assign n4167 = x112 ^ x110 ;
  assign n4168 = x114 ^ x109 ;
  assign n4171 = ~x112 & ~n4168 ;
  assign n4172 = n4171 ^ x109 ;
  assign n4173 = ~n4167 & n4172 ;
  assign n4174 = ~n4120 & n4173 ;
  assign n4175 = ~x113 & n4174 ;
  assign n4176 = ~n4166 & ~n4175 ;
  assign n4177 = ~n4155 & n4176 ;
  assign n4244 = n4243 ^ n4177 ;
  assign n4247 = n4144 & ~n4244 ;
  assign n4248 = n4247 ^ n4123 ;
  assign n4249 = n4129 & n4248 ;
  assign n4245 = n4244 ^ n4123 ;
  assign n4250 = n4249 ^ n4245 ;
  assign n4251 = n4139 ^ n4128 ;
  assign n4254 = ~n4129 & ~n4251 ;
  assign n4252 = n4251 ^ n4123 ;
  assign n4253 = ~n4134 & n4252 ;
  assign n4255 = n4254 ^ n4253 ;
  assign n4256 = n4255 ^ n4244 ;
  assign n4257 = n4256 ^ n4140 ;
  assign n4317 = ~n4257 & n4314 ;
  assign n4318 = n4317 ^ n4256 ;
  assign n4319 = n4250 & n4318 ;
  assign n4412 = n4376 ^ n4319 ;
  assign n4415 = ~n4411 & ~n4412 ;
  assign n4416 = n4415 ^ n4376 ;
  assign n4425 = n4412 ^ n4411 ;
  assign n4426 = n4425 ^ n4376 ;
  assign n4329 = n4123 & n4128 ;
  assign n4330 = n4329 ^ n4177 ;
  assign n4331 = n4244 & n4330 ;
  assign n4320 = x103 & ~n4239 ;
  assign n4321 = n4212 & n4320 ;
  assign n4322 = n4321 ^ n4212 ;
  assign n4323 = n4322 ^ n4177 ;
  assign n4332 = n4331 ^ n4323 ;
  assign n4417 = n4322 ^ n4319 ;
  assign n4422 = n4417 ^ n4335 ;
  assign n4423 = n4422 ^ n4376 ;
  assign n4424 = n4332 & n4423 ;
  assign n4427 = n4426 ^ n4424 ;
  assign n4428 = n4416 & n4427 ;
  assign n4408 = n4374 ^ n4339 ;
  assign n4409 = ~n4375 & n4408 ;
  assign n4410 = n4409 ^ n4374 ;
  assign n4336 = n4335 ^ n4332 ;
  assign n4377 = n4376 ^ n4336 ;
  assign n4378 = n4377 ^ n4319 ;
  assign n4435 = n4332 & ~n4417 ;
  assign n4436 = n4435 ^ n4319 ;
  assign n4437 = ~n4376 & n4436 ;
  assign n4438 = ~n4378 & n4437 ;
  assign n4468 = ~n4410 & ~n4438 ;
  assign n4469 = ~n4428 & n4468 ;
  assign n4470 = n4469 ^ n4428 ;
  assign n4471 = n4470 ^ n4389 ;
  assign n4474 = n4473 ^ n4471 ;
  assign n4118 = n4117 ^ n4110 ;
  assign n4379 = n4378 ^ n4118 ;
  assign n4397 = n4092 ^ n4024 ;
  assign n4315 = n4314 ^ n4256 ;
  assign n4398 = n4397 ^ n4315 ;
  assign n4399 = n4142 ^ n4129 ;
  assign n4400 = n3928 ^ n3917 ;
  assign n4401 = n4399 & n4400 ;
  assign n4402 = n4401 ^ n4397 ;
  assign n4403 = n4398 & n4402 ;
  assign n4404 = n4403 ^ n4315 ;
  assign n4405 = n4404 ^ n4378 ;
  assign n4406 = ~n4379 & ~n4405 ;
  assign n4393 = n4392 ^ n4389 ;
  assign n4394 = n4393 ^ n4382 ;
  assign n4395 = n4394 ^ n4378 ;
  assign n4407 = n4406 ^ n4395 ;
  assign n4439 = n4438 ^ n4428 ;
  assign n4440 = n4439 ^ n4410 ;
  assign n4464 = n4440 ^ n4394 ;
  assign n4465 = ~n4407 & ~n4464 ;
  assign n4466 = n4465 ^ n4440 ;
  assign n4536 = n4470 ^ n4466 ;
  assign n4537 = n4474 & n4536 ;
  assign n4538 = n4537 ^ n4470 ;
  assign n3678 = x161 & x162 ;
  assign n3675 = x162 ^ x161 ;
  assign n3689 = n3678 ^ n3675 ;
  assign n3676 = ~x159 & ~x160 ;
  assign n3665 = x160 ^ x159 ;
  assign n3677 = n3676 ^ n3665 ;
  assign n3719 = n3689 ^ n3677 ;
  assign n3683 = ~x158 & n3689 ;
  assign n3684 = n3719 ^ n3683 ;
  assign n3712 = n3676 ^ x162 ;
  assign n3690 = n3676 & ~n3678 ;
  assign n3691 = n3690 ^ n3689 ;
  assign n3692 = n3691 ^ x161 ;
  assign n3693 = n3712 ^ n3692 ;
  assign n3685 = n3683 ^ n3675 ;
  assign n3694 = n3693 ^ n3685 ;
  assign n3697 = ~n3677 & ~n3694 ;
  assign n3698 = n3697 ^ n3693 ;
  assign n3699 = ~n3684 & n3698 ;
  assign n3700 = n3699 ^ n3677 ;
  assign n3720 = n3719 ^ x157 ;
  assign n3721 = ~n3693 & n3720 ;
  assign n3715 = n3676 ^ x161 ;
  assign n3716 = n3677 & n3715 ;
  assign n3717 = ~n3712 & n3716 ;
  assign n3713 = n3712 ^ n3665 ;
  assign n3718 = n3717 ^ n3713 ;
  assign n3722 = n3718 ^ n3689 ;
  assign n3723 = n3722 ^ x158 ;
  assign n3724 = n3723 ^ n3718 ;
  assign n3725 = n3721 & n3724 ;
  assign n3726 = n3725 ^ n3722 ;
  assign n3727 = ~x158 & ~n3726 ;
  assign n3728 = n3727 ^ n3718 ;
  assign n3845 = x157 & ~n3728 ;
  assign n3846 = n3700 & n3845 ;
  assign n3608 = x153 & x154 ;
  assign n3607 = x154 ^ x153 ;
  assign n3609 = n3608 ^ n3607 ;
  assign n3610 = x156 ^ x155 ;
  assign n3605 = ~x155 & ~x156 ;
  assign n3611 = n3610 ^ n3605 ;
  assign n3614 = n3611 ^ n3608 ;
  assign n3606 = x152 & ~n3605 ;
  assign n3615 = n3608 ^ n3606 ;
  assign n3616 = ~n3614 & n3615 ;
  assign n3617 = n3616 ^ n3608 ;
  assign n3618 = n3609 & n3617 ;
  assign n3630 = x156 ^ x152 ;
  assign n3652 = x156 ^ x154 ;
  assign n3631 = ~n3630 & ~n3652 ;
  assign n3632 = n3631 ^ x153 ;
  assign n3623 = x155 ^ x153 ;
  assign n3635 = n3632 ^ n3623 ;
  assign n3636 = ~n3631 & n3635 ;
  assign n3637 = n3636 ^ n3632 ;
  assign n3656 = n3630 ^ n3607 ;
  assign n3638 = n3637 & ~n3656 ;
  assign n3639 = n3638 ^ n3632 ;
  assign n3840 = x151 & n3639 ;
  assign n3841 = ~n3618 & n3840 ;
  assign n3842 = n3841 ^ n3618 ;
  assign n3843 = n3842 ^ n3700 ;
  assign n3847 = n3846 ^ n3843 ;
  assign n3612 = ~n3609 & n3611 ;
  assign n3613 = ~n3606 & n3612 ;
  assign n3619 = n3618 ^ n3613 ;
  assign n3640 = n3639 ^ n3619 ;
  assign n3641 = ~x151 & n3640 ;
  assign n3642 = n3641 ^ n3639 ;
  assign n3643 = ~x155 & ~n3642 ;
  assign n3644 = x156 ^ x153 ;
  assign n3645 = n3644 ^ n3630 ;
  assign n3646 = n3645 ^ x156 ;
  assign n3648 = x152 & n3646 ;
  assign n3649 = n3648 ^ x156 ;
  assign n3828 = x152 ^ x151 ;
  assign n3653 = n3652 ^ n3630 ;
  assign n3654 = n3828 ^ n3653 ;
  assign n3657 = n3656 ^ x156 ;
  assign n3658 = ~n3654 & n3657 ;
  assign n3661 = n3658 ^ x153 ;
  assign n3662 = ~n3649 & ~n3661 ;
  assign n3663 = n3643 & n3662 ;
  assign n3664 = n3663 ^ n3642 ;
  assign n3666 = x160 ^ x158 ;
  assign n3667 = x162 ^ x157 ;
  assign n3670 = ~x160 & ~n3667 ;
  assign n3671 = n3670 ^ x157 ;
  assign n3672 = ~n3666 & n3671 ;
  assign n3673 = ~n3665 & n3672 ;
  assign n3674 = ~x161 & n3673 ;
  assign n3702 = n3690 ^ x158 ;
  assign n3707 = n3677 & ~n3691 ;
  assign n3708 = ~n3702 & n3707 ;
  assign n3709 = n3708 ^ n3702 ;
  assign n3710 = n3709 ^ x158 ;
  assign n3711 = n3700 & ~n3710 ;
  assign n3729 = n3728 ^ n3711 ;
  assign n3730 = ~x157 & n3729 ;
  assign n3731 = n3730 ^ n3728 ;
  assign n3732 = ~n3674 & n3731 ;
  assign n3839 = ~n3664 & n3732 ;
  assign n3877 = n3842 ^ n3839 ;
  assign n3878 = n3847 & n3877 ;
  assign n3879 = n3878 ^ n3839 ;
  assign n3738 = ~x171 & ~x172 ;
  assign n3737 = x172 ^ x171 ;
  assign n3739 = n3738 ^ n3737 ;
  assign n3735 = ~x173 & ~x174 ;
  assign n3734 = x174 ^ x173 ;
  assign n3736 = n3735 ^ n3734 ;
  assign n3740 = n3739 ^ n3736 ;
  assign n3741 = n3738 ^ x170 ;
  assign n3742 = n3741 ^ n3735 ;
  assign n3745 = n3738 ^ n3735 ;
  assign n3744 = n3735 & n3738 ;
  assign n3746 = n3745 ^ n3744 ;
  assign n3747 = n3742 & n3746 ;
  assign n3743 = n3742 ^ n3736 ;
  assign n3748 = n3747 ^ n3743 ;
  assign n3749 = n3740 & n3748 ;
  assign n3750 = n3749 ^ n3739 ;
  assign n3753 = x173 ^ x170 ;
  assign n3754 = n3753 ^ x172 ;
  assign n3755 = n3754 ^ x174 ;
  assign n3751 = x173 ^ x171 ;
  assign n3756 = n3755 ^ n3751 ;
  assign n3757 = n3756 ^ x174 ;
  assign n3758 = n3757 ^ x173 ;
  assign n3759 = n3758 ^ n3751 ;
  assign n3818 = n3737 ^ n3734 ;
  assign n3765 = n3818 ^ n3751 ;
  assign n3766 = ~n3759 & ~n3765 ;
  assign n3767 = ~x173 & n3766 ;
  assign n3770 = n3767 ^ n3766 ;
  assign n3768 = n3767 ^ n3751 ;
  assign n3769 = n3756 & n3768 ;
  assign n3771 = n3770 ^ n3769 ;
  assign n3772 = n3771 ^ x173 ;
  assign n3852 = n3772 ^ x169 ;
  assign n3810 = ~x169 & ~n3772 ;
  assign n3853 = n3852 ^ n3810 ;
  assign n3854 = n3750 & n3853 ;
  assign n3780 = x167 & x168 ;
  assign n3783 = x165 & x166 ;
  assign n3789 = n3780 & n3783 ;
  assign n3788 = n3783 ^ n3780 ;
  assign n3790 = n3789 ^ n3788 ;
  assign n3782 = x166 ^ x165 ;
  assign n3784 = n3783 ^ n3782 ;
  assign n3779 = x168 ^ x167 ;
  assign n3781 = n3780 ^ n3779 ;
  assign n3786 = n3784 ^ n3781 ;
  assign n3785 = ~n3781 & ~n3784 ;
  assign n3787 = n3786 ^ n3785 ;
  assign n3791 = n3790 ^ n3787 ;
  assign n3792 = x164 ^ x163 ;
  assign n3797 = n3792 ^ n3790 ;
  assign n3798 = n3791 & ~n3797 ;
  assign n3799 = x163 & x164 ;
  assign n3800 = ~n3789 & n3799 ;
  assign n3801 = n3800 ^ n3792 ;
  assign n3802 = n3798 & n3801 ;
  assign n3803 = n3802 ^ n3800 ;
  assign n3804 = ~n3789 & ~n3803 ;
  assign n3855 = n3854 ^ n3804 ;
  assign n3814 = n3744 ^ x169 ;
  assign n3815 = ~n3747 & ~n3814 ;
  assign n3811 = n3736 & n3739 ;
  assign n3812 = n3810 & n3811 ;
  assign n3805 = n3804 ^ n3803 ;
  assign n3793 = n3792 ^ n3781 ;
  assign n3794 = n3793 ^ n3784 ;
  assign n3795 = ~n3785 & ~n3794 ;
  assign n3796 = n3791 & ~n3795 ;
  assign n3806 = n3805 ^ n3796 ;
  assign n3807 = n3806 ^ n3799 ;
  assign n3808 = n3807 ^ n3772 ;
  assign n3776 = ~x169 & ~n3771 ;
  assign n3777 = n3776 ^ x173 ;
  assign n3778 = ~n3750 & ~n3777 ;
  assign n3809 = n3808 ^ n3778 ;
  assign n3813 = n3812 ^ n3809 ;
  assign n3816 = n3815 ^ n3813 ;
  assign n3817 = x170 ^ x169 ;
  assign n3819 = n3818 ^ n3817 ;
  assign n3820 = n3792 ^ n3782 ;
  assign n3821 = n3820 ^ n3779 ;
  assign n3822 = n3819 & n3821 ;
  assign n3849 = n3822 ^ n3807 ;
  assign n3850 = ~n3816 & n3849 ;
  assign n3851 = n3850 ^ n3807 ;
  assign n3856 = n3855 ^ n3851 ;
  assign n3848 = n3847 ^ n3839 ;
  assign n3857 = n3856 ^ n3848 ;
  assign n3823 = n3822 ^ n3816 ;
  assign n3733 = n3732 ^ n3664 ;
  assign n3824 = n3823 ^ n3733 ;
  assign n3829 = n3610 ^ n3607 ;
  assign n3830 = n3829 ^ n3828 ;
  assign n3826 = n3675 ^ n3665 ;
  assign n3825 = x158 ^ x157 ;
  assign n3827 = n3826 ^ n3825 ;
  assign n3831 = n3830 ^ n3827 ;
  assign n3832 = n3821 ^ n3819 ;
  assign n3833 = n3832 ^ n3830 ;
  assign n3834 = n3831 & n3833 ;
  assign n3835 = n3834 ^ n3830 ;
  assign n3836 = n3835 ^ n3733 ;
  assign n3837 = n3824 & ~n3836 ;
  assign n3838 = n3837 ^ n3733 ;
  assign n3871 = n3856 ^ n3838 ;
  assign n3872 = ~n3857 & ~n3871 ;
  assign n3873 = n3872 ^ n3856 ;
  assign n4490 = n3879 ^ n3873 ;
  assign n4477 = n3873 & n3879 ;
  assign n4502 = n4490 ^ n4477 ;
  assign n3466 = ~x141 & ~x142 ;
  assign n3473 = ~x143 & ~x144 ;
  assign n3474 = ~n3466 & ~n3473 ;
  assign n3467 = x142 ^ x141 ;
  assign n3468 = n3467 ^ n3466 ;
  assign n3469 = x139 & x140 ;
  assign n3470 = x144 & n3469 ;
  assign n3471 = ~n3468 & n3470 ;
  assign n3472 = n3471 ^ n3469 ;
  assign n3475 = n3474 ^ n3472 ;
  assign n3478 = x144 ^ x143 ;
  assign n3479 = n3478 ^ n3473 ;
  assign n3482 = n3468 & n3479 ;
  assign n3483 = n3482 ^ n3472 ;
  assign n3484 = n3475 & ~n3483 ;
  assign n3465 = x140 ^ x139 ;
  assign n3485 = n3484 ^ n3472 ;
  assign n3486 = ~n3465 & n3485 ;
  assign n3487 = n3484 & n3486 ;
  assign n3488 = n3487 ^ n3485 ;
  assign n3489 = n3479 ^ n3468 ;
  assign n3490 = x140 & n3474 ;
  assign n3491 = n3490 ^ n3468 ;
  assign n3492 = n3489 & ~n3491 ;
  assign n3493 = n3492 ^ n3468 ;
  assign n3494 = ~n3488 & ~n3493 ;
  assign n3495 = n3494 ^ n3488 ;
  assign n3497 = ~x147 & ~x148 ;
  assign n3504 = ~x149 & ~x150 ;
  assign n3505 = ~n3497 & ~n3504 ;
  assign n3498 = x148 ^ x147 ;
  assign n3499 = n3498 ^ n3497 ;
  assign n3500 = x145 & x146 ;
  assign n3501 = x150 & n3500 ;
  assign n3502 = ~n3499 & n3501 ;
  assign n3503 = n3502 ^ n3500 ;
  assign n3506 = n3505 ^ n3503 ;
  assign n3509 = x150 ^ x149 ;
  assign n3510 = n3509 ^ n3504 ;
  assign n3513 = n3499 & n3510 ;
  assign n3514 = n3513 ^ n3503 ;
  assign n3515 = n3506 & ~n3514 ;
  assign n3496 = x146 ^ x145 ;
  assign n3516 = n3515 ^ n3503 ;
  assign n3517 = ~n3496 & n3516 ;
  assign n3518 = n3515 & n3517 ;
  assign n3519 = n3518 ^ n3516 ;
  assign n3520 = n3510 ^ n3499 ;
  assign n3521 = x146 & n3505 ;
  assign n3522 = n3521 ^ n3499 ;
  assign n3523 = n3520 & ~n3522 ;
  assign n3524 = n3523 ^ n3499 ;
  assign n3525 = ~n3519 & ~n3524 ;
  assign n3526 = n3525 ^ n3519 ;
  assign n3889 = ~n3495 & ~n3526 ;
  assign n3527 = n3526 ^ n3495 ;
  assign n4479 = n3889 ^ n3527 ;
  assign n3549 = x149 ^ x148 ;
  assign n3553 = ~n3509 & ~n3549 ;
  assign n3548 = x147 ^ x146 ;
  assign n3550 = n3549 ^ x147 ;
  assign n3551 = n3550 ^ x150 ;
  assign n3552 = ~n3548 & n3551 ;
  assign n3554 = n3553 ^ n3552 ;
  assign n3555 = ~x145 & n3554 ;
  assign n3556 = x148 ^ x146 ;
  assign n3557 = x150 ^ x145 ;
  assign n3560 = ~x148 & ~n3557 ;
  assign n3561 = n3560 ^ x145 ;
  assign n3562 = ~n3556 & n3561 ;
  assign n3563 = ~n3498 & n3562 ;
  assign n3564 = ~x149 & n3563 ;
  assign n3565 = ~n3519 & ~n3564 ;
  assign n3566 = ~n3555 & n3565 ;
  assign n3530 = x143 ^ x142 ;
  assign n3534 = ~n3478 & ~n3530 ;
  assign n3529 = x141 ^ x140 ;
  assign n3531 = n3530 ^ x141 ;
  assign n3532 = n3531 ^ x144 ;
  assign n3533 = ~n3529 & n3532 ;
  assign n3535 = n3534 ^ n3533 ;
  assign n3536 = ~x139 & n3535 ;
  assign n3537 = x142 ^ x140 ;
  assign n3538 = x144 ^ x139 ;
  assign n3541 = ~x142 & ~n3538 ;
  assign n3542 = n3541 ^ x139 ;
  assign n3543 = ~n3537 & n3542 ;
  assign n3544 = ~n3467 & n3543 ;
  assign n3545 = ~x143 & n3544 ;
  assign n3546 = ~n3488 & ~n3545 ;
  assign n3547 = ~n3536 & n3546 ;
  assign n3567 = n3566 ^ n3547 ;
  assign n3568 = n3498 ^ n3496 ;
  assign n3569 = n3568 ^ n3509 ;
  assign n3572 = n3467 ^ n3465 ;
  assign n3573 = n3572 ^ n3478 ;
  assign n3576 = n3569 & n3573 ;
  assign n3577 = n3576 ^ n3547 ;
  assign n3578 = n3567 & ~n3577 ;
  assign n3579 = n3578 ^ n3566 ;
  assign n3580 = n3573 ^ n3569 ;
  assign n3415 = x128 ^ x127 ;
  assign n3410 = x132 ^ x131 ;
  assign n3453 = n3415 ^ n3410 ;
  assign n3418 = x130 ^ x129 ;
  assign n3454 = n3453 ^ n3418 ;
  assign n3591 = n3569 ^ n3454 ;
  assign n3345 = x136 ^ x135 ;
  assign n3344 = x134 ^ x133 ;
  assign n3455 = n3345 ^ n3344 ;
  assign n3379 = x138 ^ x137 ;
  assign n3456 = n3455 ^ n3379 ;
  assign n3592 = n3591 ^ n3456 ;
  assign n3457 = n3454 & n3456 ;
  assign n3583 = n3592 ^ n3457 ;
  assign n3584 = n3583 ^ n3569 ;
  assign n3585 = n3573 ^ n3567 ;
  assign n3586 = n3585 ^ n3569 ;
  assign n3587 = n3584 & n3586 ;
  assign n3588 = n3587 ^ n3569 ;
  assign n3589 = n3580 & ~n3588 ;
  assign n3590 = n3589 ^ n3585 ;
  assign n3409 = x131 & x132 ;
  assign n3419 = n3409 ^ x130 ;
  assign n3420 = n3418 & ~n3419 ;
  assign n3429 = n3420 ^ x129 ;
  assign n3411 = n3410 ^ n3409 ;
  assign n3414 = x128 & n3411 ;
  assign n3405 = x129 & x130 ;
  assign n3421 = n3405 & n3409 ;
  assign n3430 = ~n3414 & ~n3421 ;
  assign n3431 = n3429 & n3430 ;
  assign n3432 = n3431 ^ n3429 ;
  assign n3433 = ~x127 & n3432 ;
  assign n3412 = n3411 ^ x128 ;
  assign n3413 = n3412 ^ x127 ;
  assign n3422 = n3421 ^ n3419 ;
  assign n3423 = n3422 ^ n3420 ;
  assign n3416 = n3405 ^ x128 ;
  assign n3417 = ~n3415 & ~n3416 ;
  assign n3424 = n3423 ^ n3417 ;
  assign n3425 = ~n3414 & ~n3424 ;
  assign n3426 = n3413 & n3425 ;
  assign n3428 = n3426 ^ n3417 ;
  assign n3434 = n3433 ^ n3428 ;
  assign n3406 = x127 & x128 ;
  assign n3407 = n3405 & n3406 ;
  assign n3408 = x131 & n3407 ;
  assign n3435 = n3434 ^ n3408 ;
  assign n3436 = n3429 ^ n3423 ;
  assign n3437 = n3436 ^ n3405 ;
  assign n3438 = n3437 ^ n3429 ;
  assign n3441 = x128 & n3438 ;
  assign n3442 = n3441 ^ n3429 ;
  assign n3443 = ~n3415 & n3442 ;
  assign n3444 = n3443 ^ n3429 ;
  assign n3445 = n3444 ^ n3407 ;
  assign n3446 = ~x132 & n3445 ;
  assign n3447 = n3446 ^ n3444 ;
  assign n3448 = x131 & ~n3447 ;
  assign n3449 = n3446 & n3448 ;
  assign n3450 = n3449 ^ n3447 ;
  assign n3451 = ~n3435 & ~n3450 ;
  assign n3352 = x135 & x136 ;
  assign n3346 = x137 & x138 ;
  assign n3347 = n3346 ^ x136 ;
  assign n3348 = n3345 & ~n3347 ;
  assign n3349 = n3348 ^ x135 ;
  assign n3364 = n3352 ^ n3349 ;
  assign n3353 = n3346 & n3352 ;
  assign n3354 = n3353 ^ n3347 ;
  assign n3355 = n3354 ^ n3348 ;
  assign n3365 = n3364 ^ n3355 ;
  assign n3366 = n3365 ^ n3349 ;
  assign n3369 = x134 & n3366 ;
  assign n3370 = n3369 ^ n3349 ;
  assign n3371 = ~n3344 & n3370 ;
  assign n3356 = x134 & n3355 ;
  assign n3357 = n3356 ^ n3349 ;
  assign n3358 = ~n3344 & n3357 ;
  assign n3359 = n3358 ^ n3349 ;
  assign n3360 = ~x138 & n3359 ;
  assign n3361 = n3360 ^ x138 ;
  assign n3362 = n3361 ^ n3349 ;
  assign n3372 = n3371 ^ n3362 ;
  assign n3373 = n3372 ^ n3361 ;
  assign n3374 = n3372 ^ x138 ;
  assign n3375 = x137 & ~n3374 ;
  assign n3376 = n3373 & n3375 ;
  assign n3377 = n3376 ^ n3374 ;
  assign n3378 = ~x133 & ~n3377 ;
  assign n3380 = n3379 ^ n3346 ;
  assign n3381 = x134 & n3380 ;
  assign n3389 = ~n3355 & ~n3381 ;
  assign n3382 = n3349 & ~n3353 ;
  assign n3383 = ~n3381 & n3382 ;
  assign n3384 = n3383 ^ n3349 ;
  assign n3390 = n3389 ^ n3384 ;
  assign n3391 = n3378 & n3390 ;
  assign n3392 = n3391 ^ n3377 ;
  assign n3393 = ~x137 & ~n3392 ;
  assign n3394 = n3352 ^ x134 ;
  assign n3397 = n3345 ^ x133 ;
  assign n3398 = ~x138 & n3397 ;
  assign n3399 = n3398 ^ x133 ;
  assign n3400 = ~n3352 & n3399 ;
  assign n3401 = n3400 ^ x133 ;
  assign n3402 = ~n3394 & n3401 ;
  assign n3403 = n3393 & n3402 ;
  assign n3404 = n3403 ^ n3392 ;
  assign n3452 = n3451 ^ n3404 ;
  assign n3581 = n3456 ^ n3454 ;
  assign n3594 = ~n3581 & ~n3591 ;
  assign n3593 = ~n3573 & n3592 ;
  assign n3595 = n3594 ^ n3593 ;
  assign n3596 = n3595 ^ n3567 ;
  assign n3597 = n3596 ^ n3457 ;
  assign n3600 = ~n3452 & ~n3597 ;
  assign n3601 = n3600 ^ n3596 ;
  assign n3602 = n3590 & n3601 ;
  assign n3886 = n3579 & n3602 ;
  assign n3896 = n3886 ^ n3527 ;
  assign n3603 = n3602 ^ n3579 ;
  assign n3887 = n3886 ^ n3603 ;
  assign n3462 = ~n3377 & ~n3384 ;
  assign n3461 = ~n3432 & ~n3450 ;
  assign n3463 = n3462 ^ n3461 ;
  assign n3458 = n3457 ^ n3451 ;
  assign n3459 = n3452 & n3458 ;
  assign n3460 = n3459 ^ n3457 ;
  assign n3464 = n3463 ^ n3460 ;
  assign n3897 = n3887 ^ n3464 ;
  assign n3888 = n3464 & n3887 ;
  assign n3898 = n3897 ^ n3888 ;
  assign n3901 = n4479 ^ n3886 ;
  assign n3902 = ~n3898 & n3901 ;
  assign n3890 = n3889 ^ n3888 ;
  assign n3903 = n3902 ^ n3890 ;
  assign n3904 = n3896 & n3903 ;
  assign n3883 = n3462 ^ n3460 ;
  assign n3884 = n3463 & ~n3883 ;
  assign n3885 = n3884 ^ n3462 ;
  assign n3891 = n3890 ^ n3885 ;
  assign n3905 = n3904 ^ n3891 ;
  assign n4480 = n3885 & ~n3888 ;
  assign n4481 = n3905 & ~n4480 ;
  assign n4482 = n4479 & n4481 ;
  assign n4483 = n4482 ^ n4480 ;
  assign n3858 = n3857 ^ n3838 ;
  assign n3528 = n3527 ^ n3464 ;
  assign n3604 = n3603 ^ n3528 ;
  assign n3859 = n3858 ^ n3604 ;
  assign n3598 = n3596 ^ n3452 ;
  assign n3867 = n3858 ^ n3598 ;
  assign n3861 = n3581 ^ n3580 ;
  assign n3862 = n3832 ^ n3831 ;
  assign n3863 = n3861 & n3862 ;
  assign n3860 = n3835 ^ n3824 ;
  assign n3864 = n3863 ^ n3860 ;
  assign n3865 = n3863 ^ n3598 ;
  assign n3866 = ~n3864 & n3865 ;
  assign n3868 = n3867 ^ n3866 ;
  assign n3869 = n3859 & n3868 ;
  assign n3870 = n3869 ^ n3858 ;
  assign n4478 = n3870 & n4477 ;
  assign n3874 = n3851 ^ n3804 ;
  assign n3875 = n3855 & ~n3874 ;
  assign n3876 = n3875 ^ n3804 ;
  assign n4484 = n3876 & n4483 ;
  assign n4493 = n4490 ^ n4478 ;
  assign n4491 = n3873 ^ n3870 ;
  assign n4492 = ~n4490 & n4491 ;
  assign n4494 = n4493 ^ n4492 ;
  assign n4497 = n4484 & n4494 ;
  assign n4498 = n3905 & n4497 ;
  assign n4499 = n4498 ^ n3905 ;
  assign n4485 = n4484 ^ n3876 ;
  assign n4486 = n4485 ^ n3905 ;
  assign n4500 = n4499 ^ n4486 ;
  assign n4501 = ~n4478 & n4500 ;
  assign n4503 = ~n4483 & n4501 ;
  assign n4504 = n4502 & n4503 ;
  assign n4505 = n4504 ^ n4501 ;
  assign n3880 = n3879 ^ n3876 ;
  assign n3881 = n3880 ^ n3873 ;
  assign n4507 = ~n3881 & ~n4477 ;
  assign n4508 = ~n3870 & n4507 ;
  assign n4509 = n4508 ^ n3905 ;
  assign n4510 = ~n3905 & ~n4509 ;
  assign n4511 = ~n4480 & n4510 ;
  assign n4512 = n4511 ^ n3905 ;
  assign n4519 = n4492 ^ n3870 ;
  assign n4520 = n4483 & ~n4519 ;
  assign n4533 = n4512 & ~n4520 ;
  assign n4534 = ~n4505 & n4533 ;
  assign n4542 = n4538 ^ n4534 ;
  assign n4475 = n4474 ^ n4466 ;
  assign n4441 = n4440 ^ n4407 ;
  assign n3882 = n3881 ^ n3870 ;
  assign n3906 = n3905 ^ n3882 ;
  assign n4442 = n4441 ^ n3906 ;
  assign n4445 = n4400 ^ n4399 ;
  assign n4446 = n3862 ^ n3861 ;
  assign n4447 = n4446 ^ n4400 ;
  assign n4448 = n4445 & ~n4447 ;
  assign n4449 = n4448 ^ n4399 ;
  assign n4451 = n3860 ^ n3598 ;
  assign n4452 = n4451 ^ n3863 ;
  assign n4455 = n4449 & n4452 ;
  assign n4450 = n4449 ^ n4401 ;
  assign n4453 = n4452 ^ n4450 ;
  assign n4454 = n4398 & n4453 ;
  assign n4456 = n4455 ^ n4454 ;
  assign n4443 = n4404 ^ n4379 ;
  assign n4457 = n4456 ^ n4443 ;
  assign n4458 = n3868 ^ n3604 ;
  assign n4459 = n4458 ^ n4443 ;
  assign n4460 = n4457 & n4459 ;
  assign n4444 = n4443 ^ n4441 ;
  assign n4461 = n4460 ^ n4444 ;
  assign n4462 = n4442 & ~n4461 ;
  assign n4463 = n4462 ^ n4441 ;
  assign n4476 = n4475 ^ n4463 ;
  assign n4506 = n4480 & n4494 ;
  assign n4514 = ~n3876 & n3905 ;
  assign n4515 = n4514 ^ n4512 ;
  assign n4513 = n4512 ^ n3876 ;
  assign n4516 = n4515 ^ n4513 ;
  assign n4517 = n4506 & ~n4516 ;
  assign n4518 = n4517 ^ n4515 ;
  assign n4525 = n4477 & ~n4483 ;
  assign n4526 = n4525 ^ n4520 ;
  assign n4527 = ~n4518 & n4526 ;
  assign n4528 = n4527 ^ n4512 ;
  assign n4529 = ~n4505 & n4528 ;
  assign n4530 = n4529 ^ n4463 ;
  assign n4531 = ~n4476 & n4530 ;
  assign n4532 = n4531 ^ n4529 ;
  assign n4543 = n4542 ^ n4532 ;
  assign n5680 = n5679 ^ n4543 ;
  assign n5681 = n4529 ^ n4476 ;
  assign n5682 = n5681 ^ n5660 ;
  assign n5703 = n5627 ^ n5610 ;
  assign n5684 = n4458 ^ n4457 ;
  assign n5683 = n5624 ^ n5613 ;
  assign n5685 = n5684 ^ n5683 ;
  assign n5692 = n4450 ^ n3863 ;
  assign n5693 = n5692 ^ n4401 ;
  assign n5694 = n5693 ^ n4398 ;
  assign n5695 = n5694 ^ n4451 ;
  assign n5699 = n5695 ^ n5684 ;
  assign n5686 = n5620 ^ n5619 ;
  assign n5687 = n4446 ^ n4445 ;
  assign n5688 = n5687 ^ n5620 ;
  assign n5689 = n5686 & ~n5688 ;
  assign n5690 = n5689 ^ n5619 ;
  assign n5691 = n5690 ^ n5618 ;
  assign n5696 = n5695 ^ n5621 ;
  assign n5697 = n5696 ^ n5690 ;
  assign n5698 = n5691 & n5697 ;
  assign n5700 = n5699 ^ n5698 ;
  assign n5701 = n5685 & n5700 ;
  assign n5702 = n5701 ^ n5684 ;
  assign n5704 = n5703 ^ n5702 ;
  assign n5705 = n4461 ^ n3906 ;
  assign n5706 = n5705 ^ n5702 ;
  assign n5707 = n5704 & n5706 ;
  assign n5708 = n5707 ^ n5705 ;
  assign n5709 = n5708 ^ n5681 ;
  assign n5710 = n5682 & n5709 ;
  assign n5711 = n5710 ^ n5660 ;
  assign n5712 = n5711 ^ n4543 ;
  assign n5713 = n5680 & n5712 ;
  assign n5714 = n5713 ^ n5679 ;
  assign n4535 = n4534 ^ n4532 ;
  assign n4539 = n4538 ^ n4532 ;
  assign n4540 = ~n4535 & ~n4539 ;
  assign n4541 = n4540 ^ n4534 ;
  assign n5716 = n5714 ^ n4541 ;
  assign n8725 = n5721 ^ n5716 ;
  assign n1003 = x274 ^ x273 ;
  assign n1004 = n1003 ^ x275 ;
  assign n1005 = n1004 ^ n1003 ;
  assign n1009 = n1005 ^ x273 ;
  assign n1002 = x276 ^ x272 ;
  assign n1006 = n1005 ^ n1002 ;
  assign n1007 = n1006 ^ n1004 ;
  assign n1008 = n1007 ^ n1005 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1011 = n1010 ^ n1004 ;
  assign n1012 = n1011 ^ n1009 ;
  assign n1013 = n1012 ^ n1007 ;
  assign n1014 = n1013 ^ n1007 ;
  assign n1016 = n1004 ^ x276 ;
  assign n1017 = n1016 ^ n1009 ;
  assign n1018 = ~n1014 & ~n1017 ;
  assign n1019 = ~n1004 & n1018 ;
  assign n1022 = n1019 ^ n1018 ;
  assign n1015 = n1014 ^ n1013 ;
  assign n1020 = n1019 ^ n1009 ;
  assign n1021 = n1015 & n1020 ;
  assign n1023 = n1022 ^ n1021 ;
  assign n1024 = n1023 ^ n1005 ;
  assign n1025 = x271 & n1024 ;
  assign n1026 = x273 & x274 ;
  assign n1027 = n1026 ^ n1003 ;
  assign n1028 = ~x275 & ~x276 ;
  assign n1031 = x272 & ~n1028 ;
  assign n1034 = n1031 ^ n1026 ;
  assign n1029 = x276 ^ x275 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1035 = n1031 ^ n1030 ;
  assign n1036 = n1034 & ~n1035 ;
  assign n1037 = n1036 ^ n1031 ;
  assign n1038 = n1027 & n1037 ;
  assign n1119 = n1025 & ~n1038 ;
  assign n1067 = x278 ^ x277 ;
  assign n1066 = x282 ^ x281 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n1065 = x280 ^ x279 ;
  assign n1069 = n1068 ^ n1065 ;
  assign n1070 = x272 ^ x271 ;
  assign n1072 = n1070 ^ n1016 ;
  assign n1073 = n1069 & n1072 ;
  assign n1032 = n1030 & ~n1031 ;
  assign n1033 = ~n1027 & n1032 ;
  assign n1039 = n1038 ^ n1033 ;
  assign n1040 = n1039 ^ n1024 ;
  assign n1041 = ~x271 & n1040 ;
  assign n1042 = n1041 ^ n1024 ;
  assign n1043 = ~x275 & ~n1042 ;
  assign n1044 = x276 ^ x273 ;
  assign n1045 = n1044 ^ n1002 ;
  assign n1046 = n1045 ^ x276 ;
  assign n1048 = x272 & n1046 ;
  assign n1049 = n1048 ^ x276 ;
  assign n1052 = x276 ^ x274 ;
  assign n1053 = n1052 ^ n1002 ;
  assign n1050 = x276 ^ x271 ;
  assign n1051 = n1050 ^ n1002 ;
  assign n1054 = n1053 ^ n1051 ;
  assign n1056 = n1003 ^ n1002 ;
  assign n1057 = n1056 ^ x276 ;
  assign n1058 = ~n1054 & n1057 ;
  assign n1061 = n1058 ^ x273 ;
  assign n1062 = ~n1049 & ~n1061 ;
  assign n1063 = n1043 & n1062 ;
  assign n1064 = n1063 ^ n1042 ;
  assign n1074 = n1073 ^ n1064 ;
  assign n1083 = ~x281 & ~x282 ;
  assign n1091 = x277 & x278 ;
  assign n1096 = n1091 ^ n1067 ;
  assign n1097 = n1096 ^ x280 ;
  assign n1098 = n1096 ^ x279 ;
  assign n1099 = ~n1097 & ~n1098 ;
  assign n1100 = n1099 ^ n1096 ;
  assign n1084 = n1083 ^ n1066 ;
  assign n1101 = n1091 ^ n1084 ;
  assign n1102 = n1097 ^ n1091 ;
  assign n1103 = n1102 ^ n1098 ;
  assign n1104 = ~n1101 & n1103 ;
  assign n1105 = n1104 ^ n1096 ;
  assign n1106 = n1100 & n1105 ;
  assign n1107 = n1106 ^ n1096 ;
  assign n1108 = n1107 ^ n1091 ;
  assign n1109 = ~n1083 & n1108 ;
  assign n1075 = ~x279 & ~x280 ;
  assign n1082 = n1075 ^ n1065 ;
  assign n1085 = ~n1082 & ~n1084 ;
  assign n1092 = ~n1082 & n1091 ;
  assign n1093 = ~n1085 & n1092 ;
  assign n1110 = n1109 ^ n1093 ;
  assign n1088 = ~x278 & n1069 ;
  assign n1089 = n1082 & n1083 ;
  assign n1090 = n1088 & n1089 ;
  assign n1111 = n1110 ^ n1090 ;
  assign n1113 = n1111 ^ n1064 ;
  assign n1076 = x281 ^ x278 ;
  assign n1079 = n1066 & n1076 ;
  assign n1080 = n1079 ^ x281 ;
  assign n1081 = n1075 & ~n1080 ;
  assign n1086 = n1085 ^ n1081 ;
  assign n1087 = ~x277 & n1086 ;
  assign n1112 = n1087 & ~n1111 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1115 = ~n1074 & ~n1114 ;
  assign n1116 = n1115 ^ n1073 ;
  assign n1117 = n1116 ^ n1038 ;
  assign n1120 = n1119 ^ n1117 ;
  assign n1168 = ~x291 & ~x292 ;
  assign n1166 = ~x293 & ~x294 ;
  assign n1177 = n1168 ^ n1166 ;
  assign n1176 = n1166 & n1168 ;
  assign n1178 = n1177 ^ n1176 ;
  assign n1127 = x294 ^ x293 ;
  assign n1167 = n1166 ^ n1127 ;
  assign n1128 = x292 ^ x291 ;
  assign n1169 = n1168 ^ n1128 ;
  assign n1171 = n1167 & n1169 ;
  assign n1179 = n1178 ^ n1171 ;
  assign n1129 = x290 ^ x289 ;
  assign n1187 = n1166 ^ n1129 ;
  assign n1188 = n1187 ^ n1168 ;
  assign n1189 = ~n1176 & ~n1188 ;
  assign n1190 = ~n1179 & ~n1189 ;
  assign n1170 = n1169 ^ n1167 ;
  assign n1172 = n1171 ^ n1170 ;
  assign n1173 = x289 & x290 ;
  assign n1174 = n1172 & n1173 ;
  assign n1175 = n1174 ^ n1129 ;
  assign n1180 = n1178 ^ n1129 ;
  assign n1181 = ~n1179 & n1180 ;
  assign n1182 = n1175 & n1181 ;
  assign n1183 = n1182 ^ n1174 ;
  assign n1184 = n1172 & ~n1183 ;
  assign n1185 = n1184 ^ n1183 ;
  assign n1186 = n1185 ^ n1173 ;
  assign n1191 = n1190 ^ n1186 ;
  assign n1142 = ~x287 & ~x288 ;
  assign n1140 = ~x285 & ~x286 ;
  assign n1151 = n1142 ^ n1140 ;
  assign n1150 = n1140 & n1142 ;
  assign n1152 = n1151 ^ n1150 ;
  assign n1123 = x286 ^ x285 ;
  assign n1141 = n1140 ^ n1123 ;
  assign n1121 = x288 ^ x287 ;
  assign n1143 = n1142 ^ n1121 ;
  assign n1145 = n1141 & n1143 ;
  assign n1153 = n1152 ^ n1145 ;
  assign n1122 = x284 ^ x283 ;
  assign n1161 = n1142 ^ n1122 ;
  assign n1162 = n1161 ^ n1140 ;
  assign n1163 = ~n1150 & ~n1162 ;
  assign n1164 = ~n1153 & ~n1163 ;
  assign n1144 = n1143 ^ n1141 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1147 = x283 & x284 ;
  assign n1148 = n1146 & n1147 ;
  assign n1149 = n1148 ^ n1122 ;
  assign n1154 = n1145 ^ n1122 ;
  assign n1155 = ~n1153 & n1154 ;
  assign n1156 = n1149 & n1155 ;
  assign n1157 = n1156 ^ n1148 ;
  assign n1158 = n1146 & ~n1157 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1160 = n1159 ^ n1147 ;
  assign n1165 = n1164 ^ n1160 ;
  assign n1192 = n1191 ^ n1165 ;
  assign n1124 = n1123 ^ n1122 ;
  assign n1125 = n1124 ^ n1121 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1131 = n1130 ^ n1127 ;
  assign n1193 = n1125 & n1131 ;
  assign n1126 = n1125 ^ n1072 ;
  assign n1134 = n1131 ^ n1126 ;
  assign n1135 = ~n1069 & n1134 ;
  assign n1132 = n1131 ^ n1125 ;
  assign n1133 = ~n1126 & ~n1132 ;
  assign n1136 = n1135 ^ n1133 ;
  assign n1137 = n1136 ^ n1114 ;
  assign n1194 = n1193 ^ n1137 ;
  assign n1195 = n1192 & ~n1194 ;
  assign n1138 = n1136 ^ n1073 ;
  assign n1139 = n1137 & ~n1138 ;
  assign n1196 = n1195 ^ n1139 ;
  assign n1197 = n1196 ^ n1116 ;
  assign n1198 = n1120 & n1197 ;
  assign n1199 = n1198 ^ n1116 ;
  assign n1203 = n1184 ^ n1158 ;
  assign n1200 = n1193 ^ n1165 ;
  assign n1201 = n1192 & ~n1200 ;
  assign n1202 = n1201 ^ n1191 ;
  assign n1204 = n1203 ^ n1202 ;
  assign n1207 = n1204 ^ n1120 ;
  assign n1208 = n1207 ^ n1196 ;
  assign n1094 = n1093 ^ n1085 ;
  assign n1205 = ~n1094 & ~n1109 ;
  assign n1209 = n1208 ^ n1205 ;
  assign n1214 = n1204 & n1209 ;
  assign n1215 = n1199 & n1214 ;
  assign n1206 = n1205 ^ n1204 ;
  assign n1210 = n1209 ^ n1204 ;
  assign n1211 = ~n1206 & n1210 ;
  assign n1212 = n1211 ^ n1204 ;
  assign n1213 = ~n1199 & ~n1212 ;
  assign n1216 = n1215 ^ n1213 ;
  assign n1217 = n1202 ^ n1158 ;
  assign n1218 = n1203 & n1217 ;
  assign n1219 = n1218 ^ n1184 ;
  assign n1220 = ~n1216 & n1219 ;
  assign n1221 = n1220 ^ n1213 ;
  assign n1751 = x333 & x334 ;
  assign n1749 = x335 & x336 ;
  assign n1754 = n1751 ^ n1749 ;
  assign n1539 = x336 ^ x335 ;
  assign n1750 = n1749 ^ n1539 ;
  assign n1537 = x334 ^ x333 ;
  assign n1752 = n1751 ^ n1537 ;
  assign n1753 = n1750 & n1752 ;
  assign n1761 = x332 & n1753 ;
  assign n1762 = n1761 ^ n1749 ;
  assign n1763 = n1754 & ~n1762 ;
  assign n1764 = n1763 ^ n1751 ;
  assign n1769 = ~n1753 & ~n1754 ;
  assign n1755 = n1754 ^ n1753 ;
  assign n1773 = n1755 ^ x332 ;
  assign n1770 = n1769 & ~n1773 ;
  assign n1767 = n1773 ^ n1764 ;
  assign n1771 = n1770 ^ n1767 ;
  assign n1929 = x331 & ~n1771 ;
  assign n1930 = ~n1764 & n1929 ;
  assign n1783 = x341 & x342 ;
  assign n1781 = x339 & x340 ;
  assign n1786 = n1783 ^ n1781 ;
  assign n1544 = x340 ^ x339 ;
  assign n1782 = n1781 ^ n1544 ;
  assign n1542 = x342 ^ x341 ;
  assign n1784 = n1783 ^ n1542 ;
  assign n1785 = n1782 & n1784 ;
  assign n1793 = x338 & n1785 ;
  assign n1794 = n1793 ^ n1783 ;
  assign n1795 = n1786 & ~n1794 ;
  assign n1796 = n1795 ^ n1781 ;
  assign n1801 = ~n1785 & ~n1786 ;
  assign n1787 = n1786 ^ n1785 ;
  assign n1805 = n1787 ^ x338 ;
  assign n1802 = n1801 & ~n1805 ;
  assign n1799 = n1805 ^ n1796 ;
  assign n1803 = n1802 ^ n1799 ;
  assign n1924 = x337 & ~n1803 ;
  assign n1925 = ~n1796 & n1924 ;
  assign n1926 = n1925 ^ n1796 ;
  assign n1927 = n1926 ^ n1764 ;
  assign n1931 = n1930 ^ n1927 ;
  assign n1536 = x332 ^ x331 ;
  assign n1538 = n1537 ^ n1536 ;
  assign n1540 = n1539 ^ n1538 ;
  assign n1541 = x338 ^ x337 ;
  assign n1543 = n1542 ^ n1541 ;
  assign n1545 = n1544 ^ n1543 ;
  assign n1812 = n1540 & n1545 ;
  assign n1774 = ~x331 & ~n1773 ;
  assign n1748 = n1539 ^ n1537 ;
  assign n1756 = n1755 ^ n1748 ;
  assign n1772 = n1771 ^ n1756 ;
  assign n1775 = n1774 ^ n1772 ;
  assign n1776 = n1774 ^ n1771 ;
  assign n1777 = n1536 & n1776 ;
  assign n1778 = n1775 & n1777 ;
  assign n1779 = n1778 ^ n1776 ;
  assign n1920 = n1812 ^ n1779 ;
  assign n1806 = ~x337 & ~n1805 ;
  assign n1780 = n1544 ^ n1542 ;
  assign n1788 = n1787 ^ n1780 ;
  assign n1804 = n1803 ^ n1788 ;
  assign n1807 = n1806 ^ n1804 ;
  assign n1808 = n1806 ^ n1803 ;
  assign n1809 = n1541 & n1808 ;
  assign n1810 = n1807 & n1809 ;
  assign n1811 = n1810 ^ n1808 ;
  assign n1921 = n1811 ^ n1779 ;
  assign n1922 = n1920 & ~n1921 ;
  assign n1923 = n1922 ^ n1812 ;
  assign n1932 = n1931 ^ n1923 ;
  assign n1823 = ~x321 & ~x322 ;
  assign n1829 = ~x323 & ~x324 ;
  assign n1830 = ~n1823 & ~n1829 ;
  assign n1548 = x322 ^ x321 ;
  assign n1824 = n1823 ^ n1548 ;
  assign n1825 = x319 & x320 ;
  assign n1826 = x324 & n1825 ;
  assign n1827 = ~n1824 & n1826 ;
  assign n1828 = n1827 ^ n1825 ;
  assign n1831 = n1830 ^ n1828 ;
  assign n1550 = x324 ^ x323 ;
  assign n1834 = n1829 ^ n1550 ;
  assign n1837 = n1824 & n1834 ;
  assign n1838 = n1837 ^ n1828 ;
  assign n1839 = n1831 & ~n1838 ;
  assign n1547 = x320 ^ x319 ;
  assign n1840 = n1839 ^ n1828 ;
  assign n1841 = ~n1547 & n1840 ;
  assign n1842 = n1839 & n1841 ;
  assign n1843 = n1842 ^ n1840 ;
  assign n1911 = n1834 ^ n1824 ;
  assign n1912 = x320 & n1830 ;
  assign n1913 = n1912 ^ n1824 ;
  assign n1914 = n1911 & ~n1913 ;
  assign n1915 = n1914 ^ n1824 ;
  assign n1916 = ~n1843 & ~n1915 ;
  assign n1917 = n1916 ^ n1843 ;
  assign n1864 = ~x327 & ~x328 ;
  assign n1870 = ~x329 & ~x330 ;
  assign n1871 = ~n1864 & ~n1870 ;
  assign n1553 = x328 ^ x327 ;
  assign n1865 = n1864 ^ n1553 ;
  assign n1866 = x325 & x326 ;
  assign n1867 = x330 & n1866 ;
  assign n1868 = ~n1865 & n1867 ;
  assign n1869 = n1868 ^ n1866 ;
  assign n1872 = n1871 ^ n1869 ;
  assign n1555 = x330 ^ x329 ;
  assign n1875 = n1870 ^ n1555 ;
  assign n1878 = n1865 & n1875 ;
  assign n1879 = n1878 ^ n1869 ;
  assign n1880 = n1872 & ~n1879 ;
  assign n1552 = x326 ^ x325 ;
  assign n1881 = n1880 ^ n1869 ;
  assign n1882 = ~n1552 & n1881 ;
  assign n1883 = n1880 & n1882 ;
  assign n1884 = n1883 ^ n1881 ;
  assign n1905 = n1875 ^ n1865 ;
  assign n1906 = x326 & n1871 ;
  assign n1907 = n1906 ^ n1865 ;
  assign n1908 = n1905 & ~n1907 ;
  assign n1909 = n1908 ^ n1865 ;
  assign n1910 = ~n1884 & n1909 ;
  assign n1918 = n1917 ^ n1910 ;
  assign n1857 = x329 ^ x328 ;
  assign n1861 = ~n1555 & ~n1857 ;
  assign n1856 = x327 ^ x326 ;
  assign n1858 = n1857 ^ x327 ;
  assign n1859 = n1858 ^ x330 ;
  assign n1860 = ~n1856 & n1859 ;
  assign n1862 = n1861 ^ n1860 ;
  assign n1863 = ~x325 & n1862 ;
  assign n1885 = x328 ^ x326 ;
  assign n1886 = x330 ^ x325 ;
  assign n1889 = ~x328 & ~n1886 ;
  assign n1890 = n1889 ^ x325 ;
  assign n1891 = ~n1885 & n1890 ;
  assign n1892 = ~n1553 & n1891 ;
  assign n1893 = ~x329 & n1892 ;
  assign n1894 = ~n1884 & ~n1893 ;
  assign n1895 = ~n1863 & n1894 ;
  assign n1549 = n1548 ^ n1547 ;
  assign n1551 = n1550 ^ n1549 ;
  assign n1554 = n1553 ^ n1552 ;
  assign n1556 = n1555 ^ n1554 ;
  assign n1855 = n1551 & n1556 ;
  assign n1896 = n1895 ^ n1855 ;
  assign n1816 = x323 ^ x322 ;
  assign n1820 = ~n1550 & ~n1816 ;
  assign n1815 = x321 ^ x320 ;
  assign n1817 = n1816 ^ x321 ;
  assign n1818 = n1817 ^ x324 ;
  assign n1819 = ~n1815 & n1818 ;
  assign n1821 = n1820 ^ n1819 ;
  assign n1822 = ~x319 & n1821 ;
  assign n1844 = x322 ^ x320 ;
  assign n1845 = x324 ^ x319 ;
  assign n1848 = ~x322 & ~n1845 ;
  assign n1849 = n1848 ^ x319 ;
  assign n1850 = ~n1844 & n1849 ;
  assign n1851 = ~n1548 & n1850 ;
  assign n1852 = ~x323 & n1851 ;
  assign n1853 = ~n1843 & ~n1852 ;
  assign n1854 = ~n1822 & n1853 ;
  assign n1902 = n1855 ^ n1854 ;
  assign n1903 = n1896 & n1902 ;
  assign n1904 = n1903 ^ n1855 ;
  assign n1919 = n1918 ^ n1904 ;
  assign n1933 = n1932 ^ n1919 ;
  assign n2003 = n1917 ^ n1904 ;
  assign n2004 = ~n1918 & n2003 ;
  assign n2005 = n2004 ^ n1917 ;
  assign n1897 = n1896 ^ n1854 ;
  assign n1813 = n1812 ^ n1811 ;
  assign n1814 = n1813 ^ n1779 ;
  assign n1898 = n1897 ^ n1814 ;
  assign n1546 = n1545 ^ n1540 ;
  assign n1557 = n1556 ^ n1551 ;
  assign n1746 = n1546 & n1557 ;
  assign n1934 = n1814 ^ n1746 ;
  assign n1935 = ~n1898 & n1934 ;
  assign n1936 = n1935 ^ n1746 ;
  assign n2006 = n2005 ^ n1936 ;
  assign n2007 = n2006 ^ n1932 ;
  assign n2008 = n2007 ^ n2005 ;
  assign n2009 = n1933 & n2008 ;
  assign n2010 = n2009 ^ n2006 ;
  assign n2000 = n1926 ^ n1923 ;
  assign n2001 = n1931 & n2000 ;
  assign n2002 = n2001 ^ n1926 ;
  assign n2011 = n2010 ^ n2002 ;
  assign n1670 = ~x363 & ~x364 ;
  assign n1676 = ~x365 & ~x366 ;
  assign n1677 = ~n1670 & ~n1676 ;
  assign n1513 = x364 ^ x363 ;
  assign n1671 = n1670 ^ n1513 ;
  assign n1672 = x361 & x362 ;
  assign n1673 = x366 & n1672 ;
  assign n1674 = ~n1671 & n1673 ;
  assign n1675 = n1674 ^ n1672 ;
  assign n1678 = n1677 ^ n1675 ;
  assign n1516 = x366 ^ x365 ;
  assign n1681 = n1676 ^ n1516 ;
  assign n1684 = n1671 & n1681 ;
  assign n1685 = n1684 ^ n1675 ;
  assign n1686 = n1678 & ~n1685 ;
  assign n1514 = x362 ^ x361 ;
  assign n1687 = n1686 ^ n1675 ;
  assign n1688 = ~n1514 & n1687 ;
  assign n1689 = n1686 & n1688 ;
  assign n1690 = n1689 ^ n1687 ;
  assign n1959 = n1681 ^ n1671 ;
  assign n1960 = x362 & n1677 ;
  assign n1961 = n1960 ^ n1671 ;
  assign n1962 = n1959 & ~n1961 ;
  assign n1963 = n1962 ^ n1671 ;
  assign n1964 = ~n1690 & ~n1963 ;
  assign n1965 = n1964 ^ n1690 ;
  assign n1710 = ~x357 & ~x358 ;
  assign n1716 = ~x359 & ~x360 ;
  assign n1717 = ~n1710 & ~n1716 ;
  assign n1518 = x358 ^ x357 ;
  assign n1711 = n1710 ^ n1518 ;
  assign n1712 = x355 & x356 ;
  assign n1713 = x360 & n1712 ;
  assign n1714 = ~n1711 & n1713 ;
  assign n1715 = n1714 ^ n1712 ;
  assign n1718 = n1717 ^ n1715 ;
  assign n1521 = x360 ^ x359 ;
  assign n1721 = n1716 ^ n1521 ;
  assign n1724 = n1711 & n1721 ;
  assign n1725 = n1724 ^ n1715 ;
  assign n1726 = n1718 & ~n1725 ;
  assign n1519 = x356 ^ x355 ;
  assign n1727 = n1726 ^ n1715 ;
  assign n1728 = ~n1519 & n1727 ;
  assign n1729 = n1726 & n1728 ;
  assign n1730 = n1729 ^ n1727 ;
  assign n1953 = n1721 ^ n1711 ;
  assign n1954 = x356 & n1717 ;
  assign n1955 = n1954 ^ n1711 ;
  assign n1956 = n1953 & ~n1955 ;
  assign n1957 = n1956 ^ n1711 ;
  assign n1958 = ~n1730 & n1957 ;
  assign n1966 = n1965 ^ n1958 ;
  assign n1703 = x359 ^ x358 ;
  assign n1707 = ~n1521 & ~n1703 ;
  assign n1702 = x357 ^ x356 ;
  assign n1704 = n1703 ^ x357 ;
  assign n1705 = n1704 ^ x360 ;
  assign n1706 = ~n1702 & n1705 ;
  assign n1708 = n1707 ^ n1706 ;
  assign n1709 = ~x355 & n1708 ;
  assign n1731 = x358 ^ x356 ;
  assign n1732 = x360 ^ x355 ;
  assign n1735 = ~x358 & ~n1732 ;
  assign n1736 = n1735 ^ x355 ;
  assign n1737 = ~n1731 & n1736 ;
  assign n1738 = ~n1518 & n1737 ;
  assign n1739 = ~x359 & n1738 ;
  assign n1740 = ~n1730 & ~n1739 ;
  assign n1741 = ~n1709 & n1740 ;
  assign n1663 = x365 ^ x364 ;
  assign n1667 = ~n1516 & ~n1663 ;
  assign n1662 = x363 ^ x362 ;
  assign n1664 = n1663 ^ x363 ;
  assign n1665 = n1664 ^ x366 ;
  assign n1666 = ~n1662 & n1665 ;
  assign n1668 = n1667 ^ n1666 ;
  assign n1669 = ~x361 & n1668 ;
  assign n1691 = x364 ^ x362 ;
  assign n1692 = x366 ^ x361 ;
  assign n1695 = ~x364 & ~n1692 ;
  assign n1696 = n1695 ^ x361 ;
  assign n1697 = ~n1691 & n1696 ;
  assign n1698 = ~n1513 & n1697 ;
  assign n1699 = ~x365 & n1698 ;
  assign n1700 = ~n1690 & ~n1699 ;
  assign n1701 = ~n1669 & n1700 ;
  assign n1742 = n1741 ^ n1701 ;
  assign n1515 = n1514 ^ n1513 ;
  assign n1517 = n1516 ^ n1515 ;
  assign n1520 = n1519 ^ n1518 ;
  assign n1522 = n1521 ^ n1520 ;
  assign n1660 = n1517 & n1522 ;
  assign n1950 = n1701 ^ n1660 ;
  assign n1951 = n1742 & n1950 ;
  assign n1952 = n1951 ^ n1701 ;
  assign n1967 = n1966 ^ n1952 ;
  assign n1523 = n1522 ^ n1517 ;
  assign n1532 = x348 ^ x347 ;
  assign n1530 = x346 ^ x345 ;
  assign n1529 = x344 ^ x343 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n1527 = x354 ^ x353 ;
  assign n1525 = x352 ^ x351 ;
  assign n1524 = x350 ^ x349 ;
  assign n1526 = n1525 ^ n1524 ;
  assign n1528 = n1527 ^ n1526 ;
  assign n1534 = n1533 ^ n1528 ;
  assign n1659 = n1523 & n1534 ;
  assign n1661 = n1660 ^ n1659 ;
  assign n1743 = n1742 ^ n1661 ;
  assign n1619 = ~x349 & ~n1525 ;
  assign n1620 = x353 ^ x350 ;
  assign n1621 = ~n1527 & n1620 ;
  assign n1622 = n1621 ^ x350 ;
  assign n1623 = n1622 ^ x352 ;
  assign n1639 = ~x351 & ~x352 ;
  assign n1647 = n1639 ^ n1524 ;
  assign n1648 = ~x353 & ~n1647 ;
  assign n1640 = n1639 ^ n1525 ;
  assign n1649 = n1640 ^ x354 ;
  assign n1650 = x354 ^ x350 ;
  assign n1651 = n1649 & ~n1650 ;
  assign n1652 = n1648 & n1651 ;
  assign n1625 = x349 & x350 ;
  assign n1641 = x354 & ~n1640 ;
  assign n1642 = n1625 & n1641 ;
  assign n1624 = n1525 ^ x354 ;
  assign n1626 = n1625 ^ n1624 ;
  assign n1627 = x354 ^ x352 ;
  assign n1628 = ~n1525 & ~n1627 ;
  assign n1633 = ~x353 & ~n1628 ;
  assign n1634 = n1633 ^ n1625 ;
  assign n1635 = ~n1626 & ~n1634 ;
  assign n1636 = n1635 ^ n1628 ;
  assign n1637 = n1636 ^ n1625 ;
  assign n1643 = n1642 ^ n1637 ;
  assign n1644 = ~n1524 & n1636 ;
  assign n1645 = n1643 & n1644 ;
  assign n1646 = n1645 ^ n1643 ;
  assign n1653 = n1652 ^ n1646 ;
  assign n1654 = ~n1623 & ~n1653 ;
  assign n1655 = n1619 & n1654 ;
  assign n1656 = n1655 ^ n1653 ;
  assign n1618 = n1528 & n1533 ;
  assign n1657 = n1656 ^ n1618 ;
  assign n1566 = x345 & x346 ;
  assign n1560 = x347 & x348 ;
  assign n1561 = n1560 ^ x346 ;
  assign n1562 = n1530 & ~n1561 ;
  assign n1563 = n1562 ^ x345 ;
  assign n1578 = n1566 ^ n1563 ;
  assign n1567 = n1560 & n1566 ;
  assign n1568 = n1567 ^ n1561 ;
  assign n1569 = n1568 ^ n1562 ;
  assign n1579 = n1578 ^ n1569 ;
  assign n1580 = n1579 ^ n1563 ;
  assign n1583 = x344 & n1580 ;
  assign n1584 = n1583 ^ n1563 ;
  assign n1585 = ~n1529 & n1584 ;
  assign n1570 = x344 & n1569 ;
  assign n1571 = n1570 ^ n1563 ;
  assign n1572 = ~n1529 & n1571 ;
  assign n1573 = n1572 ^ n1563 ;
  assign n1574 = ~x348 & n1573 ;
  assign n1575 = n1574 ^ x348 ;
  assign n1576 = n1575 ^ n1563 ;
  assign n1586 = n1585 ^ n1576 ;
  assign n1587 = n1586 ^ n1575 ;
  assign n1588 = n1586 ^ x348 ;
  assign n1589 = x347 & ~n1588 ;
  assign n1590 = n1587 & n1589 ;
  assign n1591 = n1590 ^ n1588 ;
  assign n1592 = ~x343 & ~n1591 ;
  assign n1593 = n1560 ^ n1532 ;
  assign n1594 = x344 & n1593 ;
  assign n1602 = ~n1569 & ~n1594 ;
  assign n1595 = n1563 & ~n1567 ;
  assign n1596 = ~n1594 & n1595 ;
  assign n1597 = n1596 ^ n1563 ;
  assign n1603 = n1602 ^ n1597 ;
  assign n1604 = n1592 & n1603 ;
  assign n1605 = n1604 ^ n1591 ;
  assign n1606 = ~x347 & ~n1605 ;
  assign n1607 = n1566 ^ x344 ;
  assign n1610 = n1530 ^ x343 ;
  assign n1611 = ~x348 & n1610 ;
  assign n1612 = n1611 ^ x343 ;
  assign n1613 = ~n1566 & n1612 ;
  assign n1614 = n1613 ^ x343 ;
  assign n1615 = ~n1607 & n1614 ;
  assign n1616 = n1606 & n1615 ;
  assign n1617 = n1616 ^ n1605 ;
  assign n1658 = n1657 ^ n1617 ;
  assign n1947 = n1659 ^ n1658 ;
  assign n1948 = n1743 & n1947 ;
  assign n1949 = n1948 ^ n1659 ;
  assign n1968 = n1967 ^ n1949 ;
  assign n1943 = ~n1591 & ~n1597 ;
  assign n1944 = n1943 ^ n1646 ;
  assign n1941 = n1622 & ~n1640 ;
  assign n1942 = ~n1646 & n1941 ;
  assign n1945 = n1944 ^ n1942 ;
  assign n1938 = n1656 ^ n1617 ;
  assign n1939 = ~n1657 & n1938 ;
  assign n1940 = n1939 ^ n1656 ;
  assign n1946 = n1945 ^ n1940 ;
  assign n1996 = n1949 ^ n1946 ;
  assign n1997 = n1968 & n1996 ;
  assign n1998 = n1997 ^ n1946 ;
  assign n1992 = n1965 ^ n1952 ;
  assign n1993 = ~n1966 & n1992 ;
  assign n1994 = n1993 ^ n1965 ;
  assign n1989 = n1943 ^ n1940 ;
  assign n1990 = ~n1945 & n1989 ;
  assign n1991 = n1990 ^ n1943 ;
  assign n1995 = n1994 ^ n1991 ;
  assign n1999 = n1998 ^ n1995 ;
  assign n2012 = n2011 ^ n1999 ;
  assign n1969 = n1968 ^ n1946 ;
  assign n1937 = n1936 ^ n1933 ;
  assign n1970 = n1969 ^ n1937 ;
  assign n1744 = n1743 ^ n1658 ;
  assign n1535 = n1534 ^ n1523 ;
  assign n1558 = n1557 ^ n1546 ;
  assign n1559 = n1535 & n1558 ;
  assign n1745 = n1744 ^ n1559 ;
  assign n1747 = n1746 ^ n1559 ;
  assign n1899 = n1898 ^ n1747 ;
  assign n1900 = n1745 & ~n1899 ;
  assign n1901 = n1900 ^ n1744 ;
  assign n1986 = n1937 ^ n1901 ;
  assign n1987 = n1970 & n1986 ;
  assign n1988 = n1987 ^ n1969 ;
  assign n2013 = n2012 ^ n1988 ;
  assign n1971 = n1970 ^ n1901 ;
  assign n1361 = x315 & x316 ;
  assign n1460 = n1361 ^ x314 ;
  assign n1461 = ~x317 & ~n1460 ;
  assign n1236 = x314 ^ x313 ;
  assign n1237 = x316 ^ x315 ;
  assign n1355 = x317 & x318 ;
  assign n1356 = n1355 ^ x316 ;
  assign n1357 = n1237 & ~n1356 ;
  assign n1358 = n1357 ^ x315 ;
  assign n1373 = n1361 ^ n1358 ;
  assign n1362 = n1355 & n1361 ;
  assign n1363 = n1362 ^ n1356 ;
  assign n1364 = n1363 ^ n1357 ;
  assign n1374 = n1373 ^ n1364 ;
  assign n1375 = n1374 ^ n1358 ;
  assign n1378 = x314 & n1375 ;
  assign n1379 = n1378 ^ n1358 ;
  assign n1380 = ~n1236 & n1379 ;
  assign n1365 = x314 & n1364 ;
  assign n1366 = n1365 ^ n1358 ;
  assign n1367 = ~n1236 & n1366 ;
  assign n1368 = n1367 ^ n1358 ;
  assign n1369 = ~x318 & n1368 ;
  assign n1370 = n1369 ^ x318 ;
  assign n1371 = n1370 ^ n1358 ;
  assign n1381 = n1380 ^ n1371 ;
  assign n1382 = n1381 ^ n1370 ;
  assign n1383 = n1381 ^ x318 ;
  assign n1384 = x317 & ~n1383 ;
  assign n1385 = n1382 & n1384 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1387 = ~x313 & ~n1386 ;
  assign n1239 = x318 ^ x317 ;
  assign n1388 = n1355 ^ n1239 ;
  assign n1389 = x314 & n1388 ;
  assign n1397 = ~n1364 & ~n1389 ;
  assign n1390 = n1358 & ~n1362 ;
  assign n1391 = ~n1389 & n1390 ;
  assign n1392 = n1391 ^ n1358 ;
  assign n1398 = n1397 ^ n1392 ;
  assign n1399 = n1387 & n1398 ;
  assign n1400 = n1399 ^ n1386 ;
  assign n1464 = n1237 ^ x313 ;
  assign n1465 = ~x318 & n1464 ;
  assign n1466 = n1465 ^ x313 ;
  assign n1467 = ~n1361 & n1466 ;
  assign n1468 = n1467 ^ x313 ;
  assign n1469 = ~n1400 & n1468 ;
  assign n1470 = n1461 & n1469 ;
  assign n1424 = x312 ^ x308 ;
  assign n1446 = x312 ^ x310 ;
  assign n1425 = ~n1424 & ~n1446 ;
  assign n1426 = n1425 ^ x309 ;
  assign n1417 = x311 ^ x309 ;
  assign n1429 = n1426 ^ n1417 ;
  assign n1430 = ~n1425 & n1429 ;
  assign n1431 = n1430 ^ n1426 ;
  assign n1243 = x310 ^ x309 ;
  assign n1450 = n1424 ^ n1243 ;
  assign n1432 = n1431 & ~n1450 ;
  assign n1433 = n1432 ^ n1426 ;
  assign n1403 = x309 & x310 ;
  assign n1404 = n1403 ^ n1243 ;
  assign n1401 = ~x311 & ~x312 ;
  assign n1242 = x312 ^ x311 ;
  assign n1405 = n1401 ^ n1242 ;
  assign n1408 = n1405 ^ n1403 ;
  assign n1402 = x308 & ~n1401 ;
  assign n1409 = n1403 ^ n1402 ;
  assign n1410 = ~n1408 & n1409 ;
  assign n1411 = n1410 ^ n1403 ;
  assign n1412 = n1404 & n1411 ;
  assign n1406 = ~n1404 & n1405 ;
  assign n1407 = ~n1402 & n1406 ;
  assign n1413 = n1412 ^ n1407 ;
  assign n1434 = n1433 ^ n1413 ;
  assign n1435 = ~x307 & n1434 ;
  assign n1436 = n1435 ^ n1433 ;
  assign n1437 = ~x311 & ~n1436 ;
  assign n1438 = x312 ^ x309 ;
  assign n1439 = n1438 ^ n1424 ;
  assign n1440 = n1439 ^ x312 ;
  assign n1442 = x308 & n1440 ;
  assign n1443 = n1442 ^ x312 ;
  assign n1447 = n1446 ^ n1424 ;
  assign n1241 = x308 ^ x307 ;
  assign n1448 = n1447 ^ n1241 ;
  assign n1451 = n1450 ^ x312 ;
  assign n1452 = ~n1448 & n1451 ;
  assign n1455 = n1452 ^ x309 ;
  assign n1456 = ~n1443 & ~n1455 ;
  assign n1457 = n1437 & n1456 ;
  assign n1458 = n1457 ^ n1436 ;
  assign n1459 = n1458 ^ n1400 ;
  assign n1471 = n1470 ^ n1459 ;
  assign n1238 = n1237 ^ n1236 ;
  assign n1240 = n1239 ^ n1238 ;
  assign n1244 = n1243 ^ n1242 ;
  assign n1245 = n1244 ^ n1241 ;
  assign n1250 = n1240 & n1245 ;
  assign n1507 = n1458 ^ n1250 ;
  assign n1508 = ~n1471 & ~n1507 ;
  assign n1509 = n1508 ^ n1250 ;
  assign n1504 = x307 & n1433 ;
  assign n1505 = ~n1412 & n1504 ;
  assign n1506 = n1505 ^ n1412 ;
  assign n1510 = n1509 ^ n1506 ;
  assign n1256 = ~x297 & ~x298 ;
  assign n1231 = x298 ^ x297 ;
  assign n1257 = n1256 ^ n1231 ;
  assign n1255 = x299 & x300 ;
  assign n1323 = n1257 ^ n1255 ;
  assign n1232 = x300 ^ x299 ;
  assign n1324 = n1255 ^ n1232 ;
  assign n1325 = n1324 ^ x296 ;
  assign n1326 = n1325 ^ n1256 ;
  assign n1329 = n1256 & ~n1324 ;
  assign n1328 = n1324 ^ n1256 ;
  assign n1330 = n1329 ^ n1328 ;
  assign n1331 = ~n1326 & ~n1330 ;
  assign n1327 = n1326 ^ n1257 ;
  assign n1332 = n1331 ^ n1327 ;
  assign n1333 = ~n1323 & ~n1332 ;
  assign n1334 = n1333 ^ n1255 ;
  assign n1301 = x299 ^ x296 ;
  assign n1302 = n1301 ^ x298 ;
  assign n1303 = n1302 ^ x300 ;
  assign n1299 = x299 ^ x297 ;
  assign n1304 = n1303 ^ n1299 ;
  assign n1305 = n1304 ^ x300 ;
  assign n1306 = n1305 ^ x299 ;
  assign n1307 = n1306 ^ n1299 ;
  assign n1311 = n1299 ^ x298 ;
  assign n1312 = n1311 ^ x300 ;
  assign n1313 = n1312 ^ n1299 ;
  assign n1314 = ~n1307 & ~n1313 ;
  assign n1315 = ~x299 & n1314 ;
  assign n1318 = n1315 ^ n1314 ;
  assign n1316 = n1315 ^ n1299 ;
  assign n1317 = n1304 & n1316 ;
  assign n1319 = n1318 ^ n1317 ;
  assign n1320 = n1319 ^ x299 ;
  assign n1343 = x295 & n1320 ;
  assign n1496 = ~n1334 & ~n1343 ;
  assign n1276 = ~x303 & ~x304 ;
  assign n1282 = ~x305 & ~x306 ;
  assign n1283 = ~n1276 & ~n1282 ;
  assign n1226 = x304 ^ x303 ;
  assign n1277 = n1276 ^ n1226 ;
  assign n1278 = x301 & x302 ;
  assign n1279 = x306 & n1278 ;
  assign n1280 = ~n1277 & n1279 ;
  assign n1281 = n1280 ^ n1278 ;
  assign n1284 = n1283 ^ n1281 ;
  assign n1225 = x306 ^ x305 ;
  assign n1287 = n1282 ^ n1225 ;
  assign n1290 = n1277 & n1287 ;
  assign n1291 = n1290 ^ n1281 ;
  assign n1292 = n1284 & ~n1291 ;
  assign n1227 = x302 ^ x301 ;
  assign n1293 = n1292 ^ n1281 ;
  assign n1294 = ~n1227 & n1293 ;
  assign n1295 = n1292 & n1294 ;
  assign n1296 = n1295 ^ n1293 ;
  assign n1490 = n1287 ^ n1277 ;
  assign n1491 = x302 & n1283 ;
  assign n1492 = n1491 ^ n1277 ;
  assign n1493 = n1490 & ~n1492 ;
  assign n1494 = n1493 ^ n1277 ;
  assign n1495 = ~n1296 & n1494 ;
  assign n1497 = n1496 ^ n1495 ;
  assign n1351 = n1329 ^ x295 ;
  assign n1352 = ~n1331 & ~n1351 ;
  assign n1258 = ~n1255 & n1257 ;
  assign n1321 = n1320 ^ x295 ;
  assign n1344 = n1343 ^ n1321 ;
  assign n1349 = n1258 & ~n1344 ;
  assign n1335 = n1334 ^ x295 ;
  assign n1339 = ~n1319 & ~n1334 ;
  assign n1340 = n1339 ^ x299 ;
  assign n1341 = ~n1335 & ~n1340 ;
  assign n1342 = n1341 ^ n1321 ;
  assign n1345 = n1344 ^ n1342 ;
  assign n1260 = x305 ^ x304 ;
  assign n1264 = ~n1225 & ~n1260 ;
  assign n1259 = x303 ^ x302 ;
  assign n1261 = n1260 ^ x303 ;
  assign n1262 = n1261 ^ x306 ;
  assign n1263 = ~n1259 & n1262 ;
  assign n1265 = n1264 ^ n1263 ;
  assign n1266 = ~x301 & n1265 ;
  assign n1267 = x304 ^ x302 ;
  assign n1268 = x306 ^ x301 ;
  assign n1271 = ~x304 & ~n1268 ;
  assign n1272 = n1271 ^ x301 ;
  assign n1273 = ~n1267 & n1272 ;
  assign n1274 = ~n1226 & n1273 ;
  assign n1275 = ~x305 & n1274 ;
  assign n1297 = ~n1275 & ~n1296 ;
  assign n1298 = ~n1266 & n1297 ;
  assign n1346 = n1345 ^ n1298 ;
  assign n1350 = n1349 ^ n1346 ;
  assign n1353 = n1352 ^ n1350 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1229 = n1228 ^ n1225 ;
  assign n1230 = x296 ^ x295 ;
  assign n1234 = n1312 ^ n1230 ;
  assign n1252 = n1229 & n1234 ;
  assign n1498 = n1298 ^ n1252 ;
  assign n1499 = ~n1353 & n1498 ;
  assign n1500 = n1499 ^ n1298 ;
  assign n2024 = n1500 ^ n1496 ;
  assign n2025 = n1497 & ~n2024 ;
  assign n2026 = n2025 ^ n1496 ;
  assign n1501 = n1500 ^ n1497 ;
  assign n2048 = n2026 ^ n1501 ;
  assign n1489 = ~n1386 & ~n1392 ;
  assign n2044 = n2026 ^ n1489 ;
  assign n2051 = n2048 ^ n2044 ;
  assign n1235 = n1234 ^ n1229 ;
  assign n1246 = n1245 ^ n1240 ;
  assign n1247 = n1246 ^ n1229 ;
  assign n1248 = n1235 & ~n1247 ;
  assign n1249 = n1248 ^ n1234 ;
  assign n1481 = n1353 ^ n1249 ;
  assign n1485 = n1471 ^ n1252 ;
  assign n1486 = n1485 ^ n1249 ;
  assign n1487 = ~n1481 & ~n1486 ;
  assign n1482 = n1481 ^ n1252 ;
  assign n1483 = n1482 ^ n1249 ;
  assign n1484 = ~n1250 & ~n1483 ;
  assign n1488 = n1487 ^ n1484 ;
  assign n1503 = n2051 ^ n1488 ;
  assign n1511 = n1510 ^ n1503 ;
  assign n1251 = n1250 ^ n1249 ;
  assign n1354 = n1353 ^ n1251 ;
  assign n1472 = n1471 ^ n1354 ;
  assign n1222 = n1192 ^ n1136 ;
  assign n1223 = n1222 ^ n1114 ;
  assign n1473 = n1472 ^ n1223 ;
  assign n1474 = n1131 ^ n1069 ;
  assign n1475 = n1474 ^ n1126 ;
  assign n1476 = n1246 ^ n1235 ;
  assign n1477 = n1475 & n1476 ;
  assign n1478 = n1477 ^ n1223 ;
  assign n1479 = n1473 & ~n1478 ;
  assign n1224 = n1223 ^ n1209 ;
  assign n1480 = n1479 ^ n1224 ;
  assign n1512 = n1511 ^ n1480 ;
  assign n1972 = n1971 ^ n1512 ;
  assign n1976 = n1747 ^ n1744 ;
  assign n1977 = n1976 ^ n1898 ;
  assign n1982 = n1977 ^ n1971 ;
  assign n1973 = n1476 ^ n1475 ;
  assign n1974 = n1558 ^ n1535 ;
  assign n1975 = n1973 & n1974 ;
  assign n1978 = n1977 ^ n1975 ;
  assign n3267 = n1975 ^ n1477 ;
  assign n3268 = n3267 ^ n1473 ;
  assign n1981 = n1978 & ~n3268 ;
  assign n1983 = n1982 ^ n1981 ;
  assign n1984 = ~n1972 & n1983 ;
  assign n1985 = n1984 ^ n1971 ;
  assign n2014 = n2013 ^ n1985 ;
  assign n2039 = n1488 & n1501 ;
  assign n2040 = ~n1506 & ~n1509 ;
  assign n2041 = n2040 ^ n1510 ;
  assign n2042 = n2041 ^ n2026 ;
  assign n2045 = n2044 ^ n2042 ;
  assign n2046 = n2041 & n2045 ;
  assign n2047 = n2046 ^ n2042 ;
  assign n2056 = n2042 ^ n1489 ;
  assign n2049 = n2026 ^ n1488 ;
  assign n2050 = n2049 ^ n2048 ;
  assign n2052 = n2051 ^ n2026 ;
  assign n2053 = n2052 ^ n2042 ;
  assign n2054 = ~n2050 & ~n2053 ;
  assign n2057 = n2056 ^ n2054 ;
  assign n2058 = n2047 & n2057 ;
  assign n2059 = n2058 ^ n2042 ;
  assign n2060 = n2059 ^ n2026 ;
  assign n2061 = n2060 ^ n2042 ;
  assign n2062 = ~n1503 & n2040 ;
  assign n2063 = ~n2061 & n2062 ;
  assign n2064 = n2063 ^ n2061 ;
  assign n2027 = n1489 ^ n1488 ;
  assign n2021 = n1506 ^ n1501 ;
  assign n2028 = n2021 ^ n1509 ;
  assign n2029 = n2028 ^ n1488 ;
  assign n2030 = n2027 & n2029 ;
  assign n2035 = n1488 & n2030 ;
  assign n2036 = n2035 ^ n2021 ;
  assign n2037 = n1510 & ~n2036 ;
  assign n2031 = n2030 ^ n2021 ;
  assign n2032 = n2031 ^ n2026 ;
  assign n2038 = n2037 ^ n2032 ;
  assign n2065 = n2038 ^ n2026 ;
  assign n2066 = ~n2064 & n2065 ;
  assign n2067 = n2039 & n2066 ;
  assign n2068 = n2067 ^ n2038 ;
  assign n2015 = n1219 ^ n1216 ;
  assign n2016 = n2015 ^ n1209 ;
  assign n2017 = n2016 ^ n1511 ;
  assign n2018 = n2017 ^ n2015 ;
  assign n2019 = n1480 & n2018 ;
  assign n2020 = n2019 ^ n2016 ;
  assign n2069 = n2068 ^ n2020 ;
  assign n2070 = n2069 ^ n1985 ;
  assign n2071 = ~n2014 & n2070 ;
  assign n2072 = n2071 ^ n2069 ;
  assign n2073 = n1998 & n2011 ;
  assign n2074 = n2005 ^ n2002 ;
  assign n2075 = n2010 & n2074 ;
  assign n2076 = n2075 ^ n2005 ;
  assign n2077 = n2073 & n2076 ;
  assign n2078 = n2068 ^ n2015 ;
  assign n2079 = ~n2020 & ~n2078 ;
  assign n2080 = n2079 ^ n2015 ;
  assign n2081 = n2064 & ~n2080 ;
  assign n2082 = ~n2077 & n2081 ;
  assign n2083 = ~n2072 & n2082 ;
  assign n2084 = n1221 & ~n2083 ;
  assign n2087 = ~n1991 & n1994 ;
  assign n2092 = n2087 ^ n1995 ;
  assign n2093 = n1988 & n2092 ;
  assign n2105 = n2093 ^ n2011 ;
  assign n2088 = ~n1988 & n2087 ;
  assign n2091 = n2088 ^ n1995 ;
  assign n2094 = n2093 ^ n2091 ;
  assign n2095 = n2094 ^ n1988 ;
  assign n2106 = n2093 ^ n1998 ;
  assign n2107 = n2095 & ~n2106 ;
  assign n2108 = ~n2105 & n2107 ;
  assign n2109 = n2108 ^ n2093 ;
  assign n2085 = n2076 ^ n1998 ;
  assign n2086 = n2085 ^ n2011 ;
  assign n2089 = n2088 ^ n1998 ;
  assign n2090 = n2089 ^ n2011 ;
  assign n2096 = n2095 ^ n2088 ;
  assign n2097 = n2096 ^ n2076 ;
  assign n2098 = ~n2090 & ~n2097 ;
  assign n2099 = ~n2086 & n2098 ;
  assign n2100 = n2099 ^ n2088 ;
  assign n2101 = n2100 ^ n2076 ;
  assign n2102 = n2011 & n2101 ;
  assign n2103 = ~n2076 & n2102 ;
  assign n2104 = n2103 ^ n2076 ;
  assign n2111 = n2109 ^ n2104 ;
  assign n2110 = n2104 & ~n2109 ;
  assign n2112 = n2111 ^ n2110 ;
  assign n2113 = n2080 ^ n2072 ;
  assign n2114 = n2080 ^ n2064 ;
  assign n2115 = n2113 & ~n2114 ;
  assign n2116 = n2115 ^ n2080 ;
  assign n2117 = n2112 & ~n2116 ;
  assign n2118 = n2084 & ~n2117 ;
  assign n2124 = n2110 ^ n2080 ;
  assign n2125 = n2124 ^ n2064 ;
  assign n2126 = n2072 & n2125 ;
  assign n2127 = n2126 ^ n2110 ;
  assign n2128 = n2077 & ~n2095 ;
  assign n2129 = n2128 ^ n2124 ;
  assign n2130 = n2126 ^ n2125 ;
  assign n2131 = ~n2129 & n2130 ;
  assign n2132 = n2131 ^ n2124 ;
  assign n2133 = n2127 & n2132 ;
  assign n2134 = n2133 ^ n2110 ;
  assign n2135 = n2118 & ~n2134 ;
  assign n2420 = ~x375 & ~x376 ;
  assign n2426 = ~x377 & ~x378 ;
  assign n2427 = ~n2420 & ~n2426 ;
  assign n2409 = x376 ^ x375 ;
  assign n2421 = n2420 ^ n2409 ;
  assign n2422 = x373 & x374 ;
  assign n2423 = x378 & n2422 ;
  assign n2424 = ~n2421 & n2423 ;
  assign n2425 = n2424 ^ n2422 ;
  assign n2428 = n2427 ^ n2425 ;
  assign n2405 = x378 ^ x377 ;
  assign n2431 = n2426 ^ n2405 ;
  assign n2434 = n2421 & n2431 ;
  assign n2435 = n2434 ^ n2425 ;
  assign n2436 = n2428 & ~n2435 ;
  assign n2419 = x374 ^ x373 ;
  assign n2437 = n2436 ^ n2425 ;
  assign n2438 = ~n2419 & n2437 ;
  assign n2439 = n2436 & n2438 ;
  assign n2440 = n2439 ^ n2437 ;
  assign n2495 = n2431 ^ n2421 ;
  assign n2496 = x374 & n2427 ;
  assign n2497 = n2496 ^ n2421 ;
  assign n2498 = n2495 & ~n2497 ;
  assign n2499 = n2498 ^ n2421 ;
  assign n2500 = ~n2440 & ~n2499 ;
  assign n2501 = n2500 ^ n2440 ;
  assign n2444 = x371 ^ x370 ;
  assign n2448 = x372 ^ x371 ;
  assign n2449 = ~n2444 & ~n2448 ;
  assign n2443 = x369 ^ x368 ;
  assign n2445 = n2444 ^ x369 ;
  assign n2446 = n2445 ^ x372 ;
  assign n2447 = ~n2443 & n2446 ;
  assign n2450 = n2449 ^ n2447 ;
  assign n2451 = ~x367 & n2450 ;
  assign n2452 = x370 ^ x369 ;
  assign n2453 = x370 ^ x368 ;
  assign n2454 = x372 ^ x367 ;
  assign n2457 = ~x370 & ~n2454 ;
  assign n2458 = n2457 ^ x367 ;
  assign n2459 = ~n2453 & n2458 ;
  assign n2460 = ~n2452 & n2459 ;
  assign n2461 = ~x371 & n2460 ;
  assign n2463 = ~x369 & ~x370 ;
  assign n2469 = ~x371 & ~x372 ;
  assign n2470 = ~n2463 & ~n2469 ;
  assign n2464 = n2463 ^ n2452 ;
  assign n2465 = x367 & x368 ;
  assign n2466 = x372 & n2465 ;
  assign n2467 = ~n2464 & n2466 ;
  assign n2468 = n2467 ^ n2465 ;
  assign n2471 = n2470 ^ n2468 ;
  assign n2474 = n2469 ^ n2448 ;
  assign n2477 = n2464 & n2474 ;
  assign n2478 = n2477 ^ n2468 ;
  assign n2479 = n2471 & ~n2478 ;
  assign n2462 = x368 ^ x367 ;
  assign n2480 = n2479 ^ n2468 ;
  assign n2481 = ~n2462 & n2480 ;
  assign n2482 = n2479 & n2481 ;
  assign n2483 = n2482 ^ n2480 ;
  assign n2484 = ~n2461 & ~n2483 ;
  assign n2485 = ~n2451 & n2484 ;
  assign n2401 = x377 ^ x376 ;
  assign n2406 = ~n2401 & ~n2405 ;
  assign n2400 = x375 ^ x374 ;
  assign n2402 = n2401 ^ x375 ;
  assign n2403 = n2402 ^ x378 ;
  assign n2404 = ~n2400 & n2403 ;
  assign n2407 = n2406 ^ n2404 ;
  assign n2408 = ~x373 & n2407 ;
  assign n2410 = x376 ^ x374 ;
  assign n2411 = x378 ^ x373 ;
  assign n2414 = ~x376 & ~n2411 ;
  assign n2415 = n2414 ^ x373 ;
  assign n2416 = ~n2410 & n2415 ;
  assign n2417 = ~n2409 & n2416 ;
  assign n2418 = ~x377 & n2417 ;
  assign n2441 = ~n2418 & ~n2440 ;
  assign n2442 = ~n2408 & n2441 ;
  assign n2486 = n2485 ^ n2442 ;
  assign n2487 = n2419 ^ n2405 ;
  assign n2488 = n2487 ^ n2409 ;
  assign n2489 = n2462 ^ n2448 ;
  assign n2490 = n2489 ^ n2452 ;
  assign n2491 = n2488 & n2490 ;
  assign n2492 = n2491 ^ n2485 ;
  assign n2493 = n2486 & n2492 ;
  assign n2494 = n2493 ^ n2485 ;
  assign n2502 = n2501 ^ n2494 ;
  assign n2509 = x390 ^ x389 ;
  assign n2535 = x389 ^ x388 ;
  assign n2539 = ~n2509 & ~n2535 ;
  assign n2534 = x387 ^ x386 ;
  assign n2536 = n2535 ^ x387 ;
  assign n2537 = n2536 ^ x390 ;
  assign n2538 = ~n2534 & n2537 ;
  assign n2540 = n2539 ^ n2538 ;
  assign n2541 = ~x385 & n2540 ;
  assign n2510 = x388 ^ x387 ;
  assign n2542 = x388 ^ x386 ;
  assign n2543 = x390 ^ x385 ;
  assign n2546 = ~x388 & ~n2543 ;
  assign n2547 = n2546 ^ x385 ;
  assign n2548 = ~n2542 & n2547 ;
  assign n2549 = ~n2510 & n2548 ;
  assign n2550 = ~x389 & n2549 ;
  assign n2551 = ~x387 & ~x388 ;
  assign n2557 = ~x389 & ~x390 ;
  assign n2558 = ~n2551 & ~n2557 ;
  assign n2552 = n2551 ^ n2510 ;
  assign n2553 = x385 & x386 ;
  assign n2554 = x390 & n2553 ;
  assign n2555 = ~n2552 & n2554 ;
  assign n2556 = n2555 ^ n2553 ;
  assign n2559 = n2558 ^ n2556 ;
  assign n2562 = n2557 ^ n2509 ;
  assign n2565 = n2552 & n2562 ;
  assign n2566 = n2565 ^ n2556 ;
  assign n2567 = n2559 & ~n2566 ;
  assign n2511 = x386 ^ x385 ;
  assign n2568 = n2567 ^ n2556 ;
  assign n2569 = ~n2511 & n2568 ;
  assign n2570 = n2567 & n2569 ;
  assign n2571 = n2570 ^ n2568 ;
  assign n2572 = ~n2550 & ~n2571 ;
  assign n2573 = ~n2541 & n2572 ;
  assign n2519 = x383 & x384 ;
  assign n2517 = x381 & x382 ;
  assign n2525 = n2519 ^ n2517 ;
  assign n2523 = n2517 & n2519 ;
  assign n2526 = n2525 ^ n2523 ;
  assign n2516 = x379 & x380 ;
  assign n2524 = n2516 & ~n2523 ;
  assign n2527 = n2526 ^ n2524 ;
  assign n2504 = x382 ^ x381 ;
  assign n2518 = n2517 ^ n2504 ;
  assign n2506 = x384 ^ x383 ;
  assign n2520 = n2519 ^ n2506 ;
  assign n2528 = n2518 & n2520 ;
  assign n2529 = n2528 ^ n2526 ;
  assign n2505 = x380 ^ x379 ;
  assign n2530 = n2528 ^ n2505 ;
  assign n2531 = ~n2529 & ~n2530 ;
  assign n2532 = n2527 & n2531 ;
  assign n2533 = n2532 ^ n2524 ;
  assign n2574 = n2573 ^ n2533 ;
  assign n2521 = ~n2518 & ~n2520 ;
  assign n2522 = ~n2516 & n2521 ;
  assign n2575 = n2574 ^ n2522 ;
  assign n2576 = n2575 ^ n2573 ;
  assign n2583 = ~x380 & ~n2526 ;
  assign n2584 = ~n2528 & n2583 ;
  assign n2585 = n2584 ^ n2528 ;
  assign n2577 = n2528 ^ n2523 ;
  assign n2586 = n2585 ^ n2577 ;
  assign n2587 = ~x379 & n2586 ;
  assign n2588 = ~n2576 & n2587 ;
  assign n2589 = n2588 ^ n2575 ;
  assign n2512 = n2511 ^ n2510 ;
  assign n2513 = n2512 ^ n2509 ;
  assign n2507 = n2506 ^ n2505 ;
  assign n2508 = n2507 ^ n2504 ;
  assign n2514 = n2513 ^ n2508 ;
  assign n2515 = n2514 ^ n2490 ;
  assign n2590 = n2508 & n2513 ;
  assign n2591 = n2590 ^ n2589 ;
  assign n2592 = n2591 ^ n2488 ;
  assign n2593 = n2592 ^ n2514 ;
  assign n2594 = n2593 ^ n2591 ;
  assign n2595 = ~n2515 & n2594 ;
  assign n2596 = n2595 ^ n2592 ;
  assign n2597 = n2596 ^ n2486 ;
  assign n2598 = n2597 ^ n2590 ;
  assign n2503 = n2491 ^ n2486 ;
  assign n2599 = n2598 ^ n2503 ;
  assign n2601 = n2589 & n2599 ;
  assign n2602 = n2601 ^ n2590 ;
  assign n2603 = n2596 ^ n2503 ;
  assign n2604 = n2601 ^ n2599 ;
  assign n2605 = n2603 & n2604 ;
  assign n2606 = n2605 ^ n2503 ;
  assign n2607 = ~n2602 & n2606 ;
  assign n2608 = n2607 ^ n2501 ;
  assign n2609 = n2502 & n2608 ;
  assign n2610 = n2609 ^ n2501 ;
  assign n2611 = n2474 ^ n2464 ;
  assign n2612 = x368 & n2470 ;
  assign n2613 = n2612 ^ n2464 ;
  assign n2614 = n2611 & ~n2613 ;
  assign n2615 = n2614 ^ n2464 ;
  assign n2616 = ~n2483 & ~n2615 ;
  assign n2617 = n2616 ^ n2483 ;
  assign n2632 = n2617 ^ n2494 ;
  assign n2622 = n2562 ^ n2552 ;
  assign n2623 = x386 & n2558 ;
  assign n2624 = n2623 ^ n2552 ;
  assign n2625 = n2622 & ~n2624 ;
  assign n2626 = n2625 ^ n2552 ;
  assign n2627 = ~n2571 & ~n2626 ;
  assign n2628 = n2627 ^ n2571 ;
  assign n2621 = ~n2523 & ~n2533 ;
  assign n2629 = n2628 ^ n2621 ;
  assign n2618 = n2590 ^ n2573 ;
  assign n2619 = n2589 & n2618 ;
  assign n2620 = n2619 ^ n2590 ;
  assign n2630 = n2629 ^ n2620 ;
  assign n2633 = n2632 ^ n2630 ;
  assign n2634 = n2633 ^ n2608 ;
  assign n2631 = n2630 ^ n2617 ;
  assign n2635 = n2634 ^ n2617 ;
  assign n2636 = ~n2631 & ~n2635 ;
  assign n2637 = n2636 ^ n2630 ;
  assign n2641 = n2634 & ~n2637 ;
  assign n2642 = n2610 & n2641 ;
  assign n2638 = ~n2610 & n2637 ;
  assign n2649 = n2642 ^ n2638 ;
  assign n2643 = n2628 ^ n2620 ;
  assign n2644 = ~n2629 & n2643 ;
  assign n2645 = n2644 ^ n2628 ;
  assign n2650 = n2649 ^ n2645 ;
  assign n2160 = x414 ^ x413 ;
  assign n2165 = x413 ^ x410 ;
  assign n2159 = x412 ^ x411 ;
  assign n2166 = n2165 ^ n2159 ;
  assign n2167 = n2160 & n2166 ;
  assign n2168 = n2167 ^ x413 ;
  assign n2161 = n2160 ^ n2159 ;
  assign n2158 = x410 ^ x409 ;
  assign n2162 = n2161 ^ n2158 ;
  assign n2163 = x409 & ~n2162 ;
  assign n2343 = n2168 ^ n2163 ;
  assign n2170 = x411 ^ x410 ;
  assign n2171 = ~n2159 & n2170 ;
  assign n2344 = n2171 ^ x410 ;
  assign n2345 = n2344 ^ n2163 ;
  assign n2346 = n2343 & ~n2345 ;
  assign n2347 = n2346 ^ n2168 ;
  assign n2183 = ~x405 & ~x406 ;
  assign n2190 = ~x407 & ~x408 ;
  assign n2191 = ~n2183 & ~n2190 ;
  assign n2184 = x406 ^ x405 ;
  assign n2185 = n2184 ^ n2183 ;
  assign n2186 = x403 & x404 ;
  assign n2187 = x408 & n2186 ;
  assign n2188 = ~n2185 & n2187 ;
  assign n2189 = n2188 ^ n2186 ;
  assign n2192 = n2191 ^ n2189 ;
  assign n2178 = x408 ^ x407 ;
  assign n2195 = n2190 ^ n2178 ;
  assign n2198 = n2185 & n2195 ;
  assign n2199 = n2198 ^ n2189 ;
  assign n2200 = n2192 & ~n2199 ;
  assign n2182 = x404 ^ x403 ;
  assign n2201 = n2200 ^ n2189 ;
  assign n2202 = ~n2182 & n2201 ;
  assign n2203 = n2200 & n2202 ;
  assign n2204 = n2203 ^ n2201 ;
  assign n2348 = n2195 ^ n2185 ;
  assign n2349 = x404 & n2191 ;
  assign n2350 = n2349 ^ n2185 ;
  assign n2351 = n2348 & ~n2350 ;
  assign n2352 = n2351 ^ n2185 ;
  assign n2353 = ~n2204 & ~n2352 ;
  assign n2354 = n2353 ^ n2204 ;
  assign n2372 = ~n2347 & ~n2354 ;
  assign n2355 = n2354 ^ n2347 ;
  assign n2382 = n2372 ^ n2355 ;
  assign n2302 = ~x393 & ~x394 ;
  assign n2308 = ~x395 & ~x396 ;
  assign n2309 = ~n2302 & ~n2308 ;
  assign n2229 = x394 ^ x393 ;
  assign n2303 = n2302 ^ n2229 ;
  assign n2304 = x391 & x392 ;
  assign n2305 = x396 & n2304 ;
  assign n2306 = ~n2303 & n2305 ;
  assign n2307 = n2306 ^ n2304 ;
  assign n2310 = n2309 ^ n2307 ;
  assign n2232 = x396 ^ x395 ;
  assign n2313 = n2308 ^ n2232 ;
  assign n2316 = n2303 & n2313 ;
  assign n2317 = n2316 ^ n2307 ;
  assign n2318 = n2310 & ~n2317 ;
  assign n2230 = x392 ^ x391 ;
  assign n2319 = n2318 ^ n2307 ;
  assign n2320 = ~n2230 & n2319 ;
  assign n2321 = n2318 & n2320 ;
  assign n2322 = n2321 ^ n2319 ;
  assign n2361 = n2313 ^ n2303 ;
  assign n2362 = x392 & n2309 ;
  assign n2363 = n2362 ^ n2303 ;
  assign n2364 = n2361 & ~n2363 ;
  assign n2365 = n2364 ^ n2303 ;
  assign n2366 = ~n2322 & ~n2365 ;
  assign n2367 = n2366 ^ n2322 ;
  assign n2259 = x397 & x398 ;
  assign n2251 = x399 & x400 ;
  assign n2252 = x401 & x402 ;
  assign n2260 = n2251 & ~n2252 ;
  assign n2261 = ~n2259 & n2260 ;
  assign n2262 = n2261 ^ n2251 ;
  assign n2224 = x402 ^ x401 ;
  assign n2253 = n2252 ^ n2224 ;
  assign n2223 = x398 ^ x397 ;
  assign n2264 = n2259 ^ n2223 ;
  assign n2265 = n2264 ^ x400 ;
  assign n2266 = n2264 ^ x399 ;
  assign n2267 = ~n2265 & ~n2266 ;
  assign n2268 = n2267 ^ n2264 ;
  assign n2269 = n2265 ^ n2252 ;
  assign n2270 = n2269 ^ n2266 ;
  assign n2272 = n2265 ^ n2259 ;
  assign n2273 = n2272 ^ n2266 ;
  assign n2274 = ~n2270 & n2273 ;
  assign n2275 = n2274 ^ n2264 ;
  assign n2276 = n2268 & n2275 ;
  assign n2277 = n2276 ^ n2264 ;
  assign n2278 = n2277 ^ n2259 ;
  assign n2279 = n2253 & n2278 ;
  assign n2360 = ~n2262 & ~n2279 ;
  assign n2368 = n2367 ^ n2360 ;
  assign n2295 = x395 ^ x394 ;
  assign n2299 = ~n2232 & ~n2295 ;
  assign n2294 = x393 ^ x392 ;
  assign n2296 = n2295 ^ x393 ;
  assign n2297 = n2296 ^ x396 ;
  assign n2298 = ~n2294 & n2297 ;
  assign n2300 = n2299 ^ n2298 ;
  assign n2301 = ~x391 & n2300 ;
  assign n2323 = x394 ^ x392 ;
  assign n2324 = x396 ^ x391 ;
  assign n2327 = ~x394 & ~n2324 ;
  assign n2328 = n2327 ^ x391 ;
  assign n2329 = ~n2323 & n2328 ;
  assign n2330 = ~n2229 & n2329 ;
  assign n2331 = ~x395 & n2330 ;
  assign n2332 = ~n2322 & ~n2331 ;
  assign n2333 = ~n2301 & n2332 ;
  assign n2280 = n2279 ^ x397 ;
  assign n2292 = n2280 ^ n2252 ;
  assign n2226 = x400 ^ x399 ;
  assign n2225 = n2224 ^ n2223 ;
  assign n2227 = n2226 ^ n2225 ;
  assign n2282 = n2227 ^ x397 ;
  assign n2289 = ~n2227 & n2280 ;
  assign n2283 = n2251 ^ n2226 ;
  assign n2284 = ~n2252 & ~n2283 ;
  assign n2290 = n2289 ^ n2284 ;
  assign n2291 = n2282 & ~n2290 ;
  assign n2293 = n2292 ^ n2291 ;
  assign n2334 = n2333 ^ n2293 ;
  assign n2263 = n2227 & ~n2262 ;
  assign n2335 = n2334 ^ n2263 ;
  assign n2256 = ~x398 & ~n2253 ;
  assign n2257 = n2256 ^ n2252 ;
  assign n2258 = ~n2251 & n2257 ;
  assign n2336 = n2335 ^ n2258 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2233 = n2232 ^ n2231 ;
  assign n2247 = n2227 & n2233 ;
  assign n2357 = n2333 ^ n2247 ;
  assign n2358 = ~n2336 & n2357 ;
  assign n2359 = n2358 ^ n2333 ;
  assign n2369 = n2368 ^ n2359 ;
  assign n2174 = x407 ^ x406 ;
  assign n2179 = ~n2174 & ~n2178 ;
  assign n2173 = x405 ^ x404 ;
  assign n2175 = n2174 ^ x405 ;
  assign n2176 = n2175 ^ x408 ;
  assign n2177 = ~n2173 & n2176 ;
  assign n2180 = n2179 ^ n2177 ;
  assign n2181 = ~x403 & n2180 ;
  assign n2205 = x406 ^ x404 ;
  assign n2206 = x408 ^ x403 ;
  assign n2209 = ~x406 & ~n2206 ;
  assign n2210 = n2209 ^ x403 ;
  assign n2211 = ~n2205 & n2210 ;
  assign n2212 = ~n2184 & n2211 ;
  assign n2213 = ~x407 & n2212 ;
  assign n2214 = ~n2204 & ~n2213 ;
  assign n2215 = ~n2181 & n2214 ;
  assign n2164 = n2163 ^ x410 ;
  assign n2169 = n2168 ^ n2164 ;
  assign n2172 = n2171 ^ n2169 ;
  assign n2216 = n2215 ^ n2172 ;
  assign n2228 = n2227 ^ n2162 ;
  assign n2217 = n2184 ^ n2182 ;
  assign n2218 = n2217 ^ n2178 ;
  assign n2234 = n2233 ^ n2218 ;
  assign n2235 = n2234 ^ n2162 ;
  assign n2236 = n2228 & ~n2235 ;
  assign n2237 = n2236 ^ n2227 ;
  assign n2240 = n2218 & n2233 ;
  assign n2243 = ~n2237 & ~n2240 ;
  assign n2219 = n2162 & n2218 ;
  assign n2244 = n2243 ^ n2219 ;
  assign n2245 = ~n2216 & n2244 ;
  assign n2246 = n2245 ^ n2219 ;
  assign n2248 = n2240 ^ n2237 ;
  assign n2249 = n2248 ^ n2216 ;
  assign n2250 = n2249 ^ n2247 ;
  assign n2339 = n2250 & ~n2336 ;
  assign n2340 = n2339 ^ n2249 ;
  assign n2341 = ~n2246 & ~n2340 ;
  assign n2220 = n2219 ^ n2215 ;
  assign n2221 = n2216 & n2220 ;
  assign n2222 = n2221 ^ n2215 ;
  assign n2379 = n2341 ^ n2222 ;
  assign n2342 = n2222 & n2341 ;
  assign n2380 = n2379 ^ n2342 ;
  assign n2381 = ~n2369 & n2380 ;
  assign n2389 = n2382 ^ n2381 ;
  assign n2393 = n2389 ^ n2341 ;
  assign n2394 = ~n2379 & n2382 ;
  assign n2395 = n2393 & n2394 ;
  assign n2387 = n2369 & n2382 ;
  assign n2356 = n2355 ^ n2222 ;
  assign n2370 = n2369 ^ n2356 ;
  assign n2371 = n2370 ^ n2341 ;
  assign n2373 = ~n2371 & n2372 ;
  assign n2388 = n2387 ^ n2373 ;
  assign n2390 = n2389 ^ n2388 ;
  assign n2374 = n2367 ^ n2359 ;
  assign n2375 = ~n2368 & n2374 ;
  assign n2376 = n2375 ^ n2367 ;
  assign n2391 = n2390 ^ n2376 ;
  assign n2396 = n2395 ^ n2391 ;
  assign n2651 = n2650 ^ n2396 ;
  assign n2652 = n2490 ^ n2488 ;
  assign n2653 = n2652 ^ n2514 ;
  assign n2654 = n2234 ^ n2228 ;
  assign n2655 = n2653 & n2654 ;
  assign n2337 = n2336 ^ n2249 ;
  assign n2656 = n2655 ^ n2337 ;
  assign n2657 = n2597 ^ n2337 ;
  assign n2658 = ~n2656 & n2657 ;
  assign n2659 = n2658 ^ n2337 ;
  assign n2660 = n2659 ^ n2634 ;
  assign n2661 = n2634 ^ n2396 ;
  assign n2662 = n2661 ^ n2371 ;
  assign n2663 = n2662 ^ n2396 ;
  assign n2664 = n2660 & n2663 ;
  assign n2665 = n2664 ^ n2661 ;
  assign n2666 = n2651 & ~n2665 ;
  assign n2667 = n2666 ^ n2650 ;
  assign n2646 = ~n2642 & ~n2645 ;
  assign n2647 = ~n2638 & n2646 ;
  assign n2377 = ~n2373 & ~n2376 ;
  assign n2378 = ~n2342 & n2377 ;
  assign n2385 = n2378 ^ n2373 ;
  assign n2383 = n2381 & ~n2382 ;
  assign n2384 = n2378 & n2383 ;
  assign n2386 = n2385 ^ n2384 ;
  assign n2397 = n2387 & ~n2396 ;
  assign n2398 = ~n2386 & n2397 ;
  assign n2399 = n2398 ^ n2386 ;
  assign n2639 = n2638 ^ n2399 ;
  assign n2648 = n2647 ^ n2639 ;
  assign n3232 = n2667 ^ n2648 ;
  assign n3010 = ~x423 & ~x424 ;
  assign n3014 = x426 ^ x425 ;
  assign n3009 = ~x425 & ~x426 ;
  assign n3015 = n3014 ^ n3009 ;
  assign n3016 = ~n3010 & ~n3015 ;
  assign n3011 = x424 ^ x423 ;
  assign n3012 = n3011 ^ n3010 ;
  assign n3013 = ~n3009 & ~n3012 ;
  assign n3018 = n3016 ^ n3013 ;
  assign n3017 = ~n3013 & ~n3016 ;
  assign n3019 = n3018 ^ n3017 ;
  assign n3031 = x422 ^ x421 ;
  assign n3024 = n3012 ^ n3009 ;
  assign n3025 = n3024 ^ n3013 ;
  assign n3032 = n3025 ^ n3019 ;
  assign n3021 = n3015 ^ n3010 ;
  assign n3022 = n3021 ^ n3016 ;
  assign n3033 = x422 & n3022 ;
  assign n3034 = ~n3032 & n3033 ;
  assign n3035 = n3034 ^ n3017 ;
  assign n3036 = ~n3031 & ~n3035 ;
  assign n3037 = n3036 ^ n3017 ;
  assign n3102 = n3019 & n3037 ;
  assign n3049 = ~x419 & ~x420 ;
  assign n3051 = x416 ^ x415 ;
  assign n3050 = x415 & x416 ;
  assign n3052 = n3051 ^ n3050 ;
  assign n3053 = n3052 ^ x418 ;
  assign n3054 = n3052 ^ x417 ;
  assign n3055 = ~n3053 & ~n3054 ;
  assign n3056 = n3055 ^ n3052 ;
  assign n3057 = x420 ^ x419 ;
  assign n3058 = n3057 ^ n3049 ;
  assign n3059 = n3058 ^ n3050 ;
  assign n3060 = n3058 ^ n3053 ;
  assign n3061 = n3060 ^ n3054 ;
  assign n3062 = ~n3059 & n3061 ;
  assign n3063 = n3062 ^ n3052 ;
  assign n3064 = n3056 & n3063 ;
  assign n3065 = n3064 ^ n3052 ;
  assign n3066 = n3065 ^ n3050 ;
  assign n3067 = ~n3049 & n3066 ;
  assign n3070 = x417 & x418 ;
  assign n3076 = ~n3050 & n3058 ;
  assign n3077 = n3070 & n3076 ;
  assign n3078 = n3077 ^ n3070 ;
  assign n3101 = ~n3067 & ~n3078 ;
  assign n3103 = n3102 ^ n3101 ;
  assign n3068 = x418 ^ x417 ;
  assign n3069 = ~x415 & ~n3068 ;
  assign n3072 = n3068 ^ n3051 ;
  assign n3073 = ~x416 & n3072 ;
  assign n3074 = n3049 & ~n3070 ;
  assign n3075 = n3073 & n3074 ;
  assign n3079 = n3078 ^ n3075 ;
  assign n3071 = ~n3058 & n3070 ;
  assign n3080 = n3079 ^ n3071 ;
  assign n3081 = x419 ^ x418 ;
  assign n3084 = n3081 ^ x420 ;
  assign n3085 = ~x416 & n3084 ;
  assign n3086 = n3085 ^ n3081 ;
  assign n3087 = n3057 & ~n3086 ;
  assign n3088 = n3087 ^ n3081 ;
  assign n3089 = ~n3080 & ~n3088 ;
  assign n3090 = n3069 & n3089 ;
  assign n3091 = n3090 ^ n3080 ;
  assign n3092 = ~n3067 & ~n3091 ;
  assign n3020 = ~x421 & n3019 ;
  assign n3023 = n3022 ^ x422 ;
  assign n3026 = n3025 ^ x422 ;
  assign n3027 = n3023 & n3026 ;
  assign n3028 = n3027 ^ x422 ;
  assign n3029 = n3020 & n3028 ;
  assign n3030 = n3029 ^ x421 ;
  assign n3044 = ~x422 & n3010 ;
  assign n3045 = ~n3025 & n3044 ;
  assign n3046 = n3045 ^ n3025 ;
  assign n3038 = n3037 ^ n3025 ;
  assign n3047 = n3046 ^ n3038 ;
  assign n3048 = n3030 & n3047 ;
  assign n3093 = n3092 ^ n3048 ;
  assign n3094 = n3031 ^ n3014 ;
  assign n3095 = n3094 ^ n3011 ;
  assign n3096 = n3072 ^ n3057 ;
  assign n3097 = n3095 & n3096 ;
  assign n3098 = n3097 ^ n3092 ;
  assign n3099 = ~n3093 & n3098 ;
  assign n3100 = n3099 ^ n3097 ;
  assign n3104 = n3103 ^ n3100 ;
  assign n2985 = ~x427 & ~x428 ;
  assign n2987 = x430 ^ x429 ;
  assign n2986 = ~x429 & ~x430 ;
  assign n2988 = n2987 ^ n2986 ;
  assign n2989 = x432 & ~n2988 ;
  assign n2990 = ~x431 & ~x432 ;
  assign n2991 = ~n2986 & ~n2990 ;
  assign n2992 = x432 ^ x431 ;
  assign n2993 = n2992 ^ n2990 ;
  assign n2994 = n2988 & n2993 ;
  assign n2995 = ~n2991 & n2994 ;
  assign n2996 = x427 & x428 ;
  assign n2997 = ~n2995 & n2996 ;
  assign n2998 = n2997 ^ x431 ;
  assign n2999 = n2989 & n2998 ;
  assign n3000 = n2999 ^ n2997 ;
  assign n3001 = n2994 ^ n2991 ;
  assign n3002 = n3001 ^ n2995 ;
  assign n3003 = ~n3000 & n3002 ;
  assign n3006 = n2985 & n3003 ;
  assign n3004 = n3003 ^ n3000 ;
  assign n3007 = n3006 ^ n3004 ;
  assign n2965 = x436 ^ x435 ;
  assign n2964 = ~x435 & ~x436 ;
  assign n2966 = n2965 ^ n2964 ;
  assign n2962 = x438 ^ x437 ;
  assign n2961 = ~x437 & ~x438 ;
  assign n2963 = n2962 ^ n2961 ;
  assign n2967 = n2966 ^ n2963 ;
  assign n2968 = x434 ^ x433 ;
  assign n2969 = n2968 ^ n2967 ;
  assign n2975 = ~n2961 & ~n2964 ;
  assign n2970 = n2967 ^ x434 ;
  assign n2976 = n2975 ^ n2970 ;
  assign n2977 = ~n2969 & n2976 ;
  assign n2978 = n2977 ^ x433 ;
  assign n2979 = n2978 ^ n2966 ;
  assign n2980 = ~n2967 & ~n2979 ;
  assign n2982 = x433 & x434 ;
  assign n2983 = n2980 & n2982 ;
  assign n2981 = n2980 ^ n2978 ;
  assign n2984 = n2983 ^ n2981 ;
  assign n3008 = n3007 ^ n2984 ;
  assign n3105 = n3104 ^ n3008 ;
  assign n3133 = x437 ^ x434 ;
  assign n3136 = n2964 ^ x437 ;
  assign n3137 = ~n3133 & n3136 ;
  assign n3134 = n3133 ^ n2964 ;
  assign n3135 = x433 & ~n3134 ;
  assign n3138 = n3137 ^ n3135 ;
  assign n3124 = x431 ^ x428 ;
  assign n3127 = n2986 ^ x431 ;
  assign n3128 = ~n3124 & n3127 ;
  assign n3125 = n3124 ^ n2986 ;
  assign n3126 = x427 & n3125 ;
  assign n3129 = n3128 ^ n3126 ;
  assign n3108 = x428 ^ x427 ;
  assign n3109 = n3108 ^ n2987 ;
  assign n3121 = n3109 ^ x431 ;
  assign n3122 = n2988 ^ x432 ;
  assign n3123 = n3121 & n3122 ;
  assign n3130 = n3129 ^ n3123 ;
  assign n3131 = n3130 ^ x433 ;
  assign n3106 = n2968 ^ n2965 ;
  assign n3118 = n3106 ^ x437 ;
  assign n3119 = n2966 ^ x438 ;
  assign n3120 = n3118 & n3119 ;
  assign n3132 = n3131 ^ n3120 ;
  assign n3139 = n3138 ^ n3132 ;
  assign n3107 = n3106 ^ n2962 ;
  assign n3110 = n3109 ^ n2992 ;
  assign n3111 = n3107 & n3110 ;
  assign n3181 = n3130 ^ n3111 ;
  assign n3182 = n3139 & ~n3181 ;
  assign n3183 = n3182 ^ n3130 ;
  assign n3177 = n3097 ^ n3093 ;
  assign n3114 = n3110 ^ n3107 ;
  assign n3115 = n3096 ^ n3095 ;
  assign n3116 = n3114 & n3115 ;
  assign n3197 = n3116 ^ n3097 ;
  assign n3198 = n3197 ^ n3111 ;
  assign n3199 = n3198 ^ n3093 ;
  assign n3200 = n3199 ^ n3139 ;
  assign n3171 = n3200 ^ n3116 ;
  assign n3166 = n3116 ^ n3111 ;
  assign n3167 = n3166 ^ n3139 ;
  assign n3168 = n3167 ^ n3111 ;
  assign n3155 = n3168 & n3199 ;
  assign n3144 = n3116 ^ n3093 ;
  assign n3146 = n3111 ^ n3093 ;
  assign n3148 = n3171 ^ n3146 ;
  assign n3149 = n3144 & ~n3148 ;
  assign n3156 = n3155 ^ n3149 ;
  assign n3157 = n3171 ^ n3156 ;
  assign n3158 = n3155 ^ n3111 ;
  assign n3159 = n3171 ^ n3158 ;
  assign n3160 = n3157 & ~n3159 ;
  assign n3161 = n3160 & n3200 ;
  assign n3162 = n3161 ^ n3155 ;
  assign n3163 = n3168 ^ n3162 ;
  assign n3172 = n3171 ^ n3163 ;
  assign n3178 = n3177 ^ n3172 ;
  assign n3186 = n3183 ^ n3178 ;
  assign n3179 = n2984 & n3007 ;
  assign n3180 = n3178 & ~n3179 ;
  assign n3184 = n3180 & ~n3183 ;
  assign n3185 = n3184 ^ n3179 ;
  assign n3187 = n3186 ^ n3185 ;
  assign n3188 = n3187 ^ n3104 ;
  assign n3189 = n3188 ^ n3185 ;
  assign n3190 = ~n3105 & ~n3189 ;
  assign n3191 = n3190 ^ n3187 ;
  assign n2674 = x460 ^ x459 ;
  assign n2827 = x461 & x462 ;
  assign n2834 = n2827 ^ x460 ;
  assign n2835 = n2674 & ~n2834 ;
  assign n2844 = n2835 ^ x459 ;
  assign n2671 = x462 ^ x461 ;
  assign n2828 = n2827 ^ n2671 ;
  assign n2831 = x458 & n2828 ;
  assign n2823 = x459 & x460 ;
  assign n2836 = n2823 & n2827 ;
  assign n2845 = ~n2831 & ~n2836 ;
  assign n2846 = n2844 & n2845 ;
  assign n2847 = n2846 ^ n2844 ;
  assign n2672 = x458 ^ x457 ;
  assign n2837 = n2836 ^ n2834 ;
  assign n2838 = n2837 ^ n2835 ;
  assign n2851 = n2844 ^ n2838 ;
  assign n2852 = n2851 ^ n2823 ;
  assign n2853 = n2852 ^ n2844 ;
  assign n2856 = x458 & n2853 ;
  assign n2857 = n2856 ^ n2844 ;
  assign n2858 = ~n2672 & n2857 ;
  assign n2859 = n2858 ^ n2844 ;
  assign n2824 = x457 & x458 ;
  assign n2825 = n2823 & n2824 ;
  assign n2860 = n2859 ^ n2825 ;
  assign n2861 = ~x462 & n2860 ;
  assign n2862 = n2861 ^ n2859 ;
  assign n2863 = x461 & ~n2862 ;
  assign n2864 = n2861 & n2863 ;
  assign n2865 = n2864 ^ n2862 ;
  assign n2922 = ~n2847 & ~n2865 ;
  assign n2679 = x454 ^ x453 ;
  assign n2871 = x455 & x456 ;
  assign n2878 = n2871 ^ x454 ;
  assign n2879 = n2679 & ~n2878 ;
  assign n2888 = n2879 ^ x453 ;
  assign n2676 = x456 ^ x455 ;
  assign n2872 = n2871 ^ n2676 ;
  assign n2875 = x452 & n2872 ;
  assign n2867 = x453 & x454 ;
  assign n2880 = n2867 & n2871 ;
  assign n2889 = ~n2875 & ~n2880 ;
  assign n2890 = n2888 & n2889 ;
  assign n2891 = n2890 ^ n2888 ;
  assign n2892 = ~x451 & n2891 ;
  assign n2873 = n2872 ^ x452 ;
  assign n2874 = n2873 ^ x451 ;
  assign n2881 = n2880 ^ n2878 ;
  assign n2882 = n2881 ^ n2879 ;
  assign n2677 = x452 ^ x451 ;
  assign n2876 = n2867 ^ x452 ;
  assign n2877 = ~n2677 & ~n2876 ;
  assign n2883 = n2882 ^ n2877 ;
  assign n2884 = ~n2875 & ~n2883 ;
  assign n2885 = n2874 & n2884 ;
  assign n2887 = n2885 ^ n2877 ;
  assign n2893 = n2892 ^ n2887 ;
  assign n2868 = x451 & x452 ;
  assign n2869 = n2867 & n2868 ;
  assign n2870 = x455 & n2869 ;
  assign n2894 = n2893 ^ n2870 ;
  assign n2895 = n2888 ^ n2882 ;
  assign n2896 = n2895 ^ n2867 ;
  assign n2897 = n2896 ^ n2888 ;
  assign n2900 = x452 & n2897 ;
  assign n2901 = n2900 ^ n2888 ;
  assign n2902 = ~n2677 & n2901 ;
  assign n2903 = n2902 ^ n2888 ;
  assign n2904 = n2903 ^ n2869 ;
  assign n2905 = ~x456 & n2904 ;
  assign n2906 = n2905 ^ n2903 ;
  assign n2907 = x455 & ~n2906 ;
  assign n2908 = n2905 & n2907 ;
  assign n2909 = n2908 ^ n2906 ;
  assign n2910 = ~n2894 & ~n2909 ;
  assign n2848 = ~x457 & n2847 ;
  assign n2829 = n2828 ^ x458 ;
  assign n2830 = n2829 ^ x457 ;
  assign n2832 = n2823 ^ x458 ;
  assign n2833 = ~n2672 & ~n2832 ;
  assign n2839 = n2838 ^ n2833 ;
  assign n2840 = ~n2831 & ~n2839 ;
  assign n2841 = n2830 & n2840 ;
  assign n2843 = n2841 ^ n2833 ;
  assign n2849 = n2848 ^ n2843 ;
  assign n2826 = x461 & n2825 ;
  assign n2850 = n2849 ^ n2826 ;
  assign n2866 = ~n2850 & ~n2865 ;
  assign n2911 = n2910 ^ n2866 ;
  assign n2696 = x444 ^ x443 ;
  assign n2682 = x442 ^ x441 ;
  assign n2816 = n2696 ^ n2682 ;
  assign n2815 = x440 ^ x439 ;
  assign n2817 = n2816 ^ n2815 ;
  assign n2762 = x450 ^ x449 ;
  assign n2748 = x448 ^ x447 ;
  assign n2819 = n2762 ^ n2748 ;
  assign n2818 = x446 ^ x445 ;
  assign n2820 = n2819 ^ n2818 ;
  assign n2821 = n2817 & n2820 ;
  assign n2749 = x448 ^ x446 ;
  assign n2750 = x450 ^ x445 ;
  assign n2753 = ~x448 & ~n2750 ;
  assign n2754 = n2753 ^ x445 ;
  assign n2755 = ~n2749 & n2754 ;
  assign n2756 = ~n2748 & n2755 ;
  assign n2757 = ~x449 & n2756 ;
  assign n2759 = ~x447 & ~x448 ;
  assign n2793 = n2759 ^ x450 ;
  assign n2794 = n2793 ^ n2748 ;
  assign n2795 = n2794 ^ n2759 ;
  assign n2760 = n2759 ^ n2748 ;
  assign n2796 = n2748 ^ x449 ;
  assign n2797 = n2760 & ~n2796 ;
  assign n2798 = n2795 & n2797 ;
  assign n2799 = n2798 ^ n2794 ;
  assign n2758 = x449 & x450 ;
  assign n2774 = n2762 ^ n2758 ;
  assign n2801 = n2799 ^ n2774 ;
  assign n2800 = n2799 ^ x446 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2773 = ~n2758 & n2759 ;
  assign n2775 = n2774 ^ n2773 ;
  assign n2776 = n2775 ^ x449 ;
  assign n2777 = n2793 ^ n2776 ;
  assign n2803 = n2774 ^ n2760 ;
  assign n2804 = n2803 ^ x445 ;
  assign n2805 = ~n2777 & n2804 ;
  assign n2806 = n2802 & n2805 ;
  assign n2807 = n2806 ^ n2801 ;
  assign n2808 = ~x446 & ~n2807 ;
  assign n2809 = n2808 ^ n2799 ;
  assign n2768 = ~x446 & n2774 ;
  assign n2769 = n2803 ^ n2768 ;
  assign n2778 = n2777 ^ n2758 ;
  assign n2779 = n2774 ^ n2768 ;
  assign n2780 = ~n2778 & n2779 ;
  assign n2781 = n2780 ^ n2758 ;
  assign n2782 = ~n2769 & ~n2781 ;
  assign n2761 = n2760 ^ n2758 ;
  assign n2783 = n2782 ^ n2761 ;
  assign n2784 = n2783 ^ n2758 ;
  assign n2785 = n2773 ^ x446 ;
  assign n2788 = n2760 & ~n2785 ;
  assign n2789 = ~n2775 & n2788 ;
  assign n2790 = n2789 ^ n2775 ;
  assign n2791 = n2790 ^ n2774 ;
  assign n2792 = n2784 & ~n2791 ;
  assign n2810 = n2809 ^ n2792 ;
  assign n2811 = ~x445 & n2810 ;
  assign n2812 = n2811 ^ n2809 ;
  assign n2813 = ~n2757 & n2812 ;
  assign n2683 = x442 ^ x440 ;
  assign n2684 = x444 ^ x439 ;
  assign n2687 = ~x442 & ~n2684 ;
  assign n2688 = n2687 ^ x439 ;
  assign n2689 = ~n2683 & n2688 ;
  assign n2690 = ~n2682 & n2689 ;
  assign n2691 = ~x443 & n2690 ;
  assign n2693 = ~x441 & ~x442 ;
  assign n2727 = n2693 ^ x444 ;
  assign n2728 = n2727 ^ n2682 ;
  assign n2729 = n2728 ^ n2693 ;
  assign n2694 = n2693 ^ n2682 ;
  assign n2730 = n2682 ^ x443 ;
  assign n2731 = n2694 & ~n2730 ;
  assign n2732 = n2729 & n2731 ;
  assign n2733 = n2732 ^ n2728 ;
  assign n2692 = x443 & x444 ;
  assign n2708 = n2696 ^ n2692 ;
  assign n2735 = n2733 ^ n2708 ;
  assign n2734 = n2733 ^ x440 ;
  assign n2736 = n2735 ^ n2734 ;
  assign n2707 = ~n2692 & n2693 ;
  assign n2709 = n2708 ^ n2707 ;
  assign n2710 = n2709 ^ x443 ;
  assign n2711 = n2727 ^ n2710 ;
  assign n2737 = n2708 ^ n2694 ;
  assign n2738 = n2737 ^ x439 ;
  assign n2739 = ~n2711 & n2738 ;
  assign n2740 = n2736 & n2739 ;
  assign n2741 = n2740 ^ n2735 ;
  assign n2742 = ~x440 & ~n2741 ;
  assign n2743 = n2742 ^ n2733 ;
  assign n2702 = ~x440 & n2708 ;
  assign n2703 = n2737 ^ n2702 ;
  assign n2712 = n2711 ^ n2692 ;
  assign n2713 = n2708 ^ n2702 ;
  assign n2714 = ~n2712 & n2713 ;
  assign n2715 = n2714 ^ n2692 ;
  assign n2716 = ~n2703 & ~n2715 ;
  assign n2695 = n2694 ^ n2692 ;
  assign n2717 = n2716 ^ n2695 ;
  assign n2718 = n2717 ^ n2692 ;
  assign n2719 = n2707 ^ x440 ;
  assign n2722 = n2694 & ~n2719 ;
  assign n2723 = ~n2709 & n2722 ;
  assign n2724 = n2723 ^ n2709 ;
  assign n2725 = n2724 ^ n2708 ;
  assign n2726 = n2718 & ~n2725 ;
  assign n2744 = n2743 ^ n2726 ;
  assign n2745 = ~x439 & n2744 ;
  assign n2746 = n2745 ^ n2743 ;
  assign n2747 = ~n2691 & n2746 ;
  assign n2814 = n2813 ^ n2747 ;
  assign n2822 = n2821 ^ n2814 ;
  assign n2912 = n2911 ^ n2822 ;
  assign n2678 = n2677 ^ n2676 ;
  assign n2680 = n2679 ^ n2678 ;
  assign n2673 = n2672 ^ n2671 ;
  assign n2675 = n2674 ^ n2673 ;
  assign n2913 = n2680 ^ n2675 ;
  assign n2914 = n2820 ^ n2817 ;
  assign n2915 = n2913 & n2914 ;
  assign n2917 = n2915 ^ n2911 ;
  assign n2920 = n2912 & ~n2917 ;
  assign n2681 = n2675 & n2680 ;
  assign n2919 = ~n2681 & n2822 ;
  assign n2921 = n2920 ^ n2919 ;
  assign n2923 = n2922 ^ n2921 ;
  assign n2924 = ~n2891 & ~n2909 ;
  assign n2925 = n2924 ^ n2922 ;
  assign n2926 = n2923 & n2925 ;
  assign n2927 = n2926 ^ n2924 ;
  assign n2940 = n2910 ^ n2681 ;
  assign n2941 = ~n2911 & n2940 ;
  assign n2942 = n2941 ^ n2681 ;
  assign n2931 = x445 & ~n2809 ;
  assign n2937 = n2784 & n2931 ;
  assign n2932 = x439 & n2718 ;
  assign n2933 = ~n2743 & n2932 ;
  assign n2934 = n2933 ^ n2718 ;
  assign n2935 = n2934 ^ n2784 ;
  assign n2938 = n2937 ^ n2935 ;
  assign n2928 = n2821 ^ n2747 ;
  assign n2929 = ~n2814 & n2928 ;
  assign n2930 = n2929 ^ n2821 ;
  assign n2939 = n2938 ^ n2930 ;
  assign n2943 = n2942 ^ n2939 ;
  assign n2944 = n2942 ^ n2924 ;
  assign n2945 = n2944 ^ n2939 ;
  assign n2946 = n2945 ^ n2923 ;
  assign n2947 = n2946 ^ n2939 ;
  assign n2948 = n2943 & ~n2947 ;
  assign n2949 = n2948 ^ n2939 ;
  assign n2950 = n2927 & ~n2949 ;
  assign n2951 = n2934 ^ n2930 ;
  assign n2952 = ~n2938 & ~n2951 ;
  assign n2953 = n2952 ^ n2930 ;
  assign n2954 = n2939 & ~n2946 ;
  assign n2955 = ~n2927 & n2954 ;
  assign n2956 = ~n2953 & ~n2955 ;
  assign n2957 = ~n2950 & n2956 ;
  assign n2958 = n2957 ^ n2950 ;
  assign n3223 = n3185 ^ n2958 ;
  assign n3192 = n3102 ^ n3100 ;
  assign n3193 = n3103 & ~n3192 ;
  assign n3194 = n3193 ^ n3102 ;
  assign n3224 = n3223 ^ n3194 ;
  assign n3225 = n3224 ^ n2958 ;
  assign n3226 = ~n3191 & ~n3225 ;
  assign n3227 = n3226 ^ n3223 ;
  assign n3195 = n3194 ^ n3191 ;
  assign n2959 = n2955 ^ n2950 ;
  assign n2960 = n2959 ^ n2953 ;
  assign n3196 = n3195 ^ n2960 ;
  assign n3201 = n3115 ^ n3114 ;
  assign n3202 = n2914 ^ n2913 ;
  assign n3203 = n3201 & n3202 ;
  assign n3204 = n3203 ^ n3200 ;
  assign n3207 = n2821 ^ n2681 ;
  assign n3208 = n3207 ^ n2915 ;
  assign n3209 = n3208 ^ n2814 ;
  assign n3210 = n3209 ^ n2911 ;
  assign n3205 = n3186 ^ n3105 ;
  assign n3206 = n3205 ^ n3203 ;
  assign n3211 = n3210 ^ n3206 ;
  assign n3212 = n3211 ^ n3205 ;
  assign n3213 = n3204 & n3212 ;
  assign n3214 = n3213 ^ n3206 ;
  assign n3216 = n3195 ^ n2946 ;
  assign n3215 = n3205 ^ n3195 ;
  assign n3217 = n3216 ^ n3215 ;
  assign n3218 = ~n3214 & ~n3217 ;
  assign n3219 = n3218 ^ n3215 ;
  assign n3220 = ~n3196 & ~n3219 ;
  assign n3221 = n3220 ^ n3195 ;
  assign n3231 = n3227 ^ n3221 ;
  assign n3233 = n3232 ^ n3231 ;
  assign n3249 = n3219 ^ n2960 ;
  assign n3235 = n3214 ^ n2946 ;
  assign n3234 = n2660 ^ n2371 ;
  assign n3236 = n3235 ^ n3234 ;
  assign n3238 = n3210 ^ n3204 ;
  assign n3245 = n3238 ^ n3235 ;
  assign n3237 = n2656 ^ n2597 ;
  assign n3239 = n3238 ^ n3237 ;
  assign n3240 = n3202 ^ n3201 ;
  assign n3241 = n2654 ^ n2653 ;
  assign n3242 = n3240 & n3241 ;
  assign n3243 = n3242 ^ n3238 ;
  assign n3244 = n3239 & n3243 ;
  assign n3246 = n3245 ^ n3244 ;
  assign n3247 = n3236 & ~n3246 ;
  assign n3248 = n3247 ^ n3235 ;
  assign n3250 = n3249 ^ n3248 ;
  assign n3251 = n2665 ^ n2650 ;
  assign n3252 = n3251 ^ n3248 ;
  assign n3253 = n3250 & n3252 ;
  assign n3254 = n3253 ^ n3251 ;
  assign n3255 = n3254 ^ n3232 ;
  assign n3256 = ~n3233 & n3255 ;
  assign n3257 = n3256 ^ n3254 ;
  assign n3222 = n3221 ^ n2958 ;
  assign n3228 = ~n3222 & n3227 ;
  assign n3229 = n3228 ^ n3221 ;
  assign n3293 = n3257 ^ n3229 ;
  assign n2668 = n2667 ^ n2399 ;
  assign n2669 = n2648 & n2668 ;
  assign n2670 = n2669 ^ n2399 ;
  assign n3294 = n3257 ^ n2670 ;
  assign n3295 = n3293 & n3294 ;
  assign n3296 = n3295 ^ n2670 ;
  assign n3261 = n3254 ^ n3233 ;
  assign n2142 = n2128 ^ n2110 ;
  assign n3259 = n2142 ^ n2112 ;
  assign n2136 = n2072 ^ n1221 ;
  assign n2137 = n2136 ^ n2114 ;
  assign n3260 = n3259 ^ n2137 ;
  assign n3262 = n3261 ^ n3260 ;
  assign n3279 = n3246 ^ n3234 ;
  assign n3269 = n3268 ^ n1977 ;
  assign n3264 = n3241 ^ n3240 ;
  assign n3265 = n1974 ^ n1973 ;
  assign n3266 = n3264 & n3265 ;
  assign n3270 = n3269 ^ n3266 ;
  assign n5735 = n3266 ^ n3242 ;
  assign n5736 = n5735 ^ n3239 ;
  assign n3277 = n3270 & ~n5736 ;
  assign n3278 = n3277 ^ n3269 ;
  assign n3280 = n3279 ^ n3278 ;
  assign n3281 = n1983 ^ n1512 ;
  assign n3282 = n3281 ^ n3278 ;
  assign n3283 = ~n3280 & ~n3282 ;
  assign n3284 = n3283 ^ n3281 ;
  assign n3289 = n3284 ^ n3261 ;
  assign n3263 = n3251 ^ n3250 ;
  assign n3285 = n3284 ^ n3263 ;
  assign n3286 = n2069 ^ n2014 ;
  assign n3287 = n3286 ^ n3284 ;
  assign n3288 = ~n3285 & ~n3287 ;
  assign n3290 = n3289 ^ n3288 ;
  assign n3291 = n3262 & n3290 ;
  assign n3292 = n3291 ^ n3261 ;
  assign n3299 = n3296 ^ n3292 ;
  assign n3230 = n2670 & ~n3229 ;
  assign n3258 = n3230 & n3257 ;
  assign n3297 = n3292 & n3296 ;
  assign n3298 = ~n3258 & n3297 ;
  assign n3300 = n3299 ^ n3298 ;
  assign n2143 = ~n2072 & ~n2142 ;
  assign n2144 = ~n2112 & n2143 ;
  assign n2146 = ~n1221 & ~n2110 ;
  assign n2149 = ~n2072 & n2146 ;
  assign n2145 = n2143 ^ n2072 ;
  assign n2147 = n2146 ^ n2145 ;
  assign n2148 = ~n2080 & ~n2147 ;
  assign n2150 = n2149 ^ n2148 ;
  assign n2151 = n2150 ^ n2149 ;
  assign n2152 = n2144 & n2151 ;
  assign n2153 = n2152 ^ n2150 ;
  assign n3301 = n2153 ^ n2149 ;
  assign n3302 = n3301 ^ n2153 ;
  assign n3303 = n3302 ^ n1221 ;
  assign n3304 = n3303 ^ n3302 ;
  assign n3305 = n3302 ^ n2128 ;
  assign n3306 = n3305 ^ n3302 ;
  assign n3307 = ~n3304 & n3306 ;
  assign n3308 = n3307 ^ n3302 ;
  assign n3309 = n2080 & n3308 ;
  assign n3310 = n3309 ^ n3301 ;
  assign n3311 = ~n2064 & n3310 ;
  assign n3312 = n3311 ^ n2153 ;
  assign n3313 = n2080 & n2112 ;
  assign n3314 = n2146 & n3313 ;
  assign n3317 = n3314 ^ n2072 ;
  assign n3318 = n3317 ^ n3314 ;
  assign n3315 = n3314 ^ n2112 ;
  assign n3319 = n3314 ^ n2064 ;
  assign n3320 = n3319 ^ n3314 ;
  assign n3323 = n3315 & ~n3320 ;
  assign n3324 = n3318 & n3323 ;
  assign n3325 = n3324 ^ n3318 ;
  assign n3326 = n3325 ^ n3317 ;
  assign n3327 = ~n3312 & ~n3326 ;
  assign n3328 = ~n2135 & n3327 ;
  assign n3330 = n3229 ^ n2670 ;
  assign n3331 = n3330 ^ n3257 ;
  assign n2138 = n2137 ^ n2104 ;
  assign n2139 = n2137 ^ n2109 ;
  assign n2140 = n2138 & n2139 ;
  assign n2141 = n2140 ^ n2104 ;
  assign n2154 = n2064 & n2153 ;
  assign n2155 = n2141 & n2154 ;
  assign n2156 = n2155 ^ n2141 ;
  assign n2157 = ~n2135 & n2156 ;
  assign n3329 = n3258 ^ n2157 ;
  assign n3332 = n3331 ^ n3329 ;
  assign n3333 = n3332 ^ n3296 ;
  assign n3334 = ~n3328 & ~n3333 ;
  assign n3335 = n3300 & n3334 ;
  assign n5760 = ~n2135 & ~n3335 ;
  assign n5761 = n3297 ^ n2156 ;
  assign n5764 = ~n3327 & ~n5761 ;
  assign n5765 = n5764 ^ n3297 ;
  assign n5766 = ~n3258 & ~n5765 ;
  assign n5767 = n5766 ^ n2156 ;
  assign n5768 = n5760 & n5767 ;
  assign n5769 = n5768 ^ n3335 ;
  assign n5725 = n5711 ^ n5680 ;
  assign n5723 = n3328 ^ n3292 ;
  assign n5724 = n5723 ^ n3331 ;
  assign n5726 = n5725 ^ n5724 ;
  assign n5730 = n3290 ^ n3260 ;
  assign n5727 = n5708 ^ n5660 ;
  assign n5728 = n5727 ^ n5681 ;
  assign n5731 = n5730 ^ n5728 ;
  assign n5733 = n5705 ^ n5704 ;
  assign n5732 = n3286 ^ n3285 ;
  assign n5734 = n5733 ^ n5732 ;
  assign n5747 = n3281 ^ n3280 ;
  assign n5738 = n5695 ^ n5691 ;
  assign n5737 = n5736 ^ n3269 ;
  assign n5739 = n5738 ^ n5737 ;
  assign n5740 = n3265 ^ n3264 ;
  assign n5741 = n5687 ^ n5686 ;
  assign n5742 = n5740 & n5741 ;
  assign n5743 = n5742 ^ n5738 ;
  assign n5744 = ~n5739 & ~n5743 ;
  assign n5745 = n5744 ^ n5738 ;
  assign n5748 = n5747 ^ n5745 ;
  assign n5749 = n5700 ^ n5683 ;
  assign n5750 = n5749 ^ n5745 ;
  assign n5751 = n5748 & ~n5750 ;
  assign n5746 = n5745 ^ n5733 ;
  assign n5752 = n5751 ^ n5746 ;
  assign n5753 = n5734 & n5752 ;
  assign n5754 = n5753 ^ n5733 ;
  assign n5755 = n5754 ^ n5728 ;
  assign n5756 = ~n5731 & ~n5755 ;
  assign n5729 = n5728 ^ n5725 ;
  assign n5757 = n5756 ^ n5729 ;
  assign n5758 = ~n5726 & ~n5757 ;
  assign n5759 = n5758 ^ n5725 ;
  assign n5770 = n5769 ^ n5759 ;
  assign n8726 = n8725 ^ n5770 ;
  assign n6395 = x76 ^ x75 ;
  assign n6393 = x74 ^ x73 ;
  assign n6430 = n6395 ^ n6393 ;
  assign n6389 = x78 ^ x77 ;
  assign n6431 = n6430 ^ n6389 ;
  assign n6352 = x70 ^ x69 ;
  assign n6350 = x68 ^ x67 ;
  assign n6428 = n6352 ^ n6350 ;
  assign n6346 = x72 ^ x71 ;
  assign n6429 = n6428 ^ n6346 ;
  assign n6843 = n6431 ^ n6429 ;
  assign n6464 = x56 ^ x55 ;
  assign n6455 = x58 ^ x57 ;
  assign n6522 = n6464 ^ n6455 ;
  assign n6458 = x60 ^ x59 ;
  assign n6523 = n6522 ^ n6458 ;
  assign n6495 = x64 ^ x63 ;
  assign n6494 = x62 ^ x61 ;
  assign n6520 = n6495 ^ n6494 ;
  assign n6498 = x66 ^ x65 ;
  assign n6521 = n6520 ^ n6498 ;
  assign n6531 = n6523 ^ n6521 ;
  assign n6844 = n6843 ^ n6531 ;
  assign n6608 = x40 ^ x39 ;
  assign n6607 = x38 ^ x37 ;
  assign n6609 = n6608 ^ n6607 ;
  assign n6606 = x42 ^ x41 ;
  assign n6610 = n6609 ^ n6606 ;
  assign n6642 = x35 ^ x33 ;
  assign n6654 = n6642 ^ x34 ;
  assign n6655 = n6654 ^ x36 ;
  assign n6600 = x32 ^ x31 ;
  assign n6604 = n6655 ^ n6600 ;
  assign n6845 = n6610 ^ n6604 ;
  assign n6597 = x54 ^ x53 ;
  assign n6595 = x52 ^ x51 ;
  assign n6594 = x50 ^ x49 ;
  assign n6596 = n6595 ^ n6594 ;
  assign n6598 = n6597 ^ n6596 ;
  assign n6591 = x46 ^ x45 ;
  assign n6590 = x44 ^ x43 ;
  assign n6592 = n6591 ^ n6590 ;
  assign n6589 = x48 ^ x47 ;
  assign n6593 = n6592 ^ n6589 ;
  assign n6612 = n6598 ^ n6593 ;
  assign n6846 = n6845 ^ n6612 ;
  assign n6847 = n6844 & n6846 ;
  assign n6532 = n6531 ^ n6431 ;
  assign n6524 = n6521 & n6523 ;
  assign n6500 = ~x63 & ~x64 ;
  assign n6501 = n6500 ^ n6495 ;
  assign n6496 = x65 & x66 ;
  assign n6499 = n6498 ^ n6496 ;
  assign n6505 = n6501 ^ n6499 ;
  assign n6502 = n6499 & ~n6501 ;
  assign n6506 = n6505 ^ n6502 ;
  assign n6510 = n6506 ^ x62 ;
  assign n6507 = n6500 ^ n6496 ;
  assign n6497 = n6495 & n6496 ;
  assign n6508 = n6507 ^ n6497 ;
  assign n6511 = n6510 ^ n6508 ;
  assign n6512 = n6494 & ~n6511 ;
  assign n6513 = n6512 ^ x61 ;
  assign n6509 = ~n6506 & ~n6508 ;
  assign n6515 = n6513 ^ n6509 ;
  assign n6514 = ~n6509 & ~n6513 ;
  assign n6516 = n6515 ^ n6514 ;
  assign n6503 = n6502 ^ n6497 ;
  assign n6504 = n6494 & n6503 ;
  assign n6517 = n6516 ^ n6504 ;
  assign n6518 = n6517 ^ n6514 ;
  assign n6454 = ~x57 & ~x58 ;
  assign n6453 = ~x59 & ~x60 ;
  assign n6459 = n6458 ^ n6453 ;
  assign n6460 = ~n6454 & ~n6459 ;
  assign n6456 = n6455 ^ n6454 ;
  assign n6457 = ~n6453 & ~n6456 ;
  assign n6462 = n6460 ^ n6457 ;
  assign n6461 = ~n6457 & ~n6460 ;
  assign n6463 = n6462 ^ n6461 ;
  assign n6476 = ~x55 & n6463 ;
  assign n6468 = n6459 ^ n6454 ;
  assign n6469 = n6468 ^ n6460 ;
  assign n6477 = n6469 ^ x56 ;
  assign n6465 = n6456 ^ n6453 ;
  assign n6466 = n6465 ^ n6457 ;
  assign n6478 = n6466 ^ x56 ;
  assign n6479 = n6477 & n6478 ;
  assign n6480 = n6479 ^ x56 ;
  assign n6481 = n6476 & n6480 ;
  assign n6482 = n6481 ^ x55 ;
  assign n6489 = ~x56 & n6454 ;
  assign n6490 = ~n6466 & n6489 ;
  assign n6491 = n6490 ^ n6466 ;
  assign n6467 = n6466 ^ n6463 ;
  assign n6470 = x56 & n6469 ;
  assign n6471 = ~n6467 & n6470 ;
  assign n6472 = n6471 ^ n6461 ;
  assign n6473 = ~n6464 & ~n6472 ;
  assign n6474 = n6473 ^ n6461 ;
  assign n6483 = n6474 ^ n6466 ;
  assign n6492 = n6491 ^ n6483 ;
  assign n6493 = n6482 & n6492 ;
  assign n6519 = n6518 ^ n6493 ;
  assign n6529 = n6524 ^ n6519 ;
  assign n6533 = n6529 ^ n6429 ;
  assign n6534 = n6533 ^ n6531 ;
  assign n6535 = n6534 ^ n6529 ;
  assign n6536 = ~n6532 & n6535 ;
  assign n6537 = n6536 ^ n6533 ;
  assign n6385 = x77 ^ x76 ;
  assign n6390 = ~n6385 & ~n6389 ;
  assign n6384 = x75 ^ x74 ;
  assign n6386 = n6385 ^ x75 ;
  assign n6387 = n6386 ^ x78 ;
  assign n6388 = ~n6384 & n6387 ;
  assign n6391 = n6390 ^ n6388 ;
  assign n6392 = ~x73 & n6391 ;
  assign n6394 = ~x75 & ~x76 ;
  assign n6401 = ~x77 & ~x78 ;
  assign n6402 = ~n6394 & ~n6401 ;
  assign n6396 = n6395 ^ n6394 ;
  assign n6397 = x73 & x74 ;
  assign n6398 = x78 & n6397 ;
  assign n6399 = ~n6396 & n6398 ;
  assign n6400 = n6399 ^ n6397 ;
  assign n6403 = n6402 ^ n6400 ;
  assign n6406 = n6401 ^ n6389 ;
  assign n6409 = n6396 & n6406 ;
  assign n6410 = n6409 ^ n6400 ;
  assign n6411 = n6403 & ~n6410 ;
  assign n6412 = n6411 ^ n6400 ;
  assign n6413 = ~n6393 & n6412 ;
  assign n6414 = n6411 & n6413 ;
  assign n6415 = n6414 ^ n6412 ;
  assign n6416 = x76 ^ x74 ;
  assign n6417 = x78 ^ x73 ;
  assign n6420 = ~x76 & ~n6417 ;
  assign n6421 = n6420 ^ x73 ;
  assign n6422 = ~n6416 & n6421 ;
  assign n6423 = ~n6395 & n6422 ;
  assign n6424 = ~x77 & n6423 ;
  assign n6425 = ~n6415 & ~n6424 ;
  assign n6426 = ~n6392 & n6425 ;
  assign n6342 = x71 ^ x70 ;
  assign n6347 = ~n6342 & ~n6346 ;
  assign n6341 = x69 ^ x68 ;
  assign n6343 = n6342 ^ x69 ;
  assign n6344 = n6343 ^ x72 ;
  assign n6345 = ~n6341 & n6344 ;
  assign n6348 = n6347 ^ n6345 ;
  assign n6349 = ~x67 & n6348 ;
  assign n6351 = ~x69 & ~x70 ;
  assign n6358 = ~x71 & ~x72 ;
  assign n6359 = ~n6351 & ~n6358 ;
  assign n6353 = n6352 ^ n6351 ;
  assign n6354 = x67 & x68 ;
  assign n6355 = x72 & n6354 ;
  assign n6356 = ~n6353 & n6355 ;
  assign n6357 = n6356 ^ n6354 ;
  assign n6360 = n6359 ^ n6357 ;
  assign n6363 = n6358 ^ n6346 ;
  assign n6366 = n6353 & n6363 ;
  assign n6367 = n6366 ^ n6357 ;
  assign n6368 = n6360 & ~n6367 ;
  assign n6369 = n6368 ^ n6357 ;
  assign n6370 = ~n6350 & n6369 ;
  assign n6371 = n6368 & n6370 ;
  assign n6372 = n6371 ^ n6369 ;
  assign n6373 = x70 ^ x68 ;
  assign n6374 = x72 ^ x67 ;
  assign n6377 = ~x70 & ~n6374 ;
  assign n6378 = n6377 ^ x67 ;
  assign n6379 = ~n6373 & n6378 ;
  assign n6380 = ~n6352 & n6379 ;
  assign n6381 = ~x71 & n6380 ;
  assign n6382 = ~n6372 & ~n6381 ;
  assign n6383 = ~n6349 & n6382 ;
  assign n6427 = n6426 ^ n6383 ;
  assign n6538 = n6537 ^ n6427 ;
  assign n6848 = n6847 ^ n6538 ;
  assign n6740 = x53 & x54 ;
  assign n6739 = x51 & x52 ;
  assign n6741 = n6740 ^ n6739 ;
  assign n6742 = n6740 ^ n6597 ;
  assign n6743 = n6739 ^ n6595 ;
  assign n6744 = n6742 & n6743 ;
  assign n6745 = n6744 ^ n6740 ;
  assign n6746 = ~n6741 & ~n6745 ;
  assign n6691 = n6597 ^ x50 ;
  assign n6692 = n6691 ^ n6595 ;
  assign n6694 = x47 ^ x46 ;
  assign n6698 = ~n6589 & ~n6694 ;
  assign n6693 = x45 ^ x44 ;
  assign n6695 = n6694 ^ x45 ;
  assign n6696 = n6695 ^ x48 ;
  assign n6697 = ~n6693 & n6696 ;
  assign n6699 = n6698 ^ n6697 ;
  assign n6700 = ~x43 & n6699 ;
  assign n6701 = ~x45 & ~x46 ;
  assign n6707 = ~x47 & ~x48 ;
  assign n6708 = ~n6701 & ~n6707 ;
  assign n6702 = n6701 ^ n6591 ;
  assign n6703 = x43 & x44 ;
  assign n6704 = x48 & n6703 ;
  assign n6705 = ~n6702 & n6704 ;
  assign n6706 = n6705 ^ n6703 ;
  assign n6709 = n6708 ^ n6706 ;
  assign n6712 = n6707 ^ n6589 ;
  assign n6715 = n6702 & n6712 ;
  assign n6716 = n6715 ^ n6706 ;
  assign n6717 = n6709 & ~n6716 ;
  assign n6718 = n6717 ^ n6706 ;
  assign n6719 = ~n6590 & n6718 ;
  assign n6720 = n6717 & n6719 ;
  assign n6721 = n6720 ^ n6718 ;
  assign n6722 = x46 ^ x44 ;
  assign n6723 = x48 ^ x43 ;
  assign n6726 = ~x46 & ~n6723 ;
  assign n6727 = n6726 ^ x43 ;
  assign n6728 = ~n6722 & n6727 ;
  assign n6729 = ~n6591 & n6728 ;
  assign n6730 = ~x47 & n6729 ;
  assign n6731 = ~n6721 & ~n6730 ;
  assign n6732 = ~n6700 & n6731 ;
  assign n6733 = n6732 ^ x49 ;
  assign n6734 = n6733 ^ n6597 ;
  assign n6735 = n6734 ^ n6595 ;
  assign n6736 = n6735 ^ n6732 ;
  assign n6737 = ~n6692 & n6736 ;
  assign n6738 = n6737 ^ n6733 ;
  assign n6747 = n6746 ^ n6738 ;
  assign n6683 = x37 & x38 ;
  assign n6684 = n6683 ^ n6608 ;
  assign n6682 = ~x41 & ~x42 ;
  assign n6685 = n6684 ^ n6682 ;
  assign n6681 = ~x39 & ~x40 ;
  assign n6686 = n6685 ^ n6681 ;
  assign n6624 = x35 & x36 ;
  assign n6627 = ~x33 & ~x34 ;
  assign n6602 = x34 ^ x33 ;
  assign n6635 = n6627 ^ n6602 ;
  assign n6636 = ~n6624 & n6635 ;
  assign n6644 = x35 ^ x32 ;
  assign n6645 = n6644 ^ x34 ;
  assign n6646 = n6645 ^ x36 ;
  assign n6647 = n6646 ^ n6642 ;
  assign n6648 = n6647 ^ x36 ;
  assign n6649 = n6648 ^ x35 ;
  assign n6650 = n6649 ^ n6642 ;
  assign n6656 = n6655 ^ n6642 ;
  assign n6657 = ~n6650 & ~n6656 ;
  assign n6658 = ~x35 & n6657 ;
  assign n6661 = n6658 ^ n6657 ;
  assign n6659 = n6658 ^ n6642 ;
  assign n6660 = n6647 & n6659 ;
  assign n6662 = n6661 ^ n6660 ;
  assign n6663 = n6662 ^ x35 ;
  assign n6674 = x31 & n6663 ;
  assign n6664 = n6663 ^ x31 ;
  assign n6675 = n6674 ^ n6664 ;
  assign n6678 = n6636 & ~n6675 ;
  assign n6637 = n6635 ^ n6624 ;
  assign n6601 = x36 ^ x35 ;
  assign n6625 = n6624 ^ n6601 ;
  assign n6626 = n6625 ^ x32 ;
  assign n6628 = n6627 ^ n6626 ;
  assign n6638 = n6635 ^ n6628 ;
  assign n6630 = ~n6625 & n6627 ;
  assign n6629 = n6627 ^ n6625 ;
  assign n6631 = n6630 ^ n6629 ;
  assign n6632 = ~n6628 & ~n6631 ;
  assign n6639 = n6638 ^ n6632 ;
  assign n6640 = ~n6637 & ~n6639 ;
  assign n6641 = n6640 ^ n6624 ;
  assign n6665 = n6664 ^ n6641 ;
  assign n6666 = n6665 ^ n6663 ;
  assign n6670 = ~n6641 & ~n6662 ;
  assign n6671 = n6670 ^ x35 ;
  assign n6672 = ~n6666 & ~n6671 ;
  assign n6673 = n6672 ^ n6664 ;
  assign n6676 = n6675 ^ n6673 ;
  assign n6679 = n6678 ^ n6676 ;
  assign n6633 = n6630 ^ x31 ;
  assign n6634 = ~n6632 & ~n6633 ;
  assign n6680 = n6679 ^ n6634 ;
  assign n6687 = n6686 ^ n6680 ;
  assign n6622 = n6607 ^ n6606 ;
  assign n6623 = ~n6609 & n6622 ;
  assign n6688 = n6687 ^ n6623 ;
  assign n6605 = n6604 ^ n6593 ;
  assign n6611 = n6610 ^ n6605 ;
  assign n6613 = ~n6605 & ~n6612 ;
  assign n6614 = n6611 & n6613 ;
  assign n6615 = n6614 ^ n6610 ;
  assign n6618 = n6604 & n6610 ;
  assign n6619 = n6618 ^ n6613 ;
  assign n6616 = n6612 ^ n6604 ;
  assign n6617 = ~n6615 & n6616 ;
  assign n6620 = n6619 ^ n6617 ;
  assign n6621 = ~n6615 & n6620 ;
  assign n6689 = n6688 ^ n6621 ;
  assign n6748 = n6747 ^ n6689 ;
  assign n6849 = n6748 ^ n6538 ;
  assign n6850 = n6848 & ~n6849 ;
  assign n6851 = n6850 ^ n6538 ;
  assign n6811 = n6681 ^ n6608 ;
  assign n6823 = x42 & n6683 ;
  assign n6824 = ~n6811 & n6823 ;
  assign n6825 = n6824 ^ n6683 ;
  assign n6814 = ~n6681 & ~n6682 ;
  assign n6826 = n6825 ^ n6814 ;
  assign n6812 = n6682 ^ n6606 ;
  assign n6831 = n6811 & n6812 ;
  assign n6832 = n6831 ^ n6825 ;
  assign n6833 = n6826 & ~n6832 ;
  assign n6813 = n6812 ^ n6811 ;
  assign n6819 = x38 & n6814 ;
  assign n6820 = n6819 ^ n6811 ;
  assign n6821 = n6813 & n6820 ;
  assign n6822 = n6821 ^ n6812 ;
  assign n6834 = n6833 ^ n6825 ;
  assign n6835 = n6822 & n6834 ;
  assign n6836 = ~n6607 & n6835 ;
  assign n6837 = n6833 & n6836 ;
  assign n6838 = n6837 ^ n6835 ;
  assign n6839 = n6838 ^ n6822 ;
  assign n6805 = ~n6641 & ~n6674 ;
  assign n6806 = n6805 ^ n6680 ;
  assign n6807 = n6806 ^ n6618 ;
  assign n6808 = n6807 ^ n6805 ;
  assign n6809 = ~n6688 & ~n6808 ;
  assign n6810 = n6809 ^ n6806 ;
  assign n6840 = n6839 ^ n6810 ;
  assign n6599 = n6593 & n6598 ;
  assign n6800 = n6732 ^ n6599 ;
  assign n6801 = ~n6747 & n6800 ;
  assign n6802 = n6801 ^ n6732 ;
  assign n6767 = n6739 ^ x49 ;
  assign n6770 = n6767 ^ n6741 ;
  assign n6765 = n6739 ^ x50 ;
  assign n6775 = n6770 ^ n6765 ;
  assign n6766 = n6745 ^ n6741 ;
  assign n6768 = n6767 ^ n6766 ;
  assign n6776 = n6775 ^ n6768 ;
  assign n6777 = n6776 ^ n6741 ;
  assign n6779 = n6775 & n6777 ;
  assign n6772 = n6768 ^ n6741 ;
  assign n6773 = n6772 ^ n6740 ;
  assign n6774 = ~n6744 & n6773 ;
  assign n6780 = n6779 ^ n6774 ;
  assign n6781 = n6780 ^ n6772 ;
  assign n6782 = n6779 ^ n6770 ;
  assign n6783 = n6782 ^ n6772 ;
  assign n6784 = n6781 & n6783 ;
  assign n6785 = ~n6741 & n6784 ;
  assign n6786 = n6785 ^ n6779 ;
  assign n6787 = n6786 ^ n6777 ;
  assign n6795 = n6787 ^ n6739 ;
  assign n6798 = n6795 ^ n6765 ;
  assign n6759 = n6712 ^ n6702 ;
  assign n6760 = x44 & n6708 ;
  assign n6761 = n6760 ^ n6702 ;
  assign n6762 = n6759 & ~n6761 ;
  assign n6763 = n6762 ^ n6702 ;
  assign n6764 = ~n6721 & n6763 ;
  assign n6799 = n6798 ^ n6764 ;
  assign n6803 = n6802 ^ n6799 ;
  assign n6690 = n6689 ^ n6599 ;
  assign n6750 = n6690 & ~n6747 ;
  assign n6751 = n6750 ^ n6689 ;
  assign n6756 = n6620 & n6688 ;
  assign n6757 = n6756 ^ n6618 ;
  assign n6758 = ~n6751 & ~n6757 ;
  assign n6804 = n6803 ^ n6758 ;
  assign n6841 = n6840 ^ n6804 ;
  assign n6558 = n6496 & ~n6501 ;
  assign n6559 = n6517 & n6558 ;
  assign n6560 = n6559 ^ n6517 ;
  assign n6475 = n6463 & n6474 ;
  assign n6576 = n6560 ^ n6475 ;
  assign n6525 = n6524 ^ n6518 ;
  assign n6526 = n6519 & n6525 ;
  assign n6527 = n6526 ^ n6518 ;
  assign n6577 = n6576 ^ n6527 ;
  assign n6444 = n6363 ^ n6353 ;
  assign n6445 = x68 & n6359 ;
  assign n6446 = n6445 ^ n6353 ;
  assign n6447 = n6444 & ~n6446 ;
  assign n6448 = n6447 ^ n6353 ;
  assign n6449 = ~n6372 & n6448 ;
  assign n6436 = n6406 ^ n6396 ;
  assign n6437 = x74 & n6402 ;
  assign n6438 = n6437 ^ n6396 ;
  assign n6439 = n6436 & ~n6438 ;
  assign n6440 = n6439 ^ n6396 ;
  assign n6441 = ~n6415 & ~n6440 ;
  assign n6442 = n6441 ^ n6415 ;
  assign n6450 = n6449 ^ n6442 ;
  assign n6432 = n6429 & n6431 ;
  assign n6433 = n6432 ^ n6383 ;
  assign n6434 = n6427 & ~n6433 ;
  assign n6435 = n6434 ^ n6426 ;
  assign n6555 = n6450 ^ n6435 ;
  assign n6578 = n6577 ^ n6555 ;
  assign n6540 = n6432 ^ n6427 ;
  assign n6539 = n6538 ^ n6524 ;
  assign n6541 = n6540 ^ n6539 ;
  assign n6542 = ~n6519 & ~n6541 ;
  assign n6543 = n6542 ^ n6524 ;
  assign n6544 = n6540 ^ n6537 ;
  assign n6545 = n6542 ^ n6541 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = n6546 ^ n6537 ;
  assign n6548 = n6547 ^ n6544 ;
  assign n6549 = n6543 & n6548 ;
  assign n6550 = n6549 ^ n6546 ;
  assign n6551 = n6550 ^ n6540 ;
  assign n6579 = n6578 ^ n6551 ;
  assign n6842 = n6841 ^ n6579 ;
  assign n7139 = n6851 ^ n6842 ;
  assign n6961 = x22 ^ x21 ;
  assign n7096 = ~x21 & ~x22 ;
  assign n7097 = ~x23 & ~x24 ;
  assign n7098 = ~n7096 & ~n7097 ;
  assign n7099 = n7098 ^ x20 ;
  assign n7100 = n7096 ^ n6961 ;
  assign n6963 = x24 ^ x23 ;
  assign n7101 = n7097 ^ n6963 ;
  assign n7102 = n7100 & n7101 ;
  assign n7103 = n7102 ^ x20 ;
  assign n7104 = n7099 & ~n7103 ;
  assign n7105 = n7104 ^ x20 ;
  assign n7106 = x19 & ~n7105 ;
  assign n7107 = n7106 ^ x19 ;
  assign n7108 = n7107 ^ x23 ;
  assign n7109 = ~n6961 & ~n7108 ;
  assign n7110 = x22 ^ x20 ;
  assign n7111 = x24 ^ x20 ;
  assign n7112 = ~n7110 & ~n7111 ;
  assign n7113 = n7109 & n7112 ;
  assign n7114 = n7113 ^ n7108 ;
  assign n7115 = n7114 ^ x23 ;
  assign n7119 = x23 ^ x22 ;
  assign n7123 = ~n6963 & ~n7119 ;
  assign n7118 = x21 ^ x20 ;
  assign n7120 = n7119 ^ x21 ;
  assign n7121 = n7120 ^ x24 ;
  assign n7122 = ~n7118 & n7121 ;
  assign n7124 = n7123 ^ n7122 ;
  assign n7125 = ~x19 & n7124 ;
  assign n7126 = ~n7115 & n7125 ;
  assign n6957 = x28 ^ x27 ;
  assign n7053 = x28 ^ x26 ;
  assign n7054 = x30 ^ x25 ;
  assign n7057 = ~x28 & ~n7054 ;
  assign n7058 = n7057 ^ x25 ;
  assign n7059 = ~n7053 & n7058 ;
  assign n7060 = ~n6957 & n7059 ;
  assign n7061 = ~x29 & n7060 ;
  assign n7072 = ~x29 & ~x30 ;
  assign n7075 = n7072 ^ x29 ;
  assign n7076 = n7075 ^ x30 ;
  assign n7070 = x27 & x28 ;
  assign n7071 = n7070 ^ n6957 ;
  assign n7074 = ~n7071 & ~n7076 ;
  assign n7077 = n7076 ^ n7074 ;
  assign n7078 = n7072 ^ n7070 ;
  assign n7079 = n7078 ^ x25 ;
  assign n7080 = n7077 & n7079 ;
  assign n7081 = n7070 ^ x30 ;
  assign n7082 = n7081 ^ n6957 ;
  assign n6956 = x30 ^ x29 ;
  assign n7083 = n6956 & ~n7070 ;
  assign n7084 = n7082 & n7083 ;
  assign n7085 = n7084 ^ n7081 ;
  assign n7086 = n7085 ^ n7072 ;
  assign n7087 = n7086 ^ x26 ;
  assign n7088 = n7087 ^ n7085 ;
  assign n7089 = n7080 & ~n7088 ;
  assign n7090 = n7089 ^ n7086 ;
  assign n7091 = ~x26 & ~n7090 ;
  assign n7092 = n7091 ^ n7085 ;
  assign n7093 = x25 & n7092 ;
  assign n7063 = x29 ^ x28 ;
  assign n7067 = ~n6956 & ~n7063 ;
  assign n7062 = x27 ^ x26 ;
  assign n7064 = n7063 ^ x27 ;
  assign n7065 = n7064 ^ x30 ;
  assign n7066 = ~n7062 & n7065 ;
  assign n7068 = n7067 ^ n7066 ;
  assign n7069 = ~x25 & n7068 ;
  assign n7094 = n7093 ^ n7069 ;
  assign n7095 = ~n7061 & ~n7094 ;
  assign n7116 = n7115 ^ n7095 ;
  assign n7127 = n7126 ^ n7116 ;
  assign n6955 = x26 ^ x25 ;
  assign n6959 = n7065 ^ n6955 ;
  assign n6960 = x20 ^ x19 ;
  assign n6962 = n6961 ^ n6960 ;
  assign n6964 = n6963 ^ n6962 ;
  assign n7052 = n6959 & n6964 ;
  assign n7128 = n7127 ^ n7052 ;
  assign n6946 = x16 ^ x15 ;
  assign n7010 = x16 ^ x14 ;
  assign n7011 = x18 ^ x13 ;
  assign n7014 = ~x16 & ~n7011 ;
  assign n7015 = n7014 ^ x13 ;
  assign n7016 = ~n7010 & n7015 ;
  assign n7017 = ~n6946 & n7016 ;
  assign n7018 = ~x17 & n7017 ;
  assign n7028 = x15 & x16 ;
  assign n7034 = n7028 ^ n6946 ;
  assign n7035 = ~x17 & ~x18 ;
  assign n6945 = x18 ^ x17 ;
  assign n7036 = n7035 ^ n6945 ;
  assign n7037 = n7034 & ~n7036 ;
  assign n7038 = n7035 ^ n7028 ;
  assign n7039 = n7038 ^ x13 ;
  assign n7040 = ~n7037 & n7039 ;
  assign n7027 = n6946 ^ x17 ;
  assign n7029 = n7028 ^ x18 ;
  assign n7030 = n7029 ^ n6946 ;
  assign n7031 = ~n7028 & n7030 ;
  assign n7032 = ~n7027 & n7031 ;
  assign n7033 = n7032 ^ n7029 ;
  assign n7041 = n7035 ^ n7033 ;
  assign n7042 = n7041 ^ x14 ;
  assign n7043 = n7042 ^ n7033 ;
  assign n7044 = n7040 & ~n7043 ;
  assign n7045 = n7044 ^ n7041 ;
  assign n7046 = ~x14 & ~n7045 ;
  assign n7047 = n7046 ^ n7033 ;
  assign n7048 = x13 & n7047 ;
  assign n7020 = x17 ^ x16 ;
  assign n7024 = ~n6945 & ~n7020 ;
  assign n7019 = x15 ^ x14 ;
  assign n7022 = n7027 ^ x18 ;
  assign n7023 = ~n7019 & n7022 ;
  assign n7025 = n7024 ^ n7023 ;
  assign n7026 = ~x13 & n7025 ;
  assign n7049 = n7048 ^ n7026 ;
  assign n7050 = ~n7018 & ~n7049 ;
  assign n6973 = x11 & x12 ;
  assign n6952 = x12 ^ x11 ;
  assign n6975 = n6973 ^ n6952 ;
  assign n6976 = x8 & n6975 ;
  assign n6974 = n6973 ^ x10 ;
  assign n6979 = n6976 ^ n6974 ;
  assign n6980 = x9 & ~n6979 ;
  assign n6977 = n6976 ^ n6973 ;
  assign n6978 = ~n6974 & ~n6977 ;
  assign n6981 = n6980 ^ n6978 ;
  assign n6982 = ~x7 & n6981 ;
  assign n6983 = ~x9 & ~x10 ;
  assign n6950 = x10 ^ x9 ;
  assign n6984 = n6983 ^ n6950 ;
  assign n6985 = ~n6973 & n6984 ;
  assign n6990 = n6975 & ~n6983 ;
  assign n6949 = x8 ^ x7 ;
  assign n6986 = n6949 ^ x12 ;
  assign n6987 = x9 & n6986 ;
  assign n6991 = n6990 ^ n6987 ;
  assign n6992 = ~x8 & ~n6991 ;
  assign n6993 = n6992 ^ n6987 ;
  assign n6994 = x7 & ~n6993 ;
  assign n6995 = ~n6985 & n6994 ;
  assign n6996 = x7 & n6950 ;
  assign n6997 = n6976 & n6996 ;
  assign n6998 = ~n6995 & ~n6997 ;
  assign n6999 = ~x11 & ~n6996 ;
  assign n7000 = n6984 ^ x8 ;
  assign n7001 = x12 ^ x7 ;
  assign n7004 = n6984 & ~n7001 ;
  assign n7005 = n7004 ^ x7 ;
  assign n7006 = n7000 & n7005 ;
  assign n7007 = n6999 & n7006 ;
  assign n7008 = n6998 & ~n7007 ;
  assign n7009 = ~n6982 & n7008 ;
  assign n7051 = n7050 ^ n7009 ;
  assign n7129 = n7128 ^ n7051 ;
  assign n6880 = x994 ^ x993 ;
  assign n6879 = x992 ^ x991 ;
  assign n6881 = n6880 ^ n6879 ;
  assign n6878 = x996 ^ x995 ;
  assign n6882 = n6881 ^ n6878 ;
  assign n6874 = x2 ^ x1 ;
  assign n6875 = n6874 ^ x0 ;
  assign n6872 = x5 ^ x4 ;
  assign n6873 = n6872 ^ x3 ;
  assign n6876 = n6875 ^ n6873 ;
  assign n6869 = x999 ^ x998 ;
  assign n6870 = n6869 ^ x997 ;
  assign n6871 = n6870 ^ x6 ;
  assign n6877 = n6876 ^ n6871 ;
  assign n6969 = n6882 ^ n6877 ;
  assign n6965 = n6964 ^ n6959 ;
  assign n6951 = n6950 ^ n6949 ;
  assign n6953 = n6952 ^ n6951 ;
  assign n6944 = x14 ^ x13 ;
  assign n6948 = n7022 ^ n6944 ;
  assign n6954 = n6953 ^ n6948 ;
  assign n6970 = n6965 ^ n6954 ;
  assign n6971 = n6969 & n6970 ;
  assign n6966 = n6965 ^ n6953 ;
  assign n6967 = ~n6954 & n6966 ;
  assign n6968 = n6967 ^ n6965 ;
  assign n6972 = n6971 ^ n6968 ;
  assign n7130 = n7129 ^ n6972 ;
  assign n6904 = x995 ^ x994 ;
  assign n6908 = ~n6878 & ~n6904 ;
  assign n6903 = x993 ^ x992 ;
  assign n6905 = n6904 ^ x993 ;
  assign n6906 = n6905 ^ x996 ;
  assign n6907 = ~n6903 & n6906 ;
  assign n6909 = n6908 ^ n6907 ;
  assign n6910 = ~x991 & n6909 ;
  assign n6911 = ~x993 & ~x994 ;
  assign n6917 = ~x995 & ~x996 ;
  assign n6918 = ~n6911 & ~n6917 ;
  assign n6912 = n6911 ^ n6880 ;
  assign n6913 = x991 & x992 ;
  assign n6914 = x996 & n6913 ;
  assign n6915 = ~n6912 & n6914 ;
  assign n6916 = n6915 ^ n6913 ;
  assign n6919 = n6918 ^ n6916 ;
  assign n6922 = n6917 ^ n6878 ;
  assign n6925 = n6912 & n6922 ;
  assign n6926 = n6925 ^ n6916 ;
  assign n6927 = n6919 & ~n6926 ;
  assign n6928 = n6927 ^ n6916 ;
  assign n6929 = ~n6879 & n6928 ;
  assign n6930 = n6927 & n6929 ;
  assign n6931 = n6930 ^ n6928 ;
  assign n6932 = x994 ^ x992 ;
  assign n6933 = x996 ^ x991 ;
  assign n6936 = ~x994 & ~n6933 ;
  assign n6937 = n6936 ^ x991 ;
  assign n6938 = ~n6932 & n6937 ;
  assign n6939 = ~n6880 & n6938 ;
  assign n6940 = ~x995 & n6939 ;
  assign n6941 = ~n6931 & ~n6940 ;
  assign n6942 = ~n6910 & n6941 ;
  assign n6897 = x998 ^ x997 ;
  assign n6898 = ~n6869 & n6897 ;
  assign n6899 = n6898 ^ x997 ;
  assign n6885 = n6871 & n6876 ;
  assign n7160 = n6899 ^ n6885 ;
  assign n6884 = n6873 & n6875 ;
  assign n7161 = n7160 ^ n6884 ;
  assign n6889 = x1 ^ x0 ;
  assign n6890 = ~n6874 & n6889 ;
  assign n6891 = n6890 ^ x0 ;
  assign n6892 = n6891 ^ x3 ;
  assign n6893 = n6892 ^ x4 ;
  assign n6894 = n6893 ^ n6891 ;
  assign n6895 = ~n6872 & n6894 ;
  assign n6896 = n6895 ^ n6892 ;
  assign n7162 = n7161 ^ n6896 ;
  assign n7144 = n7162 ^ n6899 ;
  assign n6886 = x6 & n6870 ;
  assign n7148 = n7144 ^ n6886 ;
  assign n7198 = n7148 ^ n6899 ;
  assign n6883 = n6877 & n6882 ;
  assign n6902 = n7198 ^ n6883 ;
  assign n6943 = n6942 ^ n6902 ;
  assign n7131 = n7130 ^ n6943 ;
  assign n6868 = n6848 ^ n6748 ;
  assign n7132 = n7131 ^ n6868 ;
  assign n7133 = n6846 ^ n6844 ;
  assign n7134 = n6970 ^ n6969 ;
  assign n7135 = n7133 & n7134 ;
  assign n7136 = n7135 ^ n7131 ;
  assign n7137 = n7132 & ~n7136 ;
  assign n7138 = n7137 ^ n7131 ;
  assign n7140 = n7139 ^ n7138 ;
  assign n7305 = n6971 ^ n6943 ;
  assign n7306 = ~n7130 & n7305 ;
  assign n7307 = n7306 ^ n6971 ;
  assign n7252 = n6948 & n6953 ;
  assign n7298 = n7252 ^ n7050 ;
  assign n7299 = n7051 & n7298 ;
  assign n7300 = n7299 ^ n7050 ;
  assign n7287 = x14 & ~n7035 ;
  assign n7286 = n7048 ^ n7028 ;
  assign n7288 = n7287 ^ n7286 ;
  assign n7289 = n7037 ^ n7036 ;
  assign n7292 = ~n7028 & n7289 ;
  assign n7293 = n7292 ^ n7036 ;
  assign n7294 = n7288 & n7293 ;
  assign n7295 = n7294 ^ n7028 ;
  assign n7296 = ~n7048 & ~n7295 ;
  assign n7278 = n6984 ^ n6973 ;
  assign n7280 = n6976 & ~n6983 ;
  assign n7281 = n7280 ^ n6984 ;
  assign n7282 = ~n7278 & ~n7281 ;
  assign n7283 = n7282 ^ n6984 ;
  assign n7284 = n6998 & ~n7283 ;
  assign n7285 = n7284 ^ n6998 ;
  assign n7297 = n7296 ^ n7285 ;
  assign n7301 = n7300 ^ n7297 ;
  assign n7266 = x26 & ~n7072 ;
  assign n7265 = n7093 ^ n7070 ;
  assign n7267 = n7266 ^ n7265 ;
  assign n7271 = ~n7070 & ~n7074 ;
  assign n7272 = n7271 ^ n7076 ;
  assign n7273 = n7267 & n7272 ;
  assign n7274 = n7273 ^ n7070 ;
  assign n7275 = ~n7093 & ~n7274 ;
  assign n7259 = n7101 ^ n7100 ;
  assign n7260 = x20 & n7098 ;
  assign n7261 = n7260 ^ n7100 ;
  assign n7262 = n7259 & ~n7261 ;
  assign n7263 = n7262 ^ n7100 ;
  assign n7264 = ~n7107 & n7263 ;
  assign n7276 = n7275 ^ n7264 ;
  assign n7256 = n7095 ^ n7052 ;
  assign n7257 = ~n7127 & n7256 ;
  assign n7258 = n7257 ^ n7095 ;
  assign n7277 = n7276 ^ n7258 ;
  assign n7302 = n7301 ^ n7277 ;
  assign n7253 = n7252 ^ n6968 ;
  assign n7254 = n7051 & n7253 ;
  assign n7250 = n7051 ^ n6968 ;
  assign n7251 = ~n7128 & n7250 ;
  assign n7255 = n7254 ^ n7251 ;
  assign n7303 = n7302 ^ n7255 ;
  assign n7241 = n6922 ^ n6912 ;
  assign n7242 = x992 & n6918 ;
  assign n7243 = n7242 ^ n6912 ;
  assign n7244 = n7241 & ~n7243 ;
  assign n7245 = n7244 ^ n6912 ;
  assign n7246 = ~n6931 & ~n7245 ;
  assign n7247 = n7246 ^ n6931 ;
  assign n7238 = n6891 ^ n6884 ;
  assign n7239 = n6896 & n7238 ;
  assign n7240 = n7239 ^ n6891 ;
  assign n7248 = n7247 ^ n7240 ;
  assign n7222 = n6899 ^ n6886 ;
  assign n7227 = n7222 ^ n6884 ;
  assign n7218 = n7144 ^ n6896 ;
  assign n7219 = n7218 ^ n7162 ;
  assign n7220 = n7219 ^ n7160 ;
  assign n7203 = n7198 ^ n6896 ;
  assign n7206 = n7203 ^ n6884 ;
  assign n7207 = n7206 ^ n7144 ;
  assign n7179 = ~n7148 & n7222 ;
  assign n7180 = n7207 ^ n7179 ;
  assign n7181 = n7227 ^ n7180 ;
  assign n7182 = n7181 ^ n7162 ;
  assign n7185 = ~n6886 & n7182 ;
  assign n7186 = n7203 ^ n7144 ;
  assign n7187 = n7186 ^ n6899 ;
  assign n7189 = n7206 ^ n6899 ;
  assign n7190 = n7187 & n7189 ;
  assign n7191 = n7185 & n7190 ;
  assign n7192 = n7191 ^ n7179 ;
  assign n7193 = n7220 ^ n7192 ;
  assign n7214 = n7193 ^ n6886 ;
  assign n7215 = n7214 ^ n6884 ;
  assign n7221 = n7220 ^ n7215 ;
  assign n7232 = n7227 ^ n7221 ;
  assign n7233 = n7232 ^ n6942 ;
  assign n7234 = n7233 ^ n6883 ;
  assign n7235 = n7234 ^ n7232 ;
  assign n7236 = ~n6902 & n7235 ;
  assign n7237 = n7236 ^ n7233 ;
  assign n7249 = n7248 ^ n7237 ;
  assign n7304 = n7303 ^ n7249 ;
  assign n7308 = n7307 ^ n7304 ;
  assign n7309 = n7308 ^ n7138 ;
  assign n7310 = ~n7140 & ~n7309 ;
  assign n7311 = n7310 ^ n7308 ;
  assign n6862 = n6840 ^ n6803 ;
  assign n6863 = ~n6804 & n6862 ;
  assign n6864 = n6863 ^ n6803 ;
  assign n6858 = n6802 ^ n6798 ;
  assign n6859 = ~n6799 & n6858 ;
  assign n6860 = n6859 ^ n6798 ;
  assign n6855 = n6839 ^ n6805 ;
  assign n6856 = n6810 & n6855 ;
  assign n6857 = n6856 ^ n6805 ;
  assign n6861 = n6860 ^ n6857 ;
  assign n6865 = n6864 ^ n6861 ;
  assign n6852 = n6851 ^ n6841 ;
  assign n6853 = n6842 & n6852 ;
  assign n6854 = n6853 ^ n6851 ;
  assign n6866 = n6865 ^ n6854 ;
  assign n6528 = n6527 ^ n6475 ;
  assign n6552 = n6551 ^ n6475 ;
  assign n6553 = ~n6528 & n6552 ;
  assign n6554 = n6553 ^ n6527 ;
  assign n6584 = ~n6555 & n6579 ;
  assign n6556 = n6555 ^ n6528 ;
  assign n6557 = n6556 ^ n6551 ;
  assign n6561 = n6560 ^ n6555 ;
  assign n6562 = n6557 ^ n6475 ;
  assign n6563 = n6562 ^ n6561 ;
  assign n6564 = n6551 ^ n6528 ;
  assign n6565 = n6564 ^ n6475 ;
  assign n6566 = n6565 ^ n6561 ;
  assign n6568 = n6557 ^ n6528 ;
  assign n6569 = n6566 & n6568 ;
  assign n6570 = ~n6563 & n6569 ;
  assign n6571 = n6570 ^ n6564 ;
  assign n6572 = n6571 ^ n6557 ;
  assign n6573 = n6561 & ~n6572 ;
  assign n6574 = ~n6557 & n6573 ;
  assign n6575 = n6574 ^ n6560 ;
  assign n6585 = n6584 ^ n6575 ;
  assign n6586 = n6554 & n6585 ;
  assign n6587 = n6586 ^ n6575 ;
  assign n6443 = n6442 ^ n6435 ;
  assign n6451 = n6443 & ~n6450 ;
  assign n6452 = n6451 ^ n6442 ;
  assign n6588 = n6587 ^ n6452 ;
  assign n6867 = n6866 ^ n6588 ;
  assign n7368 = n7311 ^ n6867 ;
  assign n7315 = n7301 ^ n7255 ;
  assign n7316 = n7302 & n7315 ;
  assign n7317 = n7316 ^ n7301 ;
  assign n7312 = n7307 ^ n7303 ;
  assign n7313 = ~n7304 & n7312 ;
  assign n7314 = n7313 ^ n7307 ;
  assign n7326 = n7300 ^ n7285 ;
  assign n7327 = ~n7297 & ~n7326 ;
  assign n7328 = n7327 ^ n7300 ;
  assign n7323 = n7275 ^ n7258 ;
  assign n7324 = n7276 & ~n7323 ;
  assign n7325 = n7324 ^ n7275 ;
  assign n7318 = n7248 ^ n7232 ;
  assign n7319 = n7237 & n7318 ;
  assign n7320 = n7319 ^ n7232 ;
  assign n7321 = n7240 & n7247 ;
  assign n7369 = ~n7320 & ~n7321 ;
  assign n7381 = n7325 & n7369 ;
  assign n7382 = ~n7328 & n7381 ;
  assign n7383 = ~n7314 & n7382 ;
  assign n7322 = n7321 ^ n7320 ;
  assign n7370 = n7369 ^ n7322 ;
  assign n7371 = ~n7314 & n7370 ;
  assign n7372 = n7371 ^ n7325 ;
  assign n7373 = n7372 ^ n7328 ;
  assign n7374 = n7372 ^ n7317 ;
  assign n7375 = ~n7373 & ~n7374 ;
  assign n7376 = n7375 ^ n7372 ;
  assign n7377 = ~n7369 & ~n7376 ;
  assign n7378 = n7371 & ~n7375 ;
  assign n7379 = n7377 & n7378 ;
  assign n7380 = n7379 ^ n7377 ;
  assign n7384 = n7383 ^ n7380 ;
  assign n7385 = n7381 ^ n7371 ;
  assign n7329 = n7328 ^ n7325 ;
  assign n7330 = n7329 ^ n7322 ;
  assign n7331 = n7330 ^ n7317 ;
  assign n7332 = n7331 ^ n7314 ;
  assign n7390 = ~n7328 & ~n7332 ;
  assign n7391 = n7390 ^ n7371 ;
  assign n7392 = n7385 & ~n7391 ;
  assign n7393 = n7392 ^ n7381 ;
  assign n7394 = ~n7384 & n7393 ;
  assign n7395 = ~n7317 & n7394 ;
  assign n7396 = n7395 ^ n7384 ;
  assign n7397 = n7396 ^ n7332 ;
  assign n7398 = n7397 ^ n7311 ;
  assign n7399 = n7398 ^ n7396 ;
  assign n7400 = n7368 & ~n7399 ;
  assign n7401 = n7400 ^ n7397 ;
  assign n7459 = n7396 ^ n7380 ;
  assign n7403 = ~n6554 & n6575 ;
  assign n7405 = n6864 ^ n6857 ;
  assign n7406 = n6861 & n7405 ;
  assign n7413 = n7406 ^ n6864 ;
  assign n7407 = ~n6857 & n6860 ;
  assign n7408 = ~n6864 & n7407 ;
  assign n7409 = n7408 ^ n6861 ;
  assign n7410 = n7409 ^ n7406 ;
  assign n7414 = n7410 ^ n6854 ;
  assign n7411 = ~n6854 & n7410 ;
  assign n7415 = n7414 ^ n7411 ;
  assign n7416 = n7413 & ~n7415 ;
  assign n7449 = ~n7403 & ~n7416 ;
  assign n7443 = n7408 ^ n6588 ;
  assign n7418 = n7406 ^ n6861 ;
  assign n7402 = ~n6452 & ~n6587 ;
  assign n7404 = n7403 ^ n7402 ;
  assign n7419 = n7415 ^ n7413 ;
  assign n7420 = n7419 ^ n7416 ;
  assign n7421 = ~n6588 & ~n7420 ;
  assign n7422 = ~n7404 & n7421 ;
  assign n7423 = ~n7418 & n7422 ;
  assign n7424 = n7423 ^ n7421 ;
  assign n7444 = n7443 ^ n7424 ;
  assign n7450 = n7449 ^ n7444 ;
  assign n7451 = n6588 & ~n7450 ;
  assign n7452 = n7451 ^ n7444 ;
  assign n7412 = n7404 & n7411 ;
  assign n7417 = n7416 ^ n7403 ;
  assign n7429 = n6588 & n7417 ;
  assign n7425 = n7404 & n7408 ;
  assign n7426 = n7424 & n7425 ;
  assign n7427 = n7426 ^ n7424 ;
  assign n7430 = n7429 ^ n7427 ;
  assign n7431 = n7412 & n7430 ;
  assign n7432 = n7431 ^ n7430 ;
  assign n7442 = n7432 ^ n7380 ;
  assign n7458 = n7452 ^ n7442 ;
  assign n7460 = n7459 ^ n7458 ;
  assign n7461 = n7460 ^ n7452 ;
  assign n7462 = ~n7401 & ~n7461 ;
  assign n7463 = n7462 ^ n7458 ;
  assign n8681 = ~n7380 & n7452 ;
  assign n8682 = n7463 & n8681 ;
  assign n5826 = x952 ^ x951 ;
  assign n5821 = ~x951 & ~x952 ;
  assign n5827 = n5826 ^ n5821 ;
  assign n5820 = x950 ^ x949 ;
  assign n5828 = x949 & ~n5820 ;
  assign n5829 = x954 & n5828 ;
  assign n5830 = ~n5827 & n5829 ;
  assign n5831 = n5830 ^ n5828 ;
  assign n5822 = x954 ^ x953 ;
  assign n5823 = x953 & ~n5822 ;
  assign n5824 = n5823 ^ n5822 ;
  assign n5825 = ~n5821 & n5824 ;
  assign n5832 = n5831 ^ n5825 ;
  assign n5837 = ~n5823 & n5827 ;
  assign n5838 = n5837 ^ n5825 ;
  assign n5839 = n5832 & n5838 ;
  assign n5840 = n5839 ^ n5831 ;
  assign n5841 = n5827 ^ n5823 ;
  assign n5845 = x950 & n5825 ;
  assign n5846 = n5845 ^ n5827 ;
  assign n5847 = ~n5841 & n5846 ;
  assign n5848 = n5847 ^ n5823 ;
  assign n5849 = n5840 & ~n5848 ;
  assign n5850 = ~n5820 & n5849 ;
  assign n5851 = n5839 & n5850 ;
  assign n5852 = n5851 ^ n5849 ;
  assign n5853 = n5852 ^ n5848 ;
  assign n5792 = x946 ^ x945 ;
  assign n5787 = ~x945 & ~x946 ;
  assign n5793 = n5792 ^ n5787 ;
  assign n5786 = x944 ^ x943 ;
  assign n5794 = x943 & ~n5786 ;
  assign n5795 = x948 & n5794 ;
  assign n5796 = ~n5793 & n5795 ;
  assign n5797 = n5796 ^ n5794 ;
  assign n5788 = x948 ^ x947 ;
  assign n5789 = x947 & ~n5788 ;
  assign n5790 = n5789 ^ n5788 ;
  assign n5791 = ~n5787 & n5790 ;
  assign n5798 = n5797 ^ n5791 ;
  assign n5803 = ~n5789 & n5793 ;
  assign n5804 = n5803 ^ n5791 ;
  assign n5805 = n5798 & n5804 ;
  assign n5806 = n5805 ^ n5797 ;
  assign n5807 = n5793 ^ n5789 ;
  assign n5811 = x944 & n5791 ;
  assign n5812 = n5811 ^ n5793 ;
  assign n5813 = ~n5807 & n5812 ;
  assign n5814 = n5813 ^ n5789 ;
  assign n5815 = n5806 & ~n5814 ;
  assign n5816 = ~n5786 & n5815 ;
  assign n5817 = n5805 & n5816 ;
  assign n5818 = n5817 ^ n5815 ;
  assign n5819 = n5818 ^ n5814 ;
  assign n5855 = n5853 ^ n5819 ;
  assign n5854 = ~n5819 & ~n5853 ;
  assign n5856 = n5855 ^ n5854 ;
  assign n5877 = x961 & ~x962 ;
  assign n5879 = x966 ^ x965 ;
  assign n5878 = x965 & x966 ;
  assign n5880 = n5879 ^ n5878 ;
  assign n5881 = n5877 & n5880 ;
  assign n5882 = x964 ^ x963 ;
  assign n5883 = n5878 ^ x964 ;
  assign n5884 = n5882 & ~n5883 ;
  assign n5885 = n5884 ^ x963 ;
  assign n5886 = n5881 & n5885 ;
  assign n5887 = n5886 ^ n5877 ;
  assign n5888 = n5887 ^ x961 ;
  assign n5889 = ~x963 & ~x964 ;
  assign n5890 = n5889 ^ n5882 ;
  assign n5891 = n5882 ^ x966 ;
  assign n5892 = n5891 ^ n5889 ;
  assign n5893 = n5892 ^ x965 ;
  assign n5894 = n5892 ^ n5882 ;
  assign n5895 = ~n5893 & ~n5894 ;
  assign n5896 = n5890 & n5895 ;
  assign n5897 = n5896 ^ n5892 ;
  assign n5898 = x962 & n5897 ;
  assign n5899 = n5888 & n5898 ;
  assign n5900 = n5899 ^ n5888 ;
  assign n5901 = x962 & n5880 ;
  assign n5904 = n5901 ^ n5878 ;
  assign n6031 = n5882 ^ n5878 ;
  assign n6034 = ~n5904 & ~n6031 ;
  assign n6035 = n6034 ^ n5882 ;
  assign n6036 = ~n5889 & ~n6035 ;
  assign n6037 = ~n5900 & n6036 ;
  assign n5945 = ~x957 & ~x958 ;
  assign n5933 = x955 & ~x956 ;
  assign n5935 = x960 ^ x959 ;
  assign n5934 = x959 & x960 ;
  assign n5936 = n5935 ^ n5934 ;
  assign n5937 = n5933 & n5936 ;
  assign n5938 = x958 ^ x957 ;
  assign n5939 = n5934 ^ x958 ;
  assign n5940 = n5938 & ~n5939 ;
  assign n5941 = n5940 ^ x957 ;
  assign n5942 = n5937 & n5941 ;
  assign n5943 = n5942 ^ n5933 ;
  assign n5944 = n5943 ^ x955 ;
  assign n5946 = n5945 ^ n5938 ;
  assign n5947 = n5938 ^ x960 ;
  assign n5948 = n5947 ^ n5945 ;
  assign n5949 = n5948 ^ x959 ;
  assign n5950 = n5948 ^ n5938 ;
  assign n5951 = ~n5949 & ~n5950 ;
  assign n5952 = n5946 & n5951 ;
  assign n5953 = n5952 ^ n5948 ;
  assign n5954 = x956 & n5953 ;
  assign n5955 = n5944 & n5954 ;
  assign n5956 = n5955 ^ n5944 ;
  assign n6023 = ~n5945 & ~n5956 ;
  assign n5957 = x956 & n5936 ;
  assign n5960 = n5957 ^ n5934 ;
  assign n6024 = n5938 ^ n5934 ;
  assign n6025 = n5960 & ~n6024 ;
  assign n6026 = n6025 ^ n5934 ;
  assign n6027 = n6023 & n6026 ;
  assign n6028 = n6027 ^ n5956 ;
  assign n6029 = n6028 ^ n5900 ;
  assign n6038 = n6037 ^ n6029 ;
  assign n5961 = ~n5939 & ~n5960 ;
  assign n5958 = n5957 ^ n5939 ;
  assign n5959 = x957 & ~n5958 ;
  assign n5962 = n5961 ^ n5959 ;
  assign n5963 = ~x955 & n5962 ;
  assign n5965 = n5963 ^ n5956 ;
  assign n5966 = ~x959 & ~n5965 ;
  assign n5968 = x960 ^ x957 ;
  assign n5967 = x960 ^ x956 ;
  assign n5969 = n5968 ^ n5967 ;
  assign n5970 = n5969 ^ x960 ;
  assign n5972 = x956 & n5970 ;
  assign n5973 = n5972 ^ x960 ;
  assign n5990 = x956 ^ x955 ;
  assign n5976 = x960 ^ x958 ;
  assign n5977 = n5976 ^ n5967 ;
  assign n5978 = n5990 ^ n5977 ;
  assign n5980 = n5967 ^ n5938 ;
  assign n5981 = n5980 ^ x960 ;
  assign n5982 = ~n5978 & n5981 ;
  assign n5985 = n5982 ^ x957 ;
  assign n5986 = ~n5973 & ~n5985 ;
  assign n5987 = n5966 & n5986 ;
  assign n5988 = n5987 ^ n5965 ;
  assign n5905 = ~n5883 & ~n5904 ;
  assign n5902 = n5901 ^ n5883 ;
  assign n5903 = x963 & ~n5902 ;
  assign n5906 = n5905 ^ n5903 ;
  assign n5907 = ~x961 & n5906 ;
  assign n5909 = n5907 ^ n5900 ;
  assign n5910 = ~x965 & ~n5909 ;
  assign n5912 = x966 ^ x963 ;
  assign n5911 = x966 ^ x962 ;
  assign n5913 = n5912 ^ n5911 ;
  assign n5914 = n5913 ^ x966 ;
  assign n5916 = x962 & n5914 ;
  assign n5917 = n5916 ^ x966 ;
  assign n5994 = x962 ^ x961 ;
  assign n5920 = x966 ^ x964 ;
  assign n5921 = n5920 ^ n5911 ;
  assign n5922 = n5994 ^ n5921 ;
  assign n5924 = n5911 ^ n5882 ;
  assign n5925 = n5924 ^ x966 ;
  assign n5926 = ~n5922 & n5925 ;
  assign n5929 = n5926 ^ x963 ;
  assign n5930 = ~n5917 & ~n5929 ;
  assign n5931 = n5910 & n5930 ;
  assign n5932 = n5931 ^ n5909 ;
  assign n5989 = n5988 ^ n5932 ;
  assign n5991 = n5938 ^ n5935 ;
  assign n5992 = n5991 ^ n5990 ;
  assign n5995 = n5882 ^ n5879 ;
  assign n5996 = n5995 ^ n5994 ;
  assign n6039 = n5992 & n5996 ;
  assign n6040 = n6039 ^ n5932 ;
  assign n6041 = ~n5989 & ~n6040 ;
  assign n6042 = n6041 ^ n6039 ;
  assign n6055 = n6042 ^ n6028 ;
  assign n6056 = ~n6038 & n6055 ;
  assign n6057 = n6056 ^ n6042 ;
  assign n5866 = n5792 ^ n5786 ;
  assign n5867 = n5792 ^ n5788 ;
  assign n5868 = n5866 & n5867 ;
  assign n5863 = n5794 ^ n5789 ;
  assign n5864 = n5863 ^ n5787 ;
  assign n5860 = n5828 ^ n5823 ;
  assign n5861 = n5860 ^ n5821 ;
  assign n5857 = n5826 ^ n5820 ;
  assign n5858 = n5826 ^ n5822 ;
  assign n5859 = n5857 & n5858 ;
  assign n5862 = n5861 ^ n5859 ;
  assign n5865 = n5864 ^ n5862 ;
  assign n5869 = n5868 ^ n5865 ;
  assign n5870 = n5866 ^ n5788 ;
  assign n5871 = n5857 ^ n5822 ;
  assign n5872 = n5870 & n5871 ;
  assign n5873 = n5872 ^ n5862 ;
  assign n5874 = n5869 & ~n5873 ;
  assign n5875 = n5874 ^ n5862 ;
  assign n6044 = n5875 ^ n5855 ;
  assign n6043 = n6042 ^ n6038 ;
  assign n6045 = n6044 ^ n6043 ;
  assign n5998 = n5871 ^ n5870 ;
  assign n6008 = n5992 ^ n5871 ;
  assign n6009 = n6008 ^ n5996 ;
  assign n6001 = ~n5998 & n6009 ;
  assign n5993 = n5992 ^ n5989 ;
  assign n6006 = n6001 ^ n5993 ;
  assign n6007 = ~n5989 & ~n6006 ;
  assign n5999 = n5996 ^ n5992 ;
  assign n6011 = ~n5999 & ~n6008 ;
  assign n6010 = ~n5870 & n6009 ;
  assign n6012 = n6011 ^ n6010 ;
  assign n6013 = n6012 ^ n5989 ;
  assign n6014 = n6013 ^ n5872 ;
  assign n6015 = ~n5869 & ~n6014 ;
  assign n6016 = n6015 ^ n5872 ;
  assign n6017 = n6007 ^ n5996 ;
  assign n6018 = ~n6016 & n6017 ;
  assign n6019 = n5993 & n6018 ;
  assign n6020 = ~n6007 & n6019 ;
  assign n6021 = n6020 ^ n6018 ;
  assign n6022 = n6021 ^ n6016 ;
  assign n6046 = n6045 ^ n6022 ;
  assign n6047 = n6046 ^ n6043 ;
  assign n6052 = n5856 & n6022 ;
  assign n6053 = n6052 ^ n6046 ;
  assign n6054 = n6047 & ~n6053 ;
  assign n6058 = n6057 ^ n6054 ;
  assign n5876 = n5854 & n5875 ;
  assign n6059 = n6058 ^ n5876 ;
  assign n6060 = n5856 & ~n6059 ;
  assign n6315 = n6043 ^ n6022 ;
  assign n6316 = n6043 ^ n5875 ;
  assign n6317 = ~n6315 & ~n6316 ;
  assign n6318 = n6317 ^ n6043 ;
  assign n6319 = ~n6057 & ~n6318 ;
  assign n6322 = n6060 & ~n6319 ;
  assign n6063 = x970 ^ x969 ;
  assign n6062 = ~x969 & ~x970 ;
  assign n6064 = n6063 ^ n6062 ;
  assign n6069 = x967 & x968 ;
  assign n6070 = ~n6064 & n6069 ;
  assign n6071 = x972 & n6070 ;
  assign n6072 = n6071 ^ n6069 ;
  assign n6066 = x972 ^ x971 ;
  assign n6065 = ~x971 & ~x972 ;
  assign n6067 = n6066 ^ n6065 ;
  assign n6068 = n6064 & n6067 ;
  assign n6073 = n6072 ^ n6068 ;
  assign n6078 = ~n6062 & ~n6065 ;
  assign n6079 = n6078 ^ n6068 ;
  assign n6080 = ~n6073 & n6079 ;
  assign n6061 = x968 ^ x967 ;
  assign n6081 = n6080 ^ n6072 ;
  assign n6082 = ~n6061 & n6081 ;
  assign n6083 = n6080 & n6082 ;
  assign n6084 = n6083 ^ n6081 ;
  assign n6085 = n6067 ^ n6064 ;
  assign n6086 = n6085 ^ n6068 ;
  assign n6087 = ~n6070 & n6086 ;
  assign n6088 = ~n6084 & n6087 ;
  assign n6089 = x976 ^ x975 ;
  assign n6090 = x977 & x978 ;
  assign n6091 = n6090 ^ x976 ;
  assign n6092 = n6089 & ~n6091 ;
  assign n6093 = n6092 ^ x975 ;
  assign n6094 = x975 & x976 ;
  assign n6095 = n6090 & n6094 ;
  assign n6096 = x978 ^ x977 ;
  assign n6097 = n6096 ^ n6090 ;
  assign n6098 = x974 & n6097 ;
  assign n6099 = ~n6095 & ~n6098 ;
  assign n6100 = n6093 & n6099 ;
  assign n6101 = n6100 ^ n6093 ;
  assign n6114 = x973 & x974 ;
  assign n6115 = n6094 & n6114 ;
  assign n6102 = x974 ^ x973 ;
  assign n6103 = n6095 ^ n6091 ;
  assign n6104 = n6103 ^ n6092 ;
  assign n6105 = n6104 ^ n6093 ;
  assign n6106 = n6105 ^ n6094 ;
  assign n6107 = n6106 ^ n6093 ;
  assign n6110 = x974 & n6107 ;
  assign n6111 = n6110 ^ n6093 ;
  assign n6112 = ~n6102 & n6111 ;
  assign n6113 = n6112 ^ n6093 ;
  assign n6116 = n6115 ^ n6113 ;
  assign n6117 = ~x978 & n6116 ;
  assign n6118 = n6117 ^ n6113 ;
  assign n6119 = x977 & ~n6118 ;
  assign n6120 = n6117 & n6119 ;
  assign n6121 = n6120 ^ n6118 ;
  assign n6122 = ~n6101 & ~n6121 ;
  assign n6124 = x984 ^ x983 ;
  assign n6123 = ~x983 & ~x984 ;
  assign n6125 = n6124 ^ n6123 ;
  assign n6129 = n6125 ^ x982 ;
  assign n6126 = x981 & x982 ;
  assign n6127 = ~n6125 & n6126 ;
  assign n6141 = n6129 ^ n6127 ;
  assign n6128 = x982 ^ x981 ;
  assign n6130 = n6128 & n6129 ;
  assign n6142 = n6141 ^ n6130 ;
  assign n6204 = ~x980 & n6142 ;
  assign n6152 = x988 ^ x987 ;
  assign n6154 = x990 ^ x989 ;
  assign n6153 = ~x989 & ~x990 ;
  assign n6155 = n6154 ^ n6153 ;
  assign n6156 = n6155 ^ x988 ;
  assign n6157 = n6152 & n6156 ;
  assign n6158 = n6157 ^ x987 ;
  assign n6162 = x987 & x988 ;
  assign n6163 = ~n6155 & n6162 ;
  assign n6182 = x986 & ~n6153 ;
  assign n6183 = ~n6163 & ~n6182 ;
  assign n6184 = n6158 & n6183 ;
  assign n6185 = n6184 ^ n6158 ;
  assign n6171 = n6162 ^ x986 ;
  assign n6174 = n6152 ^ x985 ;
  assign n6175 = ~x990 & n6174 ;
  assign n6176 = n6175 ^ x985 ;
  assign n6177 = ~n6162 & n6176 ;
  assign n6178 = n6177 ^ x985 ;
  assign n6179 = ~n6171 & n6178 ;
  assign n6180 = x990 & n6179 ;
  assign n6159 = n6158 ^ n6153 ;
  assign n6160 = n6159 ^ x986 ;
  assign n6161 = n6160 ^ n6158 ;
  assign n6164 = n6163 ^ n6156 ;
  assign n6165 = n6164 ^ n6157 ;
  assign n6166 = x986 & ~n6165 ;
  assign n6167 = n6166 ^ n6158 ;
  assign n6168 = n6161 & n6167 ;
  assign n6169 = n6168 ^ n6158 ;
  assign n6170 = x985 & n6169 ;
  assign n6181 = n6180 ^ n6170 ;
  assign n6197 = n6185 ^ n6181 ;
  assign n6198 = n6185 ^ n6179 ;
  assign n6199 = ~n6197 & ~n6198 ;
  assign n6196 = x989 & n6179 ;
  assign n6200 = n6199 ^ n6196 ;
  assign n6194 = ~x985 & n6165 ;
  assign n6195 = ~n6182 & n6194 ;
  assign n6201 = n6200 ^ n6195 ;
  assign n6131 = n6130 ^ x981 ;
  assign n6132 = ~n6127 & n6131 ;
  assign n6133 = x980 & n6132 ;
  assign n6134 = ~n6123 & n6133 ;
  assign n6135 = n6134 ^ n6132 ;
  assign n6136 = n6135 ^ n6131 ;
  assign n6202 = n6201 ^ n6136 ;
  assign n6189 = n6128 ^ n6124 ;
  assign n6188 = x980 ^ x979 ;
  assign n6190 = n6189 ^ n6188 ;
  assign n6138 = n6131 ^ n6123 ;
  assign n6137 = ~n6123 & n6131 ;
  assign n6139 = n6138 ^ n6137 ;
  assign n6191 = n6190 ^ n6139 ;
  assign n6192 = n6190 ^ x979 ;
  assign n6193 = ~n6191 & n6192 ;
  assign n6203 = n6202 ^ n6193 ;
  assign n6205 = n6204 ^ n6203 ;
  assign n6206 = x986 ^ x985 ;
  assign n6207 = n6206 ^ n6152 ;
  assign n6208 = n6207 ^ n6154 ;
  assign n6209 = n6190 & n6208 ;
  assign n6210 = n6209 ^ n6201 ;
  assign n6211 = n6205 & n6210 ;
  assign n6212 = n6211 ^ n6209 ;
  assign n6186 = ~n6181 & ~n6185 ;
  assign n6147 = x979 & n6137 ;
  assign n6140 = n6139 ^ n6127 ;
  assign n6143 = x979 & ~n6142 ;
  assign n6144 = ~n6140 & n6143 ;
  assign n6148 = n6147 ^ n6144 ;
  assign n6149 = ~x980 & n6148 ;
  assign n6150 = n6149 ^ n6144 ;
  assign n6151 = ~n6136 & ~n6150 ;
  assign n6187 = n6186 ^ n6151 ;
  assign n6213 = n6212 ^ n6187 ;
  assign n6257 = ~x973 & n6101 ;
  assign n6248 = n6097 ^ x973 ;
  assign n6249 = n6248 ^ x974 ;
  assign n6250 = n6094 ^ x974 ;
  assign n6251 = ~n6102 & ~n6250 ;
  assign n6252 = n6251 ^ n6104 ;
  assign n6253 = ~n6098 & ~n6252 ;
  assign n6254 = n6249 & n6253 ;
  assign n6256 = n6254 ^ n6251 ;
  assign n6258 = n6257 ^ n6256 ;
  assign n6247 = x977 & n6115 ;
  assign n6259 = n6258 ^ n6247 ;
  assign n6260 = ~n6121 & ~n6259 ;
  assign n6229 = x971 ^ x970 ;
  assign n6233 = ~n6066 & ~n6229 ;
  assign n6228 = x969 ^ x968 ;
  assign n6230 = n6229 ^ x969 ;
  assign n6231 = n6230 ^ x972 ;
  assign n6232 = ~n6228 & n6231 ;
  assign n6234 = n6233 ^ n6232 ;
  assign n6235 = ~x967 & n6234 ;
  assign n6236 = x970 ^ x968 ;
  assign n6237 = x972 ^ x967 ;
  assign n6240 = ~x970 & ~n6237 ;
  assign n6241 = n6240 ^ x967 ;
  assign n6242 = ~n6236 & n6241 ;
  assign n6243 = ~n6063 & n6242 ;
  assign n6244 = ~x971 & n6243 ;
  assign n6245 = ~n6084 & ~n6244 ;
  assign n6246 = ~n6235 & n6245 ;
  assign n6261 = n6260 ^ n6246 ;
  assign n6215 = n6231 ^ n6061 ;
  assign n6216 = n6102 ^ n6096 ;
  assign n6217 = n6216 ^ n6089 ;
  assign n6218 = n6215 & n6217 ;
  assign n6276 = n6246 ^ n6218 ;
  assign n6277 = ~n6261 & n6276 ;
  assign n6278 = n6277 ^ n6218 ;
  assign n6275 = n6122 ^ n6088 ;
  assign n6279 = n6278 ^ n6275 ;
  assign n6280 = n6279 ^ n6213 ;
  assign n6220 = n6217 ^ n6215 ;
  assign n6221 = n6208 ^ n6190 ;
  assign n6222 = n6221 ^ n6215 ;
  assign n6223 = ~n6220 & n6222 ;
  assign n6224 = n6223 ^ n6221 ;
  assign n6225 = n6208 & ~n6224 ;
  assign n6226 = ~n6223 & n6225 ;
  assign n6227 = n6226 ^ n6224 ;
  assign n6262 = n6261 ^ n6227 ;
  assign n6219 = n6209 & n6218 ;
  assign n6265 = n6262 ^ n6219 ;
  assign n6266 = n6265 ^ n6209 ;
  assign n6267 = n6205 & n6266 ;
  assign n6268 = n6267 ^ n6209 ;
  assign n6269 = n6227 ^ n6218 ;
  assign n6272 = ~n6261 & ~n6269 ;
  assign n6273 = n6272 ^ n6218 ;
  assign n6274 = ~n6268 & ~n6273 ;
  assign n6281 = n6280 ^ n6274 ;
  assign n6282 = n6213 & ~n6281 ;
  assign n6283 = n6212 ^ n6186 ;
  assign n6284 = n6187 & ~n6283 ;
  assign n6285 = n6284 ^ n6186 ;
  assign n6286 = n6278 ^ n6122 ;
  assign n6289 = n6275 & ~n6286 ;
  assign n6290 = n6289 ^ n6122 ;
  assign n6291 = n6285 & ~n6290 ;
  assign n6292 = n6282 & n6291 ;
  assign n6293 = n6292 ^ n6285 ;
  assign n6296 = n6274 ^ n6088 ;
  assign n6301 = n6278 ^ n6274 ;
  assign n6302 = n6296 & n6301 ;
  assign n6297 = n6278 ^ n6213 ;
  assign n6298 = n6297 ^ n6285 ;
  assign n6303 = n6302 ^ n6298 ;
  assign n6294 = n6281 ^ n6122 ;
  assign n6295 = n6294 ^ n6285 ;
  assign n6304 = n6303 ^ n6295 ;
  assign n6305 = n6278 & n6304 ;
  assign n6306 = n6305 ^ n6294 ;
  assign n6307 = n6279 ^ n6274 ;
  assign n6308 = ~n6306 & ~n6307 ;
  assign n6309 = n6308 ^ n6303 ;
  assign n6310 = ~n6293 & ~n6309 ;
  assign n6311 = ~n6122 & n6310 ;
  assign n6312 = ~n6088 & n6311 ;
  assign n6313 = n6312 ^ n6310 ;
  assign n6314 = n6313 ^ n6293 ;
  assign n6320 = n6319 ^ n6314 ;
  assign n6323 = n6322 ^ n6320 ;
  assign n6325 = n6221 ^ n6220 ;
  assign n6326 = n5999 ^ n5998 ;
  assign n6327 = n6325 & n6326 ;
  assign n6324 = n6265 ^ n6205 ;
  assign n6328 = n6327 ^ n6324 ;
  assign n6329 = n6013 ^ n5869 ;
  assign n6330 = n6329 ^ n6046 ;
  assign n6331 = n6330 ^ n6324 ;
  assign n6332 = n6331 ^ n6046 ;
  assign n6333 = n6328 & n6332 ;
  assign n6334 = n6333 ^ n6330 ;
  assign n6335 = n6309 ^ n6046 ;
  assign n6336 = n6335 ^ n6281 ;
  assign n6337 = n6336 ^ n6309 ;
  assign n6338 = ~n6334 & n6337 ;
  assign n6339 = n6338 ^ n6335 ;
  assign n7363 = n6309 ^ n6059 ;
  assign n7364 = n6339 & n7363 ;
  assign n7365 = n7364 ^ n6059 ;
  assign n7439 = n7365 ^ n6314 ;
  assign n7440 = ~n6323 & n7439 ;
  assign n7366 = n7365 ^ n6323 ;
  assign n7334 = n7399 ^ n6867 ;
  assign n6340 = n6339 ^ n6059 ;
  assign n7335 = n7334 ^ n6340 ;
  assign n7353 = n6334 ^ n6281 ;
  assign n7338 = n6329 ^ n6328 ;
  assign n7344 = n7338 ^ n7135 ;
  assign n7345 = n7344 ^ n7132 ;
  assign n7336 = n6326 ^ n6325 ;
  assign n7337 = n7336 ^ n7134 ;
  assign n7339 = n7338 ^ n7133 ;
  assign n7340 = n7339 ^ n7336 ;
  assign n7341 = n7340 ^ n7338 ;
  assign n7342 = ~n7337 & n7341 ;
  assign n7343 = n7342 ^ n7339 ;
  assign n7346 = n7345 ^ n7343 ;
  assign n7347 = n7345 ^ n7135 ;
  assign n7348 = ~n7346 & n7347 ;
  assign n7349 = n7348 ^ n7344 ;
  assign n7350 = ~n7338 & n7349 ;
  assign n7351 = ~n7348 & n7350 ;
  assign n7352 = n7351 ^ n7349 ;
  assign n7354 = n7353 ^ n7352 ;
  assign n7355 = n7308 ^ n7140 ;
  assign n7358 = n7355 ^ n7352 ;
  assign n7359 = n7354 & n7358 ;
  assign n7356 = n7355 ^ n7334 ;
  assign n7360 = n7359 ^ n7356 ;
  assign n7361 = n7335 & n7360 ;
  assign n7362 = n7361 ^ n7334 ;
  assign n7367 = n7366 ^ n7362 ;
  assign n7433 = n7432 ^ n7401 ;
  assign n7434 = n7433 ^ n7362 ;
  assign n7435 = n7367 & n7434 ;
  assign n7436 = n7435 ^ n7433 ;
  assign n7437 = n7436 ^ n7365 ;
  assign n7441 = n7440 ^ n7437 ;
  assign n7464 = n7463 ^ n7436 ;
  assign n7465 = ~n7441 & ~n7464 ;
  assign n7466 = n7465 ^ n7436 ;
  assign n8680 = n7466 ^ n7463 ;
  assign n8683 = n8682 ^ n8680 ;
  assign n7725 = ~x915 & ~x916 ;
  assign n7731 = ~x917 & ~x918 ;
  assign n7732 = ~n7725 & ~n7731 ;
  assign n7724 = x913 & x914 ;
  assign n7726 = x916 ^ x915 ;
  assign n7727 = n7726 ^ n7725 ;
  assign n7728 = x918 & ~n7727 ;
  assign n7729 = n7724 & n7728 ;
  assign n7730 = n7729 ^ n7724 ;
  assign n7733 = n7732 ^ n7730 ;
  assign n7734 = x918 ^ x917 ;
  assign n7735 = n7734 ^ n7731 ;
  assign n7740 = n7727 & n7735 ;
  assign n7741 = n7740 ^ n7730 ;
  assign n7742 = n7733 & ~n7741 ;
  assign n7723 = x914 ^ x913 ;
  assign n7743 = n7742 ^ n7730 ;
  assign n7744 = ~n7723 & n7743 ;
  assign n7745 = n7742 & n7744 ;
  assign n7746 = n7745 ^ n7743 ;
  assign n7747 = n7735 ^ n7727 ;
  assign n7752 = x914 & n7732 ;
  assign n7753 = n7752 ^ n7735 ;
  assign n7754 = n7747 & n7753 ;
  assign n7755 = n7754 ^ n7727 ;
  assign n7756 = ~n7746 & n7755 ;
  assign n7800 = x917 ^ x914 ;
  assign n7803 = n7734 & n7800 ;
  assign n7804 = n7803 ^ x917 ;
  assign n7805 = n7725 & ~n7804 ;
  assign n7806 = n7805 ^ n7755 ;
  assign n7807 = ~x913 & ~n7806 ;
  assign n7808 = ~x917 & ~n7746 ;
  assign n7810 = x918 ^ x915 ;
  assign n7809 = x918 ^ x914 ;
  assign n7811 = n7810 ^ n7809 ;
  assign n7812 = n7811 ^ x918 ;
  assign n7814 = x914 & n7812 ;
  assign n7815 = n7814 ^ x918 ;
  assign n7818 = x918 ^ x916 ;
  assign n7819 = n7818 ^ n7809 ;
  assign n7820 = n7819 ^ n7723 ;
  assign n7822 = n7809 ^ n7726 ;
  assign n7823 = n7822 ^ x918 ;
  assign n7824 = ~n7820 & n7823 ;
  assign n7827 = n7824 ^ x915 ;
  assign n7828 = ~n7815 & ~n7827 ;
  assign n7829 = n7808 & n7828 ;
  assign n7830 = n7829 ^ n7746 ;
  assign n7840 = n7807 & ~n7830 ;
  assign n7759 = x911 & x912 ;
  assign n7757 = x909 & x910 ;
  assign n7760 = n7759 ^ n7757 ;
  assign n7761 = x910 ^ x909 ;
  assign n7762 = n7761 ^ n7757 ;
  assign n7763 = x912 ^ x911 ;
  assign n7764 = n7763 ^ n7759 ;
  assign n7765 = n7762 & n7764 ;
  assign n7766 = n7765 ^ n7759 ;
  assign n7836 = ~n7760 & ~n7766 ;
  assign n7831 = x908 ^ x907 ;
  assign n7832 = n7761 ^ x908 ;
  assign n7833 = n7832 ^ n7763 ;
  assign n7834 = n7831 & ~n7833 ;
  assign n7835 = n7834 ^ x907 ;
  assign n7837 = n7836 ^ n7835 ;
  assign n7838 = n7837 ^ n7830 ;
  assign n7841 = n7840 ^ n7838 ;
  assign n7842 = n7831 ^ n7763 ;
  assign n7843 = n7842 ^ n7761 ;
  assign n7844 = n7734 ^ n7723 ;
  assign n7845 = n7844 ^ n7726 ;
  assign n7846 = n7843 & n7845 ;
  assign n7847 = n7846 ^ n7837 ;
  assign n7848 = ~n7841 & ~n7847 ;
  assign n7849 = n7848 ^ n7846 ;
  assign n7768 = n7757 ^ x907 ;
  assign n7771 = n7768 ^ n7760 ;
  assign n7758 = n7757 ^ x908 ;
  assign n7776 = n7771 ^ n7758 ;
  assign n7767 = n7766 ^ n7760 ;
  assign n7769 = n7768 ^ n7767 ;
  assign n7777 = n7776 ^ n7769 ;
  assign n7778 = n7777 ^ n7760 ;
  assign n7780 = n7776 & n7778 ;
  assign n7773 = n7769 ^ n7760 ;
  assign n7774 = n7773 ^ n7759 ;
  assign n7775 = ~n7765 & n7774 ;
  assign n7781 = n7780 ^ n7775 ;
  assign n7782 = n7781 ^ n7773 ;
  assign n7783 = n7780 ^ n7771 ;
  assign n7784 = n7783 ^ n7773 ;
  assign n7785 = n7782 & n7784 ;
  assign n7786 = ~n7760 & n7785 ;
  assign n7787 = n7786 ^ n7780 ;
  assign n7788 = n7787 ^ n7778 ;
  assign n7796 = n7788 ^ n7757 ;
  assign n7799 = n7796 ^ n7758 ;
  assign n7851 = n7849 ^ n7799 ;
  assign n7850 = ~n7799 & ~n7849 ;
  assign n7852 = n7851 ^ n7850 ;
  assign n7853 = ~n7756 & ~n7852 ;
  assign n7890 = x897 & x898 ;
  assign n7889 = x899 & x900 ;
  assign n7891 = n7890 ^ n7889 ;
  assign n7856 = x900 ^ x899 ;
  assign n7892 = n7889 ^ n7856 ;
  assign n7854 = x898 ^ x897 ;
  assign n7893 = n7890 ^ n7854 ;
  assign n7894 = n7892 & n7893 ;
  assign n7895 = n7894 ^ n7890 ;
  assign n7896 = ~n7891 & ~n7895 ;
  assign n7855 = n7854 ^ x896 ;
  assign n7857 = n7856 ^ n7855 ;
  assign n7870 = x902 ^ x901 ;
  assign n7862 = ~x903 & ~x904 ;
  assign n7858 = x904 ^ x903 ;
  assign n7863 = n7862 ^ n7858 ;
  assign n7864 = x906 ^ x905 ;
  assign n7859 = x905 & x906 ;
  assign n7865 = n7864 ^ n7859 ;
  assign n7867 = ~n7863 & n7865 ;
  assign n7878 = n7859 & ~n7862 ;
  assign n7879 = ~n7867 & ~n7878 ;
  assign n7880 = n7870 & ~n7879 ;
  assign n7860 = n7859 ^ x904 ;
  assign n7861 = ~n7858 & ~n7860 ;
  assign n7871 = n7861 ^ x902 ;
  assign n7866 = n7865 ^ n7863 ;
  assign n7868 = n7867 ^ n7866 ;
  assign n7872 = n7871 ^ n7868 ;
  assign n7873 = n7870 & ~n7872 ;
  assign n7874 = n7873 ^ x901 ;
  assign n7869 = ~n7861 & ~n7868 ;
  assign n7876 = n7874 ^ n7869 ;
  assign n7875 = ~n7869 & ~n7874 ;
  assign n7877 = n7876 ^ n7875 ;
  assign n7881 = n7880 ^ n7877 ;
  assign n7882 = n7881 ^ n7875 ;
  assign n7883 = n7882 ^ x895 ;
  assign n7884 = n7883 ^ n7854 ;
  assign n7885 = n7884 ^ n7856 ;
  assign n7886 = n7885 ^ n7882 ;
  assign n7887 = ~n7857 & n7886 ;
  assign n7888 = n7887 ^ n7883 ;
  assign n7897 = n7896 ^ n7888 ;
  assign n7898 = x896 ^ x895 ;
  assign n7899 = n7898 ^ n7854 ;
  assign n7900 = n7899 ^ n7856 ;
  assign n7901 = n7870 ^ n7858 ;
  assign n7902 = n7901 ^ n7864 ;
  assign n7903 = n7900 & n7902 ;
  assign n7904 = n7903 ^ n7882 ;
  assign n7905 = n7897 & n7904 ;
  assign n7906 = n7905 ^ n7903 ;
  assign n7907 = n7878 ^ n7867 ;
  assign n7908 = n7907 ^ n7879 ;
  assign n7909 = n7881 & n7908 ;
  assign n7912 = n7889 ^ x895 ;
  assign n7915 = n7912 ^ n7891 ;
  assign n7910 = n7889 ^ x896 ;
  assign n7920 = n7915 ^ n7910 ;
  assign n7911 = n7895 ^ n7891 ;
  assign n7913 = n7912 ^ n7911 ;
  assign n7921 = n7920 ^ n7913 ;
  assign n7922 = n7921 ^ n7891 ;
  assign n7924 = n7920 & n7922 ;
  assign n7917 = n7913 ^ n7891 ;
  assign n7918 = n7917 ^ n7890 ;
  assign n7919 = ~n7894 & n7918 ;
  assign n7925 = n7924 ^ n7919 ;
  assign n7926 = n7925 ^ n7917 ;
  assign n7927 = n7924 ^ n7915 ;
  assign n7928 = n7927 ^ n7917 ;
  assign n7929 = n7926 & n7928 ;
  assign n7930 = ~n7891 & n7929 ;
  assign n7931 = n7930 ^ n7924 ;
  assign n7932 = n7931 ^ n7922 ;
  assign n7940 = n7932 ^ n7889 ;
  assign n7943 = n7940 ^ n7910 ;
  assign n7984 = n7909 & ~n7943 ;
  assign n7986 = n7756 & n7850 ;
  assign n8000 = n7984 & ~n7986 ;
  assign n8001 = ~n7906 & n8000 ;
  assign n7944 = n7943 ^ n7909 ;
  assign n7979 = n7944 ^ n7756 ;
  assign n7980 = n7979 ^ n7906 ;
  assign n7981 = n7980 ^ n7851 ;
  assign n7993 = n7986 ^ n7981 ;
  assign n7994 = n7993 ^ n7984 ;
  assign n7995 = n7994 ^ n7906 ;
  assign n7996 = n7995 ^ n7853 ;
  assign n7945 = n7851 ^ n7756 ;
  assign n7946 = n7944 & n7945 ;
  assign n7997 = n7996 ^ n7946 ;
  assign n7948 = n7902 ^ n7900 ;
  assign n7949 = n7845 ^ n7843 ;
  assign n7950 = n7949 ^ n7902 ;
  assign n7951 = n7948 & ~n7950 ;
  assign n7952 = n7951 ^ n7900 ;
  assign n7953 = n7952 ^ n7903 ;
  assign n8016 = n7953 ^ n7846 ;
  assign n8017 = n8016 ^ n7903 ;
  assign n8018 = n8017 ^ n7897 ;
  assign n8019 = n8018 ^ n7841 ;
  assign n7947 = n7846 ^ n7841 ;
  assign n7954 = n7953 ^ n7947 ;
  assign n7961 = n8019 ^ n7954 ;
  assign n7963 = n7961 ^ n7952 ;
  assign n7966 = n7953 & ~n7963 ;
  assign n7967 = n7966 ^ n7961 ;
  assign n7970 = n7966 ^ n7953 ;
  assign n7971 = ~n7841 & n7970 ;
  assign n7972 = n7971 ^ n7846 ;
  assign n7973 = n7972 ^ n7841 ;
  assign n7974 = n7967 & n7973 ;
  assign n7975 = n7974 ^ n7971 ;
  assign n7976 = n7975 ^ n7947 ;
  assign n7985 = n7984 ^ n7906 ;
  assign n7987 = n7986 ^ n7906 ;
  assign n7988 = n7985 & n7987 ;
  assign n7989 = n7988 ^ n7906 ;
  assign n7990 = n7976 & ~n7989 ;
  assign n7991 = n7990 ^ n7906 ;
  assign n7992 = n7981 & ~n7991 ;
  assign n7998 = n7997 ^ n7992 ;
  assign n7977 = n7946 & n7976 ;
  assign n7978 = n7906 & n7977 ;
  assign n7999 = n7998 ^ n7978 ;
  assign n8002 = n8001 ^ n7999 ;
  assign n8003 = ~n7853 & ~n8002 ;
  assign n8030 = n8001 ^ n7986 ;
  assign n8033 = n8003 & ~n8030 ;
  assign n7479 = x920 ^ x919 ;
  assign n7468 = ~x923 & ~x924 ;
  assign n7473 = ~x921 & ~x922 ;
  assign n7467 = x922 ^ x921 ;
  assign n7474 = n7473 ^ n7467 ;
  assign n7476 = ~n7468 & ~n7474 ;
  assign n7469 = x924 ^ x923 ;
  assign n7470 = n7469 ^ n7468 ;
  assign n7487 = ~n7470 & ~n7473 ;
  assign n7488 = ~n7476 & ~n7487 ;
  assign n7489 = n7479 & ~n7488 ;
  assign n7471 = n7470 ^ x922 ;
  assign n7472 = ~n7467 & n7471 ;
  assign n7480 = n7472 ^ x920 ;
  assign n7475 = n7474 ^ n7468 ;
  assign n7477 = n7476 ^ n7475 ;
  assign n7481 = n7480 ^ n7477 ;
  assign n7482 = n7479 & n7481 ;
  assign n7483 = n7482 ^ x919 ;
  assign n7478 = ~n7472 & n7477 ;
  assign n7485 = n7483 ^ n7478 ;
  assign n7484 = ~n7478 & ~n7483 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7490 = n7489 ^ n7486 ;
  assign n7654 = n7487 ^ n7476 ;
  assign n7655 = n7654 ^ n7488 ;
  assign n7656 = n7490 & n7655 ;
  assign n7512 = ~x927 & ~x928 ;
  assign n7518 = ~x929 & ~x930 ;
  assign n7519 = ~n7512 & ~n7518 ;
  assign n7501 = x928 ^ x927 ;
  assign n7513 = n7512 ^ n7501 ;
  assign n7514 = x925 & x926 ;
  assign n7515 = x930 & n7514 ;
  assign n7516 = ~n7513 & n7515 ;
  assign n7517 = n7516 ^ n7514 ;
  assign n7520 = n7519 ^ n7517 ;
  assign n7497 = x930 ^ x929 ;
  assign n7523 = n7518 ^ n7497 ;
  assign n7526 = n7513 & n7523 ;
  assign n7527 = n7526 ^ n7517 ;
  assign n7528 = n7520 & ~n7527 ;
  assign n7511 = x926 ^ x925 ;
  assign n7529 = n7528 ^ n7517 ;
  assign n7530 = ~n7511 & n7529 ;
  assign n7531 = n7528 & n7530 ;
  assign n7532 = n7531 ^ n7529 ;
  assign n7647 = n7523 ^ n7513 ;
  assign n7648 = x926 & n7519 ;
  assign n7649 = n7648 ^ n7513 ;
  assign n7650 = n7647 & ~n7649 ;
  assign n7651 = n7650 ^ n7513 ;
  assign n7652 = ~n7532 & ~n7651 ;
  assign n7653 = n7652 ^ n7532 ;
  assign n7657 = n7656 ^ n7653 ;
  assign n7624 = x938 ^ x937 ;
  assign n7573 = x940 ^ x939 ;
  assign n7571 = x942 ^ x941 ;
  assign n7631 = n7573 ^ n7571 ;
  assign n7569 = x941 & x942 ;
  assign n7567 = x939 & x940 ;
  assign n7577 = n7569 ^ n7567 ;
  assign n7632 = n7631 ^ n7577 ;
  assign n7572 = n7571 ^ n7569 ;
  assign n7574 = n7573 ^ n7567 ;
  assign n7575 = n7572 & n7574 ;
  assign n7633 = n7632 ^ n7575 ;
  assign n7634 = n7624 & ~n7633 ;
  assign n7586 = n7575 ^ x937 ;
  assign n7628 = n7586 & n7624 ;
  assign n7625 = n7624 ^ n7567 ;
  assign n7626 = n7625 ^ n7575 ;
  assign n7627 = ~n7577 & ~n7626 ;
  assign n7629 = n7628 ^ n7627 ;
  assign n7630 = n7629 ^ x937 ;
  assign n7636 = n7634 ^ n7630 ;
  assign n7545 = ~x933 & ~x934 ;
  assign n7549 = x936 ^ x935 ;
  assign n7544 = ~x935 & ~x936 ;
  assign n7550 = n7549 ^ n7544 ;
  assign n7551 = ~n7545 & ~n7550 ;
  assign n7546 = x934 ^ x933 ;
  assign n7547 = n7546 ^ n7545 ;
  assign n7548 = ~n7544 & ~n7547 ;
  assign n7553 = n7551 ^ n7548 ;
  assign n7552 = ~n7548 & ~n7551 ;
  assign n7554 = n7553 ^ n7552 ;
  assign n7606 = ~x931 & n7554 ;
  assign n7559 = n7550 ^ n7545 ;
  assign n7560 = n7559 ^ n7551 ;
  assign n7607 = n7560 ^ x932 ;
  assign n7556 = n7547 ^ n7544 ;
  assign n7557 = n7556 ^ n7548 ;
  assign n7608 = n7557 ^ x932 ;
  assign n7609 = n7607 & n7608 ;
  assign n7610 = n7609 ^ x932 ;
  assign n7611 = n7606 & n7610 ;
  assign n7612 = n7611 ^ x931 ;
  assign n7619 = ~x932 & n7545 ;
  assign n7620 = ~n7557 & n7619 ;
  assign n7621 = n7620 ^ n7557 ;
  assign n7555 = x932 ^ x931 ;
  assign n7558 = n7557 ^ n7554 ;
  assign n7561 = x932 & n7560 ;
  assign n7562 = ~n7558 & n7561 ;
  assign n7563 = n7562 ^ n7552 ;
  assign n7564 = ~n7555 & ~n7563 ;
  assign n7565 = n7564 ^ n7552 ;
  assign n7613 = n7565 ^ n7557 ;
  assign n7622 = n7621 ^ n7613 ;
  assign n7623 = n7612 & n7622 ;
  assign n7637 = n7636 ^ n7623 ;
  assign n7638 = n7555 ^ n7546 ;
  assign n7639 = n7638 ^ n7549 ;
  assign n7640 = n7624 ^ n7573 ;
  assign n7641 = n7640 ^ n7571 ;
  assign n7642 = n7639 & n7641 ;
  assign n7643 = n7642 ^ n7636 ;
  assign n7644 = n7637 & ~n7643 ;
  assign n7645 = n7644 ^ n7642 ;
  assign n7602 = n7577 ^ x938 ;
  assign n7603 = n7602 ^ n7569 ;
  assign n7588 = n7575 ^ n7567 ;
  assign n7570 = n7569 ^ x938 ;
  assign n7579 = n7588 ^ n7570 ;
  assign n7585 = n7579 & n7624 ;
  assign n7594 = n7624 ^ n7585 ;
  assign n7589 = n7588 ^ n7586 ;
  assign n7590 = n7589 ^ n7585 ;
  assign n7591 = ~n7577 & n7590 ;
  assign n7595 = n7594 ^ n7591 ;
  assign n7587 = n7586 ^ n7585 ;
  assign n7592 = x937 & n7591 ;
  assign n7593 = ~n7587 & n7592 ;
  assign n7596 = n7595 ^ n7593 ;
  assign n7601 = n7596 ^ n7567 ;
  assign n7604 = n7603 ^ n7601 ;
  assign n7566 = n7554 & n7565 ;
  assign n7605 = n7604 ^ n7566 ;
  assign n7646 = n7645 ^ n7605 ;
  assign n7658 = n7657 ^ n7646 ;
  assign n7493 = x929 ^ x928 ;
  assign n7498 = ~n7493 & ~n7497 ;
  assign n7492 = x927 ^ x926 ;
  assign n7494 = n7493 ^ x927 ;
  assign n7495 = n7494 ^ x930 ;
  assign n7496 = ~n7492 & n7495 ;
  assign n7499 = n7498 ^ n7496 ;
  assign n7500 = ~x925 & n7499 ;
  assign n7502 = x928 ^ x926 ;
  assign n7503 = x930 ^ x925 ;
  assign n7506 = ~x928 & ~n7503 ;
  assign n7507 = n7506 ^ x925 ;
  assign n7508 = ~n7502 & n7507 ;
  assign n7509 = ~n7501 & n7508 ;
  assign n7510 = ~x929 & n7509 ;
  assign n7533 = ~n7510 & ~n7532 ;
  assign n7534 = ~n7500 & n7533 ;
  assign n7491 = n7490 ^ n7484 ;
  assign n7535 = n7534 ^ n7491 ;
  assign n7536 = n7479 ^ n7467 ;
  assign n7537 = n7536 ^ n7469 ;
  assign n7538 = n7511 ^ n7501 ;
  assign n7539 = n7538 ^ n7497 ;
  assign n7540 = n7537 & n7539 ;
  assign n7541 = n7540 ^ n7534 ;
  assign n7542 = ~n7535 & n7541 ;
  assign n7543 = n7542 ^ n7540 ;
  assign n7659 = n7658 ^ n7543 ;
  assign n7663 = n7642 ^ n7637 ;
  assign n7665 = n7540 ^ n7535 ;
  assign n7668 = ~n7663 & n7665 ;
  assign n7660 = n7539 ^ n7537 ;
  assign n7661 = n7641 ^ n7639 ;
  assign n7662 = n7660 & n7661 ;
  assign n7664 = n7663 ^ n7540 ;
  assign n7666 = n7665 ^ n7664 ;
  assign n7667 = n7662 & ~n7666 ;
  assign n7669 = n7668 ^ n7667 ;
  assign n7670 = n7659 & n7669 ;
  assign n7671 = n7645 ^ n7604 ;
  assign n7672 = n7605 & n7671 ;
  assign n7677 = n7672 ^ n7605 ;
  assign n7675 = ~n7566 & n7604 ;
  assign n7676 = n7645 & n7675 ;
  assign n7678 = n7677 ^ n7676 ;
  assign n7679 = n7653 & ~n7678 ;
  assign n7673 = n7672 ^ n7645 ;
  assign n7680 = n7679 ^ n7673 ;
  assign n7681 = ~n7656 & n7680 ;
  assign n7674 = n7653 & n7673 ;
  assign n7682 = n7681 ^ n7674 ;
  assign n7683 = n7682 ^ n7676 ;
  assign n7684 = ~n7670 & n7683 ;
  assign n7689 = ~n7543 & n7684 ;
  assign n7690 = n7689 ^ n7669 ;
  assign n7691 = n7659 & n7690 ;
  assign n7692 = n7691 ^ n7684 ;
  assign n7693 = n7692 ^ n7670 ;
  assign n7694 = n7658 ^ n7656 ;
  assign n7695 = n7694 ^ n7679 ;
  assign n7700 = ~n7679 & ~n7695 ;
  assign n7696 = n7695 ^ n7673 ;
  assign n7701 = n7700 ^ n7696 ;
  assign n7702 = ~n7543 & n7701 ;
  assign n7703 = n7702 ^ n7696 ;
  assign n7704 = n7658 & n7703 ;
  assign n7705 = n7704 ^ n7696 ;
  assign n7706 = ~n7693 & ~n7705 ;
  assign n7707 = n7706 ^ n7670 ;
  assign n8004 = n7999 ^ n7707 ;
  assign n8006 = n7981 ^ n7976 ;
  assign n8005 = n7669 ^ n7659 ;
  assign n8007 = n8006 ^ n8005 ;
  assign n8012 = n7949 ^ n7948 ;
  assign n8013 = n7661 ^ n7660 ;
  assign n8014 = n8012 & n8013 ;
  assign n8008 = n7662 ^ n7642 ;
  assign n8009 = n8008 ^ n7540 ;
  assign n8010 = n8009 ^ n7535 ;
  assign n8011 = n8010 ^ n7637 ;
  assign n8015 = n8014 ^ n8011 ;
  assign n8020 = n8019 ^ n8006 ;
  assign n8021 = n8020 ^ n8011 ;
  assign n8022 = n8021 ^ n8006 ;
  assign n8023 = n8015 & n8022 ;
  assign n8024 = n8023 ^ n8020 ;
  assign n8025 = n8007 & ~n8024 ;
  assign n8026 = n8025 ^ n8006 ;
  assign n8027 = n8026 ^ n7999 ;
  assign n8028 = ~n8004 & n8027 ;
  assign n8029 = n8028 ^ n7707 ;
  assign n8031 = n8030 ^ n8029 ;
  assign n8034 = n8033 ^ n8031 ;
  assign n7714 = n7645 & n7653 ;
  assign n7708 = n7707 ^ n7675 ;
  assign n7709 = n7708 ^ n7692 ;
  assign n7715 = n7714 ^ n7709 ;
  assign n7716 = n7707 & n7715 ;
  assign n7717 = n7716 ^ n7709 ;
  assign n7718 = n7717 ^ n7692 ;
  assign n7720 = ~n7705 & ~n7716 ;
  assign n7721 = n7718 & n7720 ;
  assign n7722 = n7721 ^ n7717 ;
  assign n8035 = n8034 ^ n7722 ;
  assign n8320 = ~x867 & ~x868 ;
  assign n8326 = ~x869 & ~x870 ;
  assign n8327 = ~n8320 & ~n8326 ;
  assign n8309 = x868 ^ x867 ;
  assign n8321 = n8320 ^ n8309 ;
  assign n8322 = x865 & x866 ;
  assign n8323 = x870 & n8322 ;
  assign n8324 = ~n8321 & n8323 ;
  assign n8325 = n8324 ^ n8322 ;
  assign n8328 = n8327 ^ n8325 ;
  assign n8305 = x870 ^ x869 ;
  assign n8331 = n8326 ^ n8305 ;
  assign n8334 = n8321 & n8331 ;
  assign n8335 = n8334 ^ n8325 ;
  assign n8336 = n8328 & ~n8335 ;
  assign n8319 = x866 ^ x865 ;
  assign n8337 = n8336 ^ n8325 ;
  assign n8338 = ~n8319 & n8337 ;
  assign n8339 = n8336 & n8338 ;
  assign n8340 = n8339 ^ n8337 ;
  assign n8403 = n8331 ^ n8321 ;
  assign n8404 = x866 & n8327 ;
  assign n8405 = n8404 ^ n8321 ;
  assign n8406 = n8403 & ~n8405 ;
  assign n8407 = n8406 ^ n8321 ;
  assign n8408 = ~n8340 & n8407 ;
  assign n8363 = ~x861 & ~x862 ;
  assign n8369 = ~x863 & ~x864 ;
  assign n8370 = ~n8363 & ~n8369 ;
  assign n8352 = x862 ^ x861 ;
  assign n8364 = n8363 ^ n8352 ;
  assign n8365 = x859 & x860 ;
  assign n8366 = x864 & n8365 ;
  assign n8367 = ~n8364 & n8366 ;
  assign n8368 = n8367 ^ n8365 ;
  assign n8371 = n8370 ^ n8368 ;
  assign n8348 = x864 ^ x863 ;
  assign n8374 = n8369 ^ n8348 ;
  assign n8377 = n8364 & n8374 ;
  assign n8378 = n8377 ^ n8368 ;
  assign n8379 = n8371 & ~n8378 ;
  assign n8362 = x860 ^ x859 ;
  assign n8380 = n8379 ^ n8368 ;
  assign n8381 = ~n8362 & n8380 ;
  assign n8382 = n8379 & n8381 ;
  assign n8383 = n8382 ^ n8380 ;
  assign n8395 = n8374 ^ n8364 ;
  assign n8396 = x860 & n8370 ;
  assign n8397 = n8396 ^ n8364 ;
  assign n8398 = n8395 & ~n8397 ;
  assign n8399 = n8398 ^ n8364 ;
  assign n8400 = ~n8383 & ~n8399 ;
  assign n8401 = n8400 ^ n8383 ;
  assign n8409 = n8408 ^ n8401 ;
  assign n8344 = x863 ^ x862 ;
  assign n8349 = ~n8344 & ~n8348 ;
  assign n8343 = x861 ^ x860 ;
  assign n8345 = n8344 ^ x861 ;
  assign n8346 = n8345 ^ x864 ;
  assign n8347 = ~n8343 & n8346 ;
  assign n8350 = n8349 ^ n8347 ;
  assign n8351 = ~x859 & n8350 ;
  assign n8353 = x862 ^ x860 ;
  assign n8354 = x864 ^ x859 ;
  assign n8357 = ~x862 & ~n8354 ;
  assign n8358 = n8357 ^ x859 ;
  assign n8359 = ~n8353 & n8358 ;
  assign n8360 = ~n8352 & n8359 ;
  assign n8361 = ~x863 & n8360 ;
  assign n8384 = ~n8361 & ~n8383 ;
  assign n8385 = ~n8351 & n8384 ;
  assign n8301 = x869 ^ x868 ;
  assign n8306 = ~n8301 & ~n8305 ;
  assign n8300 = x867 ^ x866 ;
  assign n8302 = n8301 ^ x867 ;
  assign n8303 = n8302 ^ x870 ;
  assign n8304 = ~n8300 & n8303 ;
  assign n8307 = n8306 ^ n8304 ;
  assign n8308 = ~x865 & n8307 ;
  assign n8310 = x868 ^ x866 ;
  assign n8311 = x870 ^ x865 ;
  assign n8314 = ~x868 & ~n8311 ;
  assign n8315 = n8314 ^ x865 ;
  assign n8316 = ~n8310 & n8315 ;
  assign n8317 = ~n8309 & n8316 ;
  assign n8318 = ~x869 & n8317 ;
  assign n8341 = ~n8318 & ~n8340 ;
  assign n8342 = ~n8308 & n8341 ;
  assign n8386 = n8385 ^ n8342 ;
  assign n8387 = n8319 ^ n8309 ;
  assign n8388 = n8387 ^ n8305 ;
  assign n8389 = n8362 ^ n8352 ;
  assign n8390 = n8389 ^ n8348 ;
  assign n8391 = n8388 & n8390 ;
  assign n8392 = n8391 ^ n8342 ;
  assign n8393 = ~n8386 & n8392 ;
  assign n8394 = n8393 ^ n8391 ;
  assign n8479 = n8409 ^ n8394 ;
  assign n8420 = x858 ^ x857 ;
  assign n8418 = x856 ^ x855 ;
  assign n8417 = x854 ^ x853 ;
  assign n8419 = n8418 ^ n8417 ;
  assign n8421 = n8420 ^ n8419 ;
  assign n8415 = x852 ^ x851 ;
  assign n8413 = x850 ^ x849 ;
  assign n8412 = x848 ^ x847 ;
  assign n8414 = n8413 ^ n8412 ;
  assign n8416 = n8415 ^ n8414 ;
  assign n8422 = n8421 ^ n8416 ;
  assign n8423 = n8390 ^ n8388 ;
  assign n8424 = n8422 & n8423 ;
  assign n8425 = n8424 ^ n8391 ;
  assign n8426 = n8425 ^ n8386 ;
  assign n8452 = ~x855 & ~x856 ;
  assign n8448 = ~x857 & ~x858 ;
  assign n8454 = n8448 ^ n8420 ;
  assign n8459 = n8452 & n8454 ;
  assign n8453 = n8452 ^ n8418 ;
  assign n8467 = n8459 ^ n8453 ;
  assign n8455 = n8454 ^ x856 ;
  assign n8456 = n8418 & n8455 ;
  assign n8457 = n8456 ^ x855 ;
  assign n8458 = n8456 ^ n8455 ;
  assign n8460 = n8459 ^ n8458 ;
  assign n8461 = n8457 & ~n8460 ;
  assign n8463 = x854 & ~n8448 ;
  assign n8464 = n8461 & n8463 ;
  assign n8465 = n8464 ^ n8460 ;
  assign n8468 = n8467 ^ n8465 ;
  assign n8469 = ~x854 & ~n8468 ;
  assign n8466 = n8453 & ~n8465 ;
  assign n8470 = n8469 ^ n8466 ;
  assign n8449 = n8448 ^ n8421 ;
  assign n8450 = n8448 ^ x853 ;
  assign n8451 = ~n8449 & n8450 ;
  assign n8471 = n8470 ^ n8451 ;
  assign n8430 = x851 & x852 ;
  assign n8432 = n8430 ^ n8415 ;
  assign n8428 = x849 & x850 ;
  assign n8429 = n8428 ^ n8413 ;
  assign n8437 = n8432 ^ n8429 ;
  assign n8431 = n8430 ^ n8428 ;
  assign n8433 = n8429 & n8432 ;
  assign n8434 = n8433 ^ n8430 ;
  assign n8435 = ~n8431 & n8434 ;
  assign n8438 = n8437 ^ n8435 ;
  assign n8472 = n8471 ^ n8438 ;
  assign n8436 = n8431 ^ x848 ;
  assign n8443 = n8435 & ~n8436 ;
  assign n8439 = n8438 ^ n8436 ;
  assign n8440 = n8439 ^ n8435 ;
  assign n8445 = n8443 ^ n8440 ;
  assign n8446 = ~n8412 & n8445 ;
  assign n8473 = n8472 ^ n8446 ;
  assign n8447 = n8443 & n8446 ;
  assign n8474 = n8473 ^ n8447 ;
  assign n8427 = n8416 & n8421 ;
  assign n8475 = n8474 ^ n8427 ;
  assign n8476 = n8475 ^ n8424 ;
  assign n8477 = ~n8426 & n8476 ;
  assign n8478 = n8477 ^ n8475 ;
  assign n8480 = n8479 ^ n8478 ;
  assign n8481 = n8478 ^ n8471 ;
  assign n8482 = n8481 ^ n8427 ;
  assign n8483 = n8482 ^ n8478 ;
  assign n8484 = n8474 & n8483 ;
  assign n8485 = n8484 ^ n8481 ;
  assign n8486 = ~n8480 & ~n8485 ;
  assign n8487 = n8486 ^ n8479 ;
  assign n8402 = n8401 ^ n8394 ;
  assign n8410 = n8402 & ~n8409 ;
  assign n8411 = n8410 ^ n8401 ;
  assign n8488 = n8487 ^ n8411 ;
  assign n8522 = x853 & x854 ;
  assign n8523 = ~n8453 & n8522 ;
  assign n8524 = ~x858 & n8523 ;
  assign n8527 = x854 & n8467 ;
  assign n8528 = n8527 ^ n8457 ;
  assign n8529 = ~n8417 & n8528 ;
  assign n8530 = n8529 ^ n8457 ;
  assign n8531 = ~n8448 & n8530 ;
  assign n8532 = ~n8524 & ~n8531 ;
  assign n8533 = ~n8465 & n8532 ;
  assign n8498 = n8434 ^ n8431 ;
  assign n8491 = n8436 ^ n8428 ;
  assign n8503 = n8498 ^ n8491 ;
  assign n8494 = n8436 ^ n8434 ;
  assign n8495 = n8494 ^ x847 ;
  assign n8496 = n8495 ^ n8434 ;
  assign n8504 = n8503 ^ n8496 ;
  assign n8505 = n8504 ^ n8431 ;
  assign n8507 = n8503 & n8505 ;
  assign n8502 = ~n8436 & n8494 ;
  assign n8508 = n8507 ^ n8502 ;
  assign n8509 = n8508 ^ n8412 ;
  assign n8510 = n8507 ^ n8498 ;
  assign n8511 = n8510 ^ n8412 ;
  assign n8512 = n8509 & n8511 ;
  assign n8513 = ~n8431 & n8512 ;
  assign n8514 = n8513 ^ n8507 ;
  assign n8515 = n8514 ^ n8505 ;
  assign n8520 = n8515 ^ n8428 ;
  assign n8489 = n8436 ^ n8430 ;
  assign n8521 = n8520 ^ n8489 ;
  assign n8534 = n8533 ^ n8521 ;
  assign n8547 = n8534 ^ n8479 ;
  assign n8548 = n8547 ^ n8487 ;
  assign n8549 = n8548 ^ n8485 ;
  assign n8550 = n8549 ^ n8411 ;
  assign n8535 = n8533 ^ n8479 ;
  assign n8542 = n8479 & ~n8487 ;
  assign n8543 = n8535 & n8542 ;
  assign n8544 = n8543 ^ n8535 ;
  assign n8545 = n8544 ^ n8485 ;
  assign n8546 = n8534 & ~n8545 ;
  assign n8551 = n8550 ^ n8546 ;
  assign n8558 = n8521 & ~n8533 ;
  assign n8552 = n8551 ^ n8487 ;
  assign n8553 = n8552 ^ n8411 ;
  assign n8559 = n8558 ^ n8553 ;
  assign n8560 = n8551 & ~n8559 ;
  assign n8561 = n8560 ^ n8553 ;
  assign n8562 = n8561 ^ n8411 ;
  assign n8564 = n8488 & ~n8562 ;
  assign n8565 = n8564 ^ n8561 ;
  assign n8038 = x891 & x892 ;
  assign n8036 = x893 & x894 ;
  assign n8041 = n8038 ^ n8036 ;
  assign n8069 = n8041 ^ x890 ;
  assign n8070 = n8069 ^ n8038 ;
  assign n8040 = n8036 ^ x889 ;
  assign n8039 = n8038 ^ x890 ;
  assign n8044 = n8040 ^ n8039 ;
  assign n8045 = x894 ^ x893 ;
  assign n8046 = n8045 ^ n8036 ;
  assign n8047 = x892 ^ x891 ;
  assign n8048 = n8047 ^ n8038 ;
  assign n8049 = n8046 & n8048 ;
  assign n8050 = n8049 ^ n8038 ;
  assign n8042 = n8041 ^ n8040 ;
  assign n8051 = n8050 ^ n8042 ;
  assign n8052 = n8051 ^ n8044 ;
  assign n8053 = n8052 ^ n8041 ;
  assign n8054 = n8044 & n8053 ;
  assign n8060 = n8054 ^ n8051 ;
  assign n8056 = n8051 ^ n8040 ;
  assign n8057 = n8056 ^ n8054 ;
  assign n8058 = ~n8041 & n8057 ;
  assign n8061 = ~n8036 & n8058 ;
  assign n8062 = ~n8060 & n8061 ;
  assign n8055 = n8054 ^ n8053 ;
  assign n8059 = n8058 ^ n8055 ;
  assign n8063 = n8062 ^ n8059 ;
  assign n8068 = n8063 ^ n8036 ;
  assign n8071 = n8070 ^ n8068 ;
  assign n8076 = x886 ^ x885 ;
  assign n8075 = ~x885 & ~x886 ;
  assign n8077 = n8076 ^ n8075 ;
  assign n8073 = x888 ^ x887 ;
  assign n8072 = ~x887 & ~x888 ;
  assign n8074 = n8073 ^ n8072 ;
  assign n8078 = n8077 ^ n8074 ;
  assign n8079 = x884 ^ x883 ;
  assign n8080 = n8079 ^ n8078 ;
  assign n8086 = ~n8072 & ~n8075 ;
  assign n8081 = n8078 ^ x884 ;
  assign n8087 = n8086 ^ n8081 ;
  assign n8088 = ~n8080 & n8087 ;
  assign n8089 = n8088 ^ x883 ;
  assign n8090 = n8089 ^ n8077 ;
  assign n8091 = ~n8078 & ~n8090 ;
  assign n8093 = x883 & x884 ;
  assign n8094 = n8091 & n8093 ;
  assign n8092 = n8091 ^ n8089 ;
  assign n8095 = n8094 ^ n8092 ;
  assign n8096 = ~n8071 & ~n8095 ;
  assign n8109 = n8079 ^ n8076 ;
  assign n8110 = n8109 ^ x887 ;
  assign n8111 = n8077 ^ x888 ;
  assign n8112 = n8110 & n8111 ;
  assign n8103 = x890 ^ x889 ;
  assign n8104 = n8047 ^ x890 ;
  assign n8105 = n8104 ^ n8045 ;
  assign n8106 = n8103 & ~n8105 ;
  assign n8107 = n8106 ^ x889 ;
  assign n8102 = ~n8041 & ~n8050 ;
  assign n8108 = n8107 ^ n8102 ;
  assign n8113 = n8112 ^ n8108 ;
  assign n8097 = x887 ^ x884 ;
  assign n8100 = n8097 ^ n8075 ;
  assign n8101 = x883 & n8100 ;
  assign n8114 = n8113 ^ n8101 ;
  assign n8098 = n8075 ^ x887 ;
  assign n8099 = ~n8097 & n8098 ;
  assign n8115 = n8114 ^ n8099 ;
  assign n8116 = n8109 ^ n8073 ;
  assign n8117 = n8103 ^ n8047 ;
  assign n8118 = n8117 ^ n8045 ;
  assign n8119 = n8116 & n8118 ;
  assign n8120 = n8119 ^ n8108 ;
  assign n8121 = ~n8115 & ~n8120 ;
  assign n8122 = n8121 ^ n8119 ;
  assign n8123 = n8096 & ~n8122 ;
  assign n8127 = n8095 ^ n8071 ;
  assign n8124 = n8071 & n8122 ;
  assign n8125 = n8095 & n8124 ;
  assign n8126 = n8125 ^ n8123 ;
  assign n8128 = n8127 ^ n8126 ;
  assign n8129 = n8128 ^ n8122 ;
  assign n8131 = x879 & x880 ;
  assign n8130 = x881 & x882 ;
  assign n8132 = n8131 ^ n8130 ;
  assign n8179 = x878 ^ x877 ;
  assign n8133 = x882 ^ x881 ;
  assign n8134 = n8133 ^ n8130 ;
  assign n8135 = x880 ^ x879 ;
  assign n8136 = n8135 ^ n8131 ;
  assign n8137 = n8134 & n8136 ;
  assign n8180 = n8137 ^ n8130 ;
  assign n8147 = n8180 ^ n8132 ;
  assign n8139 = n8132 ^ x878 ;
  assign n8140 = n8139 ^ n8131 ;
  assign n8152 = n8147 ^ n8140 ;
  assign n8143 = n8180 ^ n8139 ;
  assign n8144 = n8143 ^ x877 ;
  assign n8145 = n8180 ^ n8144 ;
  assign n8153 = n8152 ^ n8145 ;
  assign n8154 = n8153 ^ n8132 ;
  assign n8156 = n8152 & n8154 ;
  assign n8151 = ~n8139 & n8143 ;
  assign n8157 = n8156 ^ n8151 ;
  assign n8158 = n8179 ^ n8157 ;
  assign n8159 = n8156 ^ n8147 ;
  assign n8160 = n8179 ^ n8159 ;
  assign n8161 = n8158 & n8160 ;
  assign n8162 = ~n8132 & n8161 ;
  assign n8163 = n8162 ^ n8156 ;
  assign n8164 = n8163 ^ n8154 ;
  assign n8169 = n8164 ^ n8130 ;
  assign n8170 = n8169 ^ n8140 ;
  assign n8196 = x874 ^ x873 ;
  assign n8173 = ~x873 & ~x874 ;
  assign n8197 = n8196 ^ n8173 ;
  assign n8198 = n8197 ^ x876 ;
  assign n8199 = x872 ^ x871 ;
  assign n8200 = n8199 ^ n8196 ;
  assign n8201 = n8200 ^ x875 ;
  assign n8202 = n8198 & n8201 ;
  assign n8181 = ~n8132 & n8180 ;
  assign n8188 = ~n8139 & n8181 ;
  assign n8182 = n8136 ^ n8134 ;
  assign n8183 = n8182 ^ n8181 ;
  assign n8184 = n8183 ^ n8139 ;
  assign n8185 = n8184 ^ n8181 ;
  assign n8189 = n8188 ^ n8185 ;
  assign n8190 = ~n8179 & n8189 ;
  assign n8193 = n8188 & n8190 ;
  assign n8191 = n8190 ^ n8183 ;
  assign n8194 = n8193 ^ n8191 ;
  assign n8171 = x875 ^ x872 ;
  assign n8174 = n8173 ^ x875 ;
  assign n8177 = ~n8171 & n8174 ;
  assign n8175 = n8174 ^ x872 ;
  assign n8176 = x871 & n8175 ;
  assign n8178 = n8177 ^ n8176 ;
  assign n8195 = n8194 ^ n8178 ;
  assign n8203 = n8202 ^ n8195 ;
  assign n8204 = n8179 ^ n8135 ;
  assign n8205 = n8204 ^ n8133 ;
  assign n8206 = x876 ^ x875 ;
  assign n8207 = n8206 ^ n8200 ;
  assign n8208 = n8205 & n8207 ;
  assign n8209 = n8208 ^ n8194 ;
  assign n8210 = n8203 & n8209 ;
  assign n8211 = n8210 ^ n8208 ;
  assign n8212 = ~n8170 & ~n8211 ;
  assign n8213 = n8129 & n8212 ;
  assign n8214 = ~n8123 & ~n8213 ;
  assign n8215 = ~x871 & ~x872 ;
  assign n8216 = x876 & ~n8197 ;
  assign n8217 = ~x875 & ~x876 ;
  assign n8218 = ~n8173 & ~n8217 ;
  assign n8219 = n8217 ^ n8206 ;
  assign n8220 = n8197 & n8219 ;
  assign n8221 = ~n8218 & n8220 ;
  assign n8222 = x871 & x872 ;
  assign n8223 = ~n8221 & n8222 ;
  assign n8224 = n8223 ^ x875 ;
  assign n8225 = n8216 & n8224 ;
  assign n8226 = n8225 ^ n8223 ;
  assign n8227 = n8220 ^ n8218 ;
  assign n8228 = n8227 ^ n8221 ;
  assign n8229 = ~n8226 & n8228 ;
  assign n8232 = n8215 & n8229 ;
  assign n8230 = n8229 ^ n8226 ;
  assign n8233 = n8232 ^ n8230 ;
  assign n8234 = n8233 ^ n8170 ;
  assign n8240 = ~n8123 & n8170 ;
  assign n8241 = n8240 ^ n8129 ;
  assign n8242 = ~n8234 & ~n8241 ;
  assign n8237 = n8129 ^ n8125 ;
  assign n8243 = n8242 ^ n8237 ;
  assign n8267 = n8207 ^ n8205 ;
  assign n8268 = n8118 ^ n8116 ;
  assign n8269 = n8268 ^ n8205 ;
  assign n8270 = ~n8267 & n8269 ;
  assign n8271 = n8270 ^ n8268 ;
  assign n8272 = n8271 ^ n8208 ;
  assign n8276 = n8203 ^ n8115 ;
  assign n8277 = n8272 & ~n8276 ;
  assign n8266 = n8119 ^ n8115 ;
  assign n8273 = n8272 ^ n8203 ;
  assign n8274 = n8273 ^ n8271 ;
  assign n8275 = n8266 & ~n8274 ;
  assign n8278 = n8277 ^ n8275 ;
  assign n8283 = n8211 & n8278 ;
  assign n8253 = n8125 & n8170 ;
  assign n8254 = n8253 ^ n8213 ;
  assign n8255 = n8254 ^ n8125 ;
  assign n8244 = n8211 ^ n8170 ;
  assign n8250 = n8126 & ~n8233 ;
  assign n8245 = n8211 ^ n8125 ;
  assign n8251 = n8250 ^ n8245 ;
  assign n8252 = ~n8244 & ~n8251 ;
  assign n8256 = n8255 ^ n8252 ;
  assign n8257 = n8233 & n8256 ;
  assign n8258 = n8257 ^ n8254 ;
  assign n8259 = n8258 ^ n8252 ;
  assign n8260 = n8254 ^ n8233 ;
  assign n8261 = n8260 ^ n8257 ;
  assign n8262 = n8258 ^ n8123 ;
  assign n8263 = ~n8261 & n8262 ;
  assign n8264 = ~n8259 & n8263 ;
  assign n8265 = n8264 ^ n8258 ;
  assign n8284 = n8283 ^ n8265 ;
  assign n8285 = n8243 & ~n8284 ;
  assign n8286 = n8170 & n8233 ;
  assign n8287 = n8285 & n8286 ;
  assign n8288 = n8287 ^ n8285 ;
  assign n8289 = n8214 & ~n8288 ;
  assign n8290 = n8234 ^ n8127 ;
  assign n8291 = n8290 ^ n8122 ;
  assign n8294 = ~n8211 & ~n8265 ;
  assign n8295 = n8294 ^ n8243 ;
  assign n8296 = ~n8278 & n8295 ;
  assign n8297 = n8296 ^ n8243 ;
  assign n8298 = n8291 & n8297 ;
  assign n8299 = n8289 & ~n8298 ;
  assign n8567 = n8565 ^ n8299 ;
  assign n8566 = ~n8299 & n8565 ;
  assign n8568 = n8567 ^ n8566 ;
  assign n8569 = n8035 & ~n8568 ;
  assign n8570 = n8268 ^ n8267 ;
  assign n8571 = n8423 ^ n8422 ;
  assign n8572 = n8570 & n8571 ;
  assign n8573 = n8572 ^ n8119 ;
  assign n8574 = n8573 ^ n8271 ;
  assign n8575 = n8574 ^ n8276 ;
  assign n8577 = n8475 ^ n8426 ;
  assign n8576 = n8547 ^ n8485 ;
  assign n8578 = n8577 ^ n8576 ;
  assign n8579 = n8578 ^ n8572 ;
  assign n8580 = n8579 ^ n8576 ;
  assign n8581 = n8575 & n8580 ;
  assign n8582 = n8581 ^ n8578 ;
  assign n8586 = n8576 ^ n8551 ;
  assign n8583 = n8291 ^ n8211 ;
  assign n8584 = n8583 ^ n8278 ;
  assign n8585 = n8584 ^ n8551 ;
  assign n8587 = n8586 ^ n8585 ;
  assign n8588 = n8582 & n8587 ;
  assign n8589 = n8588 ^ n8586 ;
  assign n8590 = ~n8285 & ~n8298 ;
  assign n8614 = n8590 ^ n8551 ;
  assign n8615 = n8589 & ~n8614 ;
  assign n8616 = n8615 ^ n8551 ;
  assign n8592 = n8027 ^ n7707 ;
  assign n8591 = n8590 ^ n8589 ;
  assign n8593 = n8592 ^ n8591 ;
  assign n8595 = n8577 ^ n8575 ;
  assign n8594 = n8019 ^ n8015 ;
  assign n8596 = n8595 ^ n8594 ;
  assign n8600 = n8571 ^ n8570 ;
  assign n8601 = n8013 ^ n8012 ;
  assign n8602 = n8600 & n8601 ;
  assign n8603 = n8602 ^ n8594 ;
  assign n8604 = ~n8596 & n8603 ;
  assign n8597 = n8584 ^ n8582 ;
  assign n8598 = n8597 ^ n8594 ;
  assign n8605 = n8604 ^ n8598 ;
  assign n8608 = n8597 ^ n8592 ;
  assign n8606 = n8024 ^ n8005 ;
  assign n8607 = n8606 ^ n8592 ;
  assign n8609 = n8608 ^ n8607 ;
  assign n8610 = n8605 & ~n8609 ;
  assign n8611 = n8610 ^ n8608 ;
  assign n8612 = n8593 & ~n8611 ;
  assign n8613 = n8612 ^ n8592 ;
  assign n8618 = n8616 ^ n8613 ;
  assign n8617 = ~n8613 & n8616 ;
  assign n8619 = n8618 ^ n8617 ;
  assign n8620 = n8569 & n8619 ;
  assign n8621 = ~n8035 & ~n8619 ;
  assign n8636 = n8568 & n8621 ;
  assign n8625 = n8566 & ~n8617 ;
  assign n8626 = n8625 ^ n8568 ;
  assign n8627 = ~n8621 & n8626 ;
  assign n8628 = n8627 ^ n8568 ;
  assign n8629 = ~n8035 & ~n8566 ;
  assign n8630 = n8617 & n8629 ;
  assign n8631 = n8029 ^ n7722 ;
  assign n8632 = n8034 & n8631 ;
  assign n8633 = n8632 ^ n7722 ;
  assign n8634 = ~n8630 & ~n8633 ;
  assign n8635 = ~n8628 & n8634 ;
  assign n8637 = n8636 ^ n8635 ;
  assign n8638 = n8637 ^ n8628 ;
  assign n8639 = ~n8620 & ~n8638 ;
  assign n8684 = n8683 ^ n8639 ;
  assign n8643 = n7463 ^ n7441 ;
  assign n8640 = n8630 ^ n8620 ;
  assign n8641 = ~n8628 & ~n8640 ;
  assign n8642 = n8641 ^ n8633 ;
  assign n8644 = n8643 ^ n8642 ;
  assign n8660 = n7360 ^ n6340 ;
  assign n8646 = n8606 ^ n8605 ;
  assign n8661 = n8660 ^ n8646 ;
  assign n8645 = n7355 ^ n7354 ;
  assign n8647 = n8646 ^ n8645 ;
  assign n8649 = n7134 ^ n7133 ;
  assign n8650 = n8649 ^ n7336 ;
  assign n8651 = n8601 ^ n8600 ;
  assign n8652 = n8650 & n8651 ;
  assign n8657 = n8652 ^ n8646 ;
  assign n8648 = n7343 ^ n7132 ;
  assign n8653 = n8652 ^ n8648 ;
  assign n8654 = n8652 ^ n8602 ;
  assign n8655 = n8654 ^ n8596 ;
  assign n8656 = n8653 & ~n8655 ;
  assign n8658 = n8657 ^ n8656 ;
  assign n8659 = n8647 & ~n8658 ;
  assign n8662 = n8661 ^ n8659 ;
  assign n8664 = n7433 ^ n7367 ;
  assign n8666 = n8664 ^ n8660 ;
  assign n8663 = n8611 ^ n8591 ;
  assign n8665 = n8664 ^ n8663 ;
  assign n8667 = n8666 ^ n8665 ;
  assign n8668 = ~n8662 & n8667 ;
  assign n8669 = n8668 ^ n8666 ;
  assign n8673 = n8664 ^ n8643 ;
  assign n8670 = n8567 ^ n8035 ;
  assign n8671 = n8670 ^ n8618 ;
  assign n8672 = n8671 ^ n8643 ;
  assign n8674 = n8673 ^ n8672 ;
  assign n8675 = ~n8669 & n8674 ;
  assign n8676 = n8675 ^ n8673 ;
  assign n8677 = n8644 & ~n8676 ;
  assign n8678 = n8677 ^ n8643 ;
  assign n8722 = n8684 ^ n8678 ;
  assign n8719 = n5757 ^ n5724 ;
  assign n8723 = n8722 ^ n8719 ;
  assign n8717 = n8676 ^ n8642 ;
  assign n8689 = n5754 ^ n5731 ;
  assign n8688 = n8671 ^ n8669 ;
  assign n8690 = n8689 ^ n8688 ;
  assign n8692 = n5752 ^ n5732 ;
  assign n8713 = n8692 ^ n8688 ;
  assign n8691 = n8663 ^ n8662 ;
  assign n8693 = n8692 ^ n8691 ;
  assign n8698 = n8655 ^ n8648 ;
  assign n8696 = n8651 ^ n8650 ;
  assign n8697 = ~n5741 & n8696 ;
  assign n8704 = n8697 ^ n5742 ;
  assign n8700 = ~n5740 & n8696 ;
  assign n8705 = n8704 ^ n8700 ;
  assign n8706 = ~n8698 & n8705 ;
  assign n8699 = n8698 ^ n8697 ;
  assign n8701 = n8700 ^ n8699 ;
  assign n8702 = ~n5739 & ~n8701 ;
  assign n8694 = n8658 ^ n8645 ;
  assign n8703 = n8702 ^ n8694 ;
  assign n8707 = n8706 ^ n8703 ;
  assign n8708 = n5749 ^ n5748 ;
  assign n8709 = n8708 ^ n8694 ;
  assign n8710 = n8707 & n8709 ;
  assign n8695 = n8694 ^ n8691 ;
  assign n8711 = n8710 ^ n8695 ;
  assign n8712 = n8693 & n8711 ;
  assign n8714 = n8713 ^ n8712 ;
  assign n8715 = n8690 & n8714 ;
  assign n8716 = n8715 ^ n8689 ;
  assign n8718 = n8717 ^ n8716 ;
  assign n8720 = n8719 ^ n8716 ;
  assign n8721 = n8718 & ~n8720 ;
  assign n8724 = n8723 ^ n8721 ;
  assign n13494 = n8726 ^ n8724 ;
  assign n11860 = x626 ^ x625 ;
  assign n11906 = ~x627 & ~x628 ;
  assign n11862 = x628 ^ x627 ;
  assign n11907 = n11906 ^ n11862 ;
  assign n11903 = x629 & x630 ;
  assign n11859 = x630 ^ x629 ;
  assign n11908 = n11903 ^ n11859 ;
  assign n11910 = ~n11907 & n11908 ;
  assign n11920 = n11903 & ~n11906 ;
  assign n11921 = ~n11910 & ~n11920 ;
  assign n11922 = n11860 & ~n11921 ;
  assign n11904 = n11903 ^ x628 ;
  assign n11905 = ~n11862 & ~n11904 ;
  assign n11913 = n11905 ^ x626 ;
  assign n11909 = n11908 ^ n11907 ;
  assign n11911 = n11910 ^ n11909 ;
  assign n11914 = n11913 ^ n11911 ;
  assign n11915 = n11860 & ~n11914 ;
  assign n11916 = n11915 ^ x625 ;
  assign n11912 = ~n11905 & ~n11911 ;
  assign n11918 = n11916 ^ n11912 ;
  assign n11917 = ~n11912 & ~n11916 ;
  assign n11919 = n11918 ^ n11917 ;
  assign n11923 = n11922 ^ n11919 ;
  assign n11924 = n11923 ^ n11917 ;
  assign n11855 = x620 ^ x619 ;
  assign n11884 = ~x621 & ~x622 ;
  assign n11857 = x622 ^ x621 ;
  assign n11885 = n11884 ^ n11857 ;
  assign n11881 = x623 & x624 ;
  assign n11854 = x624 ^ x623 ;
  assign n11886 = n11881 ^ n11854 ;
  assign n11888 = ~n11885 & n11886 ;
  assign n11898 = n11881 & ~n11884 ;
  assign n11899 = ~n11888 & ~n11898 ;
  assign n11900 = n11855 & ~n11899 ;
  assign n11882 = n11881 ^ x622 ;
  assign n11883 = ~n11857 & ~n11882 ;
  assign n11891 = n11883 ^ x620 ;
  assign n11887 = n11886 ^ n11885 ;
  assign n11889 = n11888 ^ n11887 ;
  assign n11892 = n11891 ^ n11889 ;
  assign n11893 = n11855 & ~n11892 ;
  assign n11894 = n11893 ^ x619 ;
  assign n11890 = ~n11883 & ~n11889 ;
  assign n11896 = n11894 ^ n11890 ;
  assign n11895 = ~n11890 & ~n11894 ;
  assign n11897 = n11896 ^ n11895 ;
  assign n11901 = n11900 ^ n11897 ;
  assign n11902 = n11901 ^ n11895 ;
  assign n11925 = n11924 ^ n11902 ;
  assign n11856 = n11855 ^ n11854 ;
  assign n11858 = n11857 ^ n11856 ;
  assign n11861 = n11860 ^ n11859 ;
  assign n11863 = n11862 ^ n11861 ;
  assign n11864 = n11858 & n11863 ;
  assign n12047 = n11925 ^ n11864 ;
  assign n11869 = x618 ^ x617 ;
  assign n11981 = x617 ^ x616 ;
  assign n11985 = ~n11869 & ~n11981 ;
  assign n11980 = x615 ^ x614 ;
  assign n11982 = n11981 ^ x615 ;
  assign n11983 = n11982 ^ x618 ;
  assign n11984 = ~n11980 & n11983 ;
  assign n11986 = n11985 ^ n11984 ;
  assign n11987 = ~x613 & n11986 ;
  assign n11988 = ~x615 & ~x616 ;
  assign n11994 = ~x617 & ~x618 ;
  assign n11995 = ~n11988 & ~n11994 ;
  assign n11866 = x616 ^ x615 ;
  assign n11989 = n11988 ^ n11866 ;
  assign n11990 = x613 & x614 ;
  assign n11991 = x618 & n11990 ;
  assign n11992 = ~n11989 & n11991 ;
  assign n11993 = n11992 ^ n11990 ;
  assign n11996 = n11995 ^ n11993 ;
  assign n11999 = n11994 ^ n11869 ;
  assign n12002 = n11989 & n11999 ;
  assign n12003 = n12002 ^ n11993 ;
  assign n12004 = n11996 & ~n12003 ;
  assign n11867 = x614 ^ x613 ;
  assign n12005 = n12004 ^ n11993 ;
  assign n12006 = ~n11867 & n12005 ;
  assign n12007 = n12004 & n12006 ;
  assign n12008 = n12007 ^ n12005 ;
  assign n12009 = x616 ^ x614 ;
  assign n12010 = x618 ^ x613 ;
  assign n12013 = ~x616 & ~n12010 ;
  assign n12014 = n12013 ^ x613 ;
  assign n12015 = ~n12009 & n12014 ;
  assign n12016 = ~n11866 & n12015 ;
  assign n12017 = ~x617 & n12016 ;
  assign n12018 = ~n12008 & ~n12017 ;
  assign n12019 = ~n11987 & n12018 ;
  assign n11927 = ~x609 & ~x610 ;
  assign n11872 = x610 ^ x609 ;
  assign n11936 = n11927 ^ n11872 ;
  assign n11934 = ~x611 & ~x612 ;
  assign n11874 = x612 ^ x611 ;
  assign n11935 = n11934 ^ n11874 ;
  assign n11937 = n11936 ^ n11935 ;
  assign n11938 = ~n11927 & ~n11934 ;
  assign n11943 = x608 & n11938 ;
  assign n11944 = n11943 ^ n11935 ;
  assign n11945 = n11937 & n11944 ;
  assign n11946 = n11945 ^ n11936 ;
  assign n11928 = x611 ^ x608 ;
  assign n11931 = n11874 & n11928 ;
  assign n11932 = n11931 ^ x611 ;
  assign n11933 = n11927 & ~n11932 ;
  assign n11947 = n11946 ^ n11933 ;
  assign n11948 = ~x607 & ~n11947 ;
  assign n11949 = x607 & x608 ;
  assign n11950 = x612 & ~n11936 ;
  assign n11951 = n11949 & n11950 ;
  assign n11952 = n11951 ^ n11949 ;
  assign n11953 = n11952 ^ n11938 ;
  assign n11958 = n11935 & n11936 ;
  assign n11959 = n11958 ^ n11952 ;
  assign n11960 = n11953 & ~n11959 ;
  assign n11871 = x608 ^ x607 ;
  assign n11961 = n11960 ^ n11952 ;
  assign n11962 = ~n11871 & n11961 ;
  assign n11963 = n11960 & n11962 ;
  assign n11964 = n11963 ^ n11961 ;
  assign n11873 = n11872 ^ n11871 ;
  assign n11972 = n11873 & n11934 ;
  assign n11973 = ~x608 & n11972 ;
  assign n11974 = n11973 ^ x608 ;
  assign n11965 = ~x611 & n11949 ;
  assign n11966 = n11965 ^ x608 ;
  assign n11975 = n11974 ^ n11966 ;
  assign n11976 = n11936 & n11975 ;
  assign n11977 = n11976 ^ n11965 ;
  assign n11978 = ~n11964 & ~n11977 ;
  assign n11979 = ~n11948 & n11978 ;
  assign n12020 = n12019 ^ n11979 ;
  assign n11868 = n11867 ^ n11866 ;
  assign n11870 = n11869 ^ n11868 ;
  assign n11875 = n11874 ^ n11873 ;
  assign n11879 = n11870 & n11875 ;
  assign n12050 = n12020 ^ n11879 ;
  assign n12051 = n12047 & n12050 ;
  assign n11865 = n11863 ^ n11858 ;
  assign n11876 = n11875 ^ n11870 ;
  assign n11877 = n11865 & n11876 ;
  assign n12048 = n12047 ^ n12020 ;
  assign n12049 = n11877 & n12048 ;
  assign n12052 = n12051 ^ n12049 ;
  assign n12053 = n11999 ^ n11989 ;
  assign n12054 = x614 & n11995 ;
  assign n12055 = n12054 ^ n11989 ;
  assign n12056 = n12053 & ~n12055 ;
  assign n12057 = n12056 ^ n11989 ;
  assign n12058 = ~n12008 & ~n12057 ;
  assign n12059 = n12058 ^ n12008 ;
  assign n12088 = ~n12052 & ~n12059 ;
  assign n12041 = n11979 ^ n11879 ;
  assign n12042 = ~n12020 & n12041 ;
  assign n12043 = n12042 ^ n11879 ;
  assign n12044 = n11946 & ~n11964 ;
  assign n12087 = ~n12043 & n12044 ;
  assign n12089 = n12088 ^ n12087 ;
  assign n12036 = n11920 ^ n11910 ;
  assign n12037 = n12036 ^ n11921 ;
  assign n12038 = n11923 & n12037 ;
  assign n12033 = n11898 ^ n11888 ;
  assign n12034 = n12033 ^ n11899 ;
  assign n12035 = n11901 & n12034 ;
  assign n12039 = n12038 ^ n12035 ;
  assign n12030 = n11902 ^ n11864 ;
  assign n12031 = n11925 & n12030 ;
  assign n12032 = n12031 ^ n11902 ;
  assign n12040 = n12039 ^ n12032 ;
  assign n12190 = n12087 ^ n12040 ;
  assign n12097 = ~n12089 & ~n12190 ;
  assign n12100 = n12097 ^ n12040 ;
  assign n12060 = n12059 ^ n12052 ;
  assign n12045 = n12044 ^ n12043 ;
  assign n12046 = n12045 ^ n12040 ;
  assign n12061 = n12060 ^ n12046 ;
  assign n12090 = n12089 ^ n12040 ;
  assign n12098 = n12061 & n12090 ;
  assign n12101 = n12100 ^ n12098 ;
  assign n12102 = n12038 ^ n12032 ;
  assign n12103 = n12039 & ~n12102 ;
  assign n12104 = n12103 ^ n12038 ;
  assign n12196 = n12101 & n12104 ;
  assign n12192 = ~n12040 & ~n12061 ;
  assign n12193 = n12192 ^ n12087 ;
  assign n12194 = n12089 & ~n12193 ;
  assign n12195 = n12194 ^ n12088 ;
  assign n12197 = n12196 ^ n12195 ;
  assign n12022 = n11876 ^ n11865 ;
  assign n11145 = x652 ^ x651 ;
  assign n11144 = x650 ^ x649 ;
  assign n11197 = n11145 ^ n11144 ;
  assign n11157 = x654 ^ x653 ;
  assign n11214 = n11197 ^ n11157 ;
  assign n11137 = x644 ^ x643 ;
  assign n11122 = x648 ^ x647 ;
  assign n11212 = n11137 ^ n11122 ;
  assign n11125 = x646 ^ x645 ;
  assign n11213 = n11212 ^ n11125 ;
  assign n12023 = n11214 ^ n11213 ;
  assign n11224 = x634 ^ x633 ;
  assign n11222 = x632 ^ x631 ;
  assign n11336 = n11224 ^ n11222 ;
  assign n11235 = x636 ^ x635 ;
  assign n11337 = n11336 ^ n11235 ;
  assign n11254 = x640 ^ x639 ;
  assign n11253 = x638 ^ x637 ;
  assign n11334 = n11254 ^ n11253 ;
  assign n11288 = x642 ^ x641 ;
  assign n11335 = n11334 ^ n11288 ;
  assign n11346 = n11337 ^ n11335 ;
  assign n12024 = n12023 ^ n11346 ;
  assign n12025 = n12022 & n12024 ;
  assign n12062 = n12061 ^ n12025 ;
  assign n11878 = n11877 ^ n11864 ;
  assign n11880 = n11879 ^ n11878 ;
  assign n11926 = n11925 ^ n11880 ;
  assign n12021 = n12020 ^ n11926 ;
  assign n12026 = n12025 ^ n12021 ;
  assign n11343 = n11335 ^ n11214 ;
  assign n11347 = ~n11343 & ~n11346 ;
  assign n11344 = n11343 ^ n11337 ;
  assign n11345 = ~n11213 & n11344 ;
  assign n11348 = n11347 ^ n11345 ;
  assign n11146 = ~x651 & ~x652 ;
  assign n11186 = x653 ^ x650 ;
  assign n11189 = n11157 & n11186 ;
  assign n11190 = n11189 ^ x653 ;
  assign n11191 = n11146 & ~n11190 ;
  assign n11152 = ~x653 & ~x654 ;
  assign n11158 = n11157 ^ n11152 ;
  assign n11147 = n11146 ^ n11145 ;
  assign n11168 = n11158 ^ n11147 ;
  assign n11153 = ~n11146 & ~n11152 ;
  assign n11173 = x650 & n11153 ;
  assign n11174 = n11173 ^ n11158 ;
  assign n11175 = n11168 & n11174 ;
  assign n11176 = n11175 ^ n11147 ;
  assign n11192 = n11191 ^ n11176 ;
  assign n11193 = ~x649 & ~n11192 ;
  assign n11148 = x649 & x650 ;
  assign n11149 = x654 & n11148 ;
  assign n11150 = ~n11147 & n11149 ;
  assign n11151 = n11150 ^ n11148 ;
  assign n11154 = n11153 ^ n11151 ;
  assign n11161 = n11147 & n11158 ;
  assign n11162 = n11161 ^ n11151 ;
  assign n11163 = n11154 & ~n11162 ;
  assign n11164 = n11163 ^ n11151 ;
  assign n11165 = ~n11144 & n11164 ;
  assign n11166 = n11163 & n11165 ;
  assign n11167 = n11166 ^ n11164 ;
  assign n11194 = ~x653 & n11148 ;
  assign n11200 = n11194 ^ n11152 ;
  assign n11203 = n11197 & n11200 ;
  assign n11204 = ~x650 & n11203 ;
  assign n11205 = n11204 ^ x650 ;
  assign n11195 = n11194 ^ x650 ;
  assign n11206 = n11205 ^ n11195 ;
  assign n11207 = n11147 & n11206 ;
  assign n11208 = n11207 ^ n11194 ;
  assign n11209 = ~n11167 & ~n11208 ;
  assign n11210 = ~n11193 & n11209 ;
  assign n11126 = ~x645 & ~x646 ;
  assign n11123 = ~x647 & ~x648 ;
  assign n11134 = n11126 ^ n11123 ;
  assign n11133 = n11123 & n11126 ;
  assign n11135 = n11134 ^ n11133 ;
  assign n11124 = n11123 ^ n11122 ;
  assign n11127 = n11126 ^ n11125 ;
  assign n11129 = n11124 & n11127 ;
  assign n11139 = n11135 ^ n11129 ;
  assign n11181 = n11137 ^ n11123 ;
  assign n11182 = n11181 ^ n11126 ;
  assign n11183 = ~n11133 & ~n11182 ;
  assign n11184 = ~n11139 & ~n11183 ;
  assign n11128 = n11127 ^ n11124 ;
  assign n11130 = n11129 ^ n11128 ;
  assign n11131 = x643 & x644 ;
  assign n11132 = n11130 & n11131 ;
  assign n11136 = n11135 ^ n11132 ;
  assign n11138 = n11137 ^ n11135 ;
  assign n11140 = n11138 & ~n11139 ;
  assign n11141 = ~n11136 & n11140 ;
  assign n11142 = n11141 ^ n11132 ;
  assign n11143 = n11130 & ~n11142 ;
  assign n11179 = n11143 ^ n11142 ;
  assign n11180 = n11179 ^ n11131 ;
  assign n11185 = n11184 ^ n11180 ;
  assign n11211 = n11210 ^ n11185 ;
  assign n11349 = n11348 ^ n11211 ;
  assign n11315 = x635 ^ x634 ;
  assign n11319 = ~n11235 & ~n11315 ;
  assign n11314 = x633 ^ x632 ;
  assign n11316 = n11315 ^ x633 ;
  assign n11317 = n11316 ^ x636 ;
  assign n11318 = ~n11314 & n11317 ;
  assign n11320 = n11319 ^ n11318 ;
  assign n11321 = ~x631 & n11320 ;
  assign n11223 = ~x633 & ~x634 ;
  assign n11230 = ~x635 & ~x636 ;
  assign n11231 = ~n11223 & ~n11230 ;
  assign n11225 = n11224 ^ n11223 ;
  assign n11226 = x631 & x632 ;
  assign n11227 = x636 & n11226 ;
  assign n11228 = ~n11225 & n11227 ;
  assign n11229 = n11228 ^ n11226 ;
  assign n11232 = n11231 ^ n11229 ;
  assign n11236 = n11235 ^ n11230 ;
  assign n11239 = n11225 & n11236 ;
  assign n11240 = n11239 ^ n11229 ;
  assign n11241 = n11232 & ~n11240 ;
  assign n11242 = n11241 ^ n11229 ;
  assign n11243 = ~n11222 & n11242 ;
  assign n11244 = n11241 & n11243 ;
  assign n11245 = n11244 ^ n11242 ;
  assign n11322 = x634 ^ x632 ;
  assign n11323 = x636 ^ x631 ;
  assign n11326 = ~x634 & ~n11323 ;
  assign n11327 = n11326 ^ x631 ;
  assign n11328 = ~n11322 & n11327 ;
  assign n11329 = ~n11224 & n11328 ;
  assign n11330 = ~x635 & n11329 ;
  assign n11331 = ~n11245 & ~n11330 ;
  assign n11332 = ~n11321 & n11331 ;
  assign n11261 = x639 & x640 ;
  assign n11255 = x641 & x642 ;
  assign n11256 = n11255 ^ x640 ;
  assign n11257 = n11254 & ~n11256 ;
  assign n11258 = n11257 ^ x639 ;
  assign n11273 = n11261 ^ n11258 ;
  assign n11262 = n11255 & n11261 ;
  assign n11263 = n11262 ^ n11256 ;
  assign n11264 = n11263 ^ n11257 ;
  assign n11274 = n11273 ^ n11264 ;
  assign n11275 = n11274 ^ n11258 ;
  assign n11278 = x638 & n11275 ;
  assign n11279 = n11278 ^ n11258 ;
  assign n11280 = ~n11253 & n11279 ;
  assign n11265 = x638 & n11264 ;
  assign n11266 = n11265 ^ n11258 ;
  assign n11267 = ~n11253 & n11266 ;
  assign n11268 = n11267 ^ n11258 ;
  assign n11269 = ~x642 & n11268 ;
  assign n11270 = n11269 ^ x642 ;
  assign n11271 = n11270 ^ n11258 ;
  assign n11281 = n11280 ^ n11271 ;
  assign n11282 = n11281 ^ n11270 ;
  assign n11283 = n11281 ^ x642 ;
  assign n11284 = x641 & ~n11283 ;
  assign n11285 = n11282 & n11284 ;
  assign n11286 = n11285 ^ n11283 ;
  assign n11287 = ~x637 & ~n11286 ;
  assign n11289 = n11288 ^ n11255 ;
  assign n11290 = x638 & n11289 ;
  assign n11298 = ~n11264 & ~n11290 ;
  assign n11291 = n11258 & ~n11262 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = n11292 ^ n11258 ;
  assign n11299 = n11298 ^ n11293 ;
  assign n11300 = n11287 & n11299 ;
  assign n11301 = n11300 ^ n11286 ;
  assign n11302 = ~x641 & ~n11301 ;
  assign n11303 = n11261 ^ x638 ;
  assign n11306 = n11254 ^ x637 ;
  assign n11307 = ~x642 & n11306 ;
  assign n11308 = n11307 ^ x637 ;
  assign n11309 = ~n11261 & n11308 ;
  assign n11310 = n11309 ^ x637 ;
  assign n11311 = ~n11303 & n11310 ;
  assign n11312 = n11302 & n11311 ;
  assign n11313 = n11312 ^ n11301 ;
  assign n11333 = n11332 ^ n11313 ;
  assign n12027 = n11349 ^ n11333 ;
  assign n12028 = n12027 ^ n12021 ;
  assign n12029 = n12026 & ~n12028 ;
  assign n12063 = n12062 ^ n12029 ;
  assign n12105 = n12104 ^ n12101 ;
  assign n12107 = n12105 ^ n12061 ;
  assign n11215 = n11213 & n11214 ;
  assign n11216 = n11215 ^ n11185 ;
  assign n11217 = n11211 & ~n11216 ;
  assign n11218 = n11217 ^ n11210 ;
  assign n11177 = ~n11167 & n11176 ;
  assign n11178 = n11177 ^ n11143 ;
  assign n11358 = n11218 ^ n11178 ;
  assign n11338 = n11335 & n11337 ;
  assign n11339 = n11338 ^ n11332 ;
  assign n11340 = ~n11333 & n11339 ;
  assign n11341 = n11340 ^ n11332 ;
  assign n12065 = n11358 ^ n11341 ;
  assign n11357 = ~n11286 & ~n11293 ;
  assign n11246 = n11236 ^ n11225 ;
  assign n11247 = x632 & n11231 ;
  assign n11248 = n11247 ^ n11225 ;
  assign n11249 = n11246 & ~n11248 ;
  assign n11250 = n11249 ^ n11225 ;
  assign n11251 = ~n11245 & ~n11250 ;
  assign n11252 = n11251 ^ n11245 ;
  assign n12064 = n11357 ^ n11252 ;
  assign n12066 = n12065 ^ n12064 ;
  assign n11352 = n11349 ^ n11338 ;
  assign n11353 = ~n11333 & ~n11352 ;
  assign n11350 = n11215 ^ n11211 ;
  assign n11351 = n11349 & n11350 ;
  assign n11354 = n11353 ^ n11351 ;
  assign n12067 = n12066 ^ n11354 ;
  assign n12106 = n12105 ^ n12067 ;
  assign n12108 = n12107 ^ n12106 ;
  assign n12109 = ~n12063 & n12108 ;
  assign n12110 = n12109 ^ n12107 ;
  assign n11359 = n11358 ^ n11357 ;
  assign n11360 = n11357 ^ n11341 ;
  assign n11355 = n11354 ^ n11252 ;
  assign n11361 = n11360 ^ n11355 ;
  assign n11362 = n11359 & ~n11361 ;
  assign n11219 = n11218 ^ n11143 ;
  assign n11220 = n11178 & ~n11219 ;
  assign n11221 = n11220 ^ n11143 ;
  assign n11363 = n11362 ^ n11221 ;
  assign n11342 = n11341 ^ n11252 ;
  assign n11356 = ~n11342 & ~n11355 ;
  assign n11364 = n11363 ^ n11356 ;
  assign n12185 = n12105 ^ n11364 ;
  assign n12186 = ~n12110 & ~n12185 ;
  assign n12187 = n12186 ^ n11364 ;
  assign n12198 = n12197 ^ n12187 ;
  assign n12111 = n12110 ^ n11364 ;
  assign n12068 = n12067 ^ n12063 ;
  assign n11561 = ~x591 & ~x592 ;
  assign n11391 = x592 ^ x591 ;
  assign n11801 = n11561 ^ n11391 ;
  assign n11392 = x590 ^ x589 ;
  assign n11565 = x589 & ~n11392 ;
  assign n11813 = x594 & n11565 ;
  assign n11814 = ~n11801 & n11813 ;
  assign n11815 = n11814 ^ n11565 ;
  assign n11394 = x594 ^ x593 ;
  assign n11564 = x593 & ~n11394 ;
  assign n11803 = n11564 ^ n11394 ;
  assign n11804 = ~n11561 & n11803 ;
  assign n11816 = n11815 ^ n11804 ;
  assign n11820 = ~n11564 & n11801 ;
  assign n11821 = n11820 ^ n11804 ;
  assign n11822 = n11816 & n11821 ;
  assign n11802 = n11801 ^ n11564 ;
  assign n11809 = x590 & n11804 ;
  assign n11810 = n11809 ^ n11801 ;
  assign n11811 = ~n11802 & n11810 ;
  assign n11812 = n11811 ^ n11564 ;
  assign n11823 = n11822 ^ n11815 ;
  assign n11824 = ~n11812 & n11823 ;
  assign n11825 = ~n11392 & n11824 ;
  assign n11826 = n11822 & n11825 ;
  assign n11827 = n11826 ^ n11824 ;
  assign n11828 = n11827 ^ n11812 ;
  assign n11512 = x587 & x588 ;
  assign n11387 = x588 ^ x587 ;
  assign n11538 = n11512 ^ n11387 ;
  assign n11539 = n11538 ^ x584 ;
  assign n11510 = ~x585 & ~x586 ;
  assign n11540 = n11539 ^ n11510 ;
  assign n11542 = n11538 ^ n11510 ;
  assign n11541 = n11510 & ~n11538 ;
  assign n11543 = n11542 ^ n11541 ;
  assign n11544 = ~n11540 & ~n11543 ;
  assign n11574 = n11541 ^ x583 ;
  assign n11575 = ~n11544 & ~n11574 ;
  assign n11388 = x586 ^ x585 ;
  assign n11511 = n11510 ^ n11388 ;
  assign n11513 = n11511 & ~n11512 ;
  assign n11516 = x587 ^ x584 ;
  assign n11517 = n11516 ^ x586 ;
  assign n11518 = n11517 ^ x588 ;
  assign n11514 = x587 ^ x585 ;
  assign n11519 = n11518 ^ n11514 ;
  assign n11520 = n11519 ^ x588 ;
  assign n11521 = n11520 ^ x587 ;
  assign n11522 = n11521 ^ n11514 ;
  assign n11526 = n11514 ^ x586 ;
  assign n11527 = n11526 ^ x588 ;
  assign n11528 = n11527 ^ n11514 ;
  assign n11529 = ~n11522 & ~n11528 ;
  assign n11530 = ~x587 & n11529 ;
  assign n11533 = n11530 ^ n11529 ;
  assign n11531 = n11530 ^ n11514 ;
  assign n11532 = n11519 & n11531 ;
  assign n11534 = n11533 ^ n11532 ;
  assign n11535 = n11534 ^ x587 ;
  assign n11558 = x583 & n11535 ;
  assign n11536 = n11535 ^ x583 ;
  assign n11559 = n11558 ^ n11536 ;
  assign n11572 = n11513 & ~n11559 ;
  assign n11566 = n11565 ^ n11564 ;
  assign n11393 = n11392 ^ n11391 ;
  assign n11562 = n11394 ^ n11392 ;
  assign n11563 = n11393 & ~n11562 ;
  assign n11567 = n11566 ^ n11563 ;
  assign n11568 = n11567 ^ n11561 ;
  assign n11537 = n11512 ^ n11511 ;
  assign n11545 = n11540 ^ n11512 ;
  assign n11546 = n11545 ^ n11544 ;
  assign n11547 = ~n11537 & n11546 ;
  assign n11548 = n11547 ^ n11511 ;
  assign n11549 = n11548 ^ n11536 ;
  assign n11550 = n11549 ^ n11535 ;
  assign n11554 = ~n11534 & n11548 ;
  assign n11555 = n11554 ^ x587 ;
  assign n11556 = n11550 & ~n11555 ;
  assign n11557 = n11556 ^ n11536 ;
  assign n11560 = n11559 ^ n11557 ;
  assign n11569 = n11568 ^ n11560 ;
  assign n11573 = n11572 ^ n11569 ;
  assign n11576 = n11575 ^ n11573 ;
  assign n11386 = x584 ^ x583 ;
  assign n11390 = n11527 ^ n11386 ;
  assign n11395 = n11394 ^ n11393 ;
  assign n11425 = n11390 & n11395 ;
  assign n11798 = n11568 ^ n11425 ;
  assign n11799 = n11576 & ~n11798 ;
  assign n11800 = n11799 ^ n11568 ;
  assign n12113 = n11828 ^ n11800 ;
  assign n11829 = n11548 & ~n11558 ;
  assign n12114 = n12113 ^ n11829 ;
  assign n11378 = x600 ^ x599 ;
  assign n11469 = x599 ^ x598 ;
  assign n11473 = ~n11378 & ~n11469 ;
  assign n11468 = x597 ^ x596 ;
  assign n11470 = n11469 ^ x597 ;
  assign n11471 = n11470 ^ x600 ;
  assign n11472 = ~n11468 & n11471 ;
  assign n11474 = n11473 ^ n11472 ;
  assign n11475 = ~x595 & n11474 ;
  assign n11376 = x598 ^ x597 ;
  assign n11476 = x598 ^ x596 ;
  assign n11477 = x600 ^ x595 ;
  assign n11480 = ~x598 & ~n11477 ;
  assign n11481 = n11480 ^ x595 ;
  assign n11482 = ~n11476 & n11481 ;
  assign n11483 = ~n11376 & n11482 ;
  assign n11484 = ~x599 & n11483 ;
  assign n11485 = ~x597 & ~x598 ;
  assign n11491 = ~x599 & ~x600 ;
  assign n11492 = ~n11485 & ~n11491 ;
  assign n11486 = n11485 ^ n11376 ;
  assign n11487 = x595 & x596 ;
  assign n11488 = x600 & n11487 ;
  assign n11489 = ~n11486 & n11488 ;
  assign n11490 = n11489 ^ n11487 ;
  assign n11493 = n11492 ^ n11490 ;
  assign n11496 = n11491 ^ n11378 ;
  assign n11499 = n11486 & n11496 ;
  assign n11500 = n11499 ^ n11490 ;
  assign n11501 = n11493 & ~n11500 ;
  assign n11375 = x596 ^ x595 ;
  assign n11502 = n11501 ^ n11490 ;
  assign n11503 = ~n11375 & n11502 ;
  assign n11504 = n11501 & n11503 ;
  assign n11505 = n11504 ^ n11502 ;
  assign n11506 = ~n11484 & ~n11505 ;
  assign n11507 = ~n11475 & n11506 ;
  assign n11383 = x606 ^ x605 ;
  assign n11429 = x605 ^ x604 ;
  assign n11433 = ~n11383 & ~n11429 ;
  assign n11428 = x603 ^ x602 ;
  assign n11430 = n11429 ^ x603 ;
  assign n11431 = n11430 ^ x606 ;
  assign n11432 = ~n11428 & n11431 ;
  assign n11434 = n11433 ^ n11432 ;
  assign n11435 = ~x601 & n11434 ;
  assign n11381 = x604 ^ x603 ;
  assign n11436 = x604 ^ x602 ;
  assign n11437 = x606 ^ x601 ;
  assign n11440 = ~x604 & ~n11437 ;
  assign n11441 = n11440 ^ x601 ;
  assign n11442 = ~n11436 & n11441 ;
  assign n11443 = ~n11381 & n11442 ;
  assign n11444 = ~x605 & n11443 ;
  assign n11445 = ~x603 & ~x604 ;
  assign n11451 = ~x605 & ~x606 ;
  assign n11452 = ~n11445 & ~n11451 ;
  assign n11446 = n11445 ^ n11381 ;
  assign n11447 = x601 & x602 ;
  assign n11448 = x606 & n11447 ;
  assign n11449 = ~n11446 & n11448 ;
  assign n11450 = n11449 ^ n11447 ;
  assign n11453 = n11452 ^ n11450 ;
  assign n11456 = n11451 ^ n11383 ;
  assign n11459 = n11446 & n11456 ;
  assign n11460 = n11459 ^ n11450 ;
  assign n11461 = n11453 & ~n11460 ;
  assign n11380 = x602 ^ x601 ;
  assign n11462 = n11461 ^ n11450 ;
  assign n11463 = ~n11380 & n11462 ;
  assign n11464 = n11461 & n11463 ;
  assign n11465 = n11464 ^ n11462 ;
  assign n11466 = ~n11444 & ~n11465 ;
  assign n11467 = ~n11435 & n11466 ;
  assign n11508 = n11507 ^ n11467 ;
  assign n11790 = n11508 ^ n11425 ;
  assign n11377 = n11376 ^ n11375 ;
  assign n11379 = n11378 ^ n11377 ;
  assign n11382 = n11381 ^ n11380 ;
  assign n11384 = n11383 ^ n11382 ;
  assign n11789 = n11379 & n11384 ;
  assign n11792 = n11789 ^ n11425 ;
  assign n11796 = n11790 & ~n11792 ;
  assign n11788 = n11576 ^ n11508 ;
  assign n11385 = n11384 ^ n11379 ;
  assign n11396 = n11395 ^ n11390 ;
  assign n11397 = n11396 ^ n11379 ;
  assign n11398 = n11385 & ~n11397 ;
  assign n11399 = n11398 ^ n11384 ;
  assign n11794 = n11508 ^ n11399 ;
  assign n11795 = n11788 & n11794 ;
  assign n11797 = n11796 ^ n11795 ;
  assign n12115 = n12114 ^ n11797 ;
  assign n12117 = n12115 ^ n11829 ;
  assign n11841 = n11456 ^ n11446 ;
  assign n11842 = x602 & n11452 ;
  assign n11843 = n11842 ^ n11446 ;
  assign n11844 = n11841 & ~n11843 ;
  assign n11845 = n11844 ^ n11446 ;
  assign n11846 = ~n11465 & ~n11845 ;
  assign n11847 = n11846 ^ n11465 ;
  assign n11835 = n11496 ^ n11486 ;
  assign n11836 = x596 & n11492 ;
  assign n11837 = n11836 ^ n11486 ;
  assign n11838 = n11835 & ~n11837 ;
  assign n11839 = n11838 ^ n11486 ;
  assign n11840 = ~n11505 & n11839 ;
  assign n11848 = n11847 ^ n11840 ;
  assign n11832 = n11789 ^ n11467 ;
  assign n11833 = n11508 & ~n11832 ;
  assign n11834 = n11833 ^ n11507 ;
  assign n11849 = n11848 ^ n11834 ;
  assign n12116 = n11849 ^ n11829 ;
  assign n12118 = n12117 ^ n12116 ;
  assign n11407 = x574 ^ x573 ;
  assign n11406 = x572 ^ x571 ;
  assign n11408 = n11407 ^ n11406 ;
  assign n11405 = x576 ^ x575 ;
  assign n11409 = n11408 ^ n11405 ;
  assign n11402 = x580 ^ x579 ;
  assign n11401 = x578 ^ x577 ;
  assign n11403 = n11402 ^ n11401 ;
  assign n11400 = x582 ^ x581 ;
  assign n11404 = n11403 ^ n11400 ;
  assign n11410 = n11409 ^ n11404 ;
  assign n11669 = x581 & x582 ;
  assign n11668 = x579 & x580 ;
  assign n11670 = n11669 ^ n11668 ;
  assign n11671 = n11668 ^ n11402 ;
  assign n11672 = n11669 ^ n11400 ;
  assign n11673 = n11671 & n11672 ;
  assign n11674 = n11673 ^ n11669 ;
  assign n11675 = ~n11670 & ~n11674 ;
  assign n11647 = n11402 ^ x578 ;
  assign n11648 = n11647 ^ n11400 ;
  assign n11657 = n11407 ^ x572 ;
  assign n11658 = n11657 ^ n11405 ;
  assign n11659 = n11406 & ~n11658 ;
  assign n11660 = n11659 ^ x571 ;
  assign n11650 = x575 & x576 ;
  assign n11649 = x573 & x574 ;
  assign n11651 = n11650 ^ n11649 ;
  assign n11652 = n11649 ^ n11407 ;
  assign n11653 = n11650 ^ n11405 ;
  assign n11654 = n11652 & n11653 ;
  assign n11655 = n11654 ^ n11650 ;
  assign n11656 = ~n11651 & ~n11655 ;
  assign n11661 = n11660 ^ n11656 ;
  assign n11662 = n11661 ^ x577 ;
  assign n11663 = n11662 ^ n11402 ;
  assign n11664 = n11663 ^ n11400 ;
  assign n11665 = n11664 ^ n11661 ;
  assign n11666 = ~n11648 & n11665 ;
  assign n11667 = n11666 ^ n11662 ;
  assign n11676 = n11675 ^ n11667 ;
  assign n11418 = x560 ^ x559 ;
  assign n11417 = x564 ^ x563 ;
  assign n11419 = n11418 ^ n11417 ;
  assign n11416 = x562 ^ x561 ;
  assign n11420 = n11419 ^ n11416 ;
  assign n11413 = x566 ^ x565 ;
  assign n11412 = x568 ^ x567 ;
  assign n11414 = n11413 ^ n11412 ;
  assign n11411 = x570 ^ x569 ;
  assign n11415 = n11414 ^ n11411 ;
  assign n11421 = n11420 ^ n11415 ;
  assign n11768 = n11421 ^ n11404 ;
  assign n11765 = n11415 & n11420 ;
  assign n11769 = n11768 ^ n11765 ;
  assign n11770 = n11769 ^ n11404 ;
  assign n11773 = ~n11676 & n11770 ;
  assign n11774 = n11773 ^ n11404 ;
  assign n11775 = n11410 & n11774 ;
  assign n11771 = n11676 ^ n11404 ;
  assign n11776 = n11775 ^ n11771 ;
  assign n11642 = n11415 ^ n11409 ;
  assign n11645 = ~n11410 & ~n11642 ;
  assign n11643 = n11642 ^ n11404 ;
  assign n11644 = ~n11420 & n11643 ;
  assign n11646 = n11645 ^ n11644 ;
  assign n11677 = n11676 ^ n11646 ;
  assign n11578 = x569 & x570 ;
  assign n11579 = n11578 ^ n11411 ;
  assign n11580 = ~x567 & ~x568 ;
  assign n11581 = n11580 ^ n11412 ;
  assign n11583 = n11579 & ~n11581 ;
  assign n11582 = n11581 ^ n11579 ;
  assign n11584 = n11583 ^ n11582 ;
  assign n11597 = ~x566 & n11580 ;
  assign n11598 = n11584 & n11597 ;
  assign n11586 = n11580 ^ n11578 ;
  assign n11585 = n11578 & ~n11580 ;
  assign n11587 = n11586 ^ n11585 ;
  assign n11588 = ~n11584 & ~n11587 ;
  assign n11590 = n11585 ^ n11583 ;
  assign n11589 = ~n11583 & ~n11585 ;
  assign n11591 = n11590 ^ n11589 ;
  assign n11592 = x565 & x566 ;
  assign n11593 = n11591 & n11592 ;
  assign n11594 = n11588 & n11593 ;
  assign n11595 = n11413 & ~n11589 ;
  assign n11596 = ~n11594 & ~n11595 ;
  assign n11599 = n11598 ^ n11596 ;
  assign n11600 = ~x565 & n11599 ;
  assign n11601 = n11587 ^ n11584 ;
  assign n11602 = n11591 ^ x566 ;
  assign n11603 = n11602 ^ n11587 ;
  assign n11604 = n11603 ^ n11591 ;
  assign n11605 = ~n11601 & ~n11604 ;
  assign n11606 = n11605 ^ n11602 ;
  assign n11607 = n11600 & n11606 ;
  assign n11608 = n11607 ^ n11599 ;
  assign n11609 = ~x561 & ~x562 ;
  assign n11610 = ~x563 & ~x564 ;
  assign n11611 = ~n11609 & ~n11610 ;
  assign n11612 = n11609 ^ n11416 ;
  assign n11613 = n11610 ^ n11417 ;
  assign n11615 = ~n11612 & ~n11613 ;
  assign n11614 = n11613 ^ n11612 ;
  assign n11616 = n11615 ^ n11614 ;
  assign n11617 = ~n11611 & ~n11616 ;
  assign n11618 = x559 & x560 ;
  assign n11619 = ~n11615 & n11618 ;
  assign n11620 = ~n11617 & n11619 ;
  assign n11621 = n11620 ^ n11618 ;
  assign n11633 = n11610 ^ n11609 ;
  assign n11634 = ~n11418 & ~n11616 ;
  assign n11635 = n11634 ^ n11609 ;
  assign n11636 = n11633 & n11635 ;
  assign n11637 = n11636 ^ n11609 ;
  assign n11626 = n11418 & n11611 ;
  assign n11627 = n11626 ^ n11612 ;
  assign n11631 = n11614 & n11627 ;
  assign n11628 = n11620 ^ n11613 ;
  assign n11632 = n11631 ^ n11628 ;
  assign n11639 = n11637 ^ n11632 ;
  assign n11640 = ~n11621 & ~n11639 ;
  assign n11763 = ~n11608 & n11640 ;
  assign n11641 = n11640 ^ n11608 ;
  assign n11764 = n11763 ^ n11641 ;
  assign n11784 = n11677 & n11764 ;
  assign n11785 = n11776 & n11784 ;
  assign n11779 = ~n11677 & n11763 ;
  assign n11780 = n11779 ^ n11764 ;
  assign n11781 = ~n11776 & ~n11780 ;
  assign n11782 = ~n11765 & n11781 ;
  assign n11783 = n11782 ^ n11779 ;
  assign n11786 = n11785 ^ n11783 ;
  assign n11757 = n11404 & n11409 ;
  assign n11758 = n11757 ^ n11661 ;
  assign n11759 = n11676 & ~n11758 ;
  assign n11760 = n11759 ^ n11661 ;
  assign n11720 = n11649 ^ x571 ;
  assign n11723 = n11720 ^ n11651 ;
  assign n11718 = n11649 ^ x572 ;
  assign n11728 = n11723 ^ n11718 ;
  assign n11719 = n11655 ^ n11651 ;
  assign n11721 = n11720 ^ n11719 ;
  assign n11729 = n11728 ^ n11721 ;
  assign n11730 = n11729 ^ n11651 ;
  assign n11732 = n11728 & n11730 ;
  assign n11725 = n11721 ^ n11651 ;
  assign n11726 = n11725 ^ n11650 ;
  assign n11727 = ~n11654 & n11726 ;
  assign n11733 = n11732 ^ n11727 ;
  assign n11734 = n11733 ^ n11725 ;
  assign n11735 = n11732 ^ n11723 ;
  assign n11736 = n11735 ^ n11725 ;
  assign n11737 = n11734 & n11736 ;
  assign n11738 = ~n11651 & n11737 ;
  assign n11739 = n11738 ^ n11732 ;
  assign n11740 = n11739 ^ n11730 ;
  assign n11748 = n11740 ^ n11649 ;
  assign n11751 = n11748 ^ n11718 ;
  assign n11686 = n11668 ^ x577 ;
  assign n11689 = n11686 ^ n11670 ;
  assign n11684 = n11668 ^ x578 ;
  assign n11694 = n11689 ^ n11684 ;
  assign n11685 = n11674 ^ n11670 ;
  assign n11687 = n11686 ^ n11685 ;
  assign n11695 = n11694 ^ n11687 ;
  assign n11696 = n11695 ^ n11670 ;
  assign n11698 = n11694 & n11696 ;
  assign n11691 = n11687 ^ n11670 ;
  assign n11692 = n11691 ^ n11669 ;
  assign n11693 = ~n11673 & n11692 ;
  assign n11699 = n11698 ^ n11693 ;
  assign n11700 = n11699 ^ n11691 ;
  assign n11701 = n11698 ^ n11689 ;
  assign n11702 = n11701 ^ n11691 ;
  assign n11703 = n11700 & n11702 ;
  assign n11704 = ~n11670 & n11703 ;
  assign n11705 = n11704 ^ n11698 ;
  assign n11706 = n11705 ^ n11696 ;
  assign n11714 = n11706 ^ n11668 ;
  assign n11717 = n11714 ^ n11684 ;
  assign n11752 = n11751 ^ n11717 ;
  assign n11761 = n11760 ^ n11752 ;
  assign n11682 = n11591 & n11596 ;
  assign n11683 = n11682 ^ n11632 ;
  assign n11762 = n11761 ^ n11683 ;
  assign n11787 = n11786 ^ n11762 ;
  assign n11852 = n12118 ^ n11787 ;
  assign n11422 = n11421 ^ n11410 ;
  assign n11423 = n11396 ^ n11385 ;
  assign n11424 = n11422 & n11423 ;
  assign n11426 = n11425 ^ n11424 ;
  assign n11427 = n11426 ^ n11399 ;
  assign n11509 = n11508 ^ n11427 ;
  assign n11577 = n11576 ^ n11509 ;
  assign n11678 = n11677 ^ n11641 ;
  assign n11679 = n11678 ^ n11424 ;
  assign n11680 = n11577 & n11679 ;
  assign n11681 = n11680 ^ n11424 ;
  assign n11853 = n11852 ^ n11681 ;
  assign n12069 = n12068 ^ n11853 ;
  assign n12070 = n12024 ^ n12022 ;
  assign n12071 = n11423 ^ n11422 ;
  assign n12072 = n12071 ^ n12024 ;
  assign n12073 = n12070 & ~n12072 ;
  assign n12074 = n12073 ^ n12022 ;
  assign n12075 = n12074 ^ n12028 ;
  assign n12079 = n11678 ^ n11577 ;
  assign n12080 = n12079 ^ n12028 ;
  assign n12076 = n12025 ^ n11853 ;
  assign n12077 = n12076 ^ n12028 ;
  assign n12078 = n12077 ^ n11853 ;
  assign n12081 = n12080 ^ n12078 ;
  assign n12082 = n12081 ^ n12074 ;
  assign n12083 = n12075 & ~n12082 ;
  assign n12084 = n12083 ^ n12077 ;
  assign n12085 = ~n12069 & n12084 ;
  assign n12086 = n12085 ^ n12068 ;
  assign n12112 = n12111 ^ n12086 ;
  assign n12143 = n11760 ^ n11751 ;
  assign n12144 = ~n11752 & ~n12143 ;
  assign n12145 = n12144 ^ n11760 ;
  assign n12148 = n11761 & ~n12145 ;
  assign n12149 = ~n11632 & ~n11682 ;
  assign n12150 = n12149 ^ n11632 ;
  assign n12151 = n12148 & n12150 ;
  assign n12152 = n12151 ^ n12149 ;
  assign n12146 = ~n11682 & n12145 ;
  assign n12147 = n11786 & n12146 ;
  assign n12153 = n12152 ^ n12147 ;
  assign n12158 = n12145 ^ n11761 ;
  assign n12159 = n12158 ^ n11783 ;
  assign n12160 = n12159 ^ n12145 ;
  assign n12155 = n12153 & ~n12160 ;
  assign n12156 = n12155 ^ n12146 ;
  assign n12157 = n11682 & ~n12156 ;
  assign n12164 = ~n11632 & ~n11785 ;
  assign n12165 = n12164 ^ n11786 ;
  assign n12166 = n12160 & n12165 ;
  assign n12167 = n12166 ^ n12158 ;
  assign n12174 = n11615 & n11785 ;
  assign n12175 = n11752 & n12174 ;
  assign n12176 = n12175 ^ n11752 ;
  assign n12168 = n11752 ^ n11682 ;
  assign n12177 = n12176 ^ n12168 ;
  assign n12178 = n12167 & n12177 ;
  assign n12179 = n12157 & n12178 ;
  assign n12180 = n12179 ^ n12156 ;
  assign n12140 = n11787 ^ n11681 ;
  assign n12141 = ~n11852 & n12140 ;
  assign n12134 = n11847 ^ n11834 ;
  assign n12135 = ~n11848 & n12134 ;
  assign n12136 = n12135 ^ n11847 ;
  assign n12123 = n11828 ^ n11797 ;
  assign n12124 = n12113 & ~n12123 ;
  assign n12130 = ~n11797 & n12124 ;
  assign n12125 = n12124 ^ n12116 ;
  assign n12131 = n12130 ^ n12125 ;
  assign n12132 = ~n12115 & ~n12131 ;
  assign n12133 = n12132 ^ n12125 ;
  assign n12137 = n12136 ^ n12133 ;
  assign n12138 = n12137 ^ n11787 ;
  assign n12142 = n12141 ^ n12138 ;
  assign n12181 = n12180 ^ n12142 ;
  assign n12182 = n12181 ^ n12086 ;
  assign n12183 = ~n12112 & n12182 ;
  assign n12184 = n12183 ^ n12181 ;
  assign n12199 = n12198 ^ n12184 ;
  assign n11365 = n11252 & ~n11357 ;
  assign n11366 = n11364 & n11365 ;
  assign n11367 = n11366 ^ n11364 ;
  assign n11368 = n11221 & ~n11367 ;
  assign n11369 = n11358 ^ n11354 ;
  assign n11370 = n11354 ^ n11341 ;
  assign n11371 = n11369 & n11370 ;
  assign n11372 = n11371 ^ n11354 ;
  assign n11373 = n11368 & ~n11372 ;
  assign n11374 = n11373 ^ n11367 ;
  assign n12200 = n12199 ^ n11374 ;
  assign n12235 = n12133 & ~n12136 ;
  assign n12222 = n11849 ^ n11828 ;
  assign n12223 = n12116 & ~n12222 ;
  assign n12224 = n12223 ^ n11849 ;
  assign n12229 = n12222 ^ n12116 ;
  assign n12230 = n12229 ^ n11849 ;
  assign n12225 = n11800 ^ n11797 ;
  assign n12226 = n12123 ^ n11829 ;
  assign n12227 = n12226 ^ n11849 ;
  assign n12228 = n12225 & n12227 ;
  assign n12231 = n12230 ^ n12228 ;
  assign n12232 = n12224 & ~n12231 ;
  assign n12236 = n12235 ^ n12232 ;
  assign n12215 = n12180 ^ n12137 ;
  assign n12216 = n12142 & n12215 ;
  assign n12217 = n12216 ^ n12137 ;
  assign n12201 = n12149 ^ n12145 ;
  assign n12207 = ~n11761 & ~n11783 ;
  assign n12202 = n12201 ^ n12180 ;
  assign n12208 = n12207 ^ n12202 ;
  assign n12209 = n12145 & ~n12208 ;
  assign n12210 = n12209 ^ n12202 ;
  assign n12211 = n12210 ^ n12145 ;
  assign n12212 = ~n12209 & n12211 ;
  assign n12213 = n12201 & n12212 ;
  assign n12214 = n12213 ^ n12210 ;
  assign n12218 = n12217 ^ n12214 ;
  assign n12237 = n12236 ^ n12218 ;
  assign n12238 = n12237 ^ n12187 ;
  assign n12239 = n12238 ^ n11374 ;
  assign n12240 = n12239 ^ n12238 ;
  assign n12244 = n12184 ^ n11374 ;
  assign n12245 = n12197 ^ n12184 ;
  assign n12246 = n12244 & n12245 ;
  assign n12251 = ~n12240 & n12246 ;
  assign n12252 = n12251 ^ n12238 ;
  assign n12253 = ~n12200 & ~n12252 ;
  assign n12247 = n12246 ^ n12238 ;
  assign n12242 = n12214 & ~n12217 ;
  assign n12241 = ~n12218 & n12236 ;
  assign n12243 = n12242 ^ n12241 ;
  assign n12248 = n12247 ^ n12243 ;
  assign n12254 = n12253 ^ n12248 ;
  assign n13319 = n12197 ^ n11374 ;
  assign n13320 = n13319 ^ n12184 ;
  assign n13321 = n13320 ^ n12238 ;
  assign n13444 = n12243 & ~n13321 ;
  assign n13445 = ~n12184 & n13444 ;
  assign n13446 = ~n12187 & n13445 ;
  assign n13447 = n13446 ^ n13444 ;
  assign n13448 = n13447 ^ n12243 ;
  assign n13449 = ~n12254 & ~n13448 ;
  assign n13450 = ~n11374 & n13449 ;
  assign n13451 = ~n12197 & n13450 ;
  assign n13452 = n13451 ^ n13449 ;
  assign n13453 = n13452 ^ n13448 ;
  assign n12310 = x516 ^ x515 ;
  assign n12308 = x514 ^ x513 ;
  assign n12307 = x512 ^ x511 ;
  assign n12309 = n12308 ^ n12307 ;
  assign n12311 = n12310 ^ n12309 ;
  assign n12305 = x522 ^ x521 ;
  assign n12303 = x520 ^ x519 ;
  assign n12302 = x518 ^ x517 ;
  assign n12304 = n12303 ^ n12302 ;
  assign n12306 = n12305 ^ n12304 ;
  assign n12312 = n12311 ^ n12306 ;
  assign n12321 = x534 ^ x533 ;
  assign n12319 = x532 ^ x531 ;
  assign n12318 = x530 ^ x529 ;
  assign n12320 = n12319 ^ n12318 ;
  assign n12322 = n12321 ^ n12320 ;
  assign n12316 = x528 ^ x527 ;
  assign n12314 = x526 ^ x525 ;
  assign n12313 = x524 ^ x523 ;
  assign n12315 = n12314 ^ n12313 ;
  assign n12317 = n12316 ^ n12315 ;
  assign n12323 = n12322 ^ n12317 ;
  assign n12660 = n12312 & n12323 ;
  assign n12661 = n12317 & n12322 ;
  assign n12652 = x533 & x534 ;
  assign n12651 = x531 & x532 ;
  assign n12653 = n12652 ^ n12651 ;
  assign n12654 = n12651 ^ n12319 ;
  assign n12655 = n12652 ^ n12321 ;
  assign n12656 = n12654 & n12655 ;
  assign n12657 = n12656 ^ n12652 ;
  assign n12658 = ~n12653 & ~n12657 ;
  assign n12641 = x525 & x526 ;
  assign n12640 = x527 & x528 ;
  assign n12642 = n12641 ^ n12640 ;
  assign n12643 = n12640 ^ n12316 ;
  assign n12644 = n12641 ^ n12314 ;
  assign n12645 = n12643 & n12644 ;
  assign n12646 = n12645 ^ n12641 ;
  assign n12647 = ~n12642 & ~n12646 ;
  assign n12636 = n12316 ^ x524 ;
  assign n12637 = n12636 ^ n12314 ;
  assign n12638 = n12313 & ~n12637 ;
  assign n12639 = n12638 ^ x523 ;
  assign n12648 = n12647 ^ n12639 ;
  assign n12649 = n12648 ^ x529 ;
  assign n12633 = n12321 ^ n12319 ;
  assign n12634 = n12633 ^ x530 ;
  assign n12635 = n12318 & ~n12634 ;
  assign n12650 = n12649 ^ n12635 ;
  assign n12659 = n12658 ^ n12650 ;
  assign n12864 = n12661 ^ n12659 ;
  assign n12697 = x515 & x516 ;
  assign n12698 = n12697 ^ n12310 ;
  assign n12699 = x513 & x514 ;
  assign n12700 = n12699 ^ n12308 ;
  assign n12701 = n12698 & n12700 ;
  assign n12714 = n12701 ^ x512 ;
  assign n12702 = n12699 ^ n12697 ;
  assign n12715 = n12714 ^ n12702 ;
  assign n12718 = ~n12701 & ~n12702 ;
  assign n12719 = ~n12715 & n12718 ;
  assign n12710 = x512 & n12701 ;
  assign n12711 = n12710 ^ n12699 ;
  assign n12712 = n12702 & ~n12711 ;
  assign n12713 = n12712 ^ n12697 ;
  assign n12716 = n12715 ^ n12713 ;
  assign n12720 = n12719 ^ n12716 ;
  assign n12705 = ~x511 & ~n12715 ;
  assign n12721 = n12720 ^ n12705 ;
  assign n12724 = n12310 ^ n12308 ;
  assign n12703 = n12702 ^ n12701 ;
  assign n12725 = n12724 ^ n12703 ;
  assign n12726 = n12725 ^ n12720 ;
  assign n12727 = n12726 ^ n12705 ;
  assign n12728 = n12307 & n12727 ;
  assign n12729 = n12721 & n12728 ;
  assign n12668 = x519 & x520 ;
  assign n12666 = x521 & x522 ;
  assign n12671 = n12668 ^ n12666 ;
  assign n12667 = n12666 ^ n12305 ;
  assign n12669 = n12668 ^ n12303 ;
  assign n12670 = n12667 & n12669 ;
  assign n12672 = n12671 ^ n12670 ;
  assign n12690 = n12672 ^ x518 ;
  assign n12691 = ~x517 & ~n12690 ;
  assign n12686 = ~n12670 & ~n12671 ;
  assign n12687 = n12686 & ~n12690 ;
  assign n12678 = x518 & n12670 ;
  assign n12679 = n12678 ^ n12668 ;
  assign n12680 = n12671 & ~n12679 ;
  assign n12681 = n12680 ^ n12666 ;
  assign n12684 = n12690 ^ n12681 ;
  assign n12688 = n12687 ^ n12684 ;
  assign n12665 = n12305 ^ n12303 ;
  assign n12673 = n12672 ^ n12665 ;
  assign n12689 = n12688 ^ n12673 ;
  assign n12692 = n12691 ^ n12689 ;
  assign n12693 = n12691 ^ n12688 ;
  assign n12694 = n12302 & n12693 ;
  assign n12695 = n12692 & n12694 ;
  assign n12696 = n12695 ^ n12693 ;
  assign n12722 = n12721 ^ n12696 ;
  assign n12730 = n12729 ^ n12722 ;
  assign n12865 = n12864 ^ n12730 ;
  assign n12663 = n12306 & n12311 ;
  assign n12866 = n12865 ^ n12663 ;
  assign n12867 = n12866 ^ n12660 ;
  assign n12868 = n12867 ^ n12663 ;
  assign n12869 = n12868 ^ n12864 ;
  assign n12870 = ~n12660 & ~n12869 ;
  assign n12871 = n12870 ^ n12663 ;
  assign n12874 = n12870 ^ n12869 ;
  assign n12875 = ~n12659 & ~n12874 ;
  assign n12876 = n12875 ^ n12661 ;
  assign n12877 = n12876 ^ n12659 ;
  assign n12878 = n12871 & n12877 ;
  assign n12879 = n12878 ^ n12875 ;
  assign n12880 = n12879 ^ n12864 ;
  assign n12888 = n12696 ^ n12663 ;
  assign n12889 = ~n12730 & n12888 ;
  assign n12890 = n12889 ^ n12663 ;
  assign n13211 = n12880 & n12890 ;
  assign n12931 = n12640 ^ x523 ;
  assign n12934 = n12931 ^ n12642 ;
  assign n12929 = n12640 ^ x524 ;
  assign n12939 = n12934 ^ n12929 ;
  assign n12930 = n12646 ^ n12642 ;
  assign n12932 = n12931 ^ n12930 ;
  assign n12940 = n12939 ^ n12932 ;
  assign n12941 = n12940 ^ n12642 ;
  assign n12943 = n12939 & n12941 ;
  assign n12936 = n12932 ^ n12642 ;
  assign n12937 = n12936 ^ n12641 ;
  assign n12938 = ~n12645 & n12937 ;
  assign n12944 = n12943 ^ n12938 ;
  assign n12945 = n12944 ^ n12936 ;
  assign n12946 = n12943 ^ n12934 ;
  assign n12947 = n12946 ^ n12936 ;
  assign n12948 = n12945 & n12947 ;
  assign n12949 = ~n12642 & n12948 ;
  assign n12950 = n12949 ^ n12943 ;
  assign n12951 = n12950 ^ n12941 ;
  assign n12959 = n12951 ^ n12640 ;
  assign n12962 = n12959 ^ n12929 ;
  assign n12897 = n12651 ^ x529 ;
  assign n12900 = n12897 ^ n12653 ;
  assign n12895 = n12651 ^ x530 ;
  assign n12905 = n12900 ^ n12895 ;
  assign n12896 = n12657 ^ n12653 ;
  assign n12898 = n12897 ^ n12896 ;
  assign n12906 = n12905 ^ n12898 ;
  assign n12907 = n12906 ^ n12653 ;
  assign n12909 = n12905 & n12907 ;
  assign n12902 = n12898 ^ n12653 ;
  assign n12903 = n12902 ^ n12652 ;
  assign n12904 = ~n12656 & n12903 ;
  assign n12910 = n12909 ^ n12904 ;
  assign n12911 = n12910 ^ n12902 ;
  assign n12912 = n12909 ^ n12900 ;
  assign n12913 = n12912 ^ n12902 ;
  assign n12914 = n12911 & n12913 ;
  assign n12915 = ~n12653 & n12914 ;
  assign n12916 = n12915 ^ n12909 ;
  assign n12917 = n12916 ^ n12907 ;
  assign n12925 = n12917 ^ n12651 ;
  assign n12928 = n12925 ^ n12895 ;
  assign n12963 = n12962 ^ n12928 ;
  assign n12892 = n12661 ^ n12648 ;
  assign n12893 = n12659 & ~n12892 ;
  assign n12894 = n12893 ^ n12648 ;
  assign n12964 = n12963 ^ n12894 ;
  assign n12884 = x511 & ~n12720 ;
  assign n12885 = ~n12713 & n12884 ;
  assign n12886 = n12885 ^ n12713 ;
  assign n13215 = n12964 ^ n12886 ;
  assign n12881 = x517 & ~n12688 ;
  assign n12882 = ~n12681 & n12881 ;
  assign n12883 = n12882 ^ n12681 ;
  assign n13216 = n13215 ^ n12883 ;
  assign n13217 = n13216 ^ n12886 ;
  assign n13210 = n12890 ^ n12880 ;
  assign n13212 = n13211 ^ n13210 ;
  assign n13219 = n13212 ^ n12883 ;
  assign n13221 = n13219 ^ n12886 ;
  assign n13224 = n13221 ^ n13216 ;
  assign n13227 = n13217 & n13224 ;
  assign n13229 = n13227 ^ n12883 ;
  assign n13230 = n13211 & ~n13229 ;
  assign n13235 = n13230 ^ n13227 ;
  assign n13223 = n13221 ^ n13215 ;
  assign n13231 = n13230 ^ n13223 ;
  assign n13232 = n13224 ^ n13215 ;
  assign n13233 = n13232 ^ n13217 ;
  assign n13234 = ~n13231 & n13233 ;
  assign n13236 = n13235 ^ n13234 ;
  assign n13237 = n13236 ^ n13221 ;
  assign n13238 = n13237 ^ n12883 ;
  assign n13239 = n13238 ^ n13216 ;
  assign n13207 = n12962 ^ n12894 ;
  assign n13208 = n12963 & ~n13207 ;
  assign n13209 = n13208 ^ n12962 ;
  assign n13242 = n13239 ^ n13209 ;
  assign n12887 = n12886 ^ n12883 ;
  assign n12891 = n12890 ^ n12887 ;
  assign n12965 = n12964 ^ n12891 ;
  assign n12966 = n12965 ^ n12880 ;
  assign n13243 = n13242 ^ n12966 ;
  assign n12325 = x548 ^ x547 ;
  assign n12327 = x552 ^ x551 ;
  assign n12326 = x550 ^ x549 ;
  assign n12328 = n12327 ^ n12326 ;
  assign n12828 = n12325 & n12328 ;
  assign n12816 = ~x551 & ~x552 ;
  assign n12817 = x549 & ~x550 ;
  assign n12818 = n12816 & n12817 ;
  assign n12819 = n12818 ^ x549 ;
  assign n12829 = n12828 ^ n12819 ;
  assign n12820 = x551 ^ x550 ;
  assign n12821 = ~n12327 & n12820 ;
  assign n12822 = n12821 ^ x550 ;
  assign n13026 = n12829 ^ n12822 ;
  assign n12825 = x549 & x550 ;
  assign n12826 = n12816 ^ n12327 ;
  assign n12827 = n12825 & ~n12826 ;
  assign n13027 = n13026 ^ n12827 ;
  assign n13028 = n13027 ^ n12819 ;
  assign n13029 = n13028 ^ n12827 ;
  assign n12824 = x547 & x548 ;
  assign n13014 = ~n12824 & ~n12827 ;
  assign n13008 = n12828 ^ n12827 ;
  assign n13009 = n13029 ^ n13008 ;
  assign n13015 = n13014 ^ n13009 ;
  assign n13018 = n13014 ^ n12827 ;
  assign n13019 = ~n12829 & ~n13018 ;
  assign n13020 = n13019 ^ n12819 ;
  assign n13021 = n13020 ^ n12829 ;
  assign n13022 = n13015 & ~n13021 ;
  assign n13023 = n13022 ^ n13019 ;
  assign n13024 = n13023 ^ n12827 ;
  assign n13025 = n13024 ^ n12828 ;
  assign n13030 = n13029 ^ n13025 ;
  assign n13031 = n13030 ^ n12828 ;
  assign n12330 = x554 ^ x553 ;
  assign n12791 = ~x555 & ~x556 ;
  assign n12331 = x556 ^ x555 ;
  assign n12792 = n12791 ^ n12331 ;
  assign n12788 = x557 & x558 ;
  assign n12333 = x558 ^ x557 ;
  assign n12793 = n12788 ^ n12333 ;
  assign n12794 = n12792 & ~n12793 ;
  assign n12789 = n12788 ^ x556 ;
  assign n12790 = ~n12331 & ~n12789 ;
  assign n12808 = x554 & ~n12790 ;
  assign n12809 = ~n12794 & n12808 ;
  assign n12810 = n12809 ^ n12794 ;
  assign n12800 = n12333 ^ n12331 ;
  assign n12795 = n12794 ^ n12790 ;
  assign n12801 = n12800 ^ n12795 ;
  assign n12802 = n12801 ^ n12794 ;
  assign n12811 = n12810 ^ n12802 ;
  assign n12812 = ~n12330 & n12811 ;
  assign n12813 = n12812 ^ n12801 ;
  assign n13003 = ~n12788 & n12791 ;
  assign n13004 = n13003 ^ n12790 ;
  assign n13005 = ~n12813 & ~n13004 ;
  assign n13032 = n13031 ^ n13005 ;
  assign n12830 = n12829 ^ n12827 ;
  assign n12831 = n12830 ^ n12824 ;
  assign n12823 = ~n12819 & n12822 ;
  assign n12832 = n12831 ^ n12823 ;
  assign n12814 = n12813 ^ n12790 ;
  assign n12815 = n12814 ^ n12794 ;
  assign n12833 = n12832 ^ n12815 ;
  assign n12796 = n12795 ^ x554 ;
  assign n12797 = ~n12330 & n12796 ;
  assign n12834 = n12833 ^ n12797 ;
  assign n12798 = ~n12794 & ~n12795 ;
  assign n12799 = ~n12797 & n12798 ;
  assign n12835 = n12834 ^ n12799 ;
  assign n12329 = n12328 ^ n12325 ;
  assign n12332 = n12331 ^ n12330 ;
  assign n12334 = n12333 ^ n12332 ;
  assign n12843 = n12329 & n12334 ;
  assign n12996 = n12843 ^ n12832 ;
  assign n12997 = n12835 & n12996 ;
  assign n12998 = n12997 ^ n12832 ;
  assign n13033 = n13032 ^ n12998 ;
  assign n12336 = x536 ^ x535 ;
  assign n12339 = x540 ^ x539 ;
  assign n12337 = x538 ^ x537 ;
  assign n12757 = n12339 ^ n12337 ;
  assign n12734 = x539 & x540 ;
  assign n12736 = n12734 ^ n12339 ;
  assign n12733 = x537 & x538 ;
  assign n12737 = n12733 ^ n12337 ;
  assign n12738 = n12736 & n12737 ;
  assign n12735 = n12734 ^ n12733 ;
  assign n12739 = n12738 ^ n12735 ;
  assign n12758 = n12757 ^ n12739 ;
  assign n12750 = n12738 ^ x536 ;
  assign n12751 = n12750 ^ n12735 ;
  assign n12754 = ~n12735 & ~n12738 ;
  assign n12755 = ~n12751 & n12754 ;
  assign n12746 = x536 & n12738 ;
  assign n12747 = n12746 ^ n12733 ;
  assign n12748 = n12735 & ~n12747 ;
  assign n12749 = n12748 ^ n12734 ;
  assign n12752 = n12751 ^ n12749 ;
  assign n12756 = n12755 ^ n12752 ;
  assign n12759 = n12758 ^ n12756 ;
  assign n12741 = ~x535 & ~n12751 ;
  assign n12760 = n12759 ^ n12741 ;
  assign n12761 = n12336 & n12760 ;
  assign n12762 = n12756 ^ n12741 ;
  assign n12786 = n12761 & n12762 ;
  assign n12763 = ~x545 & ~x546 ;
  assign n12764 = x543 & x544 ;
  assign n12781 = n12763 & ~n12764 ;
  assign n12782 = ~x542 & n12781 ;
  assign n12343 = x544 ^ x543 ;
  assign n12342 = x546 ^ x545 ;
  assign n12344 = n12343 ^ n12342 ;
  assign n12341 = x542 ^ x541 ;
  assign n12345 = n12344 ^ n12341 ;
  assign n12775 = n12345 ^ x541 ;
  assign n12765 = n12763 ^ n12342 ;
  assign n12767 = n12765 ^ x544 ;
  assign n12766 = n12764 & ~n12765 ;
  assign n12776 = n12767 ^ n12766 ;
  assign n12768 = n12343 & n12767 ;
  assign n12777 = n12776 ^ n12768 ;
  assign n12778 = n12777 ^ n12345 ;
  assign n12779 = n12775 & ~n12778 ;
  assign n12769 = n12768 ^ x543 ;
  assign n12770 = ~n12766 & n12769 ;
  assign n12771 = x542 & n12770 ;
  assign n12772 = ~n12763 & n12771 ;
  assign n12773 = n12772 ^ n12770 ;
  assign n12774 = n12773 ^ n12769 ;
  assign n12780 = n12779 ^ n12774 ;
  assign n12783 = n12782 ^ n12780 ;
  assign n12784 = n12783 ^ n12762 ;
  assign n12787 = n12786 ^ n12784 ;
  assign n12338 = n12337 ^ n12336 ;
  assign n12340 = n12339 ^ n12338 ;
  assign n12986 = n12340 & n12345 ;
  assign n12993 = n12986 ^ n12783 ;
  assign n12994 = n12787 & ~n12993 ;
  assign n12995 = n12994 ^ n12986 ;
  assign n13034 = n13033 ^ n12995 ;
  assign n12346 = n12345 ^ n12340 ;
  assign n12836 = n12345 ^ n12334 ;
  assign n12837 = ~n12346 & ~n12836 ;
  assign n12844 = n12843 ^ n12837 ;
  assign n12838 = n12836 ^ n12329 ;
  assign n12839 = n12837 & n12838 ;
  assign n12840 = n12839 ^ n12329 ;
  assign n12841 = n12346 ^ n12334 ;
  assign n12842 = ~n12840 & n12841 ;
  assign n12845 = n12844 ^ n12842 ;
  assign n12984 = ~n12835 & n12845 ;
  assign n12985 = n12984 ^ n12843 ;
  assign n12846 = ~n12840 & n12845 ;
  assign n12847 = n12846 ^ n12835 ;
  assign n12987 = n12986 ^ n12847 ;
  assign n12990 = n12787 & ~n12987 ;
  assign n12991 = n12990 ^ n12986 ;
  assign n12992 = ~n12985 & ~n12991 ;
  assign n13035 = n13034 ^ n12992 ;
  assign n12977 = x541 & ~n12763 ;
  assign n12978 = n12769 & n12977 ;
  assign n12974 = ~n12777 & ~n12781 ;
  assign n12975 = n12974 ^ n12766 ;
  assign n12976 = x541 & n12975 ;
  assign n12979 = n12978 ^ n12976 ;
  assign n12980 = x542 & n12979 ;
  assign n12981 = n12980 ^ n12978 ;
  assign n12982 = ~n12774 & ~n12981 ;
  assign n12967 = x535 & ~n12756 ;
  assign n12968 = ~n12749 & n12967 ;
  assign n12969 = n12968 ^ n12749 ;
  assign n12983 = n12982 ^ n12969 ;
  assign n13036 = n13035 ^ n12983 ;
  assign n13037 = n13036 ^ n12966 ;
  assign n12848 = n12847 ^ n12787 ;
  assign n12849 = n12867 ^ n12848 ;
  assign n12324 = n12323 ^ n12312 ;
  assign n12335 = n12334 ^ n12329 ;
  assign n12347 = n12346 ^ n12335 ;
  assign n12631 = n12324 & n12347 ;
  assign n12859 = n12848 ^ n12631 ;
  assign n12860 = n12849 & n12859 ;
  assign n12861 = n12860 ^ n12848 ;
  assign n13205 = n12966 ^ n12861 ;
  assign n13206 = n13037 & ~n13205 ;
  assign n13244 = n13243 ^ n13206 ;
  assign n13245 = n12992 & n13033 ;
  assign n13250 = ~n12969 & n12982 ;
  assign n13256 = n13035 & n13250 ;
  assign n13249 = ~n12995 & ~n13033 ;
  assign n13257 = n12992 & ~n13249 ;
  assign n13258 = n13256 & ~n13257 ;
  assign n13251 = n13250 ^ n12983 ;
  assign n13254 = n13249 ^ n13034 ;
  assign n13255 = n13251 & ~n13254 ;
  assign n13259 = n13258 ^ n13255 ;
  assign n13252 = ~n12992 & ~n13251 ;
  assign n13253 = n13249 & n13252 ;
  assign n13260 = n13259 ^ n13253 ;
  assign n13246 = n13031 ^ n12998 ;
  assign n13247 = n13032 & ~n13246 ;
  assign n13248 = n13247 ^ n13031 ;
  assign n13263 = n13256 ^ n13253 ;
  assign n13264 = n13248 & ~n13263 ;
  assign n13265 = n13254 ^ n13251 ;
  assign n13266 = n13257 ^ n13254 ;
  assign n13267 = ~n13265 & ~n13266 ;
  assign n13268 = n13267 ^ n13254 ;
  assign n13269 = n13264 & n13268 ;
  assign n13270 = n13269 ^ n13263 ;
  assign n13271 = ~n13260 & ~n13270 ;
  assign n13272 = n13245 & n13271 ;
  assign n13261 = n13260 ^ n13248 ;
  assign n13273 = n13272 ^ n13261 ;
  assign n13287 = n13273 ^ n13242 ;
  assign n13288 = ~n13244 & n13287 ;
  assign n13289 = n13288 ^ n13242 ;
  assign n13277 = ~n12964 & n13212 ;
  assign n13278 = n12883 & n12886 ;
  assign n13279 = n13242 & n13278 ;
  assign n13280 = n13279 ^ n13242 ;
  assign n13282 = n13209 & ~n13280 ;
  assign n13283 = n13282 ^ n13270 ;
  assign n13281 = n13280 ^ n13270 ;
  assign n13284 = n13283 ^ n13281 ;
  assign n13285 = n13277 & ~n13284 ;
  assign n13286 = n13285 ^ n13283 ;
  assign n13290 = n13289 ^ n13286 ;
  assign n12411 = x509 & x510 ;
  assign n12448 = x508 & n12411 ;
  assign n12453 = n12448 ^ x507 ;
  assign n12452 = ~x507 & ~n12448 ;
  assign n12454 = n12453 ^ n12452 ;
  assign n12455 = x505 & x506 ;
  assign n12456 = n12454 & n12455 ;
  assign n12281 = x510 ^ x509 ;
  assign n12449 = n12448 ^ n12281 ;
  assign n12412 = n12411 ^ n12281 ;
  assign n12413 = ~x508 & ~n12412 ;
  assign n12450 = n12449 ^ n12413 ;
  assign n12451 = n12450 ^ x508 ;
  assign n12457 = n12456 ^ n12451 ;
  assign n12279 = x506 ^ x505 ;
  assign n12462 = n12279 & ~n12452 ;
  assign n12458 = n12413 ^ x507 ;
  assign n12414 = ~x507 & n12413 ;
  assign n12459 = n12458 ^ n12414 ;
  assign n12463 = n12462 ^ n12459 ;
  assign n12464 = ~n12451 & ~n12463 ;
  assign n12465 = n12464 ^ n12459 ;
  assign n12466 = ~n12457 & ~n12465 ;
  assign n12467 = n12466 ^ n12456 ;
  assign n12283 = x500 ^ x499 ;
  assign n12416 = x501 & x502 ;
  assign n12284 = x502 ^ x501 ;
  assign n12417 = n12416 ^ n12284 ;
  assign n12418 = x503 & x504 ;
  assign n12286 = x504 ^ x503 ;
  assign n12419 = n12418 ^ n12286 ;
  assign n12420 = n12417 & n12419 ;
  assign n12433 = n12420 ^ x500 ;
  assign n12421 = n12418 ^ n12416 ;
  assign n12434 = n12433 ^ n12421 ;
  assign n12437 = ~n12420 & ~n12421 ;
  assign n12438 = ~n12434 & n12437 ;
  assign n12429 = x500 & n12420 ;
  assign n12430 = n12429 ^ n12418 ;
  assign n12431 = n12421 & ~n12430 ;
  assign n12432 = n12431 ^ n12416 ;
  assign n12435 = n12434 ^ n12432 ;
  assign n12439 = n12438 ^ n12435 ;
  assign n12424 = ~x499 & ~n12434 ;
  assign n12440 = n12439 ^ n12424 ;
  assign n12441 = n12286 ^ n12284 ;
  assign n12422 = n12421 ^ n12420 ;
  assign n12442 = n12441 ^ n12422 ;
  assign n12443 = n12442 ^ n12439 ;
  assign n12444 = n12443 ^ n12424 ;
  assign n12445 = n12440 & n12444 ;
  assign n12446 = n12283 & n12445 ;
  assign n12447 = n12446 ^ n12440 ;
  assign n12468 = n12467 ^ n12447 ;
  assign n12415 = ~x506 & n12414 ;
  assign n12469 = n12468 ^ n12415 ;
  assign n12475 = n12469 ^ n12447 ;
  assign n12470 = n12467 ^ n12414 ;
  assign n12471 = ~x506 & n12451 ;
  assign n12472 = ~n12459 & n12471 ;
  assign n12473 = n12472 ^ n12454 ;
  assign n12474 = ~n12470 & n12473 ;
  assign n12476 = n12475 ^ n12474 ;
  assign n12477 = ~x505 & ~n12476 ;
  assign n12478 = n12477 ^ n12469 ;
  assign n12278 = x508 ^ x507 ;
  assign n12280 = n12279 ^ n12278 ;
  assign n12282 = n12281 ^ n12280 ;
  assign n12285 = n12284 ^ n12283 ;
  assign n12287 = n12286 ^ n12285 ;
  assign n12408 = n12282 & n12287 ;
  assign n13108 = n12478 ^ n12408 ;
  assign n12296 = x492 ^ x491 ;
  assign n12295 = x490 ^ x489 ;
  assign n12297 = n12296 ^ n12295 ;
  assign n12294 = x488 ^ x487 ;
  assign n12298 = n12297 ^ n12294 ;
  assign n12291 = x496 ^ x495 ;
  assign n12290 = x494 ^ x493 ;
  assign n12292 = n12291 ^ n12290 ;
  assign n12289 = x498 ^ x497 ;
  assign n12293 = n12292 ^ n12289 ;
  assign n12299 = n12298 ^ n12293 ;
  assign n12288 = n12287 ^ n12282 ;
  assign n12405 = n12293 ^ n12288 ;
  assign n12406 = n12299 & ~n12405 ;
  assign n12407 = n12406 ^ n12298 ;
  assign n13109 = n13108 ^ n12407 ;
  assign n12352 = x491 & x492 ;
  assign n12353 = ~x489 & ~x490 ;
  assign n12354 = ~n12352 & n12353 ;
  assign n12355 = n12353 ^ n12295 ;
  assign n12356 = n12352 ^ n12296 ;
  assign n12357 = n12355 & ~n12356 ;
  assign n12358 = ~n12354 & ~n12357 ;
  assign n12360 = n12357 ^ n12354 ;
  assign n12361 = n12360 ^ n12358 ;
  assign n12359 = n12352 & ~n12355 ;
  assign n12362 = n12361 ^ n12359 ;
  assign n12363 = n12362 ^ x488 ;
  assign n12364 = ~n12294 & n12363 ;
  assign n12365 = n12358 & n12364 ;
  assign n12366 = n12364 ^ n12362 ;
  assign n12403 = n12365 & ~n12366 ;
  assign n12377 = x497 & x498 ;
  assign n12374 = x495 & x496 ;
  assign n12386 = n12377 ^ n12374 ;
  assign n12381 = ~n12374 & ~n12377 ;
  assign n12387 = n12386 ^ n12381 ;
  assign n12385 = x493 & x494 ;
  assign n12388 = n12385 & n12387 ;
  assign n12375 = n12374 ^ n12291 ;
  assign n12378 = n12377 ^ n12289 ;
  assign n12382 = n12375 & n12378 ;
  assign n12389 = n12388 ^ n12382 ;
  assign n12390 = n12381 ^ n12290 ;
  assign n12391 = n12388 ^ n12381 ;
  assign n12392 = n12390 & ~n12391 ;
  assign n12393 = n12389 & n12392 ;
  assign n12394 = n12393 ^ n12388 ;
  assign n12395 = n12387 & ~n12394 ;
  assign n12396 = n12395 ^ n12394 ;
  assign n12397 = n12396 ^ x493 ;
  assign n12383 = n12382 ^ n12290 ;
  assign n12384 = n12381 & ~n12383 ;
  assign n12398 = n12397 ^ n12384 ;
  assign n12376 = n12375 ^ x494 ;
  assign n12379 = n12378 ^ n12376 ;
  assign n12380 = n12290 & n12379 ;
  assign n12399 = n12398 ^ n12380 ;
  assign n12368 = x488 & ~n12359 ;
  assign n12369 = n12368 ^ n12297 ;
  assign n12370 = ~n12294 & n12369 ;
  assign n12371 = n12370 ^ n12297 ;
  assign n12372 = n12358 & n12371 ;
  assign n12373 = n12366 & ~n12372 ;
  assign n12400 = n12399 ^ n12373 ;
  assign n12404 = n12403 ^ n12400 ;
  assign n13110 = n13109 ^ n12404 ;
  assign n12257 = x472 ^ x471 ;
  assign n12592 = ~x473 & ~x474 ;
  assign n12256 = x474 ^ x473 ;
  assign n12593 = n12592 ^ n12256 ;
  assign n12596 = n12593 ^ x472 ;
  assign n12598 = n12257 & n12596 ;
  assign n12594 = x471 & x472 ;
  assign n12595 = ~n12593 & n12594 ;
  assign n12597 = n12596 ^ n12595 ;
  assign n12599 = n12598 ^ n12597 ;
  assign n12600 = x469 & ~n12599 ;
  assign n12601 = n12598 ^ x471 ;
  assign n12603 = ~n12592 & n12601 ;
  assign n12602 = n12601 ^ n12592 ;
  assign n12604 = n12603 ^ n12602 ;
  assign n12605 = n12604 ^ n12595 ;
  assign n12606 = n12600 & ~n12605 ;
  assign n12607 = n12606 ^ n12603 ;
  assign n12608 = x469 & ~x470 ;
  assign n12609 = n12607 & n12608 ;
  assign n12610 = n12609 ^ n12606 ;
  assign n12611 = ~x470 & n12604 ;
  assign n12612 = n12611 ^ x469 ;
  assign n12613 = x470 & ~n12592 ;
  assign n12622 = n12599 & ~n12613 ;
  assign n12614 = ~n12595 & n12601 ;
  assign n12615 = ~n12613 & n12614 ;
  assign n12616 = n12615 ^ n12601 ;
  assign n12617 = n12616 ^ n12611 ;
  assign n12623 = n12622 ^ n12617 ;
  assign n12624 = ~n12612 & ~n12623 ;
  assign n12625 = n12624 ^ x469 ;
  assign n12626 = ~n12610 & n12625 ;
  assign n12563 = x465 & x466 ;
  assign n12561 = x467 & x468 ;
  assign n12566 = n12563 ^ n12561 ;
  assign n12261 = x468 ^ x467 ;
  assign n12562 = n12561 ^ n12261 ;
  assign n12263 = x466 ^ x465 ;
  assign n12564 = n12563 ^ n12263 ;
  assign n12565 = n12562 & n12564 ;
  assign n12567 = n12566 ^ n12565 ;
  assign n12585 = n12567 ^ x464 ;
  assign n12586 = ~x463 & ~n12585 ;
  assign n12581 = ~n12565 & ~n12566 ;
  assign n12582 = n12581 & ~n12585 ;
  assign n12573 = x464 & n12565 ;
  assign n12574 = n12573 ^ n12563 ;
  assign n12575 = n12566 & ~n12574 ;
  assign n12576 = n12575 ^ n12561 ;
  assign n12579 = n12585 ^ n12576 ;
  assign n12583 = n12582 ^ n12579 ;
  assign n12560 = n12263 ^ n12261 ;
  assign n12568 = n12567 ^ n12560 ;
  assign n12584 = n12583 ^ n12568 ;
  assign n12587 = n12586 ^ n12584 ;
  assign n12260 = x464 ^ x463 ;
  assign n12588 = n12586 ^ n12583 ;
  assign n12589 = n12260 & n12588 ;
  assign n12590 = n12587 & n12589 ;
  assign n12591 = n12590 ^ n12588 ;
  assign n12627 = n12626 ^ n12591 ;
  assign n12258 = n12257 ^ n12256 ;
  assign n12255 = x470 ^ x469 ;
  assign n12259 = n12258 ^ n12255 ;
  assign n12262 = n12261 ^ n12260 ;
  assign n12264 = n12263 ^ n12262 ;
  assign n12480 = n12259 & n12264 ;
  assign n13045 = n12627 ^ n12480 ;
  assign n12269 = x480 ^ x479 ;
  assign n12267 = x478 ^ x477 ;
  assign n12266 = x476 ^ x475 ;
  assign n12268 = n12267 ^ n12266 ;
  assign n12270 = n12269 ^ n12268 ;
  assign n12273 = x482 ^ x481 ;
  assign n12272 = x484 ^ x483 ;
  assign n12274 = n12273 ^ n12272 ;
  assign n12271 = x486 ^ x485 ;
  assign n12275 = n12274 ^ n12271 ;
  assign n12483 = n12270 & n12275 ;
  assign n13046 = n13045 ^ n12483 ;
  assign n12485 = x479 & x480 ;
  assign n12486 = n12485 ^ n12269 ;
  assign n12487 = x477 & x478 ;
  assign n12488 = n12487 ^ n12267 ;
  assign n12489 = n12486 & n12488 ;
  assign n12504 = n12489 ^ x476 ;
  assign n12490 = n12487 ^ n12485 ;
  assign n12505 = n12504 ^ n12490 ;
  assign n12508 = ~n12489 & ~n12490 ;
  assign n12509 = ~n12505 & n12508 ;
  assign n12500 = x476 & n12489 ;
  assign n12501 = n12500 ^ n12487 ;
  assign n12502 = n12490 & ~n12501 ;
  assign n12503 = n12502 ^ n12485 ;
  assign n12506 = n12505 ^ n12503 ;
  assign n12510 = n12509 ^ n12506 ;
  assign n12494 = n12269 ^ n12267 ;
  assign n12491 = n12490 ^ n12489 ;
  assign n12495 = n12494 ^ n12491 ;
  assign n12511 = n12510 ^ n12495 ;
  assign n12493 = ~x475 & ~n12505 ;
  assign n12512 = n12511 ^ n12493 ;
  assign n12513 = n12266 & n12512 ;
  assign n12514 = n12510 ^ n12493 ;
  assign n12557 = n12513 & n12514 ;
  assign n12516 = x485 ^ x484 ;
  assign n12520 = ~n12271 & ~n12516 ;
  assign n12515 = x483 ^ x482 ;
  assign n12517 = n12516 ^ x483 ;
  assign n12518 = n12517 ^ x486 ;
  assign n12519 = ~n12515 & n12518 ;
  assign n12521 = n12520 ^ n12519 ;
  assign n12522 = ~x481 & n12521 ;
  assign n12523 = x484 ^ x482 ;
  assign n12524 = x486 ^ x481 ;
  assign n12527 = ~x484 & ~n12524 ;
  assign n12528 = n12527 ^ x481 ;
  assign n12529 = ~n12523 & n12528 ;
  assign n12530 = ~n12272 & n12529 ;
  assign n12531 = ~x485 & n12530 ;
  assign n12532 = ~x483 & ~x484 ;
  assign n12538 = ~x485 & ~x486 ;
  assign n12539 = ~n12532 & ~n12538 ;
  assign n12533 = n12532 ^ n12272 ;
  assign n12534 = x481 & x482 ;
  assign n12535 = x486 & n12534 ;
  assign n12536 = ~n12533 & n12535 ;
  assign n12537 = n12536 ^ n12534 ;
  assign n12540 = n12539 ^ n12537 ;
  assign n12543 = n12538 ^ n12271 ;
  assign n12546 = n12533 & n12543 ;
  assign n12547 = n12546 ^ n12537 ;
  assign n12548 = n12540 & ~n12547 ;
  assign n12549 = n12548 ^ n12537 ;
  assign n12550 = ~n12273 & n12549 ;
  assign n12551 = n12548 & n12550 ;
  assign n12552 = n12551 ^ n12549 ;
  assign n12553 = ~n12531 & ~n12552 ;
  assign n12554 = ~n12522 & n12553 ;
  assign n12555 = n12554 ^ n12514 ;
  assign n12558 = n12557 ^ n12555 ;
  assign n13047 = n13046 ^ n12558 ;
  assign n12265 = n12264 ^ n12259 ;
  assign n12276 = n12275 ^ n12270 ;
  assign n12481 = n12265 & n12276 ;
  assign n13048 = n13047 ^ n12481 ;
  assign n12629 = n13110 ^ n13048 ;
  assign n12277 = n12276 ^ n12265 ;
  assign n12300 = n12299 ^ n12288 ;
  assign n12350 = n12277 & n12300 ;
  assign n12301 = n12300 ^ n12277 ;
  assign n12348 = n12347 ^ n12324 ;
  assign n12349 = n12301 & n12348 ;
  assign n12351 = n12350 ^ n12349 ;
  assign n12630 = n12629 ^ n12351 ;
  assign n13326 = n12631 ^ n12350 ;
  assign n13327 = n13326 ^ n12349 ;
  assign n13328 = n13327 ^ n12629 ;
  assign n13329 = n13328 ^ n12849 ;
  assign n12855 = n12629 & ~n12849 ;
  assign n12856 = n13329 ^ n12855 ;
  assign n12857 = n12349 & ~n12856 ;
  assign n12858 = n12630 & ~n12857 ;
  assign n13038 = n13037 ^ n12861 ;
  assign n13039 = n13329 ^ n13038 ;
  assign n13040 = n13039 ^ n12857 ;
  assign n13041 = n13040 ^ n13038 ;
  assign n13042 = n13041 ^ n12349 ;
  assign n13043 = n12858 & n13042 ;
  assign n13044 = n13043 ^ n13040 ;
  assign n13068 = x463 & ~n12583 ;
  assign n13069 = ~n12576 & n13068 ;
  assign n13070 = n13069 ^ n12576 ;
  assign n13071 = ~n12610 & ~n12616 ;
  assign n13135 = n13070 & ~n13071 ;
  assign n13072 = n13071 ^ n13070 ;
  assign n13136 = n13135 ^ n13072 ;
  assign n13084 = n12554 ^ n12483 ;
  assign n13085 = ~n12558 & n13084 ;
  assign n13086 = n13085 ^ n12483 ;
  assign n13080 = x475 & ~n12510 ;
  assign n13081 = ~n12503 & n13080 ;
  assign n13082 = n13081 ^ n12503 ;
  assign n13074 = n12543 ^ n12533 ;
  assign n13075 = x482 & n12539 ;
  assign n13076 = n13075 ^ n12533 ;
  assign n13077 = n13074 & ~n13076 ;
  assign n13078 = n13077 ^ n12533 ;
  assign n13079 = ~n12552 & n13078 ;
  assign n13083 = n13082 ^ n13079 ;
  assign n13087 = n13086 ^ n13083 ;
  assign n13065 = n12591 ^ n12480 ;
  assign n13066 = ~n12627 & n13065 ;
  assign n13067 = n13066 ^ n12480 ;
  assign n13161 = n13087 ^ n13067 ;
  assign n13055 = n12481 & ~n12558 ;
  assign n13050 = n13047 ^ n13045 ;
  assign n13056 = n13055 ^ n13050 ;
  assign n13057 = n13048 ^ n12480 ;
  assign n13058 = n13055 ^ n12481 ;
  assign n13059 = n13057 & n13058 ;
  assign n13060 = n13059 ^ n12480 ;
  assign n13061 = n13060 ^ n13057 ;
  assign n13062 = ~n13056 & ~n13061 ;
  assign n13063 = n13062 ^ n13059 ;
  assign n13064 = n13063 ^ n13048 ;
  assign n13137 = n13087 ^ n13064 ;
  assign n13140 = n13137 ^ n13071 ;
  assign n13141 = n13140 ^ n13064 ;
  assign n13145 = n13161 ^ n13141 ;
  assign n13146 = n13145 ^ n13137 ;
  assign n13147 = ~n13072 & ~n13146 ;
  assign n13148 = n13147 ^ n13141 ;
  assign n13151 = n13147 ^ n13146 ;
  assign n13152 = n13064 & ~n13151 ;
  assign n13153 = n13152 ^ n13137 ;
  assign n13154 = ~n13148 & ~n13153 ;
  assign n13073 = n13072 ^ n13067 ;
  assign n13162 = n13073 ^ n13064 ;
  assign n13163 = n13162 ^ n13161 ;
  assign n13164 = n13161 ^ n13073 ;
  assign n13165 = n13164 ^ n13067 ;
  assign n13166 = ~n13163 & n13165 ;
  assign n13167 = n13166 ^ n13067 ;
  assign n13168 = n13067 & n13167 ;
  assign n13169 = ~n13072 & n13168 ;
  assign n13170 = n13169 ^ n13166 ;
  assign n13171 = n13170 ^ n13087 ;
  assign n13172 = n13171 ^ n13072 ;
  assign n13173 = ~n13154 & ~n13172 ;
  assign n13174 = n13136 & n13173 ;
  assign n13155 = n13086 ^ n13082 ;
  assign n13156 = ~n13083 & n13155 ;
  assign n13157 = n13156 ^ n13082 ;
  assign n13158 = n13157 ^ n13154 ;
  assign n13175 = n13174 ^ n13158 ;
  assign n13090 = n12293 & n12298 ;
  assign n13111 = n13110 ^ n13090 ;
  assign n13112 = n13111 ^ n13108 ;
  assign n13113 = ~n12404 & ~n13112 ;
  assign n13114 = n13113 ^ n13090 ;
  assign n13117 = n13113 ^ n13112 ;
  assign n13118 = n12478 & ~n13117 ;
  assign n13119 = n13118 ^ n12408 ;
  assign n13120 = n13119 ^ n12478 ;
  assign n13121 = n13114 & ~n13120 ;
  assign n13122 = n13121 ^ n13118 ;
  assign n13123 = n13122 ^ n13108 ;
  assign n13124 = n13123 ^ n12395 ;
  assign n13100 = x499 & ~n12439 ;
  assign n13101 = ~n12432 & n13100 ;
  assign n13102 = n13101 ^ n12432 ;
  assign n13099 = n12454 & ~n12467 ;
  assign n13103 = n13102 ^ n13099 ;
  assign n13096 = n12447 ^ n12408 ;
  assign n13097 = n12478 & n13096 ;
  assign n13098 = n13097 ^ n12408 ;
  assign n13104 = n13103 ^ n13098 ;
  assign n13094 = n12372 ^ n12359 ;
  assign n13091 = n13090 ^ n12399 ;
  assign n13092 = ~n12404 & n13091 ;
  assign n13093 = n13092 ^ n13090 ;
  assign n13095 = n13094 ^ n13093 ;
  assign n13105 = n13104 ^ n13095 ;
  assign n13125 = n13124 ^ n13105 ;
  assign n13176 = n13175 ^ n13125 ;
  assign n13089 = n13165 ^ n13064 ;
  assign n13177 = n13176 ^ n13089 ;
  assign n13178 = n13177 ^ n13175 ;
  assign n13127 = n13110 ^ n12350 ;
  assign n13128 = ~n12629 & ~n13127 ;
  assign n13129 = n13128 ^ n13110 ;
  assign n13130 = n13178 ^ n13129 ;
  assign n13131 = n13130 ^ n13038 ;
  assign n13132 = n13044 & ~n13131 ;
  assign n13133 = n13132 ^ n13038 ;
  assign n13291 = n13290 ^ n13133 ;
  assign n13198 = n13102 ^ n13098 ;
  assign n13199 = ~n13103 & n13198 ;
  assign n13200 = n13199 ^ n13102 ;
  assign n13181 = n13093 & n13094 ;
  assign n13184 = ~n12395 & ~n13123 ;
  assign n13187 = ~n13181 & ~n13184 ;
  assign n13188 = ~n13093 & n13104 ;
  assign n13193 = ~n13094 & n13188 ;
  assign n13182 = ~n13104 & n13125 ;
  assign n13194 = n13193 ^ n13182 ;
  assign n13195 = n13187 & n13194 ;
  assign n13196 = n13195 ^ n13182 ;
  assign n13201 = n13200 ^ n13196 ;
  assign n13183 = ~n13181 & ~n13182 ;
  assign n13185 = n13184 ^ n13124 ;
  assign n13186 = n13183 & ~n13185 ;
  assign n13197 = n13186 & ~n13196 ;
  assign n13202 = n13201 ^ n13197 ;
  assign n13134 = n13129 ^ n13089 ;
  assign n13179 = ~n13134 & n13178 ;
  assign n13180 = n13179 ^ n13176 ;
  assign n13203 = n13202 ^ n13180 ;
  assign n13204 = n13203 ^ n13133 ;
  assign n13274 = n13273 ^ n13244 ;
  assign n13275 = n13274 ^ n13133 ;
  assign n13276 = ~n13204 & ~n13275 ;
  assign n13292 = n13291 ^ n13276 ;
  assign n13314 = n13202 ^ n13175 ;
  assign n13315 = ~n13180 & n13314 ;
  assign n13316 = n13315 ^ n13202 ;
  assign n13293 = n13185 & ~n13188 ;
  assign n13294 = n13200 & n13293 ;
  assign n13295 = n13294 ^ n13185 ;
  assign n13296 = n13094 & n13295 ;
  assign n13297 = n13202 & n13296 ;
  assign n13299 = n13297 ^ n13294 ;
  assign n13300 = n13299 ^ n13200 ;
  assign n13305 = ~n13183 & n13201 ;
  assign n13308 = ~n13299 & n13305 ;
  assign n13301 = ~n13135 & ~n13175 ;
  assign n13302 = ~n13157 & ~n13301 ;
  assign n13303 = ~n13172 & n13302 ;
  assign n13304 = n13303 ^ n13301 ;
  assign n13306 = n13304 ^ n13299 ;
  assign n13309 = n13308 ^ n13306 ;
  assign n13310 = n13309 ^ n13304 ;
  assign n13311 = n13184 & ~n13310 ;
  assign n13312 = n13300 & n13311 ;
  assign n13313 = n13312 ^ n13309 ;
  assign n13317 = n13316 ^ n13313 ;
  assign n13369 = n13317 ^ n13290 ;
  assign n13370 = ~n13292 & ~n13369 ;
  assign n13371 = n13370 ^ n13290 ;
  assign n13372 = n13289 ^ n13270 ;
  assign n13373 = ~n13286 & ~n13372 ;
  assign n13374 = n13373 ^ n13270 ;
  assign n13375 = n13316 ^ n13304 ;
  assign n13376 = n13313 & n13375 ;
  assign n13377 = n13376 ^ n13316 ;
  assign n13456 = n13374 & n13377 ;
  assign n13457 = n13371 & n13456 ;
  assign n13378 = n13377 ^ n13374 ;
  assign n13458 = n13457 ^ n13378 ;
  assign n13454 = n13377 ^ n13371 ;
  assign n13455 = ~n13378 & n13454 ;
  assign n13459 = n13458 ^ n13455 ;
  assign n13318 = n13317 ^ n13292 ;
  assign n13322 = n13321 ^ n13318 ;
  assign n13362 = n13274 ^ n13204 ;
  assign n13365 = n13362 ^ n13318 ;
  assign n13360 = n12181 ^ n12112 ;
  assign n13324 = n13130 ^ n13044 ;
  assign n13323 = n12084 ^ n12068 ;
  assign n13325 = n13324 ^ n13323 ;
  assign n13332 = n12348 ^ n12301 ;
  assign n13330 = n12071 ^ n12022 ;
  assign n13333 = n13332 ^ n13330 ;
  assign n13349 = n12071 ^ n12070 ;
  assign n13334 = n13333 & n13349 ;
  assign n13335 = n13334 ^ n12071 ;
  assign n13336 = n12022 & n13335 ;
  assign n13337 = ~n13334 & n13336 ;
  assign n13338 = n13337 ^ n13335 ;
  assign n13388 = n13338 ^ n12024 ;
  assign n13389 = n13388 ^ n12070 ;
  assign n13343 = n12022 & n12071 ;
  assign n13344 = n13389 ^ n13343 ;
  assign n13345 = n13329 & n13344 ;
  assign n13346 = n13389 ^ n13345 ;
  assign n13347 = ~n12080 & n13346 ;
  assign n13348 = n13347 ^ n12080 ;
  assign n13350 = n13332 & n13349 ;
  assign n13351 = n13350 ^ n13329 ;
  assign n13352 = n12074 & n12080 ;
  assign n13353 = n13352 ^ n13329 ;
  assign n13354 = ~n13351 & n13353 ;
  assign n13355 = n13354 ^ n13329 ;
  assign n13356 = n13348 & ~n13355 ;
  assign n13357 = n13356 ^ n13324 ;
  assign n13358 = n13325 & ~n13357 ;
  assign n13359 = n13358 ^ n13324 ;
  assign n13361 = n13360 ^ n13359 ;
  assign n13363 = n13362 ^ n13359 ;
  assign n13364 = n13361 & ~n13363 ;
  assign n13366 = n13365 ^ n13364 ;
  assign n13367 = ~n13322 & n13366 ;
  assign n13368 = n13367 ^ n13321 ;
  assign n13460 = n13455 ^ n13371 ;
  assign n13462 = ~n13368 & n13460 ;
  assign n13461 = n13460 ^ n13368 ;
  assign n13463 = n13462 ^ n13461 ;
  assign n13464 = ~n13459 & ~n13463 ;
  assign n13465 = n13453 & n13464 ;
  assign n13466 = n13465 ^ n13463 ;
  assign n13467 = ~n12254 & ~n13466 ;
  assign n13468 = ~n13368 & n13459 ;
  assign n13469 = ~n13453 & ~n13457 ;
  assign n13470 = n13469 ^ n13457 ;
  assign n13471 = n13468 & n13470 ;
  assign n13472 = n13467 & ~n13471 ;
  assign n13487 = ~n13457 & ~n13462 ;
  assign n13473 = n12237 ^ n12197 ;
  assign n13474 = ~n12245 & ~n13473 ;
  assign n13475 = n13474 ^ n12197 ;
  assign n13481 = n13473 ^ n12245 ;
  assign n13482 = n13481 ^ n12197 ;
  assign n13476 = n12187 ^ n11374 ;
  assign n13477 = n12237 ^ n11374 ;
  assign n13478 = n13477 ^ n12184 ;
  assign n13479 = n13478 ^ n12197 ;
  assign n13480 = n13476 & n13479 ;
  assign n13483 = n13482 ^ n13480 ;
  assign n13484 = n13475 & n13483 ;
  assign n13488 = n13487 ^ n13484 ;
  assign n13489 = n12254 & ~n13488 ;
  assign n13490 = n13469 ^ n13453 ;
  assign n13491 = ~n13489 & n13490 ;
  assign n13492 = ~n13472 & n13491 ;
  assign n9769 = x777 & x778 ;
  assign n9767 = x779 & x780 ;
  assign n9772 = n9769 ^ n9767 ;
  assign n9776 = x780 ^ x779 ;
  assign n9777 = n9776 ^ n9767 ;
  assign n9778 = x778 ^ x777 ;
  assign n9779 = n9778 ^ n9769 ;
  assign n9780 = n9777 & n9779 ;
  assign n9781 = n9780 ^ n9769 ;
  assign n9841 = ~n9772 & ~n9781 ;
  assign n9814 = n9776 ^ x776 ;
  assign n9815 = n9814 ^ n9778 ;
  assign n9749 = x786 ^ x785 ;
  assign n9817 = x785 ^ x784 ;
  assign n9821 = ~n9749 & ~n9817 ;
  assign n9816 = x783 ^ x782 ;
  assign n9818 = n9817 ^ x783 ;
  assign n9819 = n9818 ^ x786 ;
  assign n9820 = ~n9816 & n9819 ;
  assign n9822 = n9821 ^ n9820 ;
  assign n9823 = ~x781 & n9822 ;
  assign n9737 = ~x783 & ~x784 ;
  assign n9744 = ~x785 & ~x786 ;
  assign n9745 = ~n9737 & ~n9744 ;
  assign n9738 = x784 ^ x783 ;
  assign n9739 = n9738 ^ n9737 ;
  assign n9740 = x781 & x782 ;
  assign n9741 = x786 & n9740 ;
  assign n9742 = ~n9739 & n9741 ;
  assign n9743 = n9742 ^ n9740 ;
  assign n9746 = n9745 ^ n9743 ;
  assign n9750 = n9749 ^ n9744 ;
  assign n9753 = n9739 & n9750 ;
  assign n9754 = n9753 ^ n9743 ;
  assign n9755 = n9746 & ~n9754 ;
  assign n9736 = x782 ^ x781 ;
  assign n9756 = n9755 ^ n9743 ;
  assign n9757 = ~n9736 & n9756 ;
  assign n9758 = n9755 & n9757 ;
  assign n9759 = n9758 ^ n9756 ;
  assign n9824 = x784 ^ x782 ;
  assign n9825 = x786 ^ x781 ;
  assign n9828 = ~x784 & ~n9825 ;
  assign n9829 = n9828 ^ x781 ;
  assign n9830 = ~n9824 & n9829 ;
  assign n9831 = ~n9738 & n9830 ;
  assign n9832 = ~x785 & n9831 ;
  assign n9833 = ~n9759 & ~n9832 ;
  assign n9834 = ~n9823 & n9833 ;
  assign n9835 = n9834 ^ x775 ;
  assign n9836 = n9835 ^ n9776 ;
  assign n9837 = n9836 ^ n9778 ;
  assign n9838 = n9837 ^ n9834 ;
  assign n9839 = ~n9815 & n9838 ;
  assign n9840 = n9839 ^ n9835 ;
  assign n9842 = n9841 ^ n9840 ;
  assign n9805 = x776 ^ x775 ;
  assign n9806 = n9805 ^ n9778 ;
  assign n9807 = n9806 ^ n9776 ;
  assign n9808 = n9738 ^ n9736 ;
  assign n9809 = n9808 ^ n9749 ;
  assign n9845 = n9807 & n9809 ;
  assign n9865 = n9845 ^ n9834 ;
  assign n9866 = n9842 & n9865 ;
  assign n9867 = n9866 ^ n9845 ;
  assign n9800 = n9772 ^ x776 ;
  assign n9801 = n9800 ^ n9769 ;
  assign n9771 = n9767 ^ x775 ;
  assign n9770 = n9769 ^ x776 ;
  assign n9775 = n9771 ^ n9770 ;
  assign n9773 = n9772 ^ n9771 ;
  assign n9782 = n9781 ^ n9773 ;
  assign n9783 = n9782 ^ n9775 ;
  assign n9784 = n9783 ^ n9772 ;
  assign n9785 = n9775 & n9784 ;
  assign n9791 = n9785 ^ n9782 ;
  assign n9787 = n9782 ^ n9771 ;
  assign n9788 = n9787 ^ n9785 ;
  assign n9789 = ~n9772 & n9788 ;
  assign n9792 = ~n9767 & n9789 ;
  assign n9793 = ~n9791 & n9792 ;
  assign n9786 = n9785 ^ n9784 ;
  assign n9790 = n9789 ^ n9786 ;
  assign n9794 = n9793 ^ n9790 ;
  assign n9799 = n9794 ^ n9767 ;
  assign n9802 = n9801 ^ n9799 ;
  assign n9760 = n9750 ^ n9739 ;
  assign n9761 = x782 & n9745 ;
  assign n9762 = n9761 ^ n9739 ;
  assign n9763 = n9760 & ~n9762 ;
  assign n9764 = n9763 ^ n9739 ;
  assign n9765 = ~n9759 & ~n9764 ;
  assign n9766 = n9765 ^ n9759 ;
  assign n9868 = n9802 ^ n9766 ;
  assign n9803 = ~n9766 & ~n9802 ;
  assign n9874 = n9868 ^ n9803 ;
  assign n9875 = ~n9867 & n9874 ;
  assign n9389 = ~x795 & ~x796 ;
  assign n9396 = ~x797 & ~x798 ;
  assign n9397 = ~n9389 & ~n9396 ;
  assign n9390 = x796 ^ x795 ;
  assign n9391 = n9390 ^ n9389 ;
  assign n9392 = x793 & x794 ;
  assign n9393 = x798 & n9392 ;
  assign n9394 = ~n9391 & n9393 ;
  assign n9395 = n9394 ^ n9392 ;
  assign n9398 = n9397 ^ n9395 ;
  assign n9384 = x798 ^ x797 ;
  assign n9401 = n9396 ^ n9384 ;
  assign n9404 = n9391 & n9401 ;
  assign n9405 = n9404 ^ n9395 ;
  assign n9406 = n9398 & ~n9405 ;
  assign n9388 = x794 ^ x793 ;
  assign n9407 = n9406 ^ n9395 ;
  assign n9408 = ~n9388 & n9407 ;
  assign n9409 = n9406 & n9408 ;
  assign n9410 = n9409 ^ n9407 ;
  assign n9482 = n9401 ^ n9391 ;
  assign n9483 = x794 & n9397 ;
  assign n9484 = n9483 ^ n9391 ;
  assign n9485 = n9482 & ~n9484 ;
  assign n9486 = n9485 ^ n9391 ;
  assign n9487 = ~n9410 & n9486 ;
  assign n9432 = ~x789 & ~x790 ;
  assign n9439 = ~x791 & ~x792 ;
  assign n9440 = ~n9432 & ~n9439 ;
  assign n9433 = x790 ^ x789 ;
  assign n9434 = n9433 ^ n9432 ;
  assign n9435 = x787 & x788 ;
  assign n9436 = x792 & n9435 ;
  assign n9437 = ~n9434 & n9436 ;
  assign n9438 = n9437 ^ n9435 ;
  assign n9441 = n9440 ^ n9438 ;
  assign n9427 = x792 ^ x791 ;
  assign n9444 = n9439 ^ n9427 ;
  assign n9447 = n9434 & n9444 ;
  assign n9448 = n9447 ^ n9438 ;
  assign n9449 = n9441 & ~n9448 ;
  assign n9431 = x788 ^ x787 ;
  assign n9450 = n9449 ^ n9438 ;
  assign n9451 = ~n9431 & n9450 ;
  assign n9452 = n9449 & n9451 ;
  assign n9453 = n9452 ^ n9450 ;
  assign n9474 = n9444 ^ n9434 ;
  assign n9475 = x788 & n9440 ;
  assign n9476 = n9475 ^ n9434 ;
  assign n9477 = n9474 & ~n9476 ;
  assign n9478 = n9477 ^ n9434 ;
  assign n9479 = ~n9453 & ~n9478 ;
  assign n9480 = n9479 ^ n9453 ;
  assign n9488 = n9487 ^ n9480 ;
  assign n9423 = x791 ^ x790 ;
  assign n9428 = ~n9423 & ~n9427 ;
  assign n9422 = x789 ^ x788 ;
  assign n9424 = n9423 ^ x789 ;
  assign n9425 = n9424 ^ x792 ;
  assign n9426 = ~n9422 & n9425 ;
  assign n9429 = n9428 ^ n9426 ;
  assign n9430 = ~x787 & n9429 ;
  assign n9454 = x790 ^ x788 ;
  assign n9455 = x792 ^ x787 ;
  assign n9458 = ~x790 & ~n9455 ;
  assign n9459 = n9458 ^ x787 ;
  assign n9460 = ~n9454 & n9459 ;
  assign n9461 = ~n9433 & n9460 ;
  assign n9462 = ~x791 & n9461 ;
  assign n9463 = ~n9453 & ~n9462 ;
  assign n9464 = ~n9430 & n9463 ;
  assign n9380 = x797 ^ x796 ;
  assign n9385 = ~n9380 & ~n9384 ;
  assign n9379 = x795 ^ x794 ;
  assign n9381 = n9380 ^ x795 ;
  assign n9382 = n9381 ^ x798 ;
  assign n9383 = ~n9379 & n9382 ;
  assign n9386 = n9385 ^ n9383 ;
  assign n9387 = ~x793 & n9386 ;
  assign n9411 = x796 ^ x794 ;
  assign n9412 = x798 ^ x793 ;
  assign n9415 = ~x796 & ~n9412 ;
  assign n9416 = n9415 ^ x793 ;
  assign n9417 = ~n9411 & n9416 ;
  assign n9418 = ~n9390 & n9417 ;
  assign n9419 = ~x797 & n9418 ;
  assign n9420 = ~n9410 & ~n9419 ;
  assign n9421 = ~n9387 & n9420 ;
  assign n9465 = n9464 ^ n9421 ;
  assign n9466 = n9433 ^ n9431 ;
  assign n9467 = n9466 ^ n9427 ;
  assign n9468 = n9390 ^ n9388 ;
  assign n9469 = n9468 ^ n9384 ;
  assign n9470 = n9467 & n9469 ;
  assign n9471 = n9470 ^ n9464 ;
  assign n9472 = n9465 & n9471 ;
  assign n9473 = n9472 ^ n9464 ;
  assign n9869 = n9488 ^ n9473 ;
  assign n9861 = n9842 ^ n9807 ;
  assign n9810 = n9809 ^ n9807 ;
  assign n9804 = n9469 ^ n9467 ;
  assign n9811 = n9810 ^ n9804 ;
  assign n9812 = ~n9467 & n9811 ;
  assign n9813 = n9812 ^ n9465 ;
  assign n9848 = n9842 & ~n9845 ;
  assign n9849 = n9848 ^ n9812 ;
  assign n9850 = ~n9813 & ~n9849 ;
  assign n9851 = n9850 ^ n9465 ;
  assign n9852 = ~n9469 & ~n9810 ;
  assign n9853 = n9852 ^ n9470 ;
  assign n9858 = ~n9465 & n9853 ;
  assign n9859 = n9858 ^ n9470 ;
  assign n9860 = n9851 & ~n9859 ;
  assign n9862 = ~n9810 & n9860 ;
  assign n9863 = n9861 & n9862 ;
  assign n9864 = n9863 ^ n9860 ;
  assign n9870 = n9869 ^ n9868 ;
  assign n9871 = n9870 ^ n9867 ;
  assign n9872 = n9871 ^ n9864 ;
  assign n9873 = n9803 & ~n9872 ;
  assign n9876 = ~n9864 & ~n9873 ;
  assign n9877 = n9869 & n9876 ;
  assign n9878 = n9875 & n9877 ;
  assign n9879 = n9878 ^ n9876 ;
  assign n9880 = n9879 ^ n9864 ;
  assign n9881 = n9874 ^ n9867 ;
  assign n9882 = n9881 ^ n9875 ;
  assign n9883 = ~n9864 & ~n9869 ;
  assign n9884 = ~n9882 & n9883 ;
  assign n9885 = n9884 ^ n9869 ;
  assign n9481 = n9480 ^ n9473 ;
  assign n9489 = n9481 & ~n9488 ;
  assign n9490 = n9489 ^ n9480 ;
  assign n9889 = ~n9490 & ~n9873 ;
  assign n9890 = ~n9885 & n9889 ;
  assign n9891 = ~n9875 & n9890 ;
  assign n9892 = n9891 ^ n9889 ;
  assign n9893 = n9892 ^ n9873 ;
  assign n9947 = n9880 & ~n9893 ;
  assign n9518 = x771 & x772 ;
  assign n9517 = x773 & x774 ;
  assign n9519 = n9518 ^ n9517 ;
  assign n9570 = n9517 ^ x769 ;
  assign n9573 = n9570 ^ n9519 ;
  assign n9568 = n9517 ^ x770 ;
  assign n9578 = n9573 ^ n9568 ;
  assign n9491 = x774 ^ x773 ;
  assign n9520 = n9517 ^ n9491 ;
  assign n9493 = x772 ^ x771 ;
  assign n9521 = n9518 ^ n9493 ;
  assign n9522 = n9520 & n9521 ;
  assign n9523 = n9522 ^ n9518 ;
  assign n9569 = n9523 ^ n9519 ;
  assign n9571 = n9570 ^ n9569 ;
  assign n9579 = n9578 ^ n9571 ;
  assign n9580 = n9579 ^ n9519 ;
  assign n9582 = n9578 & n9580 ;
  assign n9575 = n9571 ^ n9519 ;
  assign n9576 = n9575 ^ n9518 ;
  assign n9577 = ~n9522 & n9576 ;
  assign n9583 = n9582 ^ n9577 ;
  assign n9584 = n9583 ^ n9575 ;
  assign n9585 = n9582 ^ n9573 ;
  assign n9586 = n9585 ^ n9575 ;
  assign n9587 = n9584 & n9586 ;
  assign n9588 = ~n9519 & n9587 ;
  assign n9589 = n9588 ^ n9582 ;
  assign n9590 = n9589 ^ n9580 ;
  assign n9598 = n9590 ^ n9517 ;
  assign n9601 = n9598 ^ n9568 ;
  assign n9503 = x766 ^ x765 ;
  assign n9504 = n9503 ^ x767 ;
  assign n9565 = n9504 ^ x768 ;
  assign n9505 = x764 ^ x763 ;
  assign n9497 = ~x765 & ~x766 ;
  assign n9507 = n9503 ^ x768 ;
  assign n9530 = x768 ^ x767 ;
  assign n9538 = n9507 & n9530 ;
  assign n9539 = n9538 ^ x767 ;
  assign n9540 = ~n9497 & n9539 ;
  assign n9541 = n9540 ^ x764 ;
  assign n9542 = ~n9505 & n9541 ;
  assign n9566 = n9565 ^ n9542 ;
  assign n9550 = ~n9504 & ~n9565 ;
  assign n9551 = n9550 ^ n9542 ;
  assign n9560 = n9542 ^ x768 ;
  assign n9553 = n9566 ^ x767 ;
  assign n9552 = n9566 ^ x765 ;
  assign n9554 = n9553 ^ n9552 ;
  assign n9548 = n9566 ^ x768 ;
  assign n9555 = n9552 ^ n9548 ;
  assign n9556 = n9566 ^ n9555 ;
  assign n9557 = n9556 ^ n9542 ;
  assign n9558 = ~n9554 & ~n9557 ;
  assign n9561 = n9560 ^ n9558 ;
  assign n9562 = ~n9551 & ~n9561 ;
  assign n9567 = n9566 ^ n9562 ;
  assign n9602 = n9601 ^ n9567 ;
  assign n9524 = ~n9519 & ~n9523 ;
  assign n9492 = n9491 ^ x770 ;
  assign n9494 = n9493 ^ n9492 ;
  assign n9506 = n9505 ^ n9504 ;
  assign n9508 = n9507 ^ n9497 ;
  assign n9509 = n9506 & n9508 ;
  assign n9495 = x767 ^ x764 ;
  assign n9498 = n9497 ^ x767 ;
  assign n9501 = ~n9495 & n9498 ;
  assign n9499 = n9498 ^ x764 ;
  assign n9500 = x763 & n9499 ;
  assign n9502 = n9501 ^ n9500 ;
  assign n9510 = n9509 ^ n9502 ;
  assign n9511 = n9510 ^ x769 ;
  assign n9512 = n9511 ^ n9491 ;
  assign n9513 = n9512 ^ n9493 ;
  assign n9514 = n9513 ^ n9510 ;
  assign n9515 = ~n9494 & n9514 ;
  assign n9516 = n9515 ^ n9511 ;
  assign n9525 = n9524 ^ n9516 ;
  assign n9526 = x770 ^ x769 ;
  assign n9527 = n9526 ^ n9493 ;
  assign n9528 = n9527 ^ n9491 ;
  assign n9529 = n9505 ^ n9503 ;
  assign n9531 = n9530 ^ n9529 ;
  assign n9532 = n9528 & n9531 ;
  assign n9533 = n9532 ^ n9510 ;
  assign n9534 = ~n9525 & ~n9533 ;
  assign n9535 = n9534 ^ n9532 ;
  assign n9603 = n9602 ^ n9535 ;
  assign n9631 = x756 ^ x755 ;
  assign n9630 = ~x755 & ~x756 ;
  assign n9632 = n9631 ^ n9630 ;
  assign n9634 = ~x753 & ~x754 ;
  assign n9633 = x754 ^ x753 ;
  assign n9635 = n9634 ^ n9633 ;
  assign n9636 = n9632 & n9635 ;
  assign n9637 = ~n9630 & ~n9634 ;
  assign n9638 = n9636 & ~n9637 ;
  assign n9639 = x751 & x752 ;
  assign n9640 = ~n9638 & n9639 ;
  assign n9641 = x756 & ~n9635 ;
  assign n9642 = n9640 & n9641 ;
  assign n9643 = n9642 ^ n9640 ;
  assign n9644 = n9637 ^ n9636 ;
  assign n9645 = n9644 ^ n9638 ;
  assign n9646 = ~x752 & n9645 ;
  assign n9648 = x751 & ~n9646 ;
  assign n9647 = n9646 ^ x751 ;
  assign n9649 = n9648 ^ n9647 ;
  assign n9650 = n9649 ^ n9645 ;
  assign n9651 = n9635 ^ n9632 ;
  assign n9652 = n9651 ^ n9636 ;
  assign n9653 = ~n9650 & n9652 ;
  assign n9654 = ~n9643 & n9653 ;
  assign n9605 = x761 & x762 ;
  assign n9604 = x759 & x760 ;
  assign n9606 = n9605 ^ n9604 ;
  assign n9607 = x762 ^ x761 ;
  assign n9608 = n9607 ^ n9605 ;
  assign n9609 = x760 ^ x759 ;
  assign n9610 = n9609 ^ n9604 ;
  assign n9611 = n9608 & n9610 ;
  assign n9616 = x758 & n9611 ;
  assign n9617 = n9616 ^ n9604 ;
  assign n9618 = n9606 & ~n9617 ;
  assign n9619 = n9618 ^ n9605 ;
  assign n9624 = ~n9606 & ~n9611 ;
  assign n9657 = n9611 ^ n9606 ;
  assign n9660 = n9657 ^ x758 ;
  assign n9625 = n9624 & ~n9660 ;
  assign n9622 = n9660 ^ n9619 ;
  assign n9626 = n9625 ^ n9622 ;
  assign n9627 = x757 & ~n9626 ;
  assign n9628 = ~n9619 & n9627 ;
  assign n9629 = n9628 ^ n9619 ;
  assign n9708 = n9654 ^ n9629 ;
  assign n9712 = n9708 ^ n9603 ;
  assign n9673 = x756 ^ x752 ;
  assign n9680 = n9631 & n9673 ;
  assign n9681 = n9680 ^ x756 ;
  assign n9682 = n9634 & ~n9681 ;
  assign n9683 = n9682 ^ n9653 ;
  assign n9684 = ~n9648 & ~n9683 ;
  assign n9668 = x752 ^ x751 ;
  assign n9669 = n9668 ^ n9634 ;
  assign n9670 = ~x755 & ~n9669 ;
  assign n9671 = n9668 ^ n9633 ;
  assign n9672 = n9671 ^ x756 ;
  assign n9674 = n9672 & ~n9673 ;
  assign n9675 = n9670 & n9674 ;
  assign n9676 = n9675 ^ n9643 ;
  assign n9661 = ~x757 & ~n9660 ;
  assign n9656 = n9609 ^ n9607 ;
  assign n9658 = n9657 ^ n9656 ;
  assign n9659 = n9658 ^ n9626 ;
  assign n9662 = n9661 ^ n9659 ;
  assign n9663 = n9661 ^ n9626 ;
  assign n9664 = x758 ^ x757 ;
  assign n9665 = n9663 & n9664 ;
  assign n9666 = n9662 & n9665 ;
  assign n9667 = n9666 ^ n9663 ;
  assign n9677 = n9676 ^ n9667 ;
  assign n9686 = n9684 ^ n9677 ;
  assign n9687 = n9671 ^ n9631 ;
  assign n9688 = n9664 ^ n9609 ;
  assign n9689 = n9688 ^ n9607 ;
  assign n9690 = n9687 & n9689 ;
  assign n9691 = n9690 ^ n9667 ;
  assign n9692 = n9686 & n9691 ;
  assign n9693 = n9692 ^ n9690 ;
  assign n9713 = n9712 ^ n9693 ;
  assign n9655 = ~n9629 & n9654 ;
  assign n9938 = n9708 ^ n9655 ;
  assign n9695 = n9531 ^ n9528 ;
  assign n9696 = n9689 ^ n9687 ;
  assign n9697 = n9695 & n9696 ;
  assign n9698 = n9697 ^ n9532 ;
  assign n9699 = n9698 ^ n9690 ;
  assign n9700 = n9699 ^ n9686 ;
  assign n9701 = n9700 ^ n9525 ;
  assign n9703 = n9697 ^ n9690 ;
  assign n9706 = n9701 & n9703 ;
  assign n9702 = n9701 ^ n9690 ;
  assign n9704 = n9703 ^ n9702 ;
  assign n9705 = ~n9686 & n9704 ;
  assign n9707 = n9706 ^ n9705 ;
  assign n9937 = n9707 ^ n9655 ;
  assign n9939 = n9938 ^ n9937 ;
  assign n9719 = ~n9713 & ~n9939 ;
  assign n9694 = n9693 ^ n9655 ;
  assign n9720 = n9719 ^ n9694 ;
  assign n9723 = n9720 ^ n9693 ;
  assign n9727 = n9723 & ~n9938 ;
  assign n9728 = n9727 ^ n9720 ;
  assign n9729 = ~n9603 & n9728 ;
  assign n9730 = n9729 ^ n9720 ;
  assign n9731 = n9601 ^ n9535 ;
  assign n9732 = n9602 & n9731 ;
  assign n9733 = n9732 ^ n9601 ;
  assign n9945 = ~n9730 & n9733 ;
  assign n9940 = n9938 ^ n9694 ;
  assign n9941 = n9939 & n9940 ;
  assign n9942 = n9941 ^ n9938 ;
  assign n9943 = n9603 & n9942 ;
  assign n9944 = ~n9655 & n9943 ;
  assign n9946 = n9945 ^ n9944 ;
  assign n9948 = n9947 ^ n9946 ;
  assign n9894 = ~n9885 & n9893 ;
  assign n9886 = n9885 ^ n9880 ;
  assign n9887 = ~n9873 & ~n9886 ;
  assign n9734 = n9733 ^ n9730 ;
  assign n9735 = n9734 ^ n9490 ;
  assign n9888 = n9887 ^ n9735 ;
  assign n9895 = n9894 ^ n9888 ;
  assign n9896 = n9707 ^ n9693 ;
  assign n9897 = n9896 ^ n9712 ;
  assign n9898 = n9897 ^ n9872 ;
  assign n9908 = n9872 ^ n9701 ;
  assign n9902 = n9853 ^ n9845 ;
  assign n9903 = n9902 ^ n9812 ;
  assign n9900 = n9696 ^ n9695 ;
  assign n9901 = n9811 & n9900 ;
  assign n9904 = n9903 ^ n9901 ;
  assign n9856 = n9470 ^ n9465 ;
  assign n9899 = n9856 ^ n9842 ;
  assign n9905 = n9904 ^ n9899 ;
  assign n9906 = n9901 ^ n9701 ;
  assign n9907 = ~n9905 & ~n9906 ;
  assign n9909 = n9908 ^ n9907 ;
  assign n9910 = n9898 & n9909 ;
  assign n9911 = n9910 ^ n9872 ;
  assign n9912 = n9911 ^ n9734 ;
  assign n9913 = ~n9895 & n9912 ;
  assign n9914 = n9913 ^ n9734 ;
  assign n9121 = x842 ^ x841 ;
  assign n9130 = ~x843 & ~x844 ;
  assign n9123 = x846 ^ x845 ;
  assign n9127 = x845 & ~n9123 ;
  assign n9155 = n9127 ^ n9123 ;
  assign n9156 = ~n9130 & n9155 ;
  assign n9120 = x844 ^ x843 ;
  assign n9151 = n9130 ^ n9120 ;
  assign n9126 = x841 & ~n9121 ;
  assign n9152 = x846 & n9126 ;
  assign n9153 = ~n9151 & n9152 ;
  assign n9154 = n9153 ^ n9126 ;
  assign n9157 = n9156 ^ n9154 ;
  assign n9162 = ~n9127 & n9151 ;
  assign n9163 = n9162 ^ n9154 ;
  assign n9164 = n9157 & ~n9163 ;
  assign n9165 = ~n9121 & n9164 ;
  assign n9142 = ~x837 & ~x838 ;
  assign n9132 = x838 ^ x837 ;
  assign n9173 = n9142 ^ n9132 ;
  assign n9133 = x836 ^ x835 ;
  assign n9138 = x835 & ~n9133 ;
  assign n9185 = x840 & n9138 ;
  assign n9186 = ~n9173 & n9185 ;
  assign n9187 = n9186 ^ n9138 ;
  assign n9135 = x840 ^ x839 ;
  assign n9139 = x839 & ~n9135 ;
  assign n9175 = n9139 ^ n9135 ;
  assign n9176 = ~n9142 & n9175 ;
  assign n9188 = n9187 ^ n9176 ;
  assign n9192 = ~n9139 & n9173 ;
  assign n9193 = n9192 ^ n9176 ;
  assign n9194 = n9188 & n9193 ;
  assign n9174 = n9173 ^ n9139 ;
  assign n9181 = x836 & n9176 ;
  assign n9182 = n9181 ^ n9173 ;
  assign n9183 = ~n9174 & n9182 ;
  assign n9184 = n9183 ^ n9139 ;
  assign n9195 = n9194 ^ n9187 ;
  assign n9196 = ~n9184 & n9195 ;
  assign n9197 = ~n9133 & n9196 ;
  assign n9198 = n9194 & n9197 ;
  assign n9199 = n9198 ^ n9196 ;
  assign n9200 = n9199 ^ n9184 ;
  assign n9166 = n9164 ^ n9154 ;
  assign n9208 = n9200 ^ ~n9166 ;
  assign n9171 = x842 & n9156 ;
  assign n9172 = n9171 ^ n9151 ;
  assign n9201 = n9200 ^ n9127 ;
  assign n9202 = n9201 ^ n9151 ;
  assign n9203 = n9202 ^ n9200 ;
  assign n9204 = n9172 & ~n9203 ;
  assign n9205 = n9204 ^ n9201 ;
  assign n9209 = n9208 ^ n9205 ;
  assign n9210 = n9165 & ~n9209 ;
  assign n9211 = n9210 ^ n9208 ;
  assign n9140 = n9139 ^ n9138 ;
  assign n9134 = n9133 ^ n9132 ;
  assign n9136 = n9135 ^ n9133 ;
  assign n9137 = n9134 & ~n9136 ;
  assign n9141 = n9140 ^ n9137 ;
  assign n9143 = n9142 ^ n9141 ;
  assign n9128 = n9127 ^ n9126 ;
  assign n9122 = n9121 ^ n9120 ;
  assign n9124 = n9123 ^ n9121 ;
  assign n9125 = n9122 & ~n9124 ;
  assign n9129 = n9128 ^ n9125 ;
  assign n9131 = n9130 ^ n9129 ;
  assign n9144 = n9143 ^ n9131 ;
  assign n9145 = n9135 ^ n9134 ;
  assign n9146 = n9123 ^ n9122 ;
  assign n9147 = n9145 & n9146 ;
  assign n9148 = n9147 ^ n9131 ;
  assign n9149 = n9144 & ~n9148 ;
  assign n9150 = n9149 ^ n9131 ;
  assign n9345 = n9200 ^ n9150 ;
  assign n9346 = ~n9211 & ~n9345 ;
  assign n9347 = n9346 ^ n9200 ;
  assign n9213 = n9146 ^ n9145 ;
  assign n9222 = x834 ^ x833 ;
  assign n9220 = x830 ^ x829 ;
  assign n9219 = x832 ^ x831 ;
  assign n9221 = n9220 ^ n9219 ;
  assign n9223 = n9222 ^ n9221 ;
  assign n9217 = x828 ^ x827 ;
  assign n9215 = x826 ^ x825 ;
  assign n9214 = x824 ^ x823 ;
  assign n9216 = n9215 ^ n9214 ;
  assign n9218 = n9217 ^ n9216 ;
  assign n9224 = n9223 ^ n9218 ;
  assign n9225 = n9213 & n9224 ;
  assign n9226 = n9225 ^ n9147 ;
  assign n9227 = n9226 ^ n9144 ;
  assign n9262 = x825 & x826 ;
  assign n9263 = n9262 ^ x824 ;
  assign n9266 = n9215 ^ x823 ;
  assign n9267 = ~x828 & n9266 ;
  assign n9268 = n9267 ^ x823 ;
  assign n9269 = ~n9262 & n9268 ;
  assign n9270 = n9269 ^ x823 ;
  assign n9271 = ~n9263 & n9270 ;
  assign n9272 = ~x827 & n9271 ;
  assign n9273 = x827 & x828 ;
  assign n9274 = n9273 ^ n9217 ;
  assign n9275 = x824 & n9274 ;
  assign n9279 = n9262 & n9273 ;
  assign n9276 = n9273 ^ x826 ;
  assign n9285 = n9279 ^ n9276 ;
  assign n9277 = n9215 & ~n9276 ;
  assign n9286 = n9285 ^ n9277 ;
  assign n9289 = ~n9275 & ~n9286 ;
  assign n9278 = n9277 ^ x825 ;
  assign n9280 = n9278 & ~n9279 ;
  assign n9281 = ~n9275 & n9280 ;
  assign n9282 = n9281 ^ n9278 ;
  assign n9290 = n9289 ^ n9282 ;
  assign n9291 = ~x823 & n9290 ;
  assign n9292 = ~n9272 & ~n9291 ;
  assign n9303 = n9286 ^ n9278 ;
  assign n9304 = n9303 ^ n9262 ;
  assign n9305 = n9304 ^ n9278 ;
  assign n9308 = x824 & n9305 ;
  assign n9309 = n9308 ^ n9278 ;
  assign n9310 = ~n9214 & n9309 ;
  assign n9295 = x824 & n9286 ;
  assign n9296 = n9295 ^ n9278 ;
  assign n9297 = ~n9214 & n9296 ;
  assign n9298 = n9297 ^ n9278 ;
  assign n9299 = ~x828 & n9298 ;
  assign n9300 = n9299 ^ x828 ;
  assign n9301 = n9300 ^ n9278 ;
  assign n9311 = n9310 ^ n9301 ;
  assign n9312 = n9311 ^ n9300 ;
  assign n9313 = n9311 ^ x828 ;
  assign n9314 = x827 & ~n9313 ;
  assign n9315 = n9312 & n9314 ;
  assign n9316 = n9315 ^ n9313 ;
  assign n9317 = n9292 & ~n9316 ;
  assign n9261 = n9218 & n9223 ;
  assign n9318 = n9317 ^ n9261 ;
  assign n9228 = ~x833 & ~x834 ;
  assign n9229 = ~x831 & ~x832 ;
  assign n9232 = n9228 ^ n9222 ;
  assign n9235 = n9229 & n9232 ;
  assign n9242 = n9235 ^ x829 ;
  assign n9243 = n9235 ^ n9228 ;
  assign n9244 = n9243 ^ n9221 ;
  assign n9245 = n9242 & n9244 ;
  assign n9256 = ~n9235 & n9245 ;
  assign n9233 = n9232 ^ x832 ;
  assign n9236 = n9235 ^ n9233 ;
  assign n9234 = n9219 & n9233 ;
  assign n9237 = n9236 ^ n9234 ;
  assign n9230 = n9229 ^ n9219 ;
  assign n9231 = n9228 & n9230 ;
  assign n9238 = n9237 ^ n9231 ;
  assign n9246 = x829 & x830 ;
  assign n9247 = ~n9235 & n9246 ;
  assign n9248 = ~n9238 & n9247 ;
  assign n9239 = n9220 & ~n9228 ;
  assign n9249 = n9234 ^ x831 ;
  assign n9250 = n9239 & n9249 ;
  assign n9251 = ~n9248 & ~n9250 ;
  assign n9257 = n9256 ^ n9251 ;
  assign n9258 = ~n9228 & ~n9257 ;
  assign n9259 = n9258 ^ n9245 ;
  assign n9240 = ~x830 & ~n9239 ;
  assign n9241 = n9238 & n9240 ;
  assign n9260 = n9259 ^ n9241 ;
  assign n9319 = n9318 ^ n9260 ;
  assign n9320 = n9319 ^ n9225 ;
  assign n9321 = ~n9227 & ~n9320 ;
  assign n9322 = n9321 ^ n9319 ;
  assign n9212 = n9211 ^ n9150 ;
  assign n9324 = n9322 ^ n9212 ;
  assign n9323 = n9212 & ~n9322 ;
  assign n9325 = n9324 ^ n9323 ;
  assign n9326 = n9261 ^ n9260 ;
  assign n9327 = n9318 & n9326 ;
  assign n9328 = n9327 ^ n9317 ;
  assign n9329 = ~n9325 & n9328 ;
  assign n9330 = ~n9237 & n9251 ;
  assign n9331 = ~n9282 & ~n9316 ;
  assign n9332 = ~n9330 & ~n9331 ;
  assign n9333 = n9332 ^ n9323 ;
  assign n9334 = n9331 ^ n9330 ;
  assign n9335 = n9334 ^ n9328 ;
  assign n9336 = n9335 ^ n9324 ;
  assign n9337 = n9334 ^ n9332 ;
  assign n9338 = n9336 & n9337 ;
  assign n9341 = n9333 & n9338 ;
  assign n9342 = n9341 ^ n9332 ;
  assign n9343 = ~n9329 & ~n9342 ;
  assign n9344 = n9343 ^ n9338 ;
  assign n9354 = n9347 ^ n9344 ;
  assign n9349 = ~n9329 & ~n9332 ;
  assign n9353 = n9323 & n9349 ;
  assign n9356 = n9354 ^ n9353 ;
  assign n8834 = x810 ^ x809 ;
  assign n9010 = x809 ^ x808 ;
  assign n9014 = ~n8834 & ~n9010 ;
  assign n9009 = x807 ^ x806 ;
  assign n9011 = n9010 ^ x807 ;
  assign n9012 = n9011 ^ x810 ;
  assign n9013 = ~n9009 & n9012 ;
  assign n9015 = n9014 ^ n9013 ;
  assign n9016 = ~x805 & n9015 ;
  assign n8822 = ~x807 & ~x808 ;
  assign n8829 = ~x809 & ~x810 ;
  assign n8830 = ~n8822 & ~n8829 ;
  assign n8823 = x808 ^ x807 ;
  assign n8824 = n8823 ^ n8822 ;
  assign n8825 = x805 & x806 ;
  assign n8826 = x810 & n8825 ;
  assign n8827 = ~n8824 & n8826 ;
  assign n8828 = n8827 ^ n8825 ;
  assign n8831 = n8830 ^ n8828 ;
  assign n8835 = n8834 ^ n8829 ;
  assign n8838 = n8824 & n8835 ;
  assign n8839 = n8838 ^ n8828 ;
  assign n8840 = n8831 & ~n8839 ;
  assign n8821 = x806 ^ x805 ;
  assign n8841 = n8840 ^ n8828 ;
  assign n8842 = ~n8821 & n8841 ;
  assign n8843 = n8840 & n8842 ;
  assign n8844 = n8843 ^ n8841 ;
  assign n9017 = x808 ^ x806 ;
  assign n9018 = x810 ^ x805 ;
  assign n9021 = ~x808 & ~n9018 ;
  assign n9022 = n9021 ^ x805 ;
  assign n9023 = ~n9017 & n9022 ;
  assign n9024 = ~n8823 & n9023 ;
  assign n9025 = ~x809 & n9024 ;
  assign n9026 = ~n8844 & ~n9025 ;
  assign n9027 = ~n9016 & n9026 ;
  assign n8798 = x804 ^ x803 ;
  assign n8796 = x803 & x804 ;
  assign n8799 = n8798 ^ n8796 ;
  assign n8800 = x802 ^ x801 ;
  assign n8795 = x801 & x802 ;
  assign n8801 = n8800 ^ n8795 ;
  assign n8802 = n8799 & n8801 ;
  assign n8797 = n8796 ^ n8795 ;
  assign n8999 = n8802 ^ n8797 ;
  assign n9000 = n8999 ^ n8798 ;
  assign n9001 = n9000 ^ n8800 ;
  assign n9002 = x800 ^ x799 ;
  assign n9003 = n8999 ^ x800 ;
  assign n9004 = ~x799 & ~n9003 ;
  assign n8815 = ~n8797 & ~n8802 ;
  assign n8816 = n8815 & ~n9003 ;
  assign n8807 = x800 & n8802 ;
  assign n8808 = n8807 ^ n8795 ;
  assign n8809 = n8797 & ~n8808 ;
  assign n8810 = n8809 ^ n8796 ;
  assign n8813 = n9003 ^ n8810 ;
  assign n8817 = n8816 ^ n8813 ;
  assign n9005 = n9004 ^ n8817 ;
  assign n9006 = n9002 & n9005 ;
  assign n9007 = ~n9001 & n9006 ;
  assign n9008 = n9007 ^ n9005 ;
  assign n9028 = n9027 ^ n9008 ;
  assign n9030 = n8823 ^ n8821 ;
  assign n9031 = n9030 ^ n8834 ;
  assign n9032 = n9002 ^ n8800 ;
  assign n9033 = n9032 ^ n8798 ;
  assign n9036 = n9031 & n9033 ;
  assign n8899 = x822 ^ x821 ;
  assign n8886 = x818 ^ x817 ;
  assign n8988 = n8899 ^ n8886 ;
  assign n8888 = x820 ^ x819 ;
  assign n8989 = n8988 ^ n8888 ;
  assign n8865 = x816 ^ x815 ;
  assign n8852 = x812 ^ x811 ;
  assign n8990 = n8865 ^ n8852 ;
  assign n8855 = x814 ^ x813 ;
  assign n8991 = n8990 ^ n8855 ;
  assign n8992 = n8989 & n8991 ;
  assign n9038 = n9036 ^ n8992 ;
  assign n9029 = n8991 ^ n8989 ;
  assign n9034 = n9033 ^ n9031 ;
  assign n9035 = n9029 & n9034 ;
  assign n9039 = n9038 ^ n9035 ;
  assign n9040 = n9039 ^ n9028 ;
  assign n8854 = ~x813 & ~x814 ;
  assign n8860 = ~x815 & ~x816 ;
  assign n8861 = ~n8854 & ~n8860 ;
  assign n8853 = x811 & x812 ;
  assign n8856 = n8855 ^ n8854 ;
  assign n8857 = x816 & ~n8856 ;
  assign n8858 = n8853 & n8857 ;
  assign n8859 = n8858 ^ n8853 ;
  assign n8862 = n8861 ^ n8859 ;
  assign n8866 = n8865 ^ n8860 ;
  assign n8869 = n8856 & n8866 ;
  assign n8870 = n8869 ^ n8859 ;
  assign n8871 = n8862 & ~n8870 ;
  assign n8872 = n8871 ^ n8859 ;
  assign n8873 = ~n8852 & n8872 ;
  assign n8874 = n8871 & n8873 ;
  assign n8875 = n8874 ^ n8872 ;
  assign n8921 = ~x815 & ~n8875 ;
  assign n8923 = x816 ^ x813 ;
  assign n8922 = x816 ^ x812 ;
  assign n8924 = n8923 ^ n8922 ;
  assign n8925 = n8924 ^ x816 ;
  assign n8927 = x812 & n8925 ;
  assign n8928 = n8927 ^ x816 ;
  assign n8931 = x816 ^ x814 ;
  assign n8932 = n8931 ^ n8922 ;
  assign n8933 = n8932 ^ n8852 ;
  assign n8935 = n8922 ^ n8855 ;
  assign n8936 = n8935 ^ x816 ;
  assign n8937 = ~n8933 & n8936 ;
  assign n8940 = n8937 ^ x813 ;
  assign n8941 = ~n8928 & ~n8940 ;
  assign n8942 = n8921 & n8941 ;
  assign n8943 = n8942 ^ n8875 ;
  assign n8978 = x815 ^ x812 ;
  assign n8981 = n8865 & n8978 ;
  assign n8982 = n8981 ^ x815 ;
  assign n8983 = n8854 & ~n8982 ;
  assign n8876 = n8866 ^ n8856 ;
  assign n8881 = x812 & n8861 ;
  assign n8882 = n8881 ^ n8856 ;
  assign n8883 = n8876 & n8882 ;
  assign n8884 = n8883 ^ n8866 ;
  assign n8984 = n8983 ^ n8884 ;
  assign n8985 = ~x811 & ~n8984 ;
  assign n8986 = ~n8943 & n8985 ;
  assign n8887 = ~x819 & ~x820 ;
  assign n8894 = ~x821 & ~x822 ;
  assign n8895 = ~n8887 & ~n8894 ;
  assign n8889 = n8888 ^ n8887 ;
  assign n8890 = x817 & x818 ;
  assign n8891 = x822 & n8890 ;
  assign n8892 = ~n8889 & n8891 ;
  assign n8893 = n8892 ^ n8890 ;
  assign n8896 = n8895 ^ n8893 ;
  assign n8900 = n8899 ^ n8894 ;
  assign n8903 = n8889 & n8900 ;
  assign n8904 = n8903 ^ n8893 ;
  assign n8905 = n8896 & ~n8904 ;
  assign n8906 = n8905 ^ n8893 ;
  assign n8907 = ~n8886 & n8906 ;
  assign n8908 = n8905 & n8907 ;
  assign n8909 = n8908 ^ n8906 ;
  assign n8944 = ~x821 & ~n8909 ;
  assign n8946 = x822 ^ x819 ;
  assign n8945 = x822 ^ x818 ;
  assign n8947 = n8946 ^ n8945 ;
  assign n8948 = n8947 ^ x822 ;
  assign n8950 = x818 & n8948 ;
  assign n8951 = n8950 ^ x822 ;
  assign n8954 = x822 ^ x820 ;
  assign n8955 = n8954 ^ n8945 ;
  assign n8956 = n8955 ^ n8886 ;
  assign n8958 = n8945 ^ n8888 ;
  assign n8959 = n8958 ^ x822 ;
  assign n8960 = ~n8956 & n8959 ;
  assign n8963 = n8960 ^ x819 ;
  assign n8964 = ~n8951 & ~n8963 ;
  assign n8965 = n8944 & n8964 ;
  assign n8966 = n8965 ^ n8909 ;
  assign n8967 = x821 ^ x818 ;
  assign n8970 = n8899 & n8967 ;
  assign n8971 = n8970 ^ x821 ;
  assign n8972 = n8887 & ~n8971 ;
  assign n8910 = n8900 ^ n8889 ;
  assign n8915 = x818 & n8895 ;
  assign n8916 = n8915 ^ n8900 ;
  assign n8917 = n8910 & n8916 ;
  assign n8918 = n8917 ^ n8889 ;
  assign n8973 = n8972 ^ n8918 ;
  assign n8974 = ~x817 & ~n8973 ;
  assign n8975 = ~n8966 & n8974 ;
  assign n8976 = n8975 ^ n8966 ;
  assign n8977 = n8976 ^ n8943 ;
  assign n8987 = n8986 ^ n8977 ;
  assign n9041 = n9040 ^ n8987 ;
  assign n9042 = n8992 ^ n8987 ;
  assign n9043 = n9041 & ~n9042 ;
  assign n9037 = n9036 ^ n9035 ;
  assign n9044 = n9043 ^ n9037 ;
  assign n9045 = ~n9028 & ~n9044 ;
  assign n9046 = n9037 ^ n9008 ;
  assign n9047 = n9045 & ~n9046 ;
  assign n9048 = n9047 ^ n9043 ;
  assign n8845 = n8835 ^ n8824 ;
  assign n8846 = x806 & n8830 ;
  assign n8847 = n8846 ^ n8824 ;
  assign n8848 = n8845 & ~n8847 ;
  assign n8849 = n8848 ^ n8824 ;
  assign n8850 = ~n8844 & ~n8849 ;
  assign n8851 = n8850 ^ n8844 ;
  assign n9057 = n9048 ^ n8851 ;
  assign n9051 = n9008 & n9027 ;
  assign n9052 = n9037 & n9051 ;
  assign n9053 = ~n9041 & n9052 ;
  assign n8993 = n8992 ^ n8976 ;
  assign n8994 = ~n8987 & ~n8993 ;
  assign n8995 = n8994 ^ n8992 ;
  assign n8919 = ~n8909 & n8918 ;
  assign n8885 = ~n8875 & n8884 ;
  assign n8920 = n8919 ^ n8885 ;
  assign n9049 = n8995 ^ n8920 ;
  assign n9055 = n9053 ^ n9049 ;
  assign n9056 = n9055 ^ n9048 ;
  assign n9058 = n9057 ^ n9056 ;
  assign n9054 = n9053 ^ n9048 ;
  assign n9059 = n9058 ^ n9054 ;
  assign n8818 = x799 & ~n8817 ;
  assign n8819 = ~n8810 & n8818 ;
  assign n8820 = n8819 ^ n8810 ;
  assign n9050 = n9049 ^ n8820 ;
  assign n9060 = n9059 ^ n9050 ;
  assign n9101 = n9060 ^ n9054 ;
  assign n9102 = n9101 ^ n9049 ;
  assign n9075 = n9053 ^ n9050 ;
  assign n9076 = n9058 & n9075 ;
  assign n9077 = n9076 ^ n9058 ;
  assign n9078 = n9101 ^ n9077 ;
  assign n9369 = n8851 ^ n8820 ;
  assign n9082 = n9077 ^ n9060 ;
  assign n9370 = n9369 ^ n9049 ;
  assign n9083 = n9082 & ~n9370 ;
  assign n9084 = n9083 ^ n9076 ;
  assign n9085 = n9369 ^ n9084 ;
  assign n9086 = n9078 & n9085 ;
  assign n9087 = ~n8851 & n9086 ;
  assign n9088 = n9087 ^ n9083 ;
  assign n9089 = n9101 ^ n9088 ;
  assign n9090 = n9089 ^ n8820 ;
  assign n9091 = n9102 ^ n9090 ;
  assign n9099 = n9091 ^ n9053 ;
  assign n9100 = n9099 ^ n9055 ;
  assign n9103 = n9102 ^ n9100 ;
  assign n9104 = n9103 ^ n9048 ;
  assign n9105 = n9104 ^ n9053 ;
  assign n8996 = n8995 ^ n8919 ;
  assign n8997 = ~n8920 & ~n8996 ;
  assign n8998 = n8997 ^ n8995 ;
  assign n9106 = n9105 ^ n8998 ;
  assign n9357 = n9356 ^ n9106 ;
  assign n9361 = n9319 ^ n9227 ;
  assign n9358 = n9034 ^ n9029 ;
  assign n9359 = n9224 ^ n9213 ;
  assign n9360 = n9358 & n9359 ;
  assign n9362 = n9361 ^ n9360 ;
  assign n9365 = n9361 ^ n9041 ;
  assign n9366 = ~n9362 & ~n9365 ;
  assign n9363 = n9361 ^ n9336 ;
  assign n9367 = n9366 ^ n9363 ;
  assign n9371 = n9370 ^ n9054 ;
  assign n9372 = n9371 ^ n9106 ;
  assign n9368 = n9336 ^ n9106 ;
  assign n9373 = n9372 ^ n9368 ;
  assign n9374 = n9367 & n9373 ;
  assign n9375 = n9374 ^ n9368 ;
  assign n9376 = ~n9357 & ~n9375 ;
  assign n9377 = n9376 ^ n9106 ;
  assign n9350 = ~n9338 & n9349 ;
  assign n9348 = ~n9344 & ~n9347 ;
  assign n9351 = n9350 ^ n9348 ;
  assign n9107 = ~n9050 & ~n9054 ;
  assign n9108 = n9107 ^ n9049 ;
  assign n9109 = n9108 ^ n9053 ;
  assign n9110 = ~n8998 & ~n9109 ;
  assign n9111 = ~n9107 & n9110 ;
  assign n9112 = ~n9053 & n9111 ;
  assign n9113 = n9112 ^ n9110 ;
  assign n9114 = n9113 ^ n8998 ;
  assign n9115 = n9106 & n9114 ;
  assign n9116 = n8851 & n9115 ;
  assign n9117 = n8820 & n9116 ;
  assign n9118 = n9117 ^ n9115 ;
  assign n9119 = n9118 ^ n9114 ;
  assign n9352 = n9351 ^ n9119 ;
  assign n9378 = n9377 ^ n9352 ;
  assign n9917 = n9375 ^ n9356 ;
  assign n9916 = n9911 ^ n9895 ;
  assign n9918 = n9917 ^ n9916 ;
  assign n9921 = n9362 ^ n9041 ;
  assign n9920 = n9905 ^ n9701 ;
  assign n9922 = n9921 ^ n9920 ;
  assign n9923 = n9359 ^ n9358 ;
  assign n9924 = n9900 ^ n9811 ;
  assign n9925 = n9923 & n9924 ;
  assign n9926 = n9925 ^ n9921 ;
  assign n9927 = n9922 & ~n9926 ;
  assign n9928 = n9927 ^ n9921 ;
  assign n9933 = n9928 ^ n9917 ;
  assign n9919 = n9909 ^ n9897 ;
  assign n9929 = n9928 ^ n9919 ;
  assign n9930 = n9371 ^ n9367 ;
  assign n9931 = n9930 ^ n9928 ;
  assign n9932 = n9929 & n9931 ;
  assign n9934 = n9933 ^ n9932 ;
  assign n9935 = n9918 & ~n9934 ;
  assign n9936 = n9935 ^ n9917 ;
  assign n11092 = ~n9378 & n9936 ;
  assign n11093 = ~n9914 & n11092 ;
  assign n11094 = n11093 ^ n9914 ;
  assign n11086 = n9946 ^ n9914 ;
  assign n11095 = n11094 ^ n11086 ;
  assign n11096 = n9948 & ~n11095 ;
  assign n11097 = n11096 ^ n9947 ;
  assign n11078 = n9914 & ~n9936 ;
  assign n11098 = n9377 ^ n9351 ;
  assign n11099 = n9352 & ~n11098 ;
  assign n11100 = n11099 ^ n9377 ;
  assign n9949 = n9948 ^ n9936 ;
  assign n9915 = n9914 ^ n9378 ;
  assign n9950 = n9949 ^ n9915 ;
  assign n13430 = n9914 & n9950 ;
  assign n13426 = n9351 & ~n9377 ;
  assign n11081 = ~n9946 & ~n9947 ;
  assign n11082 = n9378 & n11081 ;
  assign n11083 = ~n9936 & n11082 ;
  assign n13427 = ~n9119 & ~n11083 ;
  assign n13428 = n13426 & n13427 ;
  assign n13429 = n13428 ^ n11083 ;
  assign n13431 = ~n11097 & ~n13429 ;
  assign n13432 = n13430 & n13431 ;
  assign n13433 = n13432 ^ n13429 ;
  assign n13434 = ~n11100 & ~n13433 ;
  assign n13435 = ~n11078 & n13434 ;
  assign n13436 = n11097 & n13435 ;
  assign n13437 = n13436 ^ n13434 ;
  assign n13438 = n13437 ^ n13433 ;
  assign n10272 = ~x701 & ~x702 ;
  assign n10256 = x702 ^ x701 ;
  assign n10273 = n10272 ^ n10256 ;
  assign n10270 = ~x699 & ~x700 ;
  assign n10257 = x700 ^ x699 ;
  assign n10271 = n10270 ^ n10257 ;
  assign n10300 = n10273 ^ n10271 ;
  assign n10301 = n10270 ^ x698 ;
  assign n10302 = n10301 ^ n10272 ;
  assign n10307 = n10302 ^ n10273 ;
  assign n10304 = n10272 ^ n10270 ;
  assign n10303 = n10270 & n10272 ;
  assign n10305 = n10304 ^ n10303 ;
  assign n10306 = n10302 & n10305 ;
  assign n10308 = n10307 ^ n10306 ;
  assign n10309 = n10300 & n10308 ;
  assign n10310 = n10309 ^ n10271 ;
  assign n10277 = x701 ^ x698 ;
  assign n10278 = n10277 ^ x700 ;
  assign n10279 = n10278 ^ x702 ;
  assign n10275 = x701 ^ x699 ;
  assign n10280 = n10279 ^ n10275 ;
  assign n10281 = n10280 ^ x702 ;
  assign n10282 = n10281 ^ x701 ;
  assign n10283 = n10282 ^ n10275 ;
  assign n10287 = n10275 ^ x700 ;
  assign n10288 = n10287 ^ x702 ;
  assign n10289 = n10288 ^ n10275 ;
  assign n10290 = ~n10283 & ~n10289 ;
  assign n10291 = ~x701 & n10290 ;
  assign n10294 = n10291 ^ n10290 ;
  assign n10292 = n10291 ^ n10275 ;
  assign n10293 = n10280 & n10292 ;
  assign n10295 = n10294 ^ n10293 ;
  assign n10296 = n10295 ^ x701 ;
  assign n10299 = n10296 ^ x697 ;
  assign n10297 = ~x697 & ~n10296 ;
  assign n10462 = n10299 ^ n10297 ;
  assign n10463 = n10310 & n10462 ;
  assign n10329 = ~x693 & ~x694 ;
  assign n10261 = x694 ^ x693 ;
  assign n10330 = n10329 ^ n10261 ;
  assign n10340 = n10330 ^ x692 ;
  assign n10341 = n10340 ^ x691 ;
  assign n10342 = ~x695 & ~x696 ;
  assign n10262 = x696 ^ x695 ;
  assign n10345 = n10342 ^ n10262 ;
  assign n10365 = n10345 ^ n10330 ;
  assign n10367 = n10365 ^ n10342 ;
  assign n10369 = n10367 ^ n10345 ;
  assign n10344 = n10369 ^ x691 ;
  assign n10348 = n10329 ^ n10262 ;
  assign n10346 = n10329 & n10345 ;
  assign n10347 = n10346 ^ n10342 ;
  assign n10349 = n10348 ^ n10347 ;
  assign n10350 = n10349 ^ n10342 ;
  assign n10351 = n10350 ^ x692 ;
  assign n10352 = ~n10344 & n10351 ;
  assign n10353 = ~n10341 & n10352 ;
  assign n10354 = n10353 ^ n10342 ;
  assign n10331 = n10261 ^ x696 ;
  assign n10332 = n10331 ^ n10329 ;
  assign n10334 = n10332 ^ n10261 ;
  assign n10335 = ~n10334 & ~n10367 ;
  assign n10336 = n10330 & n10335 ;
  assign n10337 = n10336 ^ n10332 ;
  assign n10355 = n10354 ^ n10337 ;
  assign n10356 = ~x692 & n10355 ;
  assign n10357 = n10356 ^ n10337 ;
  assign n10366 = n10365 ^ n10349 ;
  assign n10374 = ~x692 & ~n10342 ;
  assign n10375 = n10374 ^ n10342 ;
  assign n10376 = ~n10366 & ~n10375 ;
  assign n10377 = n10376 ^ n10365 ;
  assign n10378 = n10374 ^ n10262 ;
  assign n10379 = n10378 ^ n10376 ;
  assign n10380 = n10377 & ~n10379 ;
  assign n10381 = n10380 ^ n10330 ;
  assign n10459 = x691 & n10381 ;
  assign n10460 = ~n10357 & n10459 ;
  assign n10461 = n10460 ^ n10381 ;
  assign n10464 = n10463 ^ n10461 ;
  assign n10392 = n10303 ^ x697 ;
  assign n10393 = ~n10306 & ~n10392 ;
  assign n10320 = x694 ^ x692 ;
  assign n10321 = x696 ^ x691 ;
  assign n10324 = ~x694 & ~n10321 ;
  assign n10325 = n10324 ^ x691 ;
  assign n10326 = ~n10320 & n10325 ;
  assign n10327 = ~n10261 & n10326 ;
  assign n10328 = ~x695 & n10327 ;
  assign n10358 = n10342 ^ x692 ;
  assign n10359 = n10330 & n10358 ;
  assign n10360 = n10346 ^ x692 ;
  assign n10361 = n10359 & ~n10360 ;
  assign n10362 = n10361 ^ n10346 ;
  assign n10384 = ~n10362 & n10381 ;
  assign n10385 = n10384 ^ n10357 ;
  assign n10386 = ~x691 & n10385 ;
  assign n10387 = n10386 ^ n10357 ;
  assign n10388 = ~n10328 & n10387 ;
  assign n10389 = n10388 ^ n10297 ;
  assign n10311 = n10310 ^ n10299 ;
  assign n10312 = n10311 ^ n10296 ;
  assign n10316 = ~n10295 & n10310 ;
  assign n10317 = n10316 ^ x701 ;
  assign n10318 = n10312 & ~n10317 ;
  assign n10319 = n10318 ^ n10299 ;
  assign n10390 = n10389 ^ n10319 ;
  assign n10274 = n10271 & n10273 ;
  assign n10298 = n10274 & n10297 ;
  assign n10391 = n10390 ^ n10298 ;
  assign n10394 = n10393 ^ n10391 ;
  assign n10255 = x698 ^ x697 ;
  assign n10259 = n10288 ^ n10255 ;
  assign n10263 = n10262 ^ n10261 ;
  assign n10260 = x692 ^ x691 ;
  assign n10264 = n10263 ^ n10260 ;
  assign n10269 = n10259 & n10264 ;
  assign n10456 = n10388 ^ n10269 ;
  assign n10457 = n10394 & n10456 ;
  assign n10458 = n10457 ^ n10388 ;
  assign n10465 = n10464 ^ n10458 ;
  assign n10215 = x689 & x690 ;
  assign n10211 = x690 ^ x689 ;
  assign n10216 = n10215 ^ n10211 ;
  assign n10217 = ~x687 & ~x688 ;
  assign n10221 = ~n10215 & n10217 ;
  assign n10210 = x688 ^ x687 ;
  assign n10218 = n10217 ^ n10210 ;
  assign n10219 = n10215 & ~n10218 ;
  assign n10222 = n10221 ^ n10219 ;
  assign n10220 = n10215 ^ x688 ;
  assign n10223 = n10222 ^ n10220 ;
  assign n10224 = n10223 ^ x687 ;
  assign n10235 = n10216 & ~n10224 ;
  assign n10234 = n10224 ^ n10216 ;
  assign n10236 = n10235 ^ n10234 ;
  assign n10237 = ~x686 & n10236 ;
  assign n10212 = n10211 ^ n10210 ;
  assign n10209 = x686 ^ x685 ;
  assign n10213 = n10212 ^ n10209 ;
  assign n10230 = n10221 ^ n10213 ;
  assign n10231 = n10221 ^ x685 ;
  assign n10232 = ~n10230 & n10231 ;
  assign n10225 = ~n10219 & ~n10224 ;
  assign n10226 = x686 & n10225 ;
  assign n10227 = n10216 & n10226 ;
  assign n10228 = n10227 ^ n10225 ;
  assign n10229 = n10228 ^ n10224 ;
  assign n10233 = n10232 ^ n10229 ;
  assign n10238 = n10237 ^ n10233 ;
  assign n10205 = x680 ^ x679 ;
  assign n10204 = x684 ^ x683 ;
  assign n10247 = n10204 ^ x680 ;
  assign n10207 = x682 ^ x681 ;
  assign n10248 = n10247 ^ n10207 ;
  assign n10249 = n10205 & ~n10248 ;
  assign n10250 = n10249 ^ x679 ;
  assign n10240 = x683 & x684 ;
  assign n10239 = x681 & x682 ;
  assign n10241 = n10240 ^ n10239 ;
  assign n10242 = n10239 ^ n10207 ;
  assign n10243 = n10240 ^ n10204 ;
  assign n10244 = n10242 & n10243 ;
  assign n10245 = n10244 ^ n10240 ;
  assign n10246 = ~n10241 & ~n10245 ;
  assign n10251 = n10250 ^ n10246 ;
  assign n10454 = n10238 & ~n10251 ;
  assign n10421 = n10239 ^ x679 ;
  assign n10424 = n10421 ^ n10241 ;
  assign n10419 = n10239 ^ x680 ;
  assign n10429 = n10424 ^ n10419 ;
  assign n10420 = n10245 ^ n10241 ;
  assign n10422 = n10421 ^ n10420 ;
  assign n10430 = n10429 ^ n10422 ;
  assign n10431 = n10430 ^ n10241 ;
  assign n10433 = n10429 & n10431 ;
  assign n10426 = n10422 ^ n10241 ;
  assign n10427 = n10426 ^ n10240 ;
  assign n10428 = ~n10244 & n10427 ;
  assign n10434 = n10433 ^ n10428 ;
  assign n10435 = n10434 ^ n10426 ;
  assign n10436 = n10433 ^ n10424 ;
  assign n10437 = n10436 ^ n10426 ;
  assign n10438 = n10435 & n10437 ;
  assign n10439 = ~n10241 & n10438 ;
  assign n10440 = n10439 ^ n10433 ;
  assign n10441 = n10440 ^ n10431 ;
  assign n10449 = n10441 ^ n10239 ;
  assign n10452 = n10449 ^ n10419 ;
  assign n10477 = n10454 ^ n10452 ;
  assign n10206 = n10205 ^ n10204 ;
  assign n10208 = n10207 ^ n10206 ;
  assign n10214 = n10213 ^ n10208 ;
  assign n10265 = n10264 ^ n10259 ;
  assign n10266 = n10265 ^ n10213 ;
  assign n10267 = n10214 & n10266 ;
  assign n10252 = n10251 ^ n10238 ;
  assign n10253 = n10252 ^ n10213 ;
  assign n10268 = n10267 ^ n10253 ;
  assign n10395 = n10394 ^ n10269 ;
  assign n10405 = n10395 ^ n10252 ;
  assign n10406 = ~n10268 & ~n10405 ;
  assign n10407 = n10406 ^ n10252 ;
  assign n10478 = n10477 ^ n10407 ;
  assign n10412 = ~n10222 & ~n10236 ;
  assign n10413 = n10412 ^ n10235 ;
  assign n10414 = x686 & n10413 ;
  assign n10415 = n10414 ^ n10235 ;
  assign n10416 = x685 & n10415 ;
  assign n10417 = n10229 & n10416 ;
  assign n10418 = n10417 ^ n10229 ;
  assign n10479 = n10478 ^ n10418 ;
  assign n11023 = n10465 & n10479 ;
  assign n11024 = n10454 ^ n10407 ;
  assign n11025 = n10477 & n11024 ;
  assign n11026 = n11025 ^ n10452 ;
  assign n11027 = n11023 & n11026 ;
  assign n10474 = n10461 ^ n10458 ;
  assign n10475 = ~n10464 & ~n10474 ;
  assign n10476 = n10475 ^ n10458 ;
  assign n10453 = n10452 ^ n10418 ;
  assign n10480 = n10418 ^ n10407 ;
  assign n10481 = n10453 & ~n10480 ;
  assign n10488 = n10418 & n10481 ;
  assign n10482 = n10465 ^ n10454 ;
  assign n10483 = n10482 ^ n10481 ;
  assign n10489 = n10488 ^ n10483 ;
  assign n10490 = ~n10479 & ~n10489 ;
  assign n10491 = n10490 ^ n10483 ;
  assign n11022 = n10476 & n10491 ;
  assign n11028 = n11027 ^ n11022 ;
  assign n10045 = x667 & ~x668 ;
  assign n10047 = x671 & x672 ;
  assign n10046 = x672 ^ x671 ;
  assign n10048 = n10047 ^ n10046 ;
  assign n10049 = n10045 & n10048 ;
  assign n10050 = x670 ^ x669 ;
  assign n10051 = n10047 ^ x670 ;
  assign n10052 = n10050 & ~n10051 ;
  assign n10053 = n10052 ^ x669 ;
  assign n10054 = n10049 & n10053 ;
  assign n10055 = n10054 ^ n10045 ;
  assign n10056 = n10055 ^ x667 ;
  assign n10057 = ~x669 & ~x670 ;
  assign n10058 = n10057 ^ n10050 ;
  assign n10059 = n10050 ^ x672 ;
  assign n10060 = n10059 ^ n10057 ;
  assign n10061 = n10060 ^ x671 ;
  assign n10062 = n10060 ^ n10050 ;
  assign n10063 = ~n10061 & ~n10062 ;
  assign n10064 = n10058 & n10063 ;
  assign n10065 = n10064 ^ n10060 ;
  assign n10066 = x668 & n10065 ;
  assign n10067 = n10056 & n10066 ;
  assign n10068 = n10067 ^ n10056 ;
  assign n10069 = x668 & n10048 ;
  assign n10072 = n10069 ^ n10047 ;
  assign n10169 = n10050 ^ n10047 ;
  assign n10172 = ~n10072 & ~n10169 ;
  assign n10173 = n10172 ^ n10050 ;
  assign n10174 = ~n10057 & ~n10173 ;
  assign n10175 = ~n10068 & n10174 ;
  assign n10102 = ~x677 & ~x678 ;
  assign n10101 = x678 ^ x677 ;
  assign n10103 = n10102 ^ n10101 ;
  assign n10105 = x675 & x676 ;
  assign n10106 = ~n10103 & n10105 ;
  assign n10104 = n10103 ^ x676 ;
  assign n10108 = x676 ^ x675 ;
  assign n10109 = n10104 & n10108 ;
  assign n10128 = n10109 ^ x675 ;
  assign n10129 = ~n10106 & n10128 ;
  assign n10130 = x674 & n10129 ;
  assign n10131 = ~n10102 & n10130 ;
  assign n10132 = n10131 ^ n10129 ;
  assign n10133 = n10132 ^ n10128 ;
  assign n10144 = x673 & ~n10133 ;
  assign n10145 = x675 ^ x674 ;
  assign n10146 = n10145 ^ x676 ;
  assign n10147 = n10146 ^ x678 ;
  assign n10154 = n10147 ^ n10145 ;
  assign n10155 = x678 ^ x674 ;
  assign n10156 = ~n10154 & ~n10155 ;
  assign n10157 = n10156 ^ x675 ;
  assign n10148 = x677 ^ x675 ;
  assign n10160 = n10157 ^ n10148 ;
  assign n10161 = ~n10156 & n10160 ;
  assign n10162 = n10161 ^ n10157 ;
  assign n10163 = ~n10147 & n10162 ;
  assign n10164 = n10163 ^ n10157 ;
  assign n10165 = n10144 & n10164 ;
  assign n10166 = n10165 ^ n10133 ;
  assign n10167 = n10166 ^ n10068 ;
  assign n10176 = n10175 ^ n10167 ;
  assign n10114 = x677 ^ x673 ;
  assign n10115 = n10114 ^ x678 ;
  assign n10112 = x674 ^ x673 ;
  assign n10113 = n10112 ^ n10108 ;
  assign n10116 = n10115 ^ n10113 ;
  assign n10123 = ~x678 & ~n10105 ;
  assign n10124 = ~n10101 & n10123 ;
  assign n10125 = n10124 ^ n10101 ;
  assign n10126 = n10125 ^ n10113 ;
  assign n10127 = n10116 & ~n10126 ;
  assign n10134 = n10133 ^ n10127 ;
  assign n10107 = n10106 ^ n10104 ;
  assign n10110 = n10109 ^ n10107 ;
  assign n10111 = ~x674 & n10110 ;
  assign n10135 = n10134 ^ n10111 ;
  assign n10073 = ~n10051 & ~n10072 ;
  assign n10070 = n10069 ^ n10051 ;
  assign n10071 = x669 & ~n10070 ;
  assign n10074 = n10073 ^ n10071 ;
  assign n10075 = ~x667 & n10074 ;
  assign n10077 = n10075 ^ n10068 ;
  assign n10078 = ~x671 & ~n10077 ;
  assign n10080 = x672 ^ x669 ;
  assign n10079 = x672 ^ x668 ;
  assign n10081 = n10080 ^ n10079 ;
  assign n10082 = n10081 ^ x672 ;
  assign n10084 = x668 & n10082 ;
  assign n10085 = n10084 ^ x672 ;
  assign n10137 = x668 ^ x667 ;
  assign n10088 = x672 ^ x670 ;
  assign n10089 = n10088 ^ n10079 ;
  assign n10090 = n10137 ^ n10089 ;
  assign n10092 = n10079 ^ n10050 ;
  assign n10093 = n10092 ^ x672 ;
  assign n10094 = ~n10090 & n10093 ;
  assign n10097 = n10094 ^ x669 ;
  assign n10098 = ~n10085 & ~n10097 ;
  assign n10099 = n10078 & n10098 ;
  assign n10100 = n10099 ^ n10077 ;
  assign n10136 = n10135 ^ n10100 ;
  assign n10117 = n10113 ^ n10101 ;
  assign n10138 = n10050 ^ n10046 ;
  assign n10139 = n10138 ^ n10137 ;
  assign n10140 = n10117 & n10139 ;
  assign n10141 = n10140 ^ n10135 ;
  assign n10142 = n10136 & ~n10141 ;
  assign n10143 = n10142 ^ n10135 ;
  assign n10177 = n10176 ^ n10143 ;
  assign n9977 = x657 & x658 ;
  assign n9976 = x659 & x660 ;
  assign n9978 = n9977 ^ n9976 ;
  assign n10013 = n9976 ^ x655 ;
  assign n10016 = n10013 ^ n9978 ;
  assign n10011 = n9976 ^ x656 ;
  assign n10021 = n10016 ^ n10011 ;
  assign n9979 = x660 ^ x659 ;
  assign n9980 = n9979 ^ n9976 ;
  assign n9981 = x658 ^ x657 ;
  assign n9982 = n9981 ^ n9977 ;
  assign n9983 = n9980 & n9982 ;
  assign n9984 = n9983 ^ n9977 ;
  assign n10012 = n9984 ^ n9978 ;
  assign n10014 = n10013 ^ n10012 ;
  assign n10022 = n10021 ^ n10014 ;
  assign n10023 = n10022 ^ n9978 ;
  assign n10025 = n10021 & n10023 ;
  assign n10018 = n10014 ^ n9978 ;
  assign n10019 = n10018 ^ n9977 ;
  assign n10020 = ~n9983 & n10019 ;
  assign n10026 = n10025 ^ n10020 ;
  assign n10027 = n10026 ^ n10018 ;
  assign n10028 = n10025 ^ n10016 ;
  assign n10029 = n10028 ^ n10018 ;
  assign n10030 = n10027 & n10029 ;
  assign n10031 = ~n9978 & n10030 ;
  assign n10032 = n10031 ^ n10025 ;
  assign n10033 = n10032 ^ n10023 ;
  assign n10041 = n10033 ^ n9976 ;
  assign n10044 = n10041 ^ n10011 ;
  assign n10178 = n10177 ^ n10044 ;
  assign n10180 = n10139 ^ n10117 ;
  assign n9962 = x662 ^ x661 ;
  assign n9954 = x664 ^ x663 ;
  assign n10004 = n9962 ^ n9954 ;
  assign n9956 = x666 ^ x665 ;
  assign n10005 = n10004 ^ n9956 ;
  assign n9986 = x656 ^ x655 ;
  assign n10002 = n9986 ^ n9981 ;
  assign n10003 = n10002 ^ n9979 ;
  assign n10181 = n10005 ^ n10003 ;
  assign n10182 = n10181 ^ n10139 ;
  assign n10183 = n10180 & ~n10182 ;
  assign n10184 = n10183 ^ n10117 ;
  assign n10006 = n10003 & n10005 ;
  assign n10185 = n10184 ^ n10006 ;
  assign n9987 = n9981 ^ x656 ;
  assign n9988 = n9987 ^ n9979 ;
  assign n9989 = n9986 & ~n9988 ;
  assign n9990 = n9989 ^ x655 ;
  assign n9985 = ~n9978 & ~n9984 ;
  assign n9991 = n9990 ^ n9985 ;
  assign n9952 = x665 & x666 ;
  assign n9951 = ~x663 & ~x664 ;
  assign n9963 = n9952 ^ n9951 ;
  assign n9953 = ~n9951 & n9952 ;
  assign n9964 = n9963 ^ n9953 ;
  assign n9955 = n9954 ^ n9951 ;
  assign n9957 = n9956 ^ n9952 ;
  assign n9958 = ~n9955 & n9957 ;
  assign n9960 = ~n9953 & ~n9958 ;
  assign n9959 = n9958 ^ n9953 ;
  assign n9961 = n9960 ^ n9959 ;
  assign n9965 = n9964 ^ n9961 ;
  assign n9966 = n9957 ^ n9955 ;
  assign n9967 = n9966 ^ n9958 ;
  assign n9968 = x662 & ~n9967 ;
  assign n9969 = n9965 & n9968 ;
  assign n9970 = n9969 ^ n9960 ;
  assign n9971 = ~n9962 & ~n9970 ;
  assign n9972 = n9971 ^ n9960 ;
  assign n9992 = n9991 ^ n9972 ;
  assign n9974 = ~x662 & n9967 ;
  assign n9975 = n9951 & n9974 ;
  assign n9993 = n9992 ^ n9975 ;
  assign n9994 = n9993 ^ n9991 ;
  assign n9997 = n9974 ^ n9961 ;
  assign n9995 = n9957 ^ x662 ;
  assign n9996 = n9964 & n9995 ;
  assign n9998 = n9997 ^ n9996 ;
  assign n9999 = ~x661 & ~n9998 ;
  assign n10000 = n9994 & n9999 ;
  assign n10001 = n10000 ^ n9993 ;
  assign n10188 = n10185 ^ n10001 ;
  assign n10191 = n10184 & n10188 ;
  assign n10189 = n10188 ^ n10140 ;
  assign n10190 = n10136 & ~n10189 ;
  assign n10192 = n10191 ^ n10190 ;
  assign n10195 = n10192 ^ n10044 ;
  assign n10196 = ~n10178 & ~n10195 ;
  assign n10197 = n10196 ^ n10177 ;
  assign n11029 = n11028 ^ n10197 ;
  assign n10198 = n10166 ^ n10143 ;
  assign n10199 = n10176 & ~n10198 ;
  assign n10200 = n10199 ^ n10166 ;
  assign n11030 = n11029 ^ n10200 ;
  assign n10007 = n10006 ^ n9991 ;
  assign n10008 = ~n10001 & ~n10007 ;
  assign n10009 = n10008 ^ n9991 ;
  assign n10201 = n10200 ^ n10009 ;
  assign n10202 = n10201 ^ n10197 ;
  assign n9973 = n9961 & n9972 ;
  assign n10010 = n10009 ^ n9973 ;
  assign n10179 = n10178 ^ n9973 ;
  assign n10193 = n10192 ^ n10179 ;
  assign n10194 = n10010 & ~n10193 ;
  assign n10203 = n10202 ^ n10194 ;
  assign n11031 = n11030 ^ n10203 ;
  assign n11016 = ~n9973 & ~n10009 ;
  assign n11010 = n10200 ^ n10197 ;
  assign n11011 = n11010 ^ n10203 ;
  assign n11017 = n11016 ^ n11011 ;
  assign n11018 = n10203 & ~n11017 ;
  assign n11032 = n11031 ^ n11018 ;
  assign n11019 = n11010 & ~n11018 ;
  assign n11020 = n10203 ^ n10200 ;
  assign n11021 = n11019 & n11020 ;
  assign n11033 = n11032 ^ n11021 ;
  assign n10492 = n10491 ^ n10476 ;
  assign n10397 = n10188 ^ n10136 ;
  assign n10396 = n10395 ^ n10268 ;
  assign n10398 = n10397 ^ n10396 ;
  assign n10399 = n10181 ^ n10180 ;
  assign n10400 = n10265 ^ n10214 ;
  assign n10401 = n10399 & n10400 ;
  assign n10402 = n10401 ^ n10396 ;
  assign n10403 = n10398 & ~n10402 ;
  assign n10404 = n10403 ^ n10396 ;
  assign n10493 = n10492 ^ n10404 ;
  assign n10455 = n10454 ^ n10453 ;
  assign n10466 = n10465 ^ n10455 ;
  assign n10467 = n10466 ^ n10407 ;
  assign n10468 = n10467 ^ n10404 ;
  assign n10470 = n10192 ^ n10177 ;
  assign n10469 = n10044 ^ n10010 ;
  assign n10471 = n10470 ^ n10469 ;
  assign n10472 = n10471 ^ n10404 ;
  assign n10473 = ~n10468 & n10472 ;
  assign n10494 = n10493 ^ n10473 ;
  assign n11034 = n10492 ^ n10203 ;
  assign n11035 = ~n10494 & n11034 ;
  assign n11036 = n11035 ^ n10492 ;
  assign n11108 = n11036 ^ n11028 ;
  assign n11109 = ~n11033 & n11108 ;
  assign n11110 = n11109 ^ n11028 ;
  assign n10497 = x710 ^ x709 ;
  assign n10552 = ~x711 & ~x712 ;
  assign n10499 = x714 ^ x713 ;
  assign n10549 = x713 & ~n10499 ;
  assign n10670 = n10549 ^ n10499 ;
  assign n10671 = ~n10552 & n10670 ;
  assign n10496 = x712 ^ x711 ;
  assign n10666 = n10552 ^ n10496 ;
  assign n10548 = x709 & ~n10497 ;
  assign n10667 = x714 & n10548 ;
  assign n10668 = ~n10666 & n10667 ;
  assign n10669 = n10668 ^ n10548 ;
  assign n10672 = n10671 ^ n10669 ;
  assign n10677 = ~n10549 & n10666 ;
  assign n10678 = n10677 ^ n10669 ;
  assign n10679 = n10672 & ~n10678 ;
  assign n10680 = ~n10497 & n10679 ;
  assign n10560 = ~x705 & ~x706 ;
  assign n10501 = x706 ^ x705 ;
  assign n10688 = n10560 ^ n10501 ;
  assign n10502 = x704 ^ x703 ;
  assign n10556 = x703 & ~n10502 ;
  assign n10700 = x708 & n10556 ;
  assign n10701 = ~n10688 & n10700 ;
  assign n10702 = n10701 ^ n10556 ;
  assign n10504 = x708 ^ x707 ;
  assign n10557 = x707 & ~n10504 ;
  assign n10690 = n10557 ^ n10504 ;
  assign n10691 = ~n10560 & n10690 ;
  assign n10703 = n10702 ^ n10691 ;
  assign n10707 = ~n10557 & n10688 ;
  assign n10708 = n10707 ^ n10691 ;
  assign n10709 = n10703 & n10708 ;
  assign n10689 = n10688 ^ n10557 ;
  assign n10696 = x704 & n10691 ;
  assign n10697 = n10696 ^ n10688 ;
  assign n10698 = ~n10689 & n10697 ;
  assign n10699 = n10698 ^ n10557 ;
  assign n10710 = n10709 ^ n10702 ;
  assign n10711 = ~n10699 & n10710 ;
  assign n10712 = ~n10502 & n10711 ;
  assign n10713 = n10709 & n10712 ;
  assign n10714 = n10713 ^ n10711 ;
  assign n10715 = n10714 ^ n10699 ;
  assign n10681 = n10679 ^ n10669 ;
  assign n10723 = n10715 ^ ~n10681 ;
  assign n10686 = x710 & n10671 ;
  assign n10687 = n10686 ^ n10666 ;
  assign n10716 = n10715 ^ n10549 ;
  assign n10717 = n10716 ^ n10666 ;
  assign n10718 = n10717 ^ n10715 ;
  assign n10719 = n10687 & ~n10718 ;
  assign n10720 = n10719 ^ n10716 ;
  assign n10724 = n10723 ^ n10720 ;
  assign n10725 = n10680 & ~n10724 ;
  assign n10726 = n10725 ^ n10723 ;
  assign n10558 = n10557 ^ n10556 ;
  assign n10503 = n10502 ^ n10501 ;
  assign n10554 = n10504 ^ n10502 ;
  assign n10555 = n10503 & ~n10554 ;
  assign n10559 = n10558 ^ n10555 ;
  assign n10561 = n10560 ^ n10559 ;
  assign n10550 = n10549 ^ n10548 ;
  assign n10498 = n10497 ^ n10496 ;
  assign n10546 = n10499 ^ n10497 ;
  assign n10547 = n10498 & ~n10546 ;
  assign n10551 = n10550 ^ n10547 ;
  assign n10553 = n10552 ^ n10551 ;
  assign n10562 = n10561 ^ n10553 ;
  assign n10500 = n10499 ^ n10498 ;
  assign n10505 = n10504 ^ n10503 ;
  assign n10521 = n10500 & n10505 ;
  assign n10663 = n10553 ^ n10521 ;
  assign n10664 = ~n10562 & ~n10663 ;
  assign n10665 = n10664 ^ n10521 ;
  assign n10727 = n10726 ^ n10665 ;
  assign n10539 = x721 & x722 ;
  assign n10538 = ~x725 & ~x726 ;
  assign n10540 = n10539 ^ n10538 ;
  assign n10536 = ~x723 & ~x724 ;
  assign n10515 = x726 ^ x725 ;
  assign n10537 = n10536 ^ n10515 ;
  assign n10541 = n10540 ^ n10537 ;
  assign n10513 = x722 ^ x721 ;
  assign n10512 = x724 ^ x723 ;
  assign n10514 = n10513 ^ n10512 ;
  assign n10534 = n10515 ^ n10513 ;
  assign n10535 = n10514 & ~n10534 ;
  assign n10542 = n10541 ^ n10535 ;
  assign n10531 = x715 & x716 ;
  assign n10530 = ~x719 & ~x720 ;
  assign n10532 = n10531 ^ n10530 ;
  assign n10528 = ~x717 & ~x718 ;
  assign n10510 = x720 ^ x719 ;
  assign n10529 = n10528 ^ n10510 ;
  assign n10533 = n10532 ^ n10529 ;
  assign n10543 = n10542 ^ n10533 ;
  assign n10508 = x716 ^ x715 ;
  assign n10507 = x718 ^ x717 ;
  assign n10509 = n10508 ^ n10507 ;
  assign n10526 = n10510 ^ n10508 ;
  assign n10527 = n10509 & ~n10526 ;
  assign n10544 = n10543 ^ n10527 ;
  assign n10511 = n10510 ^ n10509 ;
  assign n10516 = n10515 ^ n10514 ;
  assign n10523 = n10511 & n10516 ;
  assign n10590 = n10544 ^ n10523 ;
  assign n10594 = n10562 ^ n10521 ;
  assign n10595 = n10590 & n10594 ;
  assign n10506 = n10505 ^ n10500 ;
  assign n10517 = n10516 ^ n10511 ;
  assign n10518 = n10517 ^ n10500 ;
  assign n10519 = n10506 & ~n10518 ;
  assign n10520 = n10519 ^ n10505 ;
  assign n10522 = n10521 ^ n10520 ;
  assign n10592 = n10562 ^ n10544 ;
  assign n10593 = n10522 & n10592 ;
  assign n10596 = n10595 ^ n10593 ;
  assign n10875 = n10727 ^ n10596 ;
  assign n10876 = n10715 ^ n10665 ;
  assign n10877 = ~n10726 & n10876 ;
  assign n10878 = n10877 ^ n10715 ;
  assign n10884 = ~n10596 & ~n10878 ;
  assign n10623 = n10536 ^ n10512 ;
  assign n10635 = x726 & n10539 ;
  assign n10636 = ~n10623 & n10635 ;
  assign n10637 = n10636 ^ n10539 ;
  assign n10626 = ~n10536 & ~n10538 ;
  assign n10638 = n10637 ^ n10626 ;
  assign n10624 = n10538 ^ n10515 ;
  assign n10643 = n10623 & n10624 ;
  assign n10644 = n10643 ^ n10637 ;
  assign n10645 = n10638 & ~n10644 ;
  assign n10625 = n10624 ^ n10623 ;
  assign n10631 = x722 & n10626 ;
  assign n10632 = n10631 ^ n10623 ;
  assign n10633 = n10625 & n10632 ;
  assign n10634 = n10633 ^ n10624 ;
  assign n10646 = n10645 ^ n10637 ;
  assign n10647 = n10634 & n10646 ;
  assign n10648 = ~n10513 & n10647 ;
  assign n10649 = n10645 & n10648 ;
  assign n10650 = n10649 ^ n10647 ;
  assign n10651 = n10650 ^ n10634 ;
  assign n10604 = ~n10528 & ~n10530 ;
  assign n10600 = n10528 ^ n10507 ;
  assign n10601 = x720 & n10531 ;
  assign n10602 = ~n10600 & n10601 ;
  assign n10603 = n10602 ^ n10531 ;
  assign n10605 = n10604 ^ n10603 ;
  assign n10608 = n10530 ^ n10510 ;
  assign n10611 = n10600 & n10608 ;
  assign n10612 = n10611 ^ n10603 ;
  assign n10613 = n10605 & ~n10612 ;
  assign n10614 = n10613 ^ n10603 ;
  assign n10656 = n10651 ^ ~n10614 ;
  assign n10652 = n10651 ^ n10608 ;
  assign n10615 = n10608 ^ n10600 ;
  assign n10620 = x716 & n10604 ;
  assign n10621 = n10620 ^ n10600 ;
  assign n10622 = n10615 & n10621 ;
  assign n10653 = n10652 ^ n10622 ;
  assign n10657 = n10656 ^ n10653 ;
  assign n10658 = ~n10508 & n10613 ;
  assign n10659 = n10657 & n10658 ;
  assign n10660 = n10659 ^ n10656 ;
  assign n10597 = n10542 ^ n10523 ;
  assign n10598 = n10544 & n10597 ;
  assign n10599 = n10598 ^ n10542 ;
  assign n10661 = n10660 ^ n10599 ;
  assign n10879 = n10878 ^ n10661 ;
  assign n10885 = n10884 ^ n10879 ;
  assign n10886 = n10875 & ~n10885 ;
  assign n10887 = n10886 ^ n10879 ;
  assign n10811 = ~x741 & ~x742 ;
  assign n10566 = x742 ^ x741 ;
  assign n10822 = n10811 ^ n10566 ;
  assign n10813 = ~x743 & ~x744 ;
  assign n10567 = x744 ^ x743 ;
  assign n10821 = n10813 ^ n10567 ;
  assign n10847 = n10822 ^ n10821 ;
  assign n10812 = n10811 ^ x740 ;
  assign n10814 = n10813 ^ n10812 ;
  assign n10848 = n10822 ^ n10814 ;
  assign n10816 = n10813 ^ n10811 ;
  assign n10815 = n10811 & n10813 ;
  assign n10817 = n10816 ^ n10815 ;
  assign n10818 = n10814 & n10817 ;
  assign n10849 = n10848 ^ n10818 ;
  assign n10850 = n10847 & n10849 ;
  assign n10851 = n10850 ^ n10821 ;
  assign n10826 = x743 ^ x740 ;
  assign n10827 = n10826 ^ x742 ;
  assign n10828 = n10827 ^ x744 ;
  assign n10824 = x743 ^ x741 ;
  assign n10829 = n10828 ^ n10824 ;
  assign n10830 = n10829 ^ x744 ;
  assign n10831 = n10830 ^ x743 ;
  assign n10832 = n10831 ^ n10824 ;
  assign n10836 = n10824 ^ x742 ;
  assign n10837 = n10836 ^ x744 ;
  assign n10838 = n10837 ^ n10824 ;
  assign n10839 = ~n10832 & ~n10838 ;
  assign n10840 = ~x743 & n10839 ;
  assign n10843 = n10840 ^ n10839 ;
  assign n10841 = n10840 ^ n10824 ;
  assign n10842 = n10829 & n10841 ;
  assign n10844 = n10843 ^ n10842 ;
  assign n10845 = n10844 ^ x743 ;
  assign n10861 = ~x739 & ~n10845 ;
  assign n10846 = n10845 ^ x739 ;
  assign n10943 = n10861 ^ n10846 ;
  assign n10944 = n10851 & n10943 ;
  assign n10570 = x746 ^ x745 ;
  assign n10571 = x748 ^ x747 ;
  assign n10771 = ~x749 & ~x750 ;
  assign n10573 = x750 ^ x749 ;
  assign n10774 = n10771 ^ n10573 ;
  assign n10781 = n10774 ^ x748 ;
  assign n10782 = n10571 & n10781 ;
  assign n10783 = n10782 ^ x747 ;
  assign n10765 = ~x747 & ~x748 ;
  assign n10775 = n10765 & n10774 ;
  assign n10784 = n10783 ^ n10775 ;
  assign n10766 = n10765 ^ n10571 ;
  assign n10785 = n10784 ^ n10766 ;
  assign n10786 = n10785 ^ n10783 ;
  assign n10789 = x746 & n10786 ;
  assign n10790 = n10789 ^ n10783 ;
  assign n10791 = ~n10570 & n10790 ;
  assign n10792 = n10791 ^ n10783 ;
  assign n10767 = x745 & x746 ;
  assign n10768 = ~n10766 & n10767 ;
  assign n10793 = n10792 ^ n10768 ;
  assign n10794 = ~x750 & n10793 ;
  assign n10795 = n10794 ^ n10792 ;
  assign n10796 = n10782 ^ n10781 ;
  assign n10797 = n10796 ^ n10775 ;
  assign n10798 = n10783 & ~n10797 ;
  assign n10800 = x746 & ~n10771 ;
  assign n10801 = n10798 & n10800 ;
  assign n10802 = n10801 ^ n10797 ;
  assign n10803 = ~n10795 & ~n10802 ;
  assign n10804 = x749 & n10794 ;
  assign n10805 = n10803 & n10804 ;
  assign n10806 = n10805 ^ n10803 ;
  assign n10945 = n10944 ^ n10806 ;
  assign n10823 = n10821 & n10822 ;
  assign n10864 = n10823 & n10861 ;
  assign n10852 = n10851 ^ n10846 ;
  assign n10853 = n10852 ^ n10845 ;
  assign n10857 = ~n10844 & n10851 ;
  assign n10858 = n10857 ^ x743 ;
  assign n10859 = n10853 & ~n10858 ;
  assign n10860 = n10859 ^ n10846 ;
  assign n10862 = n10861 ^ n10860 ;
  assign n10865 = n10864 ^ n10862 ;
  assign n10819 = n10815 ^ x739 ;
  assign n10820 = ~n10818 & ~n10819 ;
  assign n10866 = n10865 ^ n10820 ;
  assign n10772 = n10771 ^ x745 ;
  assign n10773 = n10772 ^ x746 ;
  assign n10777 = n10786 ^ n10772 ;
  assign n10778 = n10773 & ~n10777 ;
  assign n10779 = n10778 ^ n10775 ;
  assign n10780 = n10771 & n10779 ;
  assign n10807 = n10806 ^ n10780 ;
  assign n10867 = n10866 ^ n10807 ;
  assign n10770 = ~x745 & ~x746 ;
  assign n10809 = n10780 ^ n10779 ;
  assign n10810 = n10770 & n10809 ;
  assign n10868 = n10867 ^ n10810 ;
  assign n10769 = ~n10573 & n10768 ;
  assign n10869 = n10868 ^ n10769 ;
  assign n10565 = x740 ^ x739 ;
  assign n10569 = n10837 ^ n10565 ;
  assign n10572 = n10571 ^ n10570 ;
  assign n10574 = n10573 ^ n10572 ;
  assign n10731 = n10569 & n10574 ;
  assign n10940 = n10866 ^ n10731 ;
  assign n10941 = n10869 & n10940 ;
  assign n10942 = n10941 ^ n10866 ;
  assign n10946 = n10945 ^ n10942 ;
  assign n10906 = x733 & x734 ;
  assign n10737 = ~x735 & ~x736 ;
  assign n10577 = x736 ^ x735 ;
  assign n10760 = n10737 ^ n10577 ;
  assign n10907 = x738 & ~n10760 ;
  assign n10908 = n10906 & ~n10907 ;
  assign n10903 = ~x737 & ~x738 ;
  assign n10904 = ~n10737 & ~n10903 ;
  assign n10909 = n10908 ^ n10904 ;
  assign n10579 = x738 ^ x737 ;
  assign n10910 = n10903 ^ n10579 ;
  assign n10915 = n10760 & n10910 ;
  assign n10916 = n10915 ^ n10904 ;
  assign n10917 = n10909 & n10916 ;
  assign n10919 = n10917 ^ n10908 ;
  assign n10576 = x734 ^ x733 ;
  assign n10905 = ~n10576 & n10904 ;
  assign n10918 = n10905 & n10917 ;
  assign n10920 = n10919 ^ n10918 ;
  assign n10921 = n10910 ^ n10760 ;
  assign n10922 = x734 & n10904 ;
  assign n10923 = n10922 ^ n10760 ;
  assign n10924 = n10921 & ~n10923 ;
  assign n10925 = n10924 ^ n10760 ;
  assign n10926 = ~n10920 & ~n10925 ;
  assign n10927 = n10926 ^ n10920 ;
  assign n10953 = n10946 ^ n10927 ;
  assign n10578 = n10577 ^ n10576 ;
  assign n10759 = n10578 ^ x737 ;
  assign n10761 = n10760 ^ x738 ;
  assign n10762 = n10759 & n10761 ;
  assign n10583 = x730 ^ x729 ;
  assign n10744 = x729 ^ x728 ;
  assign n10936 = ~n10583 & n10744 ;
  assign n10582 = x732 ^ x731 ;
  assign n10584 = n10583 ^ n10582 ;
  assign n10581 = x728 ^ x727 ;
  assign n10585 = n10584 ^ n10581 ;
  assign n10750 = x727 & ~n10585 ;
  assign n10751 = n10750 ^ x728 ;
  assign n10746 = n10583 ^ x728 ;
  assign n10747 = n10746 ^ x731 ;
  assign n10748 = n10582 & n10747 ;
  assign n10749 = n10748 ^ x731 ;
  assign n10752 = n10751 ^ n10749 ;
  assign n10757 = n10936 ^ n10752 ;
  assign n10735 = x737 ^ x734 ;
  assign n10738 = n10737 ^ x737 ;
  assign n10741 = ~n10735 & n10738 ;
  assign n10739 = n10738 ^ x734 ;
  assign n10740 = x733 & n10739 ;
  assign n10742 = n10741 ^ n10740 ;
  assign n10758 = n10757 ^ n10742 ;
  assign n10763 = n10762 ^ n10758 ;
  assign n10580 = n10579 ^ n10578 ;
  assign n10733 = n10580 & n10585 ;
  assign n10900 = n10757 ^ n10733 ;
  assign n10901 = n10763 & n10900 ;
  assign n10902 = n10901 ^ n10733 ;
  assign n10954 = n10946 ^ n10902 ;
  assign n10955 = n10953 & n10954 ;
  assign n10956 = n10955 ^ n10946 ;
  assign n10928 = n10927 ^ n10902 ;
  assign n10963 = n10946 ^ n10928 ;
  assign n10930 = n10750 ^ n10749 ;
  assign n10931 = n10749 ^ x728 ;
  assign n10937 = n10936 ^ n10931 ;
  assign n10938 = n10930 & ~n10937 ;
  assign n10939 = n10938 ^ n10750 ;
  assign n10893 = n10869 ^ n10731 ;
  assign n10575 = n10574 ^ n10569 ;
  assign n10586 = n10585 ^ n10580 ;
  assign n10730 = n10575 & n10586 ;
  assign n10894 = n10893 ^ n10730 ;
  assign n10897 = n10893 ^ n10763 ;
  assign n10898 = n10894 & ~n10897 ;
  assign n10896 = ~n10733 & n10893 ;
  assign n10899 = n10898 ^ n10896 ;
  assign n10957 = n10939 ^ n10899 ;
  assign n10958 = n10939 ^ n10902 ;
  assign n10959 = n10958 ^ n10927 ;
  assign n10960 = n10959 ^ n10946 ;
  assign n10961 = ~n10957 & n10960 ;
  assign n10964 = n10963 ^ n10961 ;
  assign n10965 = ~n10956 & ~n10964 ;
  assign n10947 = n10946 ^ n10939 ;
  assign n10929 = n10928 ^ n10899 ;
  assign n10948 = n10947 ^ n10929 ;
  assign n10968 = n10927 ^ n10899 ;
  assign n10969 = n10928 & n10968 ;
  assign n10970 = n10969 ^ n10927 ;
  assign n10971 = n10946 & n10970 ;
  assign n10972 = ~n10948 & n10971 ;
  assign n10974 = n10942 ^ n10806 ;
  assign n10975 = n10945 & ~n10974 ;
  assign n10976 = n10975 ^ n10806 ;
  assign n11001 = ~n10972 & n10976 ;
  assign n11002 = ~n10965 & n11001 ;
  assign n11003 = n11002 ^ n10965 ;
  assign n10888 = n10651 ^ n10599 ;
  assign n10889 = n10660 & ~n10888 ;
  assign n10890 = n10889 ^ n10651 ;
  assign n11005 = n11003 ^ n10890 ;
  assign n11004 = n11003 ^ n10878 ;
  assign n11006 = n11005 ^ n11004 ;
  assign n11007 = ~n10887 & ~n11006 ;
  assign n11008 = n11007 ^ n11005 ;
  assign n10564 = n10517 ^ n10506 ;
  assign n10587 = n10586 ^ n10575 ;
  assign n10588 = n10564 & n10587 ;
  assign n10524 = n10523 ^ n10522 ;
  assign n10525 = n10524 ^ n10521 ;
  assign n10545 = n10544 ^ n10525 ;
  assign n10563 = n10562 ^ n10545 ;
  assign n10589 = n10588 ^ n10563 ;
  assign n10732 = n10731 ^ n10730 ;
  assign n10734 = n10733 ^ n10732 ;
  assign n10764 = n10763 ^ n10734 ;
  assign n10870 = n10869 ^ n10764 ;
  assign n10662 = n10661 ^ n10596 ;
  assign n10728 = n10727 ^ n10662 ;
  assign n10729 = n10728 ^ n10588 ;
  assign n10871 = n10870 ^ n10729 ;
  assign n10872 = n10871 ^ n10728 ;
  assign n10873 = n10589 & ~n10872 ;
  assign n10874 = n10873 ^ n10729 ;
  assign n10891 = n10890 ^ n10887 ;
  assign n10949 = n10948 ^ n10891 ;
  assign n10892 = n10891 ^ n10728 ;
  assign n10950 = n10949 ^ n10892 ;
  assign n10951 = n10874 & ~n10950 ;
  assign n10952 = n10951 ^ n10949 ;
  assign n10973 = n10972 ^ n10965 ;
  assign n10977 = n10976 ^ n10973 ;
  assign n10998 = n10977 ^ n10891 ;
  assign n10999 = ~n10952 & ~n10998 ;
  assign n11000 = n10999 ^ n10891 ;
  assign n11105 = n11003 ^ n11000 ;
  assign n11106 = n11008 & n11105 ;
  assign n11107 = n11106 ^ n11003 ;
  assign n11111 = n11110 ^ n11107 ;
  assign n13439 = n13438 ^ n11111 ;
  assign n11037 = n11036 ^ n11033 ;
  assign n11009 = n11008 ^ n11000 ;
  assign n11038 = n11037 ^ n11009 ;
  assign n10978 = n10977 ^ n10952 ;
  assign n10495 = n10494 ^ n10203 ;
  assign n10979 = n10978 ^ n10495 ;
  assign n10981 = n10471 ^ n10468 ;
  assign n10994 = n10981 ^ n10978 ;
  assign n10980 = n10948 ^ n10874 ;
  assign n10982 = n10981 ^ n10980 ;
  assign n10986 = n10870 ^ n10589 ;
  assign n10983 = n10400 ^ n10399 ;
  assign n10984 = n10587 ^ n10564 ;
  assign n10985 = n10983 & n10984 ;
  assign n10987 = n10986 ^ n10985 ;
  assign n11048 = n10985 ^ n10401 ;
  assign n11049 = n11048 ^ n10398 ;
  assign n10990 = ~n10987 & ~n11049 ;
  assign n10991 = n10990 ^ n10986 ;
  assign n10992 = n10991 ^ n10980 ;
  assign n10993 = ~n10982 & ~n10992 ;
  assign n10995 = n10994 ^ n10993 ;
  assign n10996 = n10979 & ~n10995 ;
  assign n10997 = n10996 ^ n10978 ;
  assign n11073 = n11009 ^ n10997 ;
  assign n11074 = n11038 & ~n11073 ;
  assign n11075 = n11074 ^ n11037 ;
  assign n11039 = n11038 ^ n10997 ;
  assign n11040 = n11039 ^ n9950 ;
  assign n11042 = n10995 ^ n10495 ;
  assign n11041 = n9934 ^ n9916 ;
  assign n11043 = n11042 ^ n11041 ;
  assign n11046 = n10991 ^ n10982 ;
  assign n11044 = n9930 ^ n9929 ;
  assign n11047 = n11046 ^ n11044 ;
  assign n11052 = n9924 ^ n9923 ;
  assign n11051 = n10984 ^ n10983 ;
  assign n11054 = n11052 ^ n11051 ;
  assign n11053 = ~n11051 & ~n11052 ;
  assign n11055 = n11054 ^ n11053 ;
  assign n11050 = n11049 ^ n10986 ;
  assign n11056 = n11055 ^ n11050 ;
  assign n11061 = ~n9925 & ~n11050 ;
  assign n11062 = n11061 ^ n9922 ;
  assign n11063 = n11056 & ~n11062 ;
  assign n11064 = n11063 ^ n11055 ;
  assign n11065 = n11064 ^ n11044 ;
  assign n11066 = ~n11047 & n11065 ;
  assign n11045 = n11044 ^ n11042 ;
  assign n11067 = n11066 ^ n11045 ;
  assign n11068 = ~n11043 & ~n11067 ;
  assign n11069 = n11068 ^ n11042 ;
  assign n11070 = n11069 ^ n9950 ;
  assign n11071 = ~n11040 & ~n11070 ;
  assign n11072 = n11071 ^ n11039 ;
  assign n11076 = n11075 ^ n11072 ;
  assign n11101 = n11100 ^ n9378 ;
  assign n11102 = n11101 ^ n11097 ;
  assign n11084 = n11083 ^ n11082 ;
  assign n11085 = ~n9914 & n11084 ;
  assign n11103 = n11102 ^ n11085 ;
  assign n11077 = n9948 ^ n9378 ;
  assign n11079 = n11078 ^ n9378 ;
  assign n11080 = ~n11077 & n11079 ;
  assign n11104 = n11103 ^ n11080 ;
  assign n11112 = n11111 ^ n11104 ;
  assign n11113 = n11112 ^ n11072 ;
  assign n11114 = ~n11076 & ~n11113 ;
  assign n13440 = n13439 ^ n11114 ;
  assign n11115 = n11107 ^ n11104 ;
  assign n11116 = n11111 & n11115 ;
  assign n13441 = n13440 ^ n11116 ;
  assign n13379 = n13378 ^ n13371 ;
  assign n13380 = n13379 ^ n13368 ;
  assign n13381 = n13380 ^ n12254 ;
  assign n11120 = n11111 ^ n11075 ;
  assign n11119 = n11104 ^ n11072 ;
  assign n11121 = n11120 ^ n11119 ;
  assign n13382 = n13381 ^ n11121 ;
  assign n13412 = n13366 ^ n13321 ;
  assign n13422 = n13412 ^ n11121 ;
  assign n13409 = n13362 ^ n13361 ;
  assign n13384 = n13357 ^ n13323 ;
  assign n13410 = n13409 ^ n13384 ;
  assign n13383 = n11064 ^ n11047 ;
  assign n13385 = n13384 ^ n13383 ;
  assign n13394 = n13349 ^ n13332 ;
  assign n13399 = ~n11053 & n13394 ;
  assign n13400 = n13399 ^ n9925 ;
  assign n13401 = n11055 & ~n13400 ;
  assign n11057 = n11050 ^ n9922 ;
  assign n13402 = n13401 ^ n11057 ;
  assign n13403 = n11055 ^ n9925 ;
  assign n13386 = n13350 ^ n12073 ;
  assign n13387 = n13386 ^ n13338 ;
  assign n13390 = n13389 ^ n13387 ;
  assign n13391 = n13390 ^ n12080 ;
  assign n13392 = n13391 ^ n13329 ;
  assign n13404 = n13403 ^ n13392 ;
  assign n13405 = n13404 ^ n13401 ;
  assign n13406 = ~n13402 & ~n13405 ;
  assign n13393 = n13392 ^ n13383 ;
  assign n13407 = n13406 ^ n13393 ;
  assign n13408 = n13385 & n13407 ;
  assign n13411 = n13410 ^ n13408 ;
  assign n13415 = n13412 ^ n13409 ;
  assign n13413 = n11067 ^ n11041 ;
  assign n13414 = n13413 ^ n13412 ;
  assign n13416 = n13415 ^ n13414 ;
  assign n13417 = n13411 & ~n13416 ;
  assign n13418 = n13417 ^ n13414 ;
  assign n13419 = n11069 ^ n11040 ;
  assign n13420 = n13419 ^ n13412 ;
  assign n13421 = ~n13418 & n13420 ;
  assign n13423 = n13422 ^ n13421 ;
  assign n13424 = n13382 & n13423 ;
  assign n13425 = n13424 ^ n13381 ;
  assign n13442 = n13441 ^ n13425 ;
  assign n11117 = ~n11107 & n11116 ;
  assign n11118 = n11114 & n11117 ;
  assign n13443 = n13442 ^ n11118 ;
  assign n13493 = n13492 ^ n13443 ;
  assign n13495 = n13494 ^ n13493 ;
  assign n13497 = n8719 ^ n8718 ;
  assign n13496 = n13423 ^ n13381 ;
  assign n13498 = n13497 ^ n13496 ;
  assign n13500 = n8714 ^ n8689 ;
  assign n13499 = n13419 ^ n13418 ;
  assign n13501 = n13500 ^ n13499 ;
  assign n13502 = n8711 ^ n8692 ;
  assign n13530 = n13502 ^ n13500 ;
  assign n13503 = n13413 ^ n13411 ;
  assign n13504 = n13503 ^ n13502 ;
  assign n13506 = n13407 ^ n13384 ;
  assign n13505 = n8708 ^ n8707 ;
  assign n13507 = n13506 ^ n13505 ;
  assign n13509 = n8700 ^ n5742 ;
  assign n13510 = n13509 ^ n8697 ;
  assign n13511 = n13510 ^ n8698 ;
  assign n13512 = n13511 ^ n5739 ;
  assign n13508 = n13402 ^ n13392 ;
  assign n13513 = n13512 ^ n13508 ;
  assign n13514 = n5741 ^ n5740 ;
  assign n13515 = n13514 ^ n8696 ;
  assign n13518 = n13394 ^ n11054 ;
  assign n13521 = n13515 & n13518 ;
  assign n13522 = n13521 ^ n13508 ;
  assign n13523 = ~n13513 & n13522 ;
  assign n13524 = n13523 ^ n13512 ;
  assign n13525 = n13524 ^ n13505 ;
  assign n13526 = ~n13507 & ~n13525 ;
  assign n13527 = n13526 ^ n13506 ;
  assign n13528 = n13527 ^ n13502 ;
  assign n13529 = ~n13504 & ~n13528 ;
  assign n13531 = n13530 ^ n13529 ;
  assign n13532 = ~n13501 & ~n13531 ;
  assign n13533 = n13532 ^ n13500 ;
  assign n13534 = n13533 ^ n13496 ;
  assign n13535 = ~n13498 & ~n13534 ;
  assign n13536 = n13535 ^ n13497 ;
  assign n13537 = n13536 ^ n13494 ;
  assign n13538 = ~n13495 & n13537 ;
  assign n13539 = n13538 ^ n13494 ;
  assign n5715 = n4541 & n5714 ;
  assign n5717 = n5716 ^ n5715 ;
  assign n3336 = ~n2157 & n3335 ;
  assign n3337 = ~n3258 & n3328 ;
  assign n3338 = ~n3297 & n3337 ;
  assign n3339 = n2156 & n3338 ;
  assign n3340 = n3339 ^ n3337 ;
  assign n3341 = n3340 ^ n3258 ;
  assign n3342 = n3336 & ~n3341 ;
  assign n3343 = n3342 ^ n3341 ;
  assign n5718 = n5717 ^ n3343 ;
  assign n5773 = n5769 ^ n3343 ;
  assign n5722 = n5721 ^ n3343 ;
  assign n5774 = n5773 ^ n5722 ;
  assign n5775 = n5770 & n5774 ;
  assign n5776 = n5775 ^ n5722 ;
  assign n5777 = ~n5718 & n5776 ;
  assign n5778 = n5777 ^ n5717 ;
  assign n5779 = ~n5715 & n5778 ;
  assign n5780 = n5769 ^ n5721 ;
  assign n5781 = ~n5722 & ~n5780 ;
  assign n5782 = n5770 & n5781 ;
  assign n5783 = n5782 ^ n3343 ;
  assign n5784 = n5779 & n5783 ;
  assign n5785 = n5784 ^ n5778 ;
  assign n13540 = n13539 ^ n5785 ;
  assign n8767 = ~n5759 & n5769 ;
  assign n8789 = ~n5717 & ~n8767 ;
  assign n8741 = ~n4538 & ~n5711 ;
  assign n8742 = n5721 & ~n8741 ;
  assign n8743 = ~n4534 & n8742 ;
  assign n8744 = ~n5679 & n8743 ;
  assign n8745 = n8744 ^ n8742 ;
  assign n8746 = n8745 ^ n8741 ;
  assign n8739 = n4534 & n5592 ;
  assign n8740 = n5666 & n8739 ;
  assign n8747 = n8746 ^ n8740 ;
  assign n8748 = n8746 ^ n4532 ;
  assign n8749 = n5711 ^ n4538 ;
  assign n8750 = n8749 ^ n8741 ;
  assign n8751 = n8750 ^ n8746 ;
  assign n8752 = n8751 ^ n8741 ;
  assign n8754 = ~n4534 & ~n5721 ;
  assign n8755 = n8752 & n8754 ;
  assign n8756 = n8755 ^ n8751 ;
  assign n8757 = ~n8748 & n8756 ;
  assign n8758 = n8757 ^ n8746 ;
  assign n8759 = ~n5769 & ~n8758 ;
  assign n8760 = n8746 & n8759 ;
  assign n8761 = ~n8747 & n8760 ;
  assign n8762 = n8761 ^ n8759 ;
  assign n8763 = n8762 ^ n5769 ;
  assign n8764 = n8763 ^ n5671 ;
  assign n8768 = n8767 ^ n5759 ;
  assign n8769 = n8768 ^ n5770 ;
  assign n8770 = n8769 ^ n5759 ;
  assign n8771 = n5759 ^ n4541 ;
  assign n8772 = n8771 ^ n5759 ;
  assign n8773 = ~n8770 & ~n8772 ;
  assign n8774 = n8773 ^ n5759 ;
  assign n8775 = ~n5716 & n8774 ;
  assign n8765 = n5759 ^ n5606 ;
  assign n8766 = n8765 ^ n8763 ;
  assign n8776 = n8775 ^ n8766 ;
  assign n8777 = n8763 & n8776 ;
  assign n8778 = n8777 ^ n5606 ;
  assign n8779 = n8778 ^ n8763 ;
  assign n8780 = ~n8764 & n8779 ;
  assign n8782 = n5666 & n8777 ;
  assign n8783 = n8780 & n8782 ;
  assign n8781 = n8780 ^ n8763 ;
  assign n8784 = n8783 ^ n8781 ;
  assign n8787 = n8784 ^ n3343 ;
  assign n8734 = n5769 ^ n5715 ;
  assign n8737 = n5759 & ~n8734 ;
  assign n8738 = n8737 ^ n5715 ;
  assign n8785 = ~n5721 & n8784 ;
  assign n8786 = ~n8738 & n8785 ;
  assign n8788 = n8787 ^ n8786 ;
  assign n8790 = n8788 ^ n8787 ;
  assign n8791 = n8789 & n8790 ;
  assign n8792 = n8791 ^ n8788 ;
  assign n8679 = n8678 ^ n8639 ;
  assign n8685 = ~n8679 & n8684 ;
  assign n8686 = n7466 & ~n8685 ;
  assign n8727 = n8726 ^ n8722 ;
  assign n8728 = ~n8724 & ~n8727 ;
  assign n8729 = n8728 ^ n8722 ;
  assign n8687 = n8685 ^ n8683 ;
  assign n8730 = n8729 ^ n8687 ;
  assign n8731 = n8730 ^ n8729 ;
  assign n8732 = n8686 & ~n8731 ;
  assign n8733 = n8732 ^ n8730 ;
  assign n8793 = n8792 ^ n8733 ;
  assign n8794 = n8793 ^ n5785 ;
  assign n13541 = n13540 ^ n8794 ;
  assign n13545 = ~n13466 & ~n13469 ;
  assign n13547 = ~n11075 & ~n11107 ;
  assign n13546 = n11107 ^ n11075 ;
  assign n13548 = n13547 ^ n13546 ;
  assign n13549 = n13548 ^ n13438 ;
  assign n13550 = n11104 & ~n13549 ;
  assign n13551 = n13548 & n13550 ;
  assign n13552 = n13551 ^ n13548 ;
  assign n13553 = n13552 ^ n11110 ;
  assign n13554 = n13551 ^ n13549 ;
  assign n13555 = n11119 & ~n13554 ;
  assign n13556 = n13553 & n13555 ;
  assign n13557 = n13556 ^ n13552 ;
  assign n13558 = n13438 & ~n13547 ;
  assign n13559 = n11072 & n13558 ;
  assign n13560 = n13559 ^ n13547 ;
  assign n13561 = n13559 ^ n11110 ;
  assign n13562 = n13561 ^ n13559 ;
  assign n13563 = n13559 ^ n11119 ;
  assign n13564 = ~n13562 & ~n13563 ;
  assign n13565 = ~n13560 & n13564 ;
  assign n13566 = n13565 ^ n13560 ;
  assign n13567 = n13566 ^ n13547 ;
  assign n13568 = n13557 & ~n13567 ;
  assign n13569 = n13568 ^ n13489 ;
  assign n13570 = n13569 ^ n13568 ;
  assign n13571 = n13545 & ~n13570 ;
  assign n13572 = n13571 ^ n13569 ;
  assign n13542 = n13492 ^ n13425 ;
  assign n13543 = ~n13443 & ~n13542 ;
  assign n13544 = n13543 ^ n13492 ;
  assign n13573 = n13572 ^ n13544 ;
  assign n13574 = n13573 ^ n8793 ;
  assign n13577 = n13541 & n13574 ;
  assign n13578 = n13577 ^ n8794 ;
  assign n13587 = ~n13494 & ~n13536 ;
  assign n13588 = n13536 ^ n13495 ;
  assign n13589 = n13587 & n13588 ;
  assign n13590 = n13518 ^ n13515 ;
  assign n13591 = n13518 ^ n13513 ;
  assign n13592 = ~x1000 & n13591 ;
  assign n13593 = ~n13590 & n13592 ;
  assign n13594 = n13524 ^ n13507 ;
  assign n13595 = n13506 ^ n13504 ;
  assign n13596 = n13595 ^ n13526 ;
  assign n13597 = ~n13594 & ~n13596 ;
  assign n13598 = ~n13593 & n13597 ;
  assign n13599 = n13598 ^ n13526 ;
  assign n13600 = n13599 ^ n13595 ;
  assign n13601 = n13531 ^ n13499 ;
  assign n13602 = n13533 ^ n13498 ;
  assign n13603 = ~n13601 & n13602 ;
  assign n13604 = n13600 & n13603 ;
  assign n13605 = ~n13589 & n13604 ;
  assign n13606 = n13589 ^ n13588 ;
  assign n13607 = ~n13574 & ~n13606 ;
  assign n13608 = n13607 ^ n13539 ;
  assign n13609 = n13605 & ~n13608 ;
  assign n13583 = n8792 ^ n8729 ;
  assign n13584 = ~n8733 & n13583 ;
  assign n13585 = n13584 ^ n8792 ;
  assign n13579 = n13568 ^ n13544 ;
  assign n13580 = n13572 & ~n13579 ;
  assign n13581 = n13580 ^ n13544 ;
  assign n13582 = n13581 ^ n5785 ;
  assign n13586 = n13585 ^ n13582 ;
  assign n13610 = n13609 ^ n13586 ;
  assign n13611 = n13578 & ~n13610 ;
  assign n13612 = n13611 ^ n5785 ;
  assign n13613 = n13609 ^ n13581 ;
  assign n13614 = n13585 ^ n13581 ;
  assign n13615 = ~n13613 & ~n13614 ;
  assign n13616 = n13615 ^ n13581 ;
  assign n13617 = ~n13612 & n13616 ;
  assign y0 = ~n13617 ;
endmodule
