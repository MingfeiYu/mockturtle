module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 ;
  output y0 ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2008 , n2009 , n2010 , n2011 , n2012 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2215 , n2216 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2228 , n2229 , n2232 , n2233 , n2235 , n2236 , n2237 , n2238 , n2244 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2339 , n2340 , n2342 , n2343 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2370 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2506 , n2507 , n2508 , n2509 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2529 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2555 , n2556 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2753 , n2754 , n2755 , n2756 , n2757 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2770 , n2771 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2783 , n2784 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2816 , n2817 , n2818 , n2819 , n2820 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2833 , n2834 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2846 , n2847 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2978 , n2979 , n2982 , n2983 , n2984 , n2985 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3022 , n3023 , n3024 , n3025 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3095 , n3096 , n3100 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3133 , n3134 , n3135 , n3136 , n3137 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3425 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3673 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3740 , n3741 , n3742 , n3743 , n3744 , n3747 , n3748 , n3749 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3792 , n3794 , n3795 , n3796 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3814 , n3815 , n3816 , n3817 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3859 , n3860 , n3862 , n3863 , n3864 , n3865 , n3867 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3887 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3928 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3946 , n3947 , n3948 , n3949 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3968 , n3970 , n3971 , n3973 , n3974 , n3976 , n3977 , n3978 , n3979 , n3981 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4031 , n4032 , n4033 , n4034 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4058 , n4059 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4164 , n4165 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4177 , n4178 , n4181 , n4182 , n4184 , n4185 , n4186 , n4187 , n4193 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4223 , n4224 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4236 , n4237 , n4240 , n4241 , n4243 , n4244 , n4245 , n4246 , n4252 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4838 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4941 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4967 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5049 , n5050 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5062 , n5063 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5370 , n5371 , n5372 , n5373 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5632 , n5633 , n5634 , n5635 , n5636 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5677 , n5678 , n5679 , n5680 , n5681 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5708 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5731 , n5732 , n5735 , n5736 , n5737 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6037 , n6038 , n6039 , n6040 , n6042 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6191 , n6192 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6204 , n6205 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6220 , n6221 , n6222 , n6223 , n6229 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6288 , n6289 , n6292 , n6294 , n6295 , n6296 , n6297 , n6298 , n6301 , n6302 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6588 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6609 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7041 , n7042 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7054 , n7055 , n7058 , n7059 , n7060 , n7062 , n7063 , n7064 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7259 , n7260 , n7261 , n7262 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7596 , n7597 , n7598 , n7599 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7618 , n7620 , n7621 , n7623 , n7624 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7656 , n7657 , n7658 , n7659 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7701 , n7702 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7848 , n7849 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7861 , n7862 , n7865 , n7866 , n7868 , n7869 , n7870 , n7871 , n7877 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7910 , n7911 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8028 , n8029 , n8030 , n8031 , n8032 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8084 , n8085 , n8086 , n8091 , n8092 , n8093 , n8094 , n8095 , n8098 , n8099 , n8104 , n8105 , n8106 , n8108 , n8109 , n8110 , n8113 , n8114 , n8115 , n8116 , n8117 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8153 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8177 , n8178 , n8180 , n8182 , n8184 , n8186 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8201 , n8204 , n8205 , n8208 , n8209 , n8210 , n8211 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8238 , n8239 , n8240 , n8241 , n8242 , n8244 , n8245 , n8246 , n8247 , n8248 , n8253 , n8254 , n8256 , n8258 , n8259 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8284 , n8287 , n8288 , n8289 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8348 , n8351 , n8352 , n8356 , n8359 , n8360 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8507 , n8508 , n8510 , n8512 , n8514 , n8516 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8531 , n8534 , n8535 , n8539 , n8540 , n8542 , n8544 , n8546 , n8548 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8563 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8704 , n8706 , n8707 , n8708 , n8709 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8757 , n8758 , n8759 , n8761 , n8762 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8915 , n8916 , n8917 , n8918 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9062 , n9064 , n9065 , n9066 , n9067 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9110 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9140 , n9141 , n9142 , n9143 , n9144 , n9146 , n9147 , n9148 , n9149 , n9150 , n9152 , n9157 , n9158 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9269 , n9275 , n9300 , n9301 , n9302 , n9303 , n9305 , n9306 , n9307 , n9308 , n9311 , n9312 , n9313 , n9317 , n9318 , n9319 , n9329 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9360 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9450 , n9451 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9577 , n9578 , n9579 , n9580 , n9581 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9774 , n9775 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9787 , n9788 , n9790 , n9792 , n9794 , n9796 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9811 , n9814 , n9815 , n9818 , n9819 , n9820 , n9821 , n9826 , n9831 , n9834 , n9835 , n9836 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9886 , n9887 , n9888 , n9889 , n9890 , n9893 , n9894 , n9895 , n9896 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9923 , n9924 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9995 , n9996 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10037 , n10042 , n10045 , n10046 , n10047 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10063 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10086 , n10087 , n10089 , n10091 , n10093 , n10095 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10110 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10123 , n10124 , n10125 , n10131 , n10134 , n10135 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10180 , n10181 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10217 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10445 , n10446 , n10447 , n10450 , n10452 , n10453 , n10455 , n10457 , n10459 , n10460 , n10461 , n10462 , n10463 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10561 , n10562 , n10563 , n10564 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10609 , n10610 , n10611 , n10612 , n10613 , n10619 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10631 , n10632 , n10633 , n10636 , n10637 , n10638 , n10639 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10688 , n10689 , n10690 , n10691 , n10692 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10754 , n10755 , n10756 , n10757 , n10758 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10903 , n10904 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10964 , n10965 , n10971 , n10972 , n10973 , n10975 , n10976 , n10977 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11079 , n11080 , n11081 , n11082 , n11083 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11132 , n11133 , n11139 , n11140 , n11141 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11171 , n11172 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11243 , n11244 , n11245 , n11246 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11293 , n11294 , n11295 , n11300 , n11301 , n11302 , n11303 , n11304 , n11307 , n11308 , n11309 , n11310 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11343 , n11344 , n11346 , n11351 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11402 , n11403 , n11404 , n11405 , n11406 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11424 , n11425 , n11426 , n11427 , n11428 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11496 , n11497 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11553 , n11554 , n11555 , n11556 , n11557 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11671 , n11672 , n11673 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11699 , n11702 , n11703 , n11704 , n11705 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11717 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11798 , n11799 , n11800 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11824 , n11825 , n11826 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11995 , n11997 , n11998 , n12000 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12013 , n12014 , n12015 , n12016 , n12017 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12251 , n12252 , n12253 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12600 , n12601 , n12602 , n12603 , n12604 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12765 , n12766 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12814 , n12815 , n12816 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12864 , n12865 , n12866 , n12867 , n12870 , n12871 , n12872 , n12873 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12929 , n12930 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12969 , n12970 , n12971 , n12972 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13013 , n13014 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13289 , n13290 , n13291 , n13292 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13397 , n13398 , n13399 ;
  assign n1209 = x150 ^ x149 ;
  assign n7354 = x149 ^ x148 ;
  assign n7358 = ~n1209 & ~n7354 ;
  assign n7353 = x147 ^ x146 ;
  assign n7355 = n7354 ^ x147 ;
  assign n7356 = n7355 ^ x150 ;
  assign n7357 = ~n7353 & n7356 ;
  assign n7359 = n7358 ^ n7357 ;
  assign n7360 = ~x145 & n7359 ;
  assign n1210 = x148 ^ x147 ;
  assign n7361 = ~n1210 & ~n7353 ;
  assign n7362 = x150 ^ x145 ;
  assign n7365 = ~x148 & ~n7362 ;
  assign n7366 = n7365 ^ x145 ;
  assign n7367 = n7361 & n7366 ;
  assign n7368 = ~x149 & n7367 ;
  assign n7369 = ~x147 & ~x148 ;
  assign n7372 = n7369 ^ n1210 ;
  assign n7373 = x145 & x146 ;
  assign n7374 = x150 & n7373 ;
  assign n7375 = ~n7372 & n7374 ;
  assign n7376 = n7375 ^ n7373 ;
  assign n7370 = ~x149 & ~x150 ;
  assign n7371 = ~n7369 & ~n7370 ;
  assign n7377 = n7376 ^ n7371 ;
  assign n7378 = n7370 ^ n1209 ;
  assign n7383 = n7372 & n7378 ;
  assign n7384 = n7383 ^ n7371 ;
  assign n7385 = n7377 & n7384 ;
  assign n1211 = x146 ^ x145 ;
  assign n7386 = n7385 ^ n7376 ;
  assign n7387 = ~n1211 & n7386 ;
  assign n7388 = n7385 & n7387 ;
  assign n7389 = n7388 ^ n7386 ;
  assign n7390 = ~n7368 & ~n7389 ;
  assign n7391 = ~n7360 & n7390 ;
  assign n1204 = x144 ^ x143 ;
  assign n7315 = x143 ^ x142 ;
  assign n7319 = ~n1204 & ~n7315 ;
  assign n7314 = x141 ^ x140 ;
  assign n7316 = n7315 ^ x141 ;
  assign n7317 = n7316 ^ x144 ;
  assign n7318 = ~n7314 & n7317 ;
  assign n7320 = n7319 ^ n7318 ;
  assign n7321 = ~x139 & n7320 ;
  assign n1205 = x142 ^ x141 ;
  assign n7322 = ~n1205 & ~n7314 ;
  assign n7323 = x144 ^ x139 ;
  assign n7326 = ~x142 & ~n7323 ;
  assign n7327 = n7326 ^ x139 ;
  assign n7328 = n7322 & n7327 ;
  assign n7329 = ~x143 & n7328 ;
  assign n7330 = ~x141 & ~x142 ;
  assign n7333 = n7330 ^ n1205 ;
  assign n7334 = x139 & x140 ;
  assign n7335 = x144 & n7334 ;
  assign n7336 = ~n7333 & n7335 ;
  assign n7337 = n7336 ^ n7334 ;
  assign n7331 = ~x143 & ~x144 ;
  assign n7332 = ~n7330 & ~n7331 ;
  assign n7338 = n7337 ^ n7332 ;
  assign n7339 = n7331 ^ n1204 ;
  assign n7344 = n7333 & n7339 ;
  assign n7345 = n7344 ^ n7332 ;
  assign n7346 = n7338 & n7345 ;
  assign n1206 = x140 ^ x139 ;
  assign n7347 = n7346 ^ n7337 ;
  assign n7348 = ~n1206 & n7347 ;
  assign n7349 = n7346 & n7348 ;
  assign n7350 = n7349 ^ n7347 ;
  assign n7351 = ~n7329 & ~n7350 ;
  assign n7352 = ~n7321 & n7351 ;
  assign n7392 = n7391 ^ n7352 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1208 = n1207 ^ n1204 ;
  assign n1212 = n1211 ^ n1210 ;
  assign n1213 = n1212 ^ n1209 ;
  assign n8019 = n1208 & n1213 ;
  assign n8020 = n8019 ^ n7352 ;
  assign n8021 = n7392 & ~n8020 ;
  assign n8022 = n8021 ^ n7391 ;
  assign n1214 = n1213 ^ n1208 ;
  assign n1195 = x134 ^ x133 ;
  assign n1194 = x136 ^ x135 ;
  assign n1196 = n1195 ^ n1194 ;
  assign n1193 = x138 ^ x137 ;
  assign n1197 = n1196 ^ n1193 ;
  assign n1200 = x128 ^ x127 ;
  assign n1199 = x132 ^ x131 ;
  assign n1201 = n1200 ^ n1199 ;
  assign n1198 = x130 ^ x129 ;
  assign n1202 = n1201 ^ n1198 ;
  assign n7994 = n1197 & n1202 ;
  assign n8023 = n7994 ^ n1208 ;
  assign n1203 = n1202 ^ n1197 ;
  assign n8024 = n8023 ^ n1203 ;
  assign n8025 = n8024 ^ n1208 ;
  assign n8028 = ~n7392 & n8025 ;
  assign n8029 = n8028 ^ n1208 ;
  assign n8030 = n1214 & n8029 ;
  assign n8026 = n7392 ^ n1208 ;
  assign n8031 = n8030 ^ n8026 ;
  assign n7261 = x135 & x136 ;
  assign n7262 = n7261 ^ x134 ;
  assign n7265 = n1194 ^ x133 ;
  assign n7266 = ~x138 & n7265 ;
  assign n7267 = n7266 ^ x133 ;
  assign n7268 = ~n7261 & n7267 ;
  assign n7269 = n7268 ^ x133 ;
  assign n7270 = ~n7262 & n7269 ;
  assign n7271 = ~x137 & n7270 ;
  assign n7272 = x137 & x138 ;
  assign n7273 = n7272 ^ n1193 ;
  assign n7278 = n7261 & n7272 ;
  assign n7274 = n7272 ^ x136 ;
  assign n7279 = n7278 ^ n7274 ;
  assign n7275 = n1194 & ~n7274 ;
  assign n7280 = n7279 ^ n7275 ;
  assign n7276 = n7275 ^ x135 ;
  assign n7277 = n7276 ^ n7261 ;
  assign n7281 = n7280 ^ n7277 ;
  assign n7282 = n7281 ^ n7276 ;
  assign n7285 = x134 & n7282 ;
  assign n7286 = n7285 ^ n7276 ;
  assign n7287 = ~n1195 & n7286 ;
  assign n7288 = n7287 ^ n7276 ;
  assign n7289 = n7273 & n7288 ;
  assign n7290 = x133 & x134 ;
  assign n7291 = ~x138 & n7261 ;
  assign n7292 = n7290 & n7291 ;
  assign n7293 = ~n7289 & ~n7292 ;
  assign n7294 = ~x133 & n7293 ;
  assign n7295 = x134 & n7273 ;
  assign n7303 = ~n7280 & ~n7295 ;
  assign n7296 = n7276 & ~n7278 ;
  assign n7297 = ~n7295 & n7296 ;
  assign n7298 = n7297 ^ n7276 ;
  assign n7304 = n7303 ^ n7298 ;
  assign n7305 = n7294 & n7304 ;
  assign n7306 = n7305 ^ n7293 ;
  assign n7307 = ~n7271 & n7306 ;
  assign n7222 = x129 & x130 ;
  assign n7243 = x127 & x128 ;
  assign n7244 = n7222 & n7243 ;
  assign n7245 = x131 & n7244 ;
  assign n7216 = x131 & x132 ;
  assign n7220 = n7216 ^ n1199 ;
  assign n7221 = x128 & n7220 ;
  assign n7228 = n7220 ^ x127 ;
  assign n7229 = n7228 ^ x128 ;
  assign n7230 = ~n7221 & n7229 ;
  assign n7223 = n7216 & n7222 ;
  assign n7217 = n7216 ^ x130 ;
  assign n7231 = n7223 ^ n7217 ;
  assign n7218 = n1198 & ~n7217 ;
  assign n7232 = n7231 ^ n7218 ;
  assign n7233 = n7232 ^ x128 ;
  assign n7234 = n7233 ^ n7222 ;
  assign n7235 = n7234 ^ n7232 ;
  assign n7238 = ~n1200 & ~n7235 ;
  assign n7239 = n7238 ^ n7232 ;
  assign n7240 = ~n7230 & ~n7239 ;
  assign n7241 = n7240 ^ n7232 ;
  assign n7219 = n7218 ^ x129 ;
  assign n7224 = ~n7221 & ~n7223 ;
  assign n7225 = n7219 & n7224 ;
  assign n7226 = n7225 ^ n7219 ;
  assign n7227 = ~x127 & n7226 ;
  assign n7242 = n7241 ^ n7227 ;
  assign n7246 = n7245 ^ n7242 ;
  assign n7257 = ~x132 & n7244 ;
  assign n7247 = n7232 ^ n7219 ;
  assign n7248 = n7247 ^ n7222 ;
  assign n7249 = n7248 ^ n7219 ;
  assign n7252 = x128 & n7249 ;
  assign n7253 = n7252 ^ n7219 ;
  assign n7254 = ~n1200 & n7253 ;
  assign n7255 = n7254 ^ n7219 ;
  assign n7256 = n7220 & n7255 ;
  assign n7259 = n7257 ^ n7256 ;
  assign n7260 = n7246 & ~n7259 ;
  assign n7308 = n7307 ^ n7260 ;
  assign n7309 = n1208 ^ n1202 ;
  assign n7312 = ~n1203 & ~n7309 ;
  assign n7310 = n7309 ^ n1197 ;
  assign n7311 = ~n1213 & n7310 ;
  assign n7313 = n7312 ^ n7311 ;
  assign n7393 = n7392 ^ n7313 ;
  assign n8032 = n7994 ^ n7393 ;
  assign n8035 = ~n7308 & ~n8032 ;
  assign n8036 = n8035 ^ n7994 ;
  assign n8037 = n8031 & ~n8036 ;
  assign n11814 = n8022 & n8037 ;
  assign n8006 = n7378 ^ n7372 ;
  assign n8007 = x146 & n7371 ;
  assign n8008 = n8007 ^ n7372 ;
  assign n8009 = n8006 & ~n8008 ;
  assign n8010 = n8009 ^ n7372 ;
  assign n8011 = ~n7389 & ~n8010 ;
  assign n8012 = n8011 ^ n7389 ;
  assign n7999 = n7339 ^ n7333 ;
  assign n8000 = x140 & n7332 ;
  assign n8001 = n8000 ^ n7333 ;
  assign n8002 = n7999 & ~n8001 ;
  assign n8003 = n8002 ^ n7333 ;
  assign n8004 = ~n7350 & ~n8003 ;
  assign n8005 = n8004 ^ n7350 ;
  assign n8013 = n8012 ^ n8005 ;
  assign n11824 = n11814 ^ n8013 ;
  assign n8038 = n8037 ^ n8022 ;
  assign n11815 = n11814 ^ n8038 ;
  assign n7995 = n7994 ^ n7307 ;
  assign n7996 = n7308 & n7995 ;
  assign n7997 = n7996 ^ n7307 ;
  assign n7992 = n7293 & ~n7298 ;
  assign n7991 = ~n7226 & ~n7259 ;
  assign n7993 = n7992 ^ n7991 ;
  assign n7998 = n7997 ^ n7993 ;
  assign n11825 = n11815 ^ n7998 ;
  assign n11816 = n7998 & n11815 ;
  assign n11826 = n11825 ^ n11816 ;
  assign n11817 = ~n8005 & ~n8012 ;
  assign n12589 = n11817 ^ n8013 ;
  assign n11829 = n12589 ^ n11814 ;
  assign n11830 = ~n11826 & n11829 ;
  assign n11818 = n11817 ^ n11816 ;
  assign n11831 = n11830 ^ n11818 ;
  assign n11832 = n11824 & n11831 ;
  assign n11811 = n7997 ^ n7992 ;
  assign n11812 = ~n7993 & ~n11811 ;
  assign n11813 = n11812 ^ n7997 ;
  assign n11819 = n11818 ^ n11813 ;
  assign n11833 = n11832 ^ n11819 ;
  assign n12590 = ~n11813 & ~n11816 ;
  assign n7075 = ~x155 & ~x156 ;
  assign n1234 = x156 ^ x155 ;
  assign n7077 = n7075 ^ n1234 ;
  assign n7076 = x152 & ~n7075 ;
  assign n7081 = n7077 ^ n7076 ;
  assign n7078 = n7077 ^ x154 ;
  assign n7964 = n7078 ^ x153 ;
  assign n7965 = n7081 & n7964 ;
  assign n1233 = x154 ^ x153 ;
  assign n7966 = n7965 ^ n1233 ;
  assign n7967 = ~x154 & ~n7966 ;
  assign n7968 = ~n7965 & n7967 ;
  assign n7969 = n7968 ^ n7966 ;
  assign n7060 = n1233 ^ x155 ;
  assign n7062 = x155 ^ x153 ;
  assign n7036 = x156 ^ x154 ;
  assign n7037 = x156 ^ x152 ;
  assign n7059 = ~n7036 & ~n7037 ;
  assign n7063 = n7062 ^ n7059 ;
  assign n7064 = n7063 ^ x154 ;
  assign n7067 = ~n7060 & ~n7064 ;
  assign n7068 = n7067 ^ x154 ;
  assign n7069 = n7063 ^ x155 ;
  assign n7070 = n7069 ^ n7037 ;
  assign n7071 = n7070 ^ n7060 ;
  assign n7072 = n7071 ^ n7063 ;
  assign n7073 = ~n7068 & ~n7072 ;
  assign n7074 = n7073 ^ n7069 ;
  assign n7970 = x151 & n7074 ;
  assign n7971 = n7969 & n7970 ;
  assign n7972 = n7971 ^ n7969 ;
  assign n7090 = x157 & ~x158 ;
  assign n7091 = x162 ^ x159 ;
  assign n7092 = x161 ^ x160 ;
  assign n7093 = n7092 ^ x162 ;
  assign n7094 = n7091 & ~n7093 ;
  assign n7095 = n7094 ^ x162 ;
  assign n7096 = n7090 & ~n7095 ;
  assign n7100 = n7096 ^ x157 ;
  assign n7097 = n7096 ^ n7090 ;
  assign n7098 = ~x160 & ~x161 ;
  assign n7099 = n7097 & n7098 ;
  assign n7101 = n7100 ^ n7099 ;
  assign n1229 = x160 ^ x159 ;
  assign n7102 = x161 ^ x159 ;
  assign n7103 = ~n1229 & n7102 ;
  assign n1228 = x162 ^ x161 ;
  assign n7104 = n7103 ^ n1228 ;
  assign n7105 = n7104 ^ n1229 ;
  assign n7110 = x162 & ~n7103 ;
  assign n7111 = n7105 & n7110 ;
  assign n7112 = n7111 ^ n7105 ;
  assign n7113 = n7112 ^ n1229 ;
  assign n7114 = x158 & ~n7113 ;
  assign n7115 = n7101 & ~n7114 ;
  assign n7116 = x159 ^ x158 ;
  assign n7954 = x160 ^ x158 ;
  assign n7955 = n7116 & n7954 ;
  assign n7956 = n7955 ^ x158 ;
  assign n7960 = n1229 ^ x158 ;
  assign n7117 = n7092 ^ x159 ;
  assign n7957 = n7117 ^ x158 ;
  assign n7958 = ~n1228 & n7957 ;
  assign n7961 = n7960 ^ n7958 ;
  assign n7962 = n7956 & n7961 ;
  assign n7963 = ~n7115 & ~n7962 ;
  assign n7973 = n7972 ^ n7963 ;
  assign n7038 = n7037 ^ n7036 ;
  assign n7039 = n7038 ^ x156 ;
  assign n7041 = x152 & n7039 ;
  assign n7042 = n7041 ^ x156 ;
  assign n7045 = x156 ^ x153 ;
  assign n7046 = n7045 ^ n7037 ;
  assign n1232 = x152 ^ x151 ;
  assign n7047 = n7046 ^ n1232 ;
  assign n7048 = n7038 ^ n1232 ;
  assign n7049 = n7048 ^ n7037 ;
  assign n7050 = n7049 ^ x156 ;
  assign n7051 = ~n7047 & n7050 ;
  assign n7054 = n7051 ^ x154 ;
  assign n7055 = ~n7042 & ~n7054 ;
  assign n7058 = ~x155 & n7055 ;
  assign n7082 = n7078 & n7081 ;
  assign n7079 = n7078 ^ n7076 ;
  assign n7080 = x153 & n7079 ;
  assign n7083 = n7082 ^ n7080 ;
  assign n7084 = n7083 ^ n7074 ;
  assign n7087 = x151 & n7084 ;
  assign n7088 = n7087 ^ n7083 ;
  assign n7089 = ~n7058 & ~n7088 ;
  assign n7120 = ~n1228 & ~n7092 ;
  assign n7118 = n7117 ^ x162 ;
  assign n7119 = ~n7116 & n7118 ;
  assign n7121 = n7120 ^ n7119 ;
  assign n7122 = ~x157 & n7121 ;
  assign n7123 = ~n7115 & ~n7122 ;
  assign n7124 = ~n1229 & ~n7116 ;
  assign n7125 = x162 ^ x157 ;
  assign n7128 = ~x160 & ~n7125 ;
  assign n7129 = n7128 ^ x157 ;
  assign n7130 = n7124 & n7129 ;
  assign n7131 = ~x161 & n7130 ;
  assign n7132 = n7123 & ~n7131 ;
  assign n7974 = n7089 & n7132 ;
  assign n11840 = n7974 ^ n7972 ;
  assign n11841 = n7973 & ~n11840 ;
  assign n11842 = n11841 ^ n7972 ;
  assign n7135 = ~x171 & ~x172 ;
  assign n1217 = x172 ^ x171 ;
  assign n7146 = n7135 ^ n1217 ;
  assign n7137 = ~x173 & ~x174 ;
  assign n1218 = x174 ^ x173 ;
  assign n7145 = n7137 ^ n1218 ;
  assign n7147 = n7146 ^ n7145 ;
  assign n7136 = n7135 ^ x170 ;
  assign n7138 = n7137 ^ n7136 ;
  assign n7148 = n7145 ^ n7138 ;
  assign n7140 = n7137 ^ n7135 ;
  assign n7139 = n7135 & n7137 ;
  assign n7141 = n7140 ^ n7139 ;
  assign n7142 = n7138 & n7141 ;
  assign n7149 = n7148 ^ n7142 ;
  assign n7150 = n7147 & n7149 ;
  assign n7151 = n7150 ^ n7146 ;
  assign n7154 = x173 ^ x170 ;
  assign n7155 = n7154 ^ x172 ;
  assign n7156 = n7155 ^ x174 ;
  assign n7152 = x173 ^ x171 ;
  assign n7157 = n7156 ^ n7152 ;
  assign n7158 = n7157 ^ x174 ;
  assign n7159 = n7158 ^ x173 ;
  assign n7160 = n7159 ^ n7152 ;
  assign n7164 = n7152 ^ x172 ;
  assign n7165 = n7164 ^ x174 ;
  assign n7166 = n7165 ^ n7152 ;
  assign n7167 = ~n7160 & ~n7166 ;
  assign n7168 = ~x173 & n7167 ;
  assign n7171 = n7168 ^ n7167 ;
  assign n7169 = n7168 ^ n7152 ;
  assign n7170 = n7157 & n7169 ;
  assign n7172 = n7171 ^ n7170 ;
  assign n7173 = n7172 ^ x173 ;
  assign n7979 = n7173 ^ x169 ;
  assign n7209 = ~x169 & ~n7173 ;
  assign n7980 = n7979 ^ n7209 ;
  assign n7981 = n7151 & n7980 ;
  assign n7180 = x167 & x168 ;
  assign n7182 = x165 & x166 ;
  assign n7188 = n7180 & n7182 ;
  assign n7187 = n7182 ^ n7180 ;
  assign n7189 = n7188 ^ n7187 ;
  assign n1221 = x166 ^ x165 ;
  assign n7183 = n7182 ^ n1221 ;
  assign n1224 = x168 ^ x167 ;
  assign n7181 = n7180 ^ n1224 ;
  assign n7185 = n7183 ^ n7181 ;
  assign n7184 = ~n7181 & ~n7183 ;
  assign n7186 = n7185 ^ n7184 ;
  assign n7190 = n7189 ^ n7186 ;
  assign n1222 = x164 ^ x163 ;
  assign n7195 = n7189 ^ n1222 ;
  assign n7196 = n7190 & ~n7195 ;
  assign n7197 = x163 & x164 ;
  assign n7198 = ~n7188 & n7197 ;
  assign n7199 = n7198 ^ n1222 ;
  assign n7200 = n7196 & n7199 ;
  assign n7201 = n7200 ^ n7198 ;
  assign n7202 = ~n7188 & ~n7201 ;
  assign n7982 = n7981 ^ n7202 ;
  assign n7208 = n7145 & n7146 ;
  assign n7210 = n7208 & n7209 ;
  assign n7203 = n7202 ^ n7201 ;
  assign n7191 = n7181 ^ n1222 ;
  assign n7192 = n7191 ^ n7183 ;
  assign n7193 = ~n7184 & ~n7192 ;
  assign n7194 = n7190 & ~n7193 ;
  assign n7204 = n7203 ^ n7194 ;
  assign n7205 = n7204 ^ n7197 ;
  assign n7206 = n7205 ^ n7173 ;
  assign n7177 = ~x169 & ~n7172 ;
  assign n7178 = n7177 ^ x173 ;
  assign n7179 = ~n7151 & ~n7178 ;
  assign n7207 = n7206 ^ n7179 ;
  assign n7211 = n7210 ^ n7207 ;
  assign n7143 = n7139 ^ x169 ;
  assign n7144 = ~n7142 & ~n7143 ;
  assign n7212 = n7211 ^ n7144 ;
  assign n1216 = x170 ^ x169 ;
  assign n1220 = n7165 ^ n1216 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1225 = n1224 ^ n1223 ;
  assign n7134 = n1220 & n1225 ;
  assign n7976 = n7205 ^ n7134 ;
  assign n7977 = ~n7212 & n7976 ;
  assign n7978 = n7977 ^ n7205 ;
  assign n11837 = n7981 ^ n7978 ;
  assign n11838 = n7982 & n11837 ;
  assign n11839 = n11838 ^ n7202 ;
  assign n11843 = n11842 ^ n11839 ;
  assign n7983 = n7982 ^ n7978 ;
  assign n7975 = n7974 ^ n7973 ;
  assign n7984 = n7983 ^ n7975 ;
  assign n7213 = n7212 ^ n7134 ;
  assign n7133 = n7132 ^ n7089 ;
  assign n7214 = n7213 ^ n7133 ;
  assign n1235 = n1234 ^ n1233 ;
  assign n1236 = n1235 ^ n1232 ;
  assign n1227 = x158 ^ x157 ;
  assign n1231 = n7118 ^ n1227 ;
  assign n1237 = n1236 ^ n1231 ;
  assign n1226 = n1225 ^ n1220 ;
  assign n7033 = n1236 ^ n1226 ;
  assign n7034 = n1237 & n7033 ;
  assign n7035 = n7034 ^ n1236 ;
  assign n7951 = n7133 ^ n7035 ;
  assign n7952 = ~n7214 & n7951 ;
  assign n7953 = n7952 ^ n7133 ;
  assign n11834 = n7983 ^ n7953 ;
  assign n11835 = n7984 & n11834 ;
  assign n11836 = n11835 ^ n7983 ;
  assign n11844 = n11843 ^ n11836 ;
  assign n7394 = n7393 ^ n7308 ;
  assign n7215 = n7214 ^ n7035 ;
  assign n7395 = n7394 ^ n7215 ;
  assign n7985 = n7984 ^ n7953 ;
  assign n7986 = n7985 ^ n7394 ;
  assign n1215 = n1214 ^ n1203 ;
  assign n1238 = n1237 ^ n1226 ;
  assign n6706 = n1215 & n1238 ;
  assign n7987 = n7986 ^ n6706 ;
  assign n7988 = n7987 ^ n7985 ;
  assign n7989 = n7395 & ~n7988 ;
  assign n7990 = n7989 ^ n7986 ;
  assign n8014 = n8013 ^ n7998 ;
  assign n8039 = n8038 ^ n8014 ;
  assign n11845 = n8039 ^ n7985 ;
  assign n11846 = ~n7990 & n11845 ;
  assign n11847 = n11846 ^ n7985 ;
  assign n12587 = n11836 & ~n11842 ;
  assign n12617 = ~n11847 & ~n12587 ;
  assign n12618 = n11844 & n12617 ;
  assign n12619 = n12618 ^ n12590 ;
  assign n12620 = ~n12590 & ~n12619 ;
  assign n12621 = n11833 & n12620 ;
  assign n12622 = n12621 ^ n11833 ;
  assign n12600 = n11842 ^ n11836 ;
  assign n12612 = n12600 ^ n12587 ;
  assign n12591 = ~n11833 & ~n12590 ;
  assign n12592 = n12589 & n12591 ;
  assign n12593 = n12592 ^ n12590 ;
  assign n12588 = n11847 & n12587 ;
  assign n12594 = n11839 & n12593 ;
  assign n12602 = n11847 ^ n11836 ;
  assign n12603 = n12600 & n12602 ;
  assign n12601 = n12600 ^ n12588 ;
  assign n12604 = n12603 ^ n12601 ;
  assign n12607 = ~n11833 & ~n12604 ;
  assign n12608 = n12594 & n12607 ;
  assign n12609 = n12608 ^ n12594 ;
  assign n12610 = n12609 ^ n11839 ;
  assign n12611 = ~n12588 & n12610 ;
  assign n12613 = ~n12593 & n12611 ;
  assign n12614 = ~n12612 & n12613 ;
  assign n12615 = n12614 ^ n12611 ;
  assign n12629 = n12603 ^ n11847 ;
  assign n12630 = n12593 & ~n12629 ;
  assign n12836 = ~n12615 & ~n12630 ;
  assign n12837 = ~n12622 & n12836 ;
  assign n7434 = x237 & x238 ;
  assign n7433 = x239 & x240 ;
  assign n7441 = n7434 ^ n7433 ;
  assign n7435 = ~n7433 & ~n7434 ;
  assign n7442 = n7441 ^ n7435 ;
  assign n7443 = x235 & x236 ;
  assign n7444 = n7442 & n7443 ;
  assign n1340 = x240 ^ x239 ;
  assign n7436 = n7433 ^ n1340 ;
  assign n1343 = x238 ^ x237 ;
  assign n7437 = n7434 ^ n1343 ;
  assign n7438 = n7436 & n7437 ;
  assign n7445 = n7444 ^ n7438 ;
  assign n1341 = x236 ^ x235 ;
  assign n7446 = n7435 ^ n1341 ;
  assign n7447 = n7444 ^ n7435 ;
  assign n7448 = n7446 & ~n7447 ;
  assign n7449 = n7445 & n7448 ;
  assign n7450 = n7449 ^ n7444 ;
  assign n7451 = n7442 & ~n7450 ;
  assign n7405 = x243 & x244 ;
  assign n7404 = x245 & x246 ;
  assign n7413 = n7405 ^ n7404 ;
  assign n7406 = ~n7404 & ~n7405 ;
  assign n7414 = n7413 ^ n7406 ;
  assign n7415 = x241 & x242 ;
  assign n7416 = n7414 & n7415 ;
  assign n1338 = x244 ^ x243 ;
  assign n7408 = n7405 ^ n1338 ;
  assign n1336 = x246 ^ x245 ;
  assign n7407 = n7404 ^ n1336 ;
  assign n7410 = n7408 ^ n7407 ;
  assign n7409 = ~n7407 & ~n7408 ;
  assign n7411 = n7410 ^ n7409 ;
  assign n7420 = n7416 ^ n7411 ;
  assign n7421 = n7416 ^ n7406 ;
  assign n7412 = n7411 ^ n7406 ;
  assign n1335 = x242 ^ x241 ;
  assign n7417 = n7416 ^ n1335 ;
  assign n7418 = ~n7412 & ~n7417 ;
  assign n7422 = n7421 ^ n7418 ;
  assign n7423 = ~n7420 & n7422 ;
  assign n7424 = n7423 ^ n7411 ;
  assign n8297 = n7414 & n7424 ;
  assign n11871 = ~n7451 & ~n8297 ;
  assign n7419 = n7406 & n7418 ;
  assign n7425 = n7409 ^ x241 ;
  assign n7426 = n7425 ^ n7424 ;
  assign n7427 = n7414 ^ x242 ;
  assign n7428 = ~n7409 & ~n7427 ;
  assign n7429 = n7428 ^ x242 ;
  assign n7430 = n7426 & n7429 ;
  assign n7431 = n7430 ^ n7409 ;
  assign n7432 = n7424 & ~n7431 ;
  assign n7461 = n7419 & n7432 ;
  assign n7455 = n7436 ^ x236 ;
  assign n7456 = n7455 ^ n7437 ;
  assign n7457 = n1341 & n7456 ;
  assign n7452 = n7450 ^ x235 ;
  assign n7453 = n7452 ^ n7451 ;
  assign n7439 = n7438 ^ n1341 ;
  assign n7440 = n7435 & ~n7439 ;
  assign n7454 = n7453 ^ n7440 ;
  assign n7458 = n7457 ^ n7454 ;
  assign n7459 = n7458 ^ n7432 ;
  assign n7462 = n7461 ^ n7459 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1339 = n1338 ^ n1337 ;
  assign n1342 = n1341 ^ n1340 ;
  assign n1344 = n1343 ^ n1342 ;
  assign n7403 = n1339 & n1344 ;
  assign n8294 = n7458 ^ n7403 ;
  assign n8295 = n7462 & n8294 ;
  assign n8296 = n8295 ^ n7458 ;
  assign n7486 = x227 & x228 ;
  assign n7485 = x225 & x226 ;
  assign n7487 = n7486 ^ n7485 ;
  assign n1351 = x226 ^ x225 ;
  assign n7488 = n7485 ^ n1351 ;
  assign n1353 = x228 ^ x227 ;
  assign n7489 = n7486 ^ n1353 ;
  assign n7490 = n7488 & n7489 ;
  assign n7491 = n7490 ^ n7485 ;
  assign n7492 = ~n7487 & ~n7491 ;
  assign n7464 = n1353 ^ x224 ;
  assign n7465 = n7464 ^ n1351 ;
  assign n1347 = x230 ^ x229 ;
  assign n1348 = x234 ^ x233 ;
  assign n7474 = n1348 ^ x230 ;
  assign n1346 = x232 ^ x231 ;
  assign n7475 = n7474 ^ n1346 ;
  assign n7476 = n1347 & ~n7475 ;
  assign n7477 = n7476 ^ x229 ;
  assign n7467 = x233 & x234 ;
  assign n7466 = x231 & x232 ;
  assign n7468 = n7467 ^ n7466 ;
  assign n7469 = n7466 ^ n1346 ;
  assign n7470 = n7467 ^ n1348 ;
  assign n7471 = n7469 & n7470 ;
  assign n7472 = n7471 ^ n7466 ;
  assign n7473 = ~n7468 & ~n7472 ;
  assign n7478 = n7477 ^ n7473 ;
  assign n7479 = n7478 ^ x223 ;
  assign n7480 = n7479 ^ n1353 ;
  assign n7481 = n7480 ^ n1351 ;
  assign n7482 = n7481 ^ n7478 ;
  assign n7483 = ~n7465 & n7482 ;
  assign n7484 = n7483 ^ n7479 ;
  assign n7493 = n7492 ^ n7484 ;
  assign n1349 = n1348 ^ n1347 ;
  assign n1350 = n1349 ^ n1346 ;
  assign n1352 = x224 ^ x223 ;
  assign n1354 = n1353 ^ n1352 ;
  assign n1355 = n1354 ^ n1351 ;
  assign n7494 = n1350 & n1355 ;
  assign n8324 = n7494 ^ n7478 ;
  assign n8325 = ~n7493 & ~n8324 ;
  assign n8326 = n8325 ^ n7494 ;
  assign n8300 = n7490 ^ x224 ;
  assign n8301 = n7487 ^ x223 ;
  assign n8302 = n8301 ^ n7490 ;
  assign n8303 = n8300 & ~n8302 ;
  assign n8304 = n8303 ^ n7491 ;
  assign n8305 = ~n7487 & n8304 ;
  assign n8306 = x223 & n8305 ;
  assign n8307 = n8303 ^ n7490 ;
  assign n8308 = n8307 ^ n8305 ;
  assign n8322 = n8306 & ~n8308 ;
  assign n8309 = n7471 ^ x230 ;
  assign n8310 = n7468 ^ x229 ;
  assign n8311 = n8310 ^ n7471 ;
  assign n8312 = n8309 & ~n8311 ;
  assign n8315 = n8312 ^ n7471 ;
  assign n8313 = n8312 ^ n7472 ;
  assign n8314 = ~n7468 & n8313 ;
  assign n8316 = n8315 ^ n8314 ;
  assign n8317 = x229 & n8314 ;
  assign n8318 = ~n8316 & n8317 ;
  assign n8319 = n8318 ^ n8316 ;
  assign n8320 = n8319 ^ n8308 ;
  assign n8323 = n8322 ^ n8320 ;
  assign n8327 = n8326 ^ n8323 ;
  assign n7495 = n7494 ^ n7493 ;
  assign n7463 = n7462 ^ n7403 ;
  assign n7496 = n7495 ^ n7463 ;
  assign n1345 = n1344 ^ n1339 ;
  assign n1356 = n1355 ^ n1350 ;
  assign n7401 = n1345 & n1356 ;
  assign n8329 = n7463 ^ n7401 ;
  assign n8330 = ~n7496 & n8329 ;
  assign n8331 = n8330 ^ n7401 ;
  assign n8298 = n8297 ^ n7451 ;
  assign n8299 = n8298 ^ n8296 ;
  assign n8328 = n8327 ^ n8299 ;
  assign n8332 = n8331 ^ n8328 ;
  assign n11873 = ~n8327 & ~n8332 ;
  assign n11874 = ~n8296 & n11873 ;
  assign n11875 = n11874 ^ n8332 ;
  assign n11876 = ~n11871 & n11875 ;
  assign n11872 = n11871 ^ n8298 ;
  assign n11877 = n11876 ^ n11872 ;
  assign n11878 = n11876 ^ n8327 ;
  assign n11879 = ~n11877 & n11878 ;
  assign n11880 = n11879 ^ n8327 ;
  assign n11886 = n11880 ^ n11876 ;
  assign n11883 = n8326 ^ n8319 ;
  assign n11884 = n8323 & n11883 ;
  assign n11885 = n11884 ^ n8319 ;
  assign n11887 = n11886 ^ n11885 ;
  assign n11881 = ~n8331 & n11880 ;
  assign n11882 = ~n8296 & n11881 ;
  assign n11888 = n11887 ^ n11882 ;
  assign n12548 = ~n11871 & ~n11888 ;
  assign n12549 = n11875 & ~n11885 ;
  assign n12550 = ~n12548 & n12549 ;
  assign n12551 = n12550 ^ n12548 ;
  assign n7582 = x249 & x250 ;
  assign n7580 = x251 & x252 ;
  assign n7585 = n7582 ^ n7580 ;
  assign n1361 = x252 ^ x251 ;
  assign n7581 = n7580 ^ n1361 ;
  assign n1359 = x250 ^ x249 ;
  assign n7583 = n7582 ^ n1359 ;
  assign n7584 = n7581 & n7583 ;
  assign n8227 = n7584 ^ n7582 ;
  assign n7596 = n7584 ^ x248 ;
  assign n8209 = n7580 ^ x247 ;
  assign n8210 = n8209 ^ n7585 ;
  assign n8208 = n7580 ^ x248 ;
  assign n8211 = n8210 ^ n8208 ;
  assign n8225 = n7596 & n8211 ;
  assign n8228 = n8227 ^ n8225 ;
  assign n8229 = ~n7585 & n8228 ;
  assign n8231 = n7584 & n8209 ;
  assign n8232 = n8229 & n8231 ;
  assign n8226 = n8225 ^ n7596 ;
  assign n8230 = n8229 ^ n8226 ;
  assign n8233 = n8232 ^ n8230 ;
  assign n8238 = n8233 ^ n7580 ;
  assign n8239 = n8238 ^ n8208 ;
  assign n7602 = x257 & x258 ;
  assign n7601 = x255 & x256 ;
  assign n7603 = n7602 ^ n7601 ;
  assign n1363 = x254 ^ x253 ;
  assign n8201 = n7602 ^ x254 ;
  assign n1366 = x258 ^ x257 ;
  assign n7604 = n7602 ^ n1366 ;
  assign n1364 = x256 ^ x255 ;
  assign n7605 = n7601 ^ n1364 ;
  assign n7606 = n7604 & n7605 ;
  assign n7607 = n7606 ^ n7602 ;
  assign n8180 = n7607 ^ n7603 ;
  assign n8186 = n8201 ^ n8180 ;
  assign n8190 = n1363 & n8186 ;
  assign n8184 = n7602 & ~n7606 ;
  assign n8191 = n8190 ^ n8184 ;
  assign n8177 = n7602 ^ x253 ;
  assign n8178 = n8177 ^ n7607 ;
  assign n8182 = n8178 ^ n7603 ;
  assign n8192 = n8191 ^ n8182 ;
  assign n8193 = n8190 ^ n8180 ;
  assign n8194 = n8193 ^ n8182 ;
  assign n8195 = n8192 & n8194 ;
  assign n8196 = ~n7603 & n8195 ;
  assign n8197 = n8196 ^ n8190 ;
  assign n8198 = n8197 ^ n1363 ;
  assign n8204 = n8198 ^ n7602 ;
  assign n8205 = n8204 ^ n8201 ;
  assign n8240 = n8239 ^ n8205 ;
  assign n1371 = x266 ^ x265 ;
  assign n1370 = x268 ^ x267 ;
  assign n1372 = n1371 ^ n1370 ;
  assign n1369 = x270 ^ x269 ;
  assign n1373 = n1372 ^ n1369 ;
  assign n1376 = x262 ^ x261 ;
  assign n1375 = x260 ^ x259 ;
  assign n1377 = n1376 ^ n1375 ;
  assign n1374 = x264 ^ x263 ;
  assign n1378 = n1377 ^ n1374 ;
  assign n8158 = n1373 & n1378 ;
  assign n7541 = x269 ^ x268 ;
  assign n7545 = ~n1369 & ~n7541 ;
  assign n7540 = x267 ^ x266 ;
  assign n7542 = n7541 ^ x267 ;
  assign n7543 = n7542 ^ x270 ;
  assign n7544 = ~n7540 & n7543 ;
  assign n7546 = n7545 ^ n7544 ;
  assign n7547 = ~x265 & n7546 ;
  assign n7548 = ~n1370 & ~n7540 ;
  assign n7549 = x270 ^ x265 ;
  assign n7552 = ~x268 & ~n7549 ;
  assign n7553 = n7552 ^ x265 ;
  assign n7554 = n7548 & n7553 ;
  assign n7555 = ~x269 & n7554 ;
  assign n7556 = ~x267 & ~x268 ;
  assign n7559 = n7556 ^ n1370 ;
  assign n7560 = x265 & x266 ;
  assign n7561 = x270 & n7560 ;
  assign n7562 = ~n7559 & n7561 ;
  assign n7563 = n7562 ^ n7560 ;
  assign n7557 = ~x269 & ~x270 ;
  assign n7558 = ~n7556 & ~n7557 ;
  assign n7564 = n7563 ^ n7558 ;
  assign n7565 = n7557 ^ n1369 ;
  assign n7570 = n7559 & n7565 ;
  assign n7571 = n7570 ^ n7558 ;
  assign n7572 = n7564 & n7571 ;
  assign n7573 = n7572 ^ n7563 ;
  assign n7574 = ~n1371 & n7573 ;
  assign n7575 = n7572 & n7574 ;
  assign n7576 = n7575 ^ n7573 ;
  assign n7577 = ~n7555 & ~n7576 ;
  assign n7578 = ~n7547 & n7577 ;
  assign n7499 = ~x263 & ~x264 ;
  assign n7502 = n7499 ^ n1374 ;
  assign n7498 = x261 & x262 ;
  assign n7504 = x259 & x260 ;
  assign n7505 = n7498 & ~n7504 ;
  assign n7506 = n7502 & n7505 ;
  assign n7507 = n7506 ^ n7498 ;
  assign n7503 = n7498 & ~n7502 ;
  assign n7508 = n7507 ^ n7503 ;
  assign n7497 = ~x260 & n1377 ;
  assign n7500 = ~n7498 & n7499 ;
  assign n7501 = n7497 & n7500 ;
  assign n7509 = n7508 ^ n7501 ;
  assign n7510 = n7498 ^ n1376 ;
  assign n7511 = n7502 & ~n7510 ;
  assign n7519 = x260 & n7511 ;
  assign n7520 = ~n7499 & n7519 ;
  assign n7521 = n7520 ^ n7499 ;
  assign n7512 = n7511 ^ n7503 ;
  assign n7513 = n7512 ^ n7499 ;
  assign n7522 = n7521 ^ n7513 ;
  assign n7523 = ~x259 & n7522 ;
  assign n7524 = ~n7509 & ~n7523 ;
  assign n7525 = n7504 ^ n1375 ;
  assign n7526 = n7525 ^ x262 ;
  assign n7527 = n7525 ^ x261 ;
  assign n7528 = ~n7526 & ~n7527 ;
  assign n7529 = n7528 ^ n7525 ;
  assign n7530 = n7504 ^ n7502 ;
  assign n7531 = n7526 ^ n7502 ;
  assign n7532 = n7531 ^ n7527 ;
  assign n7533 = ~n7530 & n7532 ;
  assign n7534 = n7533 ^ n7525 ;
  assign n7535 = n7529 & n7534 ;
  assign n7536 = n7535 ^ n7525 ;
  assign n7537 = n7536 ^ n7504 ;
  assign n7538 = ~n7499 & n7537 ;
  assign n7539 = n7524 & ~n7538 ;
  assign n7579 = n7578 ^ n7539 ;
  assign n8248 = n8158 ^ n7579 ;
  assign n1379 = n1378 ^ n1373 ;
  assign n1365 = n1364 ^ n1363 ;
  assign n1367 = n1366 ^ n1365 ;
  assign n1358 = x248 ^ x247 ;
  assign n1360 = n1359 ^ n1358 ;
  assign n1362 = n1361 ^ n1360 ;
  assign n1368 = n1367 ^ n1362 ;
  assign n7628 = n1373 ^ n1368 ;
  assign n7629 = n1379 & ~n7628 ;
  assign n7630 = n7629 ^ n1378 ;
  assign n8288 = n8248 ^ n7630 ;
  assign n7631 = n1362 & n1367 ;
  assign n7590 = n7584 ^ n7580 ;
  assign n7591 = n7590 ^ n1358 ;
  assign n7592 = ~n7585 & ~n7591 ;
  assign n7586 = n1361 ^ n1359 ;
  assign n7587 = n7586 ^ n7585 ;
  assign n7588 = n7587 ^ x248 ;
  assign n7589 = n7588 ^ n7584 ;
  assign n7593 = n7592 ^ n7589 ;
  assign n7594 = n7593 ^ n7588 ;
  assign n7597 = n7596 ^ n7588 ;
  assign n7598 = n7594 & ~n7597 ;
  assign n7599 = n7598 ^ n7588 ;
  assign n7626 = n1358 & n7599 ;
  assign n7623 = n7592 ^ x247 ;
  assign n7615 = n7606 ^ x254 ;
  assign n7608 = n7607 ^ n1363 ;
  assign n7609 = ~n7603 & ~n7608 ;
  assign n7610 = n7609 ^ n7606 ;
  assign n7611 = n1366 ^ n1364 ;
  assign n7612 = n7611 ^ n7603 ;
  assign n7613 = n7612 ^ n7609 ;
  assign n7614 = ~n7610 & ~n7613 ;
  assign n7616 = n7615 ^ n7614 ;
  assign n7620 = n1363 & ~n7616 ;
  assign n7618 = n7609 ^ x253 ;
  assign n7621 = n7620 ^ n7618 ;
  assign n7624 = n7623 ^ n7621 ;
  assign n7627 = n7626 ^ n7624 ;
  assign n8244 = n7631 ^ n7627 ;
  assign n8245 = n8244 ^ n7579 ;
  assign n8246 = n8245 ^ n7630 ;
  assign n8287 = n8245 ^ n8158 ;
  assign n8289 = n8288 ^ n8287 ;
  assign n8265 = n8288 & n8289 ;
  assign n8247 = n8246 ^ n8158 ;
  assign n8253 = n8247 ^ n8245 ;
  assign n8254 = n8253 ^ n7631 ;
  assign n8256 = n8158 ^ n7631 ;
  assign n8258 = n8287 ^ n8256 ;
  assign n8259 = ~n8254 & n8258 ;
  assign n8266 = n8265 ^ n8259 ;
  assign n8267 = n8287 ^ n8266 ;
  assign n8268 = n8265 ^ n8158 ;
  assign n8269 = n8287 ^ n8268 ;
  assign n8270 = n8267 & ~n8269 ;
  assign n8271 = n8246 & n8270 ;
  assign n8272 = n8271 ^ n8265 ;
  assign n8284 = n8288 ^ n8272 ;
  assign n8291 = n8284 ^ n7579 ;
  assign n8292 = n8291 ^ n8158 ;
  assign n8171 = n7631 ^ n7621 ;
  assign n8172 = ~n7627 & ~n8171 ;
  assign n8173 = n8172 ^ n7631 ;
  assign n8241 = n8240 ^ n8173 ;
  assign n11857 = n8292 ^ n8241 ;
  assign n8159 = n8158 ^ n7539 ;
  assign n8160 = n7579 & ~n8159 ;
  assign n8161 = n8160 ^ n7578 ;
  assign n11858 = n8241 ^ n8161 ;
  assign n11859 = n11857 & ~n11858 ;
  assign n11860 = n11859 ^ n8292 ;
  assign n11861 = n11860 ^ n8239 ;
  assign n11862 = n11861 ^ n8173 ;
  assign n11863 = n11862 ^ n11860 ;
  assign n11864 = n8240 & n11863 ;
  assign n11865 = n11864 ^ n11861 ;
  assign n8168 = ~n7507 & ~n7538 ;
  assign n8162 = n7565 ^ n7559 ;
  assign n8163 = x266 & n7558 ;
  assign n8164 = n8163 ^ n7559 ;
  assign n8165 = n8162 & ~n8164 ;
  assign n8166 = n8165 ^ n7559 ;
  assign n8167 = ~n7576 & n8166 ;
  assign n8169 = n8168 ^ n8167 ;
  assign n8170 = n8169 ^ n8161 ;
  assign n8242 = n8241 ^ n8170 ;
  assign n8293 = n8292 ^ n8242 ;
  assign n11866 = n8293 ^ n8168 ;
  assign n11867 = n8169 & n11866 ;
  assign n11868 = n11867 ^ n8168 ;
  assign n12545 = n11868 ^ n11860 ;
  assign n12546 = ~n11865 & ~n12545 ;
  assign n12547 = n12546 ^ n11868 ;
  assign n12552 = n12551 ^ n12547 ;
  assign n11869 = n11868 ^ n11865 ;
  assign n8333 = n8332 ^ n8293 ;
  assign n7635 = n8246 ^ n7496 ;
  assign n1357 = n1356 ^ n1345 ;
  assign n1380 = n1379 ^ n1368 ;
  assign n7400 = n1357 & n1380 ;
  assign n8153 = n7496 ^ n7400 ;
  assign n8156 = n7635 & ~n8153 ;
  assign n8155 = ~n7401 & n8246 ;
  assign n8157 = n8156 ^ n8155 ;
  assign n11854 = n8293 ^ n8157 ;
  assign n11855 = n8333 & ~n11854 ;
  assign n11856 = n11855 ^ n8332 ;
  assign n11870 = n11869 ^ n11856 ;
  assign n12542 = n11888 ^ n11856 ;
  assign n12543 = n11870 & ~n12542 ;
  assign n12544 = n12543 ^ n11888 ;
  assign n12553 = n12552 ^ n12544 ;
  assign n7711 = ~x189 & ~x190 ;
  assign n1324 = x190 ^ x189 ;
  assign n7720 = n7711 ^ n1324 ;
  assign n7709 = ~x191 & ~x192 ;
  assign n1323 = x192 ^ x191 ;
  assign n7719 = n7709 ^ n1323 ;
  assign n7721 = n7720 ^ n7719 ;
  assign n7710 = n7709 ^ x188 ;
  assign n7712 = n7711 ^ n7710 ;
  assign n7722 = n7719 ^ n7712 ;
  assign n7714 = n7711 ^ n7709 ;
  assign n7713 = n7709 & n7711 ;
  assign n7715 = n7714 ^ n7713 ;
  assign n7716 = n7712 & n7715 ;
  assign n7723 = n7722 ^ n7716 ;
  assign n7724 = n7721 & n7723 ;
  assign n7725 = n7724 ^ n7720 ;
  assign n7728 = x191 ^ x188 ;
  assign n7729 = n7728 ^ x190 ;
  assign n7730 = n7729 ^ x192 ;
  assign n7726 = x191 ^ x189 ;
  assign n7731 = n7730 ^ n7726 ;
  assign n7732 = n7731 ^ x192 ;
  assign n7733 = n7732 ^ x191 ;
  assign n7734 = n7733 ^ n7726 ;
  assign n7738 = n7726 ^ x190 ;
  assign n7739 = n7738 ^ x192 ;
  assign n7740 = n7739 ^ n7726 ;
  assign n7741 = ~n7734 & ~n7740 ;
  assign n7742 = ~x191 & n7741 ;
  assign n7745 = n7742 ^ n7741 ;
  assign n7743 = n7742 ^ n7726 ;
  assign n7744 = n7731 & n7743 ;
  assign n7746 = n7745 ^ n7744 ;
  assign n7747 = n7746 ^ x191 ;
  assign n8456 = n7747 ^ x187 ;
  assign n7783 = ~x187 & ~n7747 ;
  assign n8457 = n8456 ^ n7783 ;
  assign n8458 = n7725 & n8457 ;
  assign n7754 = x195 & x196 ;
  assign n7756 = x197 & x198 ;
  assign n7762 = n7754 & n7756 ;
  assign n7761 = n7756 ^ n7754 ;
  assign n7763 = n7762 ^ n7761 ;
  assign n1327 = x198 ^ x197 ;
  assign n7757 = n7756 ^ n1327 ;
  assign n1330 = x196 ^ x195 ;
  assign n7755 = n7754 ^ n1330 ;
  assign n7759 = n7757 ^ n7755 ;
  assign n7758 = ~n7755 & ~n7757 ;
  assign n7760 = n7759 ^ n7758 ;
  assign n7764 = n7763 ^ n7760 ;
  assign n1328 = x194 ^ x193 ;
  assign n7769 = n7763 ^ n1328 ;
  assign n7770 = n7764 & ~n7769 ;
  assign n7771 = x193 & x194 ;
  assign n7772 = ~n7762 & n7771 ;
  assign n7773 = n7772 ^ n7763 ;
  assign n7774 = n7770 & n7773 ;
  assign n7775 = n7774 ^ n7772 ;
  assign n7776 = ~n7762 & ~n7775 ;
  assign n8459 = n8458 ^ n7776 ;
  assign n7782 = n7719 & n7720 ;
  assign n7784 = n7782 & n7783 ;
  assign n7777 = n7776 ^ n7775 ;
  assign n7765 = n7755 ^ n1328 ;
  assign n7766 = n7765 ^ n7757 ;
  assign n7767 = ~n7758 & ~n7766 ;
  assign n7768 = n7764 & ~n7767 ;
  assign n7778 = n7777 ^ n7768 ;
  assign n7779 = n7778 ^ n7771 ;
  assign n7780 = n7779 ^ n7747 ;
  assign n7751 = ~x187 & ~n7746 ;
  assign n7752 = n7751 ^ x191 ;
  assign n7753 = ~n7725 & ~n7752 ;
  assign n7781 = n7780 ^ n7753 ;
  assign n7785 = n7784 ^ n7781 ;
  assign n7717 = n7713 ^ x187 ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7786 = n7785 ^ n7718 ;
  assign n1322 = x188 ^ x187 ;
  assign n1326 = n7739 ^ n1322 ;
  assign n1329 = n1328 ^ n1327 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n7708 = n1326 & n1331 ;
  assign n8453 = n7779 ^ n7708 ;
  assign n8454 = ~n7786 & n8453 ;
  assign n8455 = n8454 ^ n7779 ;
  assign n11921 = n8458 ^ n8455 ;
  assign n11922 = n8459 & n11921 ;
  assign n11923 = n11922 ^ n7776 ;
  assign n8460 = n8459 ^ n8455 ;
  assign n7641 = x179 & x180 ;
  assign n7640 = x177 & x178 ;
  assign n7642 = n7641 ^ n7640 ;
  assign n1314 = x180 ^ x179 ;
  assign n7645 = n7641 ^ n1314 ;
  assign n1312 = x178 ^ x177 ;
  assign n7646 = n7640 ^ n1312 ;
  assign n7647 = n7645 & n7646 ;
  assign n7648 = n7647 ^ x176 ;
  assign n8441 = n7647 ^ x175 ;
  assign n8442 = n8441 ^ n7642 ;
  assign n8443 = n7648 & n8442 ;
  assign n8444 = n8443 ^ x176 ;
  assign n8445 = n8444 ^ n7640 ;
  assign n8446 = n7642 & ~n8445 ;
  assign n8447 = n8446 ^ n7641 ;
  assign n8448 = x175 & n8444 ;
  assign n8449 = ~n8447 & n8448 ;
  assign n8450 = n8449 ^ n8447 ;
  assign n11913 = n8460 ^ n8450 ;
  assign n1311 = x176 ^ x175 ;
  assign n7650 = n7647 ^ n7641 ;
  assign n7651 = n7650 ^ n1311 ;
  assign n7652 = ~n7642 & ~n7651 ;
  assign n7643 = n1314 ^ n1312 ;
  assign n7644 = n7643 ^ n7642 ;
  assign n7649 = n7648 ^ n7644 ;
  assign n7653 = n7652 ^ n7649 ;
  assign n7654 = n7653 ^ n7648 ;
  assign n7656 = n7644 ^ x176 ;
  assign n7657 = n7656 ^ n7648 ;
  assign n7658 = ~n7654 & ~n7657 ;
  assign n7659 = n7658 ^ n7648 ;
  assign n7704 = n1311 & ~n7659 ;
  assign n7701 = n7652 ^ x175 ;
  assign n1319 = x186 ^ x185 ;
  assign n7662 = x185 ^ x184 ;
  assign n7666 = ~n1319 & ~n7662 ;
  assign n7661 = x183 ^ x182 ;
  assign n7663 = n7662 ^ x183 ;
  assign n7664 = n7663 ^ x186 ;
  assign n7665 = ~n7661 & n7664 ;
  assign n7667 = n7666 ^ n7665 ;
  assign n7668 = ~x181 & n7667 ;
  assign n1317 = x184 ^ x183 ;
  assign n7669 = ~n1317 & ~n7661 ;
  assign n7670 = x186 ^ x181 ;
  assign n7673 = ~x184 & ~n7670 ;
  assign n7674 = n7673 ^ x181 ;
  assign n7675 = n7669 & n7674 ;
  assign n7676 = ~x185 & n7675 ;
  assign n7677 = ~x183 & ~x184 ;
  assign n7680 = n7677 ^ n1317 ;
  assign n7681 = x181 & x182 ;
  assign n7682 = x186 & n7681 ;
  assign n7683 = ~n7680 & n7682 ;
  assign n7684 = n7683 ^ n7681 ;
  assign n7678 = ~x185 & ~x186 ;
  assign n7679 = ~n7677 & ~n7678 ;
  assign n7685 = n7684 ^ n7679 ;
  assign n7686 = n7678 ^ n1319 ;
  assign n7691 = n7680 & n7686 ;
  assign n7692 = n7691 ^ n7679 ;
  assign n7693 = n7685 & n7692 ;
  assign n1316 = x182 ^ x181 ;
  assign n7694 = n7693 ^ n7684 ;
  assign n7695 = ~n1316 & n7694 ;
  assign n7696 = n7693 & n7695 ;
  assign n7697 = n7696 ^ n7694 ;
  assign n7698 = ~n7676 & ~n7697 ;
  assign n7699 = ~n7668 & n7698 ;
  assign n7702 = n7701 ^ n7699 ;
  assign n7705 = n7704 ^ n7702 ;
  assign n1313 = n1312 ^ n1311 ;
  assign n1315 = n1314 ^ n1313 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1320 = n1319 ^ n1318 ;
  assign n7706 = n1315 & n1320 ;
  assign n8431 = n7706 ^ n7699 ;
  assign n8432 = ~n7705 & n8431 ;
  assign n8433 = n8432 ^ n7699 ;
  assign n11914 = n8450 ^ n8433 ;
  assign n11915 = n11913 & ~n11914 ;
  assign n11916 = n11915 ^ n8460 ;
  assign n7787 = n7786 ^ n7708 ;
  assign n7707 = n7706 ^ n7705 ;
  assign n7788 = n7787 ^ n7707 ;
  assign n1321 = n1320 ^ n1315 ;
  assign n1332 = n1331 ^ n1326 ;
  assign n8335 = n1321 & n1332 ;
  assign n8462 = n8335 ^ n7787 ;
  assign n8463 = n7788 & ~n8462 ;
  assign n8464 = n8463 ^ n7787 ;
  assign n8434 = n7686 ^ n7680 ;
  assign n8435 = x182 & n7679 ;
  assign n8436 = n8435 ^ n7680 ;
  assign n8437 = n8434 & ~n8436 ;
  assign n8438 = n8437 ^ n7680 ;
  assign n8439 = ~n7697 & ~n8438 ;
  assign n8440 = n8439 ^ n7697 ;
  assign n11909 = n8464 ^ n8440 ;
  assign n8451 = n8450 ^ n8440 ;
  assign n8452 = n8451 ^ n8433 ;
  assign n8461 = n8460 ^ n8452 ;
  assign n8465 = n8464 ^ n8461 ;
  assign n11910 = n8465 ^ n8440 ;
  assign n11911 = ~n11909 & ~n11910 ;
  assign n11912 = n11911 ^ n8464 ;
  assign n11917 = n11916 ^ n11912 ;
  assign n11924 = n11923 ^ n11917 ;
  assign n7790 = x213 & x214 ;
  assign n1299 = x214 ^ x213 ;
  assign n7793 = n7790 ^ n1299 ;
  assign n7791 = x215 & x216 ;
  assign n1301 = x216 ^ x215 ;
  assign n7794 = n7791 ^ n1301 ;
  assign n7795 = n7793 & n7794 ;
  assign n8398 = n7795 ^ x212 ;
  assign n7792 = n7791 ^ n7790 ;
  assign n8399 = n7792 ^ x211 ;
  assign n8400 = n8399 ^ n7795 ;
  assign n8401 = n8398 & ~n8400 ;
  assign n8404 = n8401 ^ n7795 ;
  assign n7796 = n7795 ^ n7790 ;
  assign n8402 = n8401 ^ n7796 ;
  assign n8403 = ~n7792 & n8402 ;
  assign n8405 = n8404 ^ n8403 ;
  assign n8406 = x211 & n8403 ;
  assign n8407 = ~n8405 & n8406 ;
  assign n8408 = n8407 ^ n8405 ;
  assign n7819 = ~x219 & ~x220 ;
  assign n1304 = x220 ^ x219 ;
  assign n7822 = n7819 ^ n1304 ;
  assign n7823 = x217 & x218 ;
  assign n7824 = x222 & n7823 ;
  assign n7825 = ~n7822 & n7824 ;
  assign n7826 = n7825 ^ n7823 ;
  assign n7820 = ~x221 & ~x222 ;
  assign n7821 = ~n7819 & ~n7820 ;
  assign n7827 = n7826 ^ n7821 ;
  assign n1305 = x222 ^ x221 ;
  assign n7828 = n7820 ^ n1305 ;
  assign n7833 = n7822 & n7828 ;
  assign n7834 = n7833 ^ n7821 ;
  assign n7835 = n7827 & n7834 ;
  assign n1306 = x218 ^ x217 ;
  assign n7836 = n7835 ^ n7826 ;
  assign n7837 = ~n1306 & n7836 ;
  assign n7838 = n7835 & n7837 ;
  assign n7839 = n7838 ^ n7836 ;
  assign n8392 = n7828 ^ n7822 ;
  assign n8393 = x218 & n7821 ;
  assign n8394 = n8393 ^ n7822 ;
  assign n8395 = n8392 & ~n8394 ;
  assign n8396 = n8395 ^ n7822 ;
  assign n8397 = ~n7839 & n8396 ;
  assign n8409 = n8408 ^ n8397 ;
  assign n7804 = x221 ^ x220 ;
  assign n7808 = ~n1305 & ~n7804 ;
  assign n7803 = x219 ^ x218 ;
  assign n7805 = n7804 ^ x219 ;
  assign n7806 = n7805 ^ x222 ;
  assign n7807 = ~n7803 & n7806 ;
  assign n7809 = n7808 ^ n7807 ;
  assign n7810 = ~x217 & n7809 ;
  assign n7811 = ~n1304 & ~n7803 ;
  assign n7812 = x222 ^ x217 ;
  assign n7815 = ~x220 & ~n7812 ;
  assign n7816 = n7815 ^ x217 ;
  assign n7817 = n7811 & n7816 ;
  assign n7818 = ~x221 & n7817 ;
  assign n7840 = ~n7818 & ~n7839 ;
  assign n7841 = ~n7810 & n7840 ;
  assign n1300 = x212 ^ x211 ;
  assign n7798 = n1301 ^ x212 ;
  assign n7799 = n7798 ^ n1299 ;
  assign n7800 = n1300 & ~n7799 ;
  assign n7801 = n7800 ^ x211 ;
  assign n7797 = ~n7792 & ~n7796 ;
  assign n7802 = n7801 ^ n7797 ;
  assign n7842 = n7841 ^ n7802 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1303 = n1302 ^ n1299 ;
  assign n1307 = n1306 ^ n1305 ;
  assign n1308 = n1307 ^ n1304 ;
  assign n7931 = n1303 & n1308 ;
  assign n8389 = n7931 ^ n7802 ;
  assign n8390 = n7842 & ~n8389 ;
  assign n8391 = n8390 ^ n7931 ;
  assign n11905 = n8408 ^ n8391 ;
  assign n11906 = ~n8409 & n11905 ;
  assign n11907 = n11906 ^ n8408 ;
  assign n7868 = x203 ^ x200 ;
  assign n7869 = n7868 ^ x202 ;
  assign n7870 = n7869 ^ x204 ;
  assign n7866 = x203 ^ x201 ;
  assign n7871 = n7870 ^ n7866 ;
  assign n7843 = x204 ^ x202 ;
  assign n7844 = x204 ^ x200 ;
  assign n7845 = n7844 ^ n7843 ;
  assign n7877 = ~n7843 & ~n7845 ;
  assign n7881 = n7877 ^ x201 ;
  assign n7882 = n7881 ^ n7866 ;
  assign n7883 = n7877 & n7882 ;
  assign n7884 = n7883 ^ n7866 ;
  assign n7885 = ~n7871 & n7884 ;
  assign n7886 = n7885 ^ n7881 ;
  assign n8423 = x199 & n7886 ;
  assign n7887 = ~x203 & ~x204 ;
  assign n1290 = x204 ^ x203 ;
  assign n7889 = n7887 ^ n1290 ;
  assign n7888 = x200 & ~n7887 ;
  assign n7893 = n7889 ^ n7888 ;
  assign n8414 = n7888 ^ x202 ;
  assign n8415 = n8414 ^ x201 ;
  assign n8416 = n7893 & ~n8415 ;
  assign n1289 = x202 ^ x201 ;
  assign n8417 = n8416 ^ n1289 ;
  assign n8420 = ~x202 & ~n8416 ;
  assign n8421 = ~n8417 & n8420 ;
  assign n1294 = x206 ^ x205 ;
  assign n7902 = x209 & x210 ;
  assign n1293 = x210 ^ x209 ;
  assign n7903 = n7902 ^ n1293 ;
  assign n7904 = n1294 & n7903 ;
  assign n1295 = x208 ^ x207 ;
  assign n7905 = n1295 ^ x205 ;
  assign n7910 = x207 & x208 ;
  assign n7911 = ~n7903 & ~n7910 ;
  assign n7914 = ~x206 & n7911 ;
  assign n7906 = n7902 ^ x208 ;
  assign n7907 = ~x205 & ~n7906 ;
  assign n7915 = n7914 ^ n7907 ;
  assign n7916 = n7905 & n7915 ;
  assign n7917 = n7916 ^ n7907 ;
  assign n7918 = ~n7904 & n7917 ;
  assign n7920 = ~n1295 & ~n7906 ;
  assign n7924 = n7920 ^ n7906 ;
  assign n7925 = n7924 ^ x207 ;
  assign n7926 = n7904 & ~n7925 ;
  assign n7919 = x205 & x206 ;
  assign n7921 = ~n7911 & ~n7920 ;
  assign n7922 = n7919 & n7921 ;
  assign n7927 = n7926 ^ n7922 ;
  assign n7928 = ~n7918 & ~n7927 ;
  assign n7846 = n7845 ^ x204 ;
  assign n7848 = x200 & n7846 ;
  assign n7849 = n7848 ^ x204 ;
  assign n7852 = x204 ^ x201 ;
  assign n7853 = n7852 ^ n7844 ;
  assign n1288 = x200 ^ x199 ;
  assign n7854 = n7853 ^ n1288 ;
  assign n7855 = n7845 ^ n1288 ;
  assign n7856 = n7855 ^ n7844 ;
  assign n7857 = n7856 ^ x204 ;
  assign n7858 = ~n7854 & n7857 ;
  assign n7861 = n7858 ^ x202 ;
  assign n7862 = ~n7849 & ~n7861 ;
  assign n7865 = ~x203 & n7862 ;
  assign n7890 = n7889 ^ x202 ;
  assign n7894 = n7890 & n7893 ;
  assign n7891 = n7890 ^ n7888 ;
  assign n7892 = x201 & n7891 ;
  assign n7895 = n7894 ^ n7892 ;
  assign n7896 = n7895 ^ n7886 ;
  assign n7899 = x199 & n7896 ;
  assign n7900 = n7899 ^ n7895 ;
  assign n7901 = ~n7865 & ~n7900 ;
  assign n7929 = n7928 ^ n7901 ;
  assign n1291 = n1290 ^ n1289 ;
  assign n1292 = n1291 ^ n1288 ;
  assign n1296 = n1295 ^ n1294 ;
  assign n1297 = n1296 ^ n1293 ;
  assign n7930 = n1292 & n1297 ;
  assign n8411 = n7930 ^ n7928 ;
  assign n8412 = ~n7929 & n8411 ;
  assign n8413 = n8412 ^ n7930 ;
  assign n8418 = n8417 ^ n8413 ;
  assign n8422 = n8421 ^ n8418 ;
  assign n8424 = n8422 ^ n8413 ;
  assign n8425 = n8423 & n8424 ;
  assign n8426 = n8425 ^ n8422 ;
  assign n8410 = n8409 ^ n8391 ;
  assign n8427 = n8426 ^ n8410 ;
  assign n8351 = n7930 ^ n7929 ;
  assign n8348 = n7931 ^ n7842 ;
  assign n8352 = n8351 ^ n8348 ;
  assign n8367 = n8352 ^ n7929 ;
  assign n8359 = n8352 ^ n7930 ;
  assign n1298 = n1297 ^ n1292 ;
  assign n1309 = n1308 ^ n1303 ;
  assign n7932 = n1298 & n1309 ;
  assign n8356 = n7932 ^ n7930 ;
  assign n8360 = n8359 ^ n8356 ;
  assign n8368 = n8367 ^ n8360 ;
  assign n8369 = ~n7929 & n8368 ;
  assign n8378 = n8369 ^ n8368 ;
  assign n8372 = n8369 ^ n8351 ;
  assign n8373 = n8348 ^ n7932 ;
  assign n8374 = n8373 ^ n8369 ;
  assign n8375 = n8372 & n8374 ;
  assign n8379 = n8378 ^ n8375 ;
  assign n8370 = n8369 ^ n7931 ;
  assign n8371 = n8369 ^ n7842 ;
  assign n8376 = ~n8371 & n8375 ;
  assign n8377 = ~n8370 & n8376 ;
  assign n8380 = n8379 ^ n8377 ;
  assign n8381 = n8380 ^ n8351 ;
  assign n8382 = n8381 ^ n8356 ;
  assign n8385 = n8382 ^ n7929 ;
  assign n8386 = n8385 ^ n8348 ;
  assign n8387 = n8386 ^ n7930 ;
  assign n8388 = n8387 ^ n8348 ;
  assign n8428 = n8427 ^ n8388 ;
  assign n8341 = n7902 & n7910 ;
  assign n8342 = ~n7927 & n8341 ;
  assign n8343 = n8342 ^ n7927 ;
  assign n8429 = n8428 ^ n8343 ;
  assign n11893 = n8429 ^ n8410 ;
  assign n11896 = n8413 ^ n8388 ;
  assign n11897 = n8426 & n11896 ;
  assign n11898 = n11897 ^ n8388 ;
  assign n11899 = n11898 ^ n8410 ;
  assign n11900 = n11899 ^ n8429 ;
  assign n11901 = n8343 & n11900 ;
  assign n11902 = n11901 ^ n8429 ;
  assign n11903 = n11893 & n11902 ;
  assign n11904 = n11903 ^ n11899 ;
  assign n11908 = n11907 ^ n11904 ;
  assign n11925 = n11924 ^ n11908 ;
  assign n1333 = n1332 ^ n1321 ;
  assign n1310 = n1309 ^ n1298 ;
  assign n7637 = n1321 ^ n1310 ;
  assign n7638 = n1333 & ~n7637 ;
  assign n7639 = n7638 ^ n1332 ;
  assign n8339 = n7639 & ~n8360 ;
  assign n8336 = n8360 ^ n8335 ;
  assign n8337 = n8336 ^ n7639 ;
  assign n8338 = n7788 & ~n8337 ;
  assign n8340 = n8339 ^ n8338 ;
  assign n8430 = n8429 ^ n8340 ;
  assign n11890 = n8465 ^ n8429 ;
  assign n11891 = ~n8430 & ~n11890 ;
  assign n11892 = n11891 ^ n8465 ;
  assign n11926 = n11925 ^ n11892 ;
  assign n11889 = n11888 ^ n11870 ;
  assign n11927 = n11926 ^ n11889 ;
  assign n8466 = n8465 ^ n8430 ;
  assign n8334 = n8333 ^ n8157 ;
  assign n8467 = n8466 ^ n8334 ;
  assign n7789 = n7788 ^ n7639 ;
  assign n7937 = n8360 ^ n7789 ;
  assign n7402 = n7401 ^ n7400 ;
  assign n7636 = n7635 ^ n7402 ;
  assign n7938 = n7937 ^ n7636 ;
  assign n1334 = n1333 ^ n1310 ;
  assign n1381 = n1380 ^ n1357 ;
  assign n7947 = n1334 & n1381 ;
  assign n8149 = n7947 ^ n7636 ;
  assign n8150 = ~n7938 & ~n8149 ;
  assign n8151 = n8150 ^ n7937 ;
  assign n11928 = n8466 ^ n8151 ;
  assign n11929 = ~n8467 & n11928 ;
  assign n11930 = n11929 ^ n8466 ;
  assign n12539 = n11930 ^ n11926 ;
  assign n12540 = ~n11927 & ~n12539 ;
  assign n12541 = n12540 ^ n11930 ;
  assign n12562 = n11924 ^ n11892 ;
  assign n12563 = ~n11925 & ~n12562 ;
  assign n12564 = n12563 ^ n11924 ;
  assign n12555 = n11912 & ~n11916 ;
  assign n12554 = ~n11917 & n11923 ;
  assign n12556 = n12555 ^ n12554 ;
  assign n12559 = ~n11904 & n11907 ;
  assign n12557 = ~n8410 & ~n8429 ;
  assign n12558 = n11898 & n12557 ;
  assign n12560 = n12559 ^ n12558 ;
  assign n12840 = ~n12556 & n12560 ;
  assign n12844 = ~n12564 & ~n12840 ;
  assign n12842 = n12840 ^ n12556 ;
  assign n12843 = n12842 ^ n12560 ;
  assign n12847 = n12844 ^ n12843 ;
  assign n12845 = ~n12843 & ~n12844 ;
  assign n12848 = n12847 ^ n12845 ;
  assign n12841 = n12840 ^ n12564 ;
  assign n12846 = n12845 ^ n12841 ;
  assign n12849 = n12848 ^ n12846 ;
  assign n12850 = n12547 ^ n12544 ;
  assign n12851 = n12552 & ~n12850 ;
  assign n12852 = n12851 ^ n12551 ;
  assign n12853 = n12849 & n12852 ;
  assign n12854 = ~n12541 & n12853 ;
  assign n12855 = ~n12553 & n12854 ;
  assign n12856 = n12855 ^ n12853 ;
  assign n12857 = n12856 ^ n12849 ;
  assign n12858 = n12857 ^ n12564 ;
  assign n12561 = n12560 ^ n12556 ;
  assign n12565 = n12564 ^ n12561 ;
  assign n12566 = n12565 ^ n12553 ;
  assign n12567 = n12566 ^ n12541 ;
  assign n12876 = ~n12567 & ~n12840 ;
  assign n12859 = ~n12547 & ~n12551 ;
  assign n12870 = n12842 & n12859 ;
  assign n12860 = ~n12556 & n12558 ;
  assign n12861 = ~n12547 & n12860 ;
  assign n12862 = n12861 ^ n12556 ;
  assign n12864 = ~n12551 & n12560 ;
  assign n12865 = ~n12862 & n12864 ;
  assign n12866 = n12865 ^ n12861 ;
  assign n12867 = n12866 ^ n12840 ;
  assign n12871 = n12870 ^ n12867 ;
  assign n12872 = ~n12544 & n12871 ;
  assign n12873 = n12872 ^ n12866 ;
  assign n12877 = n12876 ^ n12873 ;
  assign n12878 = n12857 & n12877 ;
  assign n12879 = n12878 ^ n12873 ;
  assign n12880 = n12858 & n12879 ;
  assign n12881 = n12880 ^ n12857 ;
  assign n12882 = n12848 ^ n12553 ;
  assign n12883 = ~n12845 & ~n12882 ;
  assign n12884 = n12848 ^ n12541 ;
  assign n12885 = n12883 & ~n12884 ;
  assign n12886 = n12885 ^ n12848 ;
  assign n12887 = n12886 ^ n12852 ;
  assign n12888 = n12887 ^ n12886 ;
  assign n12889 = ~n12541 & n12848 ;
  assign n12890 = n12889 ^ n12886 ;
  assign n12891 = ~n12888 & ~n12890 ;
  assign n12892 = n12891 ^ n12886 ;
  assign n12893 = ~n12881 & ~n12892 ;
  assign n12894 = n12893 ^ n12881 ;
  assign n13142 = ~n12881 & n12886 ;
  assign n13143 = n12852 & n13142 ;
  assign n13144 = n13143 ^ n12886 ;
  assign n11931 = n11930 ^ n11927 ;
  assign n6981 = x95 & x96 ;
  assign n1259 = x96 ^ x95 ;
  assign n6982 = n6981 ^ n1259 ;
  assign n6983 = x91 & x92 ;
  assign n1257 = x92 ^ x91 ;
  assign n6984 = n6983 ^ n1257 ;
  assign n6985 = n6984 ^ x94 ;
  assign n6986 = n6984 ^ x93 ;
  assign n6987 = ~n6985 & ~n6986 ;
  assign n6988 = n6987 ^ n6984 ;
  assign n6989 = n6983 ^ n6981 ;
  assign n6990 = n6985 ^ n6983 ;
  assign n6991 = n6990 ^ n6986 ;
  assign n6992 = n6989 & n6991 ;
  assign n6993 = n6992 ^ n6984 ;
  assign n6994 = n6988 & n6993 ;
  assign n6995 = n6994 ^ n6984 ;
  assign n6996 = n6995 ^ n6983 ;
  assign n6997 = n6982 & n6996 ;
  assign n1256 = x94 ^ x93 ;
  assign n6998 = x95 ^ x94 ;
  assign n7001 = n6998 ^ x96 ;
  assign n7002 = ~x92 & n7001 ;
  assign n7003 = n7002 ^ n6998 ;
  assign n7004 = n1259 & ~n7003 ;
  assign n7005 = n7004 ^ n6998 ;
  assign n7006 = ~n1256 & ~n7005 ;
  assign n7007 = ~x91 & n7006 ;
  assign n7008 = x93 & x94 ;
  assign n7020 = ~n6981 & ~n6983 ;
  assign n7021 = n7008 & n7020 ;
  assign n7022 = n7021 ^ n7008 ;
  assign n7023 = n7022 ^ n6981 ;
  assign n1258 = n1257 ^ n1256 ;
  assign n7015 = ~x92 & ~n6982 ;
  assign n7016 = n1258 & n7015 ;
  assign n7017 = n7016 ^ n1258 ;
  assign n7009 = n6981 ^ n1258 ;
  assign n7018 = n7017 ^ n7009 ;
  assign n7019 = ~n7008 & n7018 ;
  assign n7024 = n7023 ^ n7019 ;
  assign n7025 = ~n7007 & ~n7024 ;
  assign n7026 = ~n6997 & n7025 ;
  assign n6935 = x101 & x102 ;
  assign n1254 = x102 ^ x101 ;
  assign n6936 = n6935 ^ n1254 ;
  assign n6937 = x97 & x98 ;
  assign n1252 = x98 ^ x97 ;
  assign n6938 = n6937 ^ n1252 ;
  assign n6939 = n6938 ^ x100 ;
  assign n6940 = n6938 ^ x99 ;
  assign n6941 = ~n6939 & ~n6940 ;
  assign n6942 = n6941 ^ n6938 ;
  assign n6943 = n6937 ^ n6935 ;
  assign n6944 = n6939 ^ n6937 ;
  assign n6945 = n6944 ^ n6940 ;
  assign n6946 = n6943 & n6945 ;
  assign n6947 = n6946 ^ n6938 ;
  assign n6948 = n6942 & n6947 ;
  assign n6949 = n6948 ^ n6938 ;
  assign n6950 = n6949 ^ n6937 ;
  assign n6951 = n6936 & n6950 ;
  assign n1251 = x100 ^ x99 ;
  assign n6952 = x101 ^ x100 ;
  assign n6955 = n6952 ^ x102 ;
  assign n6956 = ~x98 & n6955 ;
  assign n6957 = n6956 ^ n6952 ;
  assign n6958 = n1254 & ~n6957 ;
  assign n6959 = n6958 ^ n6952 ;
  assign n6960 = ~n1251 & ~n6959 ;
  assign n6961 = ~x97 & n6960 ;
  assign n6962 = x99 & x100 ;
  assign n6974 = ~n6935 & ~n6937 ;
  assign n6975 = n6962 & n6974 ;
  assign n6976 = n6975 ^ n6962 ;
  assign n6977 = n6976 ^ n6935 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n6969 = ~x98 & ~n6936 ;
  assign n6970 = n1253 & n6969 ;
  assign n6971 = n6970 ^ n1253 ;
  assign n6963 = n6935 ^ n1253 ;
  assign n6972 = n6971 ^ n6963 ;
  assign n6973 = ~n6962 & n6972 ;
  assign n6978 = n6977 ^ n6973 ;
  assign n6979 = ~n6961 & ~n6978 ;
  assign n6980 = ~n6951 & n6979 ;
  assign n7027 = n7026 ^ n6980 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n1255 = n1254 ^ n1253 ;
  assign n1261 = n1260 ^ n1255 ;
  assign n1247 = x82 ^ x81 ;
  assign n1246 = x84 ^ x83 ;
  assign n1248 = n1247 ^ n1246 ;
  assign n1245 = x80 ^ x79 ;
  assign n1249 = n1248 ^ n1245 ;
  assign n1243 = x90 ^ x89 ;
  assign n1241 = x88 ^ x87 ;
  assign n1240 = x86 ^ x85 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1244 = n1243 ^ n1242 ;
  assign n1250 = n1249 ^ n1244 ;
  assign n6929 = n1260 ^ n1250 ;
  assign n6930 = ~n1261 & n6929 ;
  assign n6931 = n6930 ^ n1250 ;
  assign n6932 = n1249 & ~n6931 ;
  assign n6933 = ~n6930 & n6932 ;
  assign n6934 = n6933 ^ n6931 ;
  assign n7028 = n7027 ^ n6934 ;
  assign n6926 = n1255 & n1260 ;
  assign n6927 = n1244 & n1249 ;
  assign n6928 = n6926 & n6927 ;
  assign n7029 = n7028 ^ n6928 ;
  assign n6890 = ~x83 & ~x84 ;
  assign n6891 = n6890 ^ n1246 ;
  assign n6892 = n6891 ^ x82 ;
  assign n6893 = n1247 & n6892 ;
  assign n6894 = n6893 ^ x81 ;
  assign n6896 = ~n6890 & n6894 ;
  assign n6895 = n6894 ^ n6890 ;
  assign n6897 = n6896 ^ n6895 ;
  assign n6898 = ~x80 & n6897 ;
  assign n6899 = x81 & x82 ;
  assign n6900 = n6899 ^ n1247 ;
  assign n6901 = n6898 & ~n6900 ;
  assign n6913 = x80 & ~n6890 ;
  assign n6912 = ~n6891 & n6899 ;
  assign n6902 = n6893 ^ n6892 ;
  assign n6919 = n6912 ^ n6902 ;
  assign n6920 = ~n6913 & n6919 ;
  assign n6914 = n6894 & ~n6913 ;
  assign n6915 = ~n6912 & n6914 ;
  assign n6916 = n6915 ^ n6894 ;
  assign n6911 = n6901 ^ n6898 ;
  assign n6917 = n6916 ^ n6911 ;
  assign n6907 = ~n6897 & ~n6902 ;
  assign n6908 = n6907 ^ n6896 ;
  assign n6909 = x80 & n6908 ;
  assign n6910 = n6909 ^ n6896 ;
  assign n6918 = n6917 ^ n6910 ;
  assign n6921 = n6920 ^ n6918 ;
  assign n6922 = ~x79 & n6921 ;
  assign n6923 = n6922 ^ n6910 ;
  assign n6924 = ~n6901 & ~n6923 ;
  assign n6849 = ~x89 & ~x90 ;
  assign n6850 = n6849 ^ n1243 ;
  assign n6851 = ~x87 & ~x88 ;
  assign n6852 = n6851 ^ n1241 ;
  assign n6854 = ~n6850 & ~n6852 ;
  assign n6853 = n6852 ^ n6850 ;
  assign n6855 = n6854 ^ n6853 ;
  assign n6856 = ~n6849 & ~n6851 ;
  assign n6861 = ~x86 & ~n6856 ;
  assign n6862 = ~n6855 & n6861 ;
  assign n6863 = n6862 ^ n6855 ;
  assign n6864 = n6863 ^ n6853 ;
  assign n6865 = ~x85 & n6864 ;
  assign n6866 = x85 & x86 ;
  assign n6885 = n6849 & n6851 ;
  assign n6886 = ~n6866 & n6885 ;
  assign n6887 = n6886 ^ n6866 ;
  assign n6867 = n6866 ^ n6856 ;
  assign n6868 = n6867 ^ n6852 ;
  assign n6869 = n6866 ^ n6853 ;
  assign n6870 = n6869 ^ n1240 ;
  assign n6871 = ~n6856 & n6870 ;
  assign n6872 = n6871 ^ n6870 ;
  assign n6873 = ~n6868 & n6872 ;
  assign n6874 = n6873 ^ n6867 ;
  assign n6875 = n6871 ^ n1240 ;
  assign n6876 = n6875 ^ n6873 ;
  assign n6877 = n6874 & n6876 ;
  assign n6888 = n6887 ^ n6877 ;
  assign n6889 = ~n6865 & ~n6888 ;
  assign n6925 = n6924 ^ n6889 ;
  assign n7030 = n7029 ^ n6925 ;
  assign n6766 = ~x111 & ~x112 ;
  assign n6768 = ~x113 & ~x114 ;
  assign n6774 = ~n6766 & ~n6768 ;
  assign n1280 = x112 ^ x111 ;
  assign n1279 = x114 ^ x113 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n6767 = n6766 ^ n1280 ;
  assign n6769 = n6768 ^ n1279 ;
  assign n6770 = n6767 & n6769 ;
  assign n6771 = n6770 ^ x110 ;
  assign n6772 = ~n1281 & ~n6771 ;
  assign n6773 = n6772 ^ x110 ;
  assign n6775 = n6774 ^ n6773 ;
  assign n6821 = x111 ^ x110 ;
  assign n6822 = ~n1280 & ~n6821 ;
  assign n6823 = x114 ^ x109 ;
  assign n6826 = ~x112 & ~n6823 ;
  assign n6827 = n6826 ^ x109 ;
  assign n6828 = n6822 & n6827 ;
  assign n6829 = ~x113 & n6828 ;
  assign n6830 = n6774 ^ n6770 ;
  assign n6831 = x109 & x110 ;
  assign n6832 = x114 & ~n6767 ;
  assign n6833 = n6831 & n6832 ;
  assign n6834 = n6833 ^ n6831 ;
  assign n6835 = n6834 ^ n6770 ;
  assign n6836 = n6830 & ~n6835 ;
  assign n1282 = x110 ^ x109 ;
  assign n6837 = n6836 ^ n6834 ;
  assign n6838 = ~n1282 & n6837 ;
  assign n6839 = n6836 & n6838 ;
  assign n6840 = n6839 ^ n6837 ;
  assign n6841 = ~n6829 & ~n6840 ;
  assign n6844 = ~x109 & n6841 ;
  assign n6845 = ~n6775 & n6844 ;
  assign n6776 = x103 & ~x104 ;
  assign n6803 = x107 ^ x106 ;
  assign n6778 = x108 ^ x105 ;
  assign n6804 = n6803 ^ n6778 ;
  assign n6777 = n6804 ^ x105 ;
  assign n6781 = n6777 & n6778 ;
  assign n6782 = n6781 ^ x105 ;
  assign n6783 = n6776 & ~n6782 ;
  assign n6785 = n6783 ^ n6776 ;
  assign n6786 = ~x106 & ~x107 ;
  assign n6787 = n6785 & n6786 ;
  assign n6784 = n6783 ^ x103 ;
  assign n6788 = n6787 ^ n6784 ;
  assign n1276 = x106 ^ x105 ;
  assign n6789 = x107 ^ x105 ;
  assign n6790 = ~n1276 & n6789 ;
  assign n1275 = x108 ^ x107 ;
  assign n6791 = n6790 ^ n1275 ;
  assign n6792 = n6791 ^ n1276 ;
  assign n6797 = x108 & ~n6790 ;
  assign n6798 = n6792 & n6797 ;
  assign n6799 = n6798 ^ n6792 ;
  assign n6800 = n6799 ^ n1276 ;
  assign n6801 = x104 & ~n6800 ;
  assign n6802 = n6788 & ~n6801 ;
  assign n6807 = x105 ^ x104 ;
  assign n6808 = n6804 & ~n6807 ;
  assign n6806 = ~n1275 & ~n6803 ;
  assign n6809 = n6808 ^ n6806 ;
  assign n6810 = ~x103 & n6809 ;
  assign n6811 = ~n6802 & ~n6810 ;
  assign n6812 = ~n1276 & ~n6807 ;
  assign n6813 = x108 ^ x103 ;
  assign n6816 = ~x106 & ~n6813 ;
  assign n6817 = n6816 ^ x103 ;
  assign n6818 = n6812 & n6817 ;
  assign n6819 = ~x107 & n6818 ;
  assign n6820 = n6811 & ~n6819 ;
  assign n6842 = n6841 ^ n6820 ;
  assign n6846 = n6845 ^ n6842 ;
  assign n1271 = x120 ^ x119 ;
  assign n1269 = x116 ^ x115 ;
  assign n1268 = x118 ^ x117 ;
  assign n1270 = n1269 ^ n1268 ;
  assign n1272 = n1271 ^ n1270 ;
  assign n1266 = x124 ^ x123 ;
  assign n1264 = x126 ^ x125 ;
  assign n1263 = x122 ^ x121 ;
  assign n1265 = n1264 ^ n1263 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1273 = n1272 ^ n1267 ;
  assign n1274 = x104 ^ x103 ;
  assign n1278 = n6804 ^ n1274 ;
  assign n6761 = n1278 ^ n1272 ;
  assign n6764 = ~n1273 & ~n6761 ;
  assign n1283 = n1282 ^ n1281 ;
  assign n6762 = n6761 ^ n1267 ;
  assign n6763 = ~n1283 & n6762 ;
  assign n6765 = n6764 ^ n6763 ;
  assign n6847 = n6846 ^ n6765 ;
  assign n6710 = x125 & x126 ;
  assign n6709 = x123 & x124 ;
  assign n6753 = n6709 ^ n1266 ;
  assign n6754 = ~n6710 & ~n6753 ;
  assign n6711 = n6710 ^ n1264 ;
  assign n6717 = x121 & x122 ;
  assign n6723 = n6717 ^ n1263 ;
  assign n6724 = n6723 ^ x124 ;
  assign n6725 = n6723 ^ x123 ;
  assign n6726 = ~n6724 & ~n6725 ;
  assign n6727 = n6726 ^ n6723 ;
  assign n6728 = n6717 ^ n6710 ;
  assign n6729 = n6724 ^ n6717 ;
  assign n6730 = n6729 ^ n6725 ;
  assign n6731 = n6728 & n6730 ;
  assign n6732 = n6731 ^ n6723 ;
  assign n6733 = n6727 & n6732 ;
  assign n6734 = n6733 ^ n6723 ;
  assign n6735 = n6734 ^ n6717 ;
  assign n6736 = n6711 & n6735 ;
  assign n6752 = ~n1267 & ~n6736 ;
  assign n6755 = n6754 ^ n6752 ;
  assign n6756 = n1267 ^ x121 ;
  assign n6757 = ~n6755 & n6756 ;
  assign n6746 = n1271 ^ x116 ;
  assign n6747 = n6746 ^ n1268 ;
  assign n6748 = n1269 & ~n6747 ;
  assign n6749 = n6748 ^ x115 ;
  assign n6739 = x119 & x120 ;
  assign n6738 = x117 & x118 ;
  assign n6740 = n6739 ^ n6738 ;
  assign n6741 = n6738 ^ n1268 ;
  assign n6742 = n6739 ^ n1271 ;
  assign n6743 = n6741 & n6742 ;
  assign n6744 = n6743 ^ n6738 ;
  assign n6745 = ~n6740 & ~n6744 ;
  assign n6750 = n6749 ^ n6745 ;
  assign n6722 = n6710 ^ x121 ;
  assign n6737 = n6736 ^ n6722 ;
  assign n6751 = n6750 ^ n6737 ;
  assign n6758 = n6757 ^ n6751 ;
  assign n6718 = n6709 & ~n6710 ;
  assign n6719 = ~n6717 & n6718 ;
  assign n6720 = n6719 ^ n6709 ;
  assign n6721 = n1267 & ~n6720 ;
  assign n6759 = n6758 ^ n6721 ;
  assign n6714 = x122 & ~n6711 ;
  assign n6715 = n6714 ^ n1264 ;
  assign n6716 = ~n6709 & ~n6715 ;
  assign n6760 = n6759 ^ n6716 ;
  assign n6848 = n6847 ^ n6760 ;
  assign n7031 = n7030 ^ n6848 ;
  assign n1284 = n1283 ^ n1278 ;
  assign n1285 = n1284 ^ n1273 ;
  assign n1262 = n1261 ^ n1250 ;
  assign n1286 = n1285 ^ n1262 ;
  assign n1239 = n1238 ^ n1215 ;
  assign n6701 = n1262 ^ n1239 ;
  assign n6702 = n1286 & ~n6701 ;
  assign n6703 = n6702 ^ n1285 ;
  assign n8140 = n7031 ^ n6703 ;
  assign n8141 = n7395 ^ n6706 ;
  assign n8142 = n8141 ^ n6703 ;
  assign n8143 = ~n8140 & ~n8142 ;
  assign n8115 = n6773 & n6774 ;
  assign n8116 = ~n6840 & n8115 ;
  assign n8117 = n8116 ^ n6840 ;
  assign n8095 = x106 ^ x104 ;
  assign n8098 = n6807 & n8095 ;
  assign n8099 = n8098 ^ x104 ;
  assign n8108 = n1276 ^ x104 ;
  assign n8104 = n6803 ^ x105 ;
  assign n8105 = n8104 ^ x104 ;
  assign n8106 = ~n1275 & n8105 ;
  assign n8109 = n8108 ^ n8106 ;
  assign n8110 = n8099 & n8109 ;
  assign n8113 = ~n6802 & ~n8110 ;
  assign n11783 = n8117 ^ n8113 ;
  assign n8091 = n1278 & n1283 ;
  assign n8092 = n8091 ^ n6820 ;
  assign n8093 = n6846 & n8092 ;
  assign n8094 = n8093 ^ n6820 ;
  assign n11784 = n11783 ^ n8094 ;
  assign n8071 = n1267 & n1272 ;
  assign n8132 = n8071 ^ n6750 ;
  assign n8133 = n6760 & ~n8132 ;
  assign n8134 = n8133 ^ n6750 ;
  assign n8120 = n6743 ^ x116 ;
  assign n8121 = n6740 ^ x115 ;
  assign n8122 = n8121 ^ n6743 ;
  assign n8123 = n8120 & ~n8122 ;
  assign n8126 = n8123 ^ n6743 ;
  assign n8124 = n8123 ^ n6744 ;
  assign n8125 = ~n6740 & n8124 ;
  assign n8127 = n8126 ^ n8125 ;
  assign n8128 = x115 & n8125 ;
  assign n8129 = ~n8127 & n8128 ;
  assign n8130 = n8129 ^ n8127 ;
  assign n8119 = ~n6720 & ~n6736 ;
  assign n8131 = n8130 ^ n8119 ;
  assign n8135 = n8134 ^ n8131 ;
  assign n8136 = n11784 ^ n8135 ;
  assign n8072 = n8071 ^ n1278 ;
  assign n8073 = n8072 ^ n1273 ;
  assign n8074 = n8073 ^ n1278 ;
  assign n8075 = n6846 ^ n1283 ;
  assign n8076 = n8075 ^ n1278 ;
  assign n8077 = n8074 & n8076 ;
  assign n8078 = n8077 ^ n1278 ;
  assign n8079 = n1284 & ~n8078 ;
  assign n8080 = n8079 ^ n8075 ;
  assign n8081 = n8071 ^ n6847 ;
  assign n8084 = ~n6760 & ~n8081 ;
  assign n8085 = n8084 ^ n8071 ;
  assign n8086 = n8080 & ~n8085 ;
  assign n8137 = n8136 ^ n8086 ;
  assign n8067 = ~n6997 & ~n7022 ;
  assign n8066 = ~n6951 & ~n6976 ;
  assign n8068 = n8067 ^ n8066 ;
  assign n8063 = n7026 ^ n6926 ;
  assign n8064 = n7027 & n8063 ;
  assign n8065 = n8064 ^ n7026 ;
  assign n8069 = n8068 ^ n8065 ;
  assign n6878 = n6877 ^ n6866 ;
  assign n8059 = ~n6854 & ~n6878 ;
  assign n8056 = x79 & ~n6916 ;
  assign n8057 = n6910 & n8056 ;
  assign n8058 = n8057 ^ n6916 ;
  assign n8060 = n8059 ^ n8058 ;
  assign n8053 = n6927 ^ n6924 ;
  assign n8054 = ~n6925 & n8053 ;
  assign n8055 = n8054 ^ n6927 ;
  assign n8061 = n8060 ^ n8055 ;
  assign n8045 = n6934 ^ n6926 ;
  assign n8046 = ~n7027 & ~n8045 ;
  assign n8047 = n8046 ^ n6926 ;
  assign n8048 = n7029 ^ n6927 ;
  assign n8050 = n6925 & n8048 ;
  assign n8051 = n8050 ^ n7029 ;
  assign n8052 = ~n8047 & ~n8051 ;
  assign n8062 = n8061 ^ n8052 ;
  assign n8070 = n8069 ^ n8062 ;
  assign n8138 = n8137 ^ n8070 ;
  assign n6704 = n1262 & n1285 ;
  assign n8042 = n7030 ^ n6704 ;
  assign n8043 = ~n7031 & n8042 ;
  assign n8044 = n8043 ^ n7030 ;
  assign n8139 = n8138 ^ n8044 ;
  assign n8144 = n8143 ^ n8139 ;
  assign n8041 = ~n6704 & ~n7031 ;
  assign n8145 = n8144 ^ n8041 ;
  assign n8040 = n8039 ^ n7990 ;
  assign n8146 = n8145 ^ n8040 ;
  assign n6705 = n6704 ^ n6703 ;
  assign n6707 = n6706 ^ n6705 ;
  assign n6708 = n6707 ^ n6704 ;
  assign n7032 = n7031 ^ n6708 ;
  assign n7396 = n7395 ^ n7032 ;
  assign n8147 = n8146 ^ n7396 ;
  assign n1382 = n1381 ^ n1334 ;
  assign n1287 = n1286 ^ n1239 ;
  assign n7397 = n1334 ^ n1287 ;
  assign n7398 = n1382 & ~n7397 ;
  assign n7399 = n7398 ^ n1381 ;
  assign n7939 = n7938 ^ n7399 ;
  assign n7948 = n7947 ^ n7396 ;
  assign n7949 = n7948 ^ n7399 ;
  assign n7950 = n7939 & ~n7949 ;
  assign n8148 = n8147 ^ n7950 ;
  assign n8468 = n8467 ^ n8151 ;
  assign n11851 = n8468 ^ n8146 ;
  assign n11852 = ~n8148 & ~n11851 ;
  assign n11853 = n11852 ^ n8468 ;
  assign n11932 = n11931 ^ n11853 ;
  assign n11848 = n11847 ^ n11844 ;
  assign n11849 = n11848 ^ n11833 ;
  assign n11791 = n8135 ^ n8113 ;
  assign n11792 = n8135 ^ n8117 ;
  assign n11793 = ~n11791 & n11792 ;
  assign n11794 = n11793 ^ n8135 ;
  assign n11798 = n11783 ^ n8135 ;
  assign n11795 = n8094 ^ n8086 ;
  assign n11796 = ~n8136 & ~n11795 ;
  assign n11799 = n11798 ^ n11796 ;
  assign n11800 = ~n11794 & n11799 ;
  assign n11785 = n11784 ^ n8086 ;
  assign n11786 = n8135 & ~n11785 ;
  assign n8114 = n8113 ^ n8094 ;
  assign n11787 = n8113 ^ n8086 ;
  assign n11788 = ~n8114 & ~n11787 ;
  assign n11789 = n11788 ^ n8113 ;
  assign n11790 = n11786 & ~n11789 ;
  assign n11803 = n11800 ^ n11790 ;
  assign n11780 = n8134 ^ n8130 ;
  assign n11781 = n8131 & ~n11780 ;
  assign n11782 = n11781 ^ n8134 ;
  assign n11804 = n11803 ^ n11782 ;
  assign n11777 = n8137 ^ n8044 ;
  assign n11778 = n8138 & ~n11777 ;
  assign n11771 = n8067 ^ n8065 ;
  assign n11772 = n8068 & ~n11771 ;
  assign n11773 = n11772 ^ n8067 ;
  assign n11760 = ~n8055 & ~n8058 ;
  assign n11761 = ~n8052 & n8059 ;
  assign n11767 = ~n11760 & ~n11761 ;
  assign n11763 = ~n8062 & ~n8069 ;
  assign n11768 = n11763 ^ n8062 ;
  assign n11769 = n11767 & ~n11768 ;
  assign n11762 = n11761 ^ n11760 ;
  assign n11764 = n11763 ^ n11760 ;
  assign n11765 = n11762 & ~n11764 ;
  assign n11766 = n11765 ^ n11761 ;
  assign n11770 = n11769 ^ n11766 ;
  assign n11774 = n11773 ^ n11770 ;
  assign n11775 = n11774 ^ n8137 ;
  assign n11779 = n11778 ^ n11775 ;
  assign n11805 = n11804 ^ n11779 ;
  assign n11806 = n11805 ^ n8139 ;
  assign n11807 = n11806 ^ n8040 ;
  assign n11808 = n11807 ^ n11805 ;
  assign n11809 = n8145 & ~n11808 ;
  assign n11810 = n11809 ^ n11806 ;
  assign n11850 = n11849 ^ n11810 ;
  assign n12568 = n11853 ^ n11850 ;
  assign n12569 = n11932 & n12568 ;
  assign n12570 = n12569 ^ n11850 ;
  assign n12571 = n12570 ^ n12567 ;
  assign n12616 = n12590 & ~n12604 ;
  assign n12624 = ~n11833 & ~n11839 ;
  assign n12625 = n12624 ^ n12622 ;
  assign n12623 = n12622 ^ n11839 ;
  assign n12626 = n12625 ^ n12623 ;
  assign n12627 = n12616 & ~n12626 ;
  assign n12628 = n12627 ^ n12625 ;
  assign n12635 = n12587 & ~n12593 ;
  assign n12636 = n12635 ^ n12630 ;
  assign n12637 = n12628 & n12636 ;
  assign n12638 = n12637 ^ n12622 ;
  assign n12639 = ~n12615 & ~n12638 ;
  assign n12583 = n11849 ^ n11805 ;
  assign n12584 = ~n11810 & n12583 ;
  assign n12585 = n12584 ^ n11805 ;
  assign n12579 = n11804 ^ n11774 ;
  assign n12580 = ~n11779 & n12579 ;
  assign n12581 = n12580 ^ n11774 ;
  assign n12574 = n11782 & ~n11800 ;
  assign n12575 = ~n11790 & n12574 ;
  assign n12576 = n12575 ^ n11800 ;
  assign n12577 = n12576 ^ n11766 ;
  assign n12572 = ~n11769 & n11773 ;
  assign n12573 = ~n11766 & n12572 ;
  assign n12578 = n12577 ^ n12573 ;
  assign n12582 = n12581 ^ n12578 ;
  assign n12586 = n12585 ^ n12582 ;
  assign n12640 = n12639 ^ n12586 ;
  assign n12827 = n12640 ^ n12570 ;
  assign n12828 = n12571 & n12827 ;
  assign n12829 = n12828 ^ n12640 ;
  assign n12833 = n12581 ^ n12576 ;
  assign n12834 = ~n12578 & ~n12833 ;
  assign n12835 = n12834 ^ n12581 ;
  assign n13269 = n12829 & n12835 ;
  assign n13270 = n13144 & ~n13269 ;
  assign n13271 = n12894 & n13270 ;
  assign n13272 = ~n12837 & n13271 ;
  assign n13273 = n13272 ^ n13270 ;
  assign n13274 = n13273 ^ n13269 ;
  assign n12830 = n12639 ^ n12585 ;
  assign n12831 = n12586 & n12830 ;
  assign n12832 = n12831 ^ n12639 ;
  assign n13275 = n13274 ^ n12832 ;
  assign n13276 = n12835 ^ n12829 ;
  assign n13277 = n13276 ^ n13269 ;
  assign n13278 = n13277 ^ n13274 ;
  assign n13289 = n13278 ^ n13144 ;
  assign n13290 = n13289 ^ n13278 ;
  assign n13291 = n13278 ^ n12837 ;
  assign n13292 = n13291 ^ n13278 ;
  assign n13295 = n13277 & ~n13292 ;
  assign n13296 = ~n13290 & n13295 ;
  assign n13297 = n13296 ^ n13290 ;
  assign n13298 = n13297 ^ n13289 ;
  assign n13299 = ~n13275 & n13298 ;
  assign n13300 = n13299 ^ n13274 ;
  assign n5823 = ~x375 & ~x376 ;
  assign n1010 = x376 ^ x375 ;
  assign n5826 = n5823 ^ n1010 ;
  assign n5827 = x373 & x374 ;
  assign n5828 = x378 & n5827 ;
  assign n5829 = ~n5826 & n5828 ;
  assign n5830 = n5829 ^ n5827 ;
  assign n5824 = ~x377 & ~x378 ;
  assign n5825 = ~n5823 & ~n5824 ;
  assign n5831 = n5830 ^ n5825 ;
  assign n1008 = x378 ^ x377 ;
  assign n5832 = n5824 ^ n1008 ;
  assign n5837 = n5826 & n5832 ;
  assign n5838 = n5837 ^ n5825 ;
  assign n5839 = n5831 & n5838 ;
  assign n1007 = x374 ^ x373 ;
  assign n5840 = n5839 ^ n5830 ;
  assign n5841 = ~n1007 & n5840 ;
  assign n5842 = n5839 & n5841 ;
  assign n5843 = n5842 ^ n5840 ;
  assign n8879 = n5832 ^ n5826 ;
  assign n8880 = x374 & n5825 ;
  assign n8881 = n8880 ^ n5826 ;
  assign n8882 = n8879 & ~n8881 ;
  assign n8883 = n8882 ^ n5826 ;
  assign n8884 = ~n5843 & ~n8883 ;
  assign n8885 = n8884 ^ n5843 ;
  assign n1013 = x390 ^ x389 ;
  assign n5765 = x389 ^ x388 ;
  assign n5769 = ~n1013 & ~n5765 ;
  assign n5764 = x387 ^ x386 ;
  assign n5766 = n5765 ^ x387 ;
  assign n5767 = n5766 ^ x390 ;
  assign n5768 = ~n5764 & n5767 ;
  assign n5770 = n5769 ^ n5768 ;
  assign n5771 = ~x385 & n5770 ;
  assign n1014 = x388 ^ x387 ;
  assign n5772 = ~n1014 & ~n5764 ;
  assign n5773 = x390 ^ x385 ;
  assign n5776 = ~x388 & ~n5773 ;
  assign n5777 = n5776 ^ x385 ;
  assign n5778 = n5772 & n5777 ;
  assign n5779 = ~x389 & n5778 ;
  assign n5780 = ~x387 & ~x388 ;
  assign n5783 = n5780 ^ n1014 ;
  assign n5784 = x385 & x386 ;
  assign n5785 = x390 & n5784 ;
  assign n5786 = ~n5783 & n5785 ;
  assign n5787 = n5786 ^ n5784 ;
  assign n5781 = ~x389 & ~x390 ;
  assign n5782 = ~n5780 & ~n5781 ;
  assign n5788 = n5787 ^ n5782 ;
  assign n5789 = n5781 ^ n1013 ;
  assign n5794 = n5783 & n5789 ;
  assign n5795 = n5794 ^ n5782 ;
  assign n5796 = n5788 & n5795 ;
  assign n1015 = x386 ^ x385 ;
  assign n5797 = n5796 ^ n5787 ;
  assign n5798 = ~n1015 & n5797 ;
  assign n5799 = n5796 & n5798 ;
  assign n5800 = n5799 ^ n5797 ;
  assign n5801 = ~n5779 & ~n5800 ;
  assign n5802 = ~n5771 & n5801 ;
  assign n5727 = x383 & x384 ;
  assign n5726 = x381 & x382 ;
  assign n5731 = n5727 ^ n5726 ;
  assign n5728 = n5726 & n5727 ;
  assign n5732 = n5731 ^ n5728 ;
  assign n1018 = x382 ^ x381 ;
  assign n5735 = n5726 ^ n1018 ;
  assign n1019 = x384 ^ x383 ;
  assign n5736 = n5727 ^ n1019 ;
  assign n5737 = n5735 & n5736 ;
  assign n5740 = ~n5732 & ~n5737 ;
  assign n5741 = ~x380 & n5740 ;
  assign n5742 = n5741 ^ x380 ;
  assign n5729 = n5728 ^ x380 ;
  assign n5743 = n5742 ^ n5729 ;
  assign n5744 = ~x379 & n5743 ;
  assign n5748 = x379 & x380 ;
  assign n5759 = ~n5735 & ~n5736 ;
  assign n5760 = ~n5748 & n5759 ;
  assign n5761 = n5760 ^ n5748 ;
  assign n5745 = n5737 ^ n5732 ;
  assign n1020 = x380 ^ x379 ;
  assign n5746 = n5737 ^ n1020 ;
  assign n5747 = ~n5745 & ~n5746 ;
  assign n5749 = ~n5728 & n5748 ;
  assign n5750 = n5749 ^ n5732 ;
  assign n5751 = n5747 & n5750 ;
  assign n5752 = n5751 ^ n5749 ;
  assign n5753 = n5752 ^ n5748 ;
  assign n5762 = n5761 ^ n5753 ;
  assign n5763 = ~n5744 & ~n5762 ;
  assign n5803 = n5802 ^ n5763 ;
  assign n1005 = x370 ^ x369 ;
  assign n1003 = x372 ^ x371 ;
  assign n1002 = x368 ^ x367 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1009 = n1008 ^ n1007 ;
  assign n1011 = n1010 ^ n1009 ;
  assign n8867 = n1006 & n1011 ;
  assign n5847 = x371 ^ x370 ;
  assign n5851 = ~n1003 & ~n5847 ;
  assign n5846 = x369 ^ x368 ;
  assign n5848 = n5847 ^ x369 ;
  assign n5849 = n5848 ^ x372 ;
  assign n5850 = ~n5846 & n5849 ;
  assign n5852 = n5851 ^ n5850 ;
  assign n5853 = ~x367 & n5852 ;
  assign n5854 = ~n1005 & ~n5846 ;
  assign n5855 = x372 ^ x367 ;
  assign n5858 = ~x370 & ~n5855 ;
  assign n5859 = n5858 ^ x367 ;
  assign n5860 = n5854 & n5859 ;
  assign n5861 = ~x371 & n5860 ;
  assign n5862 = ~x369 & ~x370 ;
  assign n5865 = n5862 ^ n1005 ;
  assign n5866 = x367 & x368 ;
  assign n5867 = x372 & n5866 ;
  assign n5868 = ~n5865 & n5867 ;
  assign n5869 = n5868 ^ n5866 ;
  assign n5863 = ~x371 & ~x372 ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5870 = n5869 ^ n5864 ;
  assign n5871 = n5863 ^ n1003 ;
  assign n5876 = n5865 & n5871 ;
  assign n5877 = n5876 ^ n5864 ;
  assign n5878 = n5870 & n5877 ;
  assign n5879 = n5878 ^ n5869 ;
  assign n5880 = ~n1002 & n5879 ;
  assign n5881 = n5878 & n5880 ;
  assign n5882 = n5881 ^ n5879 ;
  assign n5883 = ~n5861 & ~n5882 ;
  assign n5884 = ~n5853 & n5883 ;
  assign n5808 = x377 ^ x376 ;
  assign n5812 = ~n1008 & ~n5808 ;
  assign n5807 = x375 ^ x374 ;
  assign n5809 = n5808 ^ x375 ;
  assign n5810 = n5809 ^ x378 ;
  assign n5811 = ~n5807 & n5810 ;
  assign n5813 = n5812 ^ n5811 ;
  assign n5814 = ~x373 & n5813 ;
  assign n5815 = ~n1010 & ~n5807 ;
  assign n5816 = x378 ^ x373 ;
  assign n5819 = ~x376 & ~n5816 ;
  assign n5820 = n5819 ^ x373 ;
  assign n5821 = n5815 & n5820 ;
  assign n5822 = ~x377 & n5821 ;
  assign n5844 = ~n5822 & ~n5843 ;
  assign n5845 = ~n5814 & n5844 ;
  assign n5885 = n5884 ^ n5845 ;
  assign n8868 = n8867 ^ n5885 ;
  assign n1016 = n1015 ^ n1014 ;
  assign n1017 = n1016 ^ n1013 ;
  assign n1021 = n1020 ^ n1019 ;
  assign n1022 = n1021 ^ n1018 ;
  assign n5804 = n1017 & n1022 ;
  assign n8869 = n8868 ^ n5804 ;
  assign n1012 = n1011 ^ n1006 ;
  assign n5805 = n5804 ^ n5803 ;
  assign n1023 = n1022 ^ n1017 ;
  assign n5806 = n5805 ^ n1023 ;
  assign n5886 = n5885 ^ n5806 ;
  assign n5887 = n5886 ^ n1006 ;
  assign n5888 = n5887 ^ n5805 ;
  assign n5889 = n5888 ^ n5885 ;
  assign n5890 = ~n1012 & n5889 ;
  assign n5891 = n5890 ^ n5886 ;
  assign n8870 = n8869 ^ n5891 ;
  assign n8872 = ~n5803 & ~n8870 ;
  assign n8873 = n8872 ^ n5804 ;
  assign n8874 = n8867 ^ n5891 ;
  assign n8875 = n8872 ^ n8870 ;
  assign n8876 = n8874 & ~n8875 ;
  assign n8877 = n8876 ^ n5891 ;
  assign n8878 = ~n8873 & ~n8877 ;
  assign n8886 = n8885 ^ n8878 ;
  assign n8887 = n8867 ^ n5884 ;
  assign n8888 = n5885 & n8887 ;
  assign n8889 = n8888 ^ n5884 ;
  assign n12103 = n8889 ^ n8885 ;
  assign n12104 = n8886 & n12103 ;
  assign n12105 = n12104 ^ n8885 ;
  assign n8902 = n5789 ^ n5783 ;
  assign n8903 = x386 & n5782 ;
  assign n8904 = n8903 ^ n5783 ;
  assign n8905 = n8902 & ~n8904 ;
  assign n8906 = n8905 ^ n5783 ;
  assign n8907 = ~n5800 & ~n8906 ;
  assign n8908 = n8907 ^ n5800 ;
  assign n8901 = ~n5728 & ~n5752 ;
  assign n8909 = n8908 ^ n8901 ;
  assign n8898 = n5804 ^ n5802 ;
  assign n8899 = ~n5803 & n8898 ;
  assign n8900 = n8899 ^ n5804 ;
  assign n8910 = n8909 ^ n8900 ;
  assign n8890 = n5871 ^ n5865 ;
  assign n8891 = x368 & n5864 ;
  assign n8892 = n8891 ^ n5865 ;
  assign n8893 = n8890 & ~n8892 ;
  assign n8894 = n8893 ^ n5865 ;
  assign n8895 = ~n5882 & ~n8894 ;
  assign n8896 = n8895 ^ n5882 ;
  assign n12106 = n8910 ^ n8896 ;
  assign n8897 = n8896 ^ n8889 ;
  assign n8911 = n8910 ^ n8897 ;
  assign n8912 = n8911 ^ n8886 ;
  assign n12107 = n8912 ^ n8896 ;
  assign n12108 = ~n12106 & ~n12107 ;
  assign n12109 = n12108 ^ n8910 ;
  assign n12110 = ~n12105 & n12109 ;
  assign n12100 = n8908 ^ n8900 ;
  assign n12101 = ~n8909 & n12100 ;
  assign n12102 = n12101 ^ n8908 ;
  assign n12111 = n8912 & n12105 ;
  assign n12112 = ~n12109 & n12111 ;
  assign n12668 = ~n12102 & ~n12112 ;
  assign n12669 = ~n12110 & n12668 ;
  assign n5921 = ~x393 & ~x394 ;
  assign n1038 = x394 ^ x393 ;
  assign n5924 = n5921 ^ n1038 ;
  assign n5925 = x391 & x392 ;
  assign n5926 = x396 & n5925 ;
  assign n5927 = ~n5924 & n5926 ;
  assign n5928 = n5927 ^ n5925 ;
  assign n5922 = ~x395 & ~x396 ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5929 = n5928 ^ n5923 ;
  assign n1036 = x396 ^ x395 ;
  assign n5930 = n5922 ^ n1036 ;
  assign n5935 = n5924 & n5930 ;
  assign n5936 = n5935 ^ n5923 ;
  assign n5937 = n5929 & n5936 ;
  assign n1037 = x392 ^ x391 ;
  assign n5938 = n5937 ^ n5928 ;
  assign n5939 = ~n1037 & n5938 ;
  assign n5940 = n5937 & n5939 ;
  assign n5941 = n5940 ^ n5938 ;
  assign n8937 = n5930 ^ n5924 ;
  assign n8938 = x392 & n5923 ;
  assign n8939 = n8938 ^ n5924 ;
  assign n8940 = n8937 & ~n8939 ;
  assign n8941 = n8940 ^ n5924 ;
  assign n8942 = ~n5941 & ~n8941 ;
  assign n8943 = n8942 ^ n5941 ;
  assign n5900 = x397 & x398 ;
  assign n5892 = x399 & x400 ;
  assign n5893 = x401 & x402 ;
  assign n5901 = n5892 & ~n5893 ;
  assign n5902 = ~n5900 & n5901 ;
  assign n5903 = n5902 ^ n5892 ;
  assign n1025 = x402 ^ x401 ;
  assign n5894 = n5893 ^ n1025 ;
  assign n1026 = x398 ^ x397 ;
  assign n5945 = n5900 ^ n1026 ;
  assign n5946 = n5945 ^ x400 ;
  assign n5947 = n5945 ^ x399 ;
  assign n5948 = ~n5946 & ~n5947 ;
  assign n5949 = n5948 ^ n5945 ;
  assign n5950 = n5900 ^ n5893 ;
  assign n5951 = n5946 ^ n5900 ;
  assign n5952 = n5951 ^ n5947 ;
  assign n5953 = n5950 & n5952 ;
  assign n5954 = n5953 ^ n5945 ;
  assign n5955 = n5949 & n5954 ;
  assign n5956 = n5955 ^ n5945 ;
  assign n5957 = n5956 ^ n5900 ;
  assign n5958 = n5894 & n5957 ;
  assign n8936 = ~n5903 & ~n5958 ;
  assign n8944 = n8943 ^ n8936 ;
  assign n1028 = x400 ^ x399 ;
  assign n5962 = n5892 ^ n1028 ;
  assign n5963 = ~n5893 & ~n5962 ;
  assign n1027 = n1026 ^ n1025 ;
  assign n1029 = n1028 ^ n1027 ;
  assign n5961 = ~n1029 & ~n5958 ;
  assign n5964 = n5963 ^ n5961 ;
  assign n5965 = n1029 ^ x397 ;
  assign n5966 = ~n5964 & n5965 ;
  assign n5944 = n5893 ^ x397 ;
  assign n5959 = n5958 ^ n5944 ;
  assign n5906 = x395 ^ x394 ;
  assign n5910 = ~n1036 & ~n5906 ;
  assign n5905 = x393 ^ x392 ;
  assign n5907 = n5906 ^ x393 ;
  assign n5908 = n5907 ^ x396 ;
  assign n5909 = ~n5905 & n5908 ;
  assign n5911 = n5910 ^ n5909 ;
  assign n5912 = ~x391 & n5911 ;
  assign n5913 = ~n1038 & ~n5905 ;
  assign n5914 = x396 ^ x391 ;
  assign n5917 = ~x394 & ~n5914 ;
  assign n5918 = n5917 ^ x391 ;
  assign n5919 = n5913 & n5918 ;
  assign n5920 = ~x395 & n5919 ;
  assign n5942 = ~n5920 & ~n5941 ;
  assign n5943 = ~n5912 & n5942 ;
  assign n5960 = n5959 ^ n5943 ;
  assign n5967 = n5966 ^ n5960 ;
  assign n5904 = n1029 & ~n5903 ;
  assign n5968 = n5967 ^ n5904 ;
  assign n5897 = x398 & ~n5894 ;
  assign n5898 = n5897 ^ n1025 ;
  assign n5899 = ~n5892 & ~n5898 ;
  assign n5969 = n5968 ^ n5899 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1040 = n1039 ^ n1036 ;
  assign n8927 = n1029 & n1040 ;
  assign n8933 = n8927 ^ n5943 ;
  assign n8934 = ~n5969 & n8933 ;
  assign n8935 = n8934 ^ n5943 ;
  assign n12085 = n8943 ^ n8935 ;
  assign n12086 = ~n8944 & n12085 ;
  assign n12087 = n12086 ^ n8943 ;
  assign n1041 = x408 ^ x407 ;
  assign n5983 = x407 ^ x406 ;
  assign n5987 = ~n1041 & ~n5983 ;
  assign n5982 = x405 ^ x404 ;
  assign n5984 = n5983 ^ x405 ;
  assign n5985 = n5984 ^ x408 ;
  assign n5986 = ~n5982 & n5985 ;
  assign n5988 = n5987 ^ n5986 ;
  assign n5989 = ~x403 & n5988 ;
  assign n1042 = x406 ^ x405 ;
  assign n5990 = ~n1042 & ~n5982 ;
  assign n5991 = x408 ^ x403 ;
  assign n5994 = ~x406 & ~n5991 ;
  assign n5995 = n5994 ^ x403 ;
  assign n5996 = n5990 & n5995 ;
  assign n5997 = ~x407 & n5996 ;
  assign n5998 = ~x405 & ~x406 ;
  assign n6001 = n5998 ^ n1042 ;
  assign n6002 = x403 & x404 ;
  assign n6003 = x408 & n6002 ;
  assign n6004 = ~n6001 & n6003 ;
  assign n6005 = n6004 ^ n6002 ;
  assign n5999 = ~x407 & ~x408 ;
  assign n6000 = ~n5998 & ~n5999 ;
  assign n6006 = n6005 ^ n6000 ;
  assign n6007 = n5999 ^ n1041 ;
  assign n6012 = n6001 & n6007 ;
  assign n6013 = n6012 ^ n6000 ;
  assign n6014 = n6006 & n6013 ;
  assign n1043 = x404 ^ x403 ;
  assign n6015 = n6014 ^ n6005 ;
  assign n6016 = ~n1043 & n6015 ;
  assign n6017 = n6014 & n6016 ;
  assign n6018 = n6017 ^ n6015 ;
  assign n6019 = ~n5997 & ~n6018 ;
  assign n6020 = ~n5989 & n6019 ;
  assign n1032 = x412 ^ x411 ;
  assign n1031 = x414 ^ x413 ;
  assign n5970 = n1032 ^ x413 ;
  assign n5971 = n5970 ^ x410 ;
  assign n5972 = n1031 & n5971 ;
  assign n5973 = n5972 ^ x413 ;
  assign n8955 = n5973 ^ x410 ;
  assign n8954 = n5973 ^ x412 ;
  assign n8956 = n8955 ^ n8954 ;
  assign n5980 = ~n1032 & n8956 ;
  assign n1033 = n1032 ^ n1031 ;
  assign n1030 = x410 ^ x409 ;
  assign n1034 = n1033 ^ n1030 ;
  assign n5974 = x409 & ~n1034 ;
  assign n5975 = n5974 ^ x410 ;
  assign n5976 = n5975 ^ n5973 ;
  assign n5981 = n5980 ^ n5976 ;
  assign n6021 = n6020 ^ n5981 ;
  assign n1035 = n1034 ^ n1029 ;
  assign n1044 = n1043 ^ n1042 ;
  assign n1045 = n1044 ^ n1041 ;
  assign n1046 = n1045 ^ n1040 ;
  assign n6022 = n1046 ^ n1034 ;
  assign n6023 = ~n1035 & n6022 ;
  assign n6024 = n6023 ^ n1046 ;
  assign n6025 = n1040 & n1045 ;
  assign n8923 = ~n6024 & ~n6025 ;
  assign n8918 = n1034 & n1045 ;
  assign n8924 = n8923 ^ n8918 ;
  assign n8925 = ~n6021 & n8924 ;
  assign n8926 = n8925 ^ n8918 ;
  assign n6026 = n6025 ^ n6024 ;
  assign n6027 = n6026 ^ n6021 ;
  assign n8928 = n8927 ^ n6027 ;
  assign n8930 = ~n5969 & n8928 ;
  assign n8931 = n8930 ^ n6027 ;
  assign n8932 = ~n8926 & ~n8931 ;
  assign n8964 = n8918 ^ n5981 ;
  assign n8965 = n8918 ^ n6020 ;
  assign n8966 = ~n8964 & n8965 ;
  assign n8967 = n8966 ^ n6020 ;
  assign n12077 = n8932 & n8967 ;
  assign n8953 = n5974 ^ n5973 ;
  assign n8959 = n1032 & n8956 ;
  assign n8960 = n8959 ^ n8954 ;
  assign n8961 = n8953 & ~n8960 ;
  assign n8962 = n8961 ^ n5974 ;
  assign n8946 = n6007 ^ n6001 ;
  assign n8947 = x404 & n6000 ;
  assign n8948 = n8947 ^ n6001 ;
  assign n8949 = n8946 & ~n8948 ;
  assign n8950 = n8949 ^ n6001 ;
  assign n8951 = ~n6018 & ~n8950 ;
  assign n8952 = n8951 ^ n6018 ;
  assign n8963 = n8962 ^ n8952 ;
  assign n8968 = n8967 ^ n8963 ;
  assign n8945 = n8944 ^ n8935 ;
  assign n8969 = n8968 ^ n8945 ;
  assign n8970 = n8969 ^ n8932 ;
  assign n12081 = ~n8952 & ~n8962 ;
  assign n12088 = ~n8970 & n12081 ;
  assign n12657 = ~n12077 & ~n12088 ;
  assign n12658 = ~n12087 & n12657 ;
  assign n12076 = n8967 ^ n8932 ;
  assign n12078 = n12077 ^ n12076 ;
  assign n12079 = ~n8945 & n12078 ;
  assign n12082 = n12081 ^ n8963 ;
  assign n12660 = n12079 & ~n12082 ;
  assign n12661 = n12658 & n12660 ;
  assign n12659 = n12658 ^ n12088 ;
  assign n12662 = n12661 ^ n12659 ;
  assign n12089 = n8945 & n12082 ;
  assign n12091 = n12082 ^ n12079 ;
  assign n12090 = n12089 ^ n12088 ;
  assign n12092 = n12091 ^ n12090 ;
  assign n12093 = n12092 ^ n12087 ;
  assign n12080 = n12079 ^ n8967 ;
  assign n12083 = ~n12080 & n12082 ;
  assign n12084 = ~n12076 & n12083 ;
  assign n12094 = n12093 ^ n12084 ;
  assign n12663 = n12089 & ~n12094 ;
  assign n12664 = ~n12662 & n12663 ;
  assign n12665 = n12664 ^ n12662 ;
  assign n12666 = n12665 ^ n12110 ;
  assign n12670 = n12669 ^ n12666 ;
  assign n1024 = n1023 ^ n1012 ;
  assign n1047 = n1046 ^ n1035 ;
  assign n6029 = n1024 & n1047 ;
  assign n6028 = n6027 ^ n5969 ;
  assign n6030 = n6029 ^ n6028 ;
  assign n8915 = n6028 ^ n5891 ;
  assign n8916 = ~n6030 & ~n8915 ;
  assign n8913 = n8912 ^ n6028 ;
  assign n8917 = n8916 ^ n8913 ;
  assign n12096 = n12094 ^ n8912 ;
  assign n12095 = n12094 ^ n8970 ;
  assign n12097 = n12096 ^ n12095 ;
  assign n12098 = n8917 & n12097 ;
  assign n12099 = n12098 ^ n12096 ;
  assign n12113 = n12112 ^ n12110 ;
  assign n12114 = n12113 ^ n12102 ;
  assign n12671 = n12114 ^ n12094 ;
  assign n12672 = n12099 & n12671 ;
  assign n12673 = n12672 ^ n12094 ;
  assign n12905 = n12673 ^ n12665 ;
  assign n12906 = n12670 & n12905 ;
  assign n12907 = n12906 ^ n12665 ;
  assign n5422 = ~x423 & ~x424 ;
  assign n5421 = ~x425 & ~x426 ;
  assign n1050 = x426 ^ x425 ;
  assign n5425 = n5421 ^ n1050 ;
  assign n5426 = ~n5422 & ~n5425 ;
  assign n1049 = x424 ^ x423 ;
  assign n5423 = n5422 ^ n1049 ;
  assign n5424 = ~n5421 & ~n5423 ;
  assign n5428 = n5426 ^ n5424 ;
  assign n5427 = ~n5424 & ~n5426 ;
  assign n5429 = n5428 ^ n5427 ;
  assign n1051 = x422 ^ x421 ;
  assign n5431 = n5423 ^ n5421 ;
  assign n5432 = n5431 ^ n5424 ;
  assign n5441 = n5432 ^ n5429 ;
  assign n5434 = n5425 ^ n5422 ;
  assign n5435 = n5434 ^ n5426 ;
  assign n5442 = x422 & n5435 ;
  assign n5443 = ~n5441 & n5442 ;
  assign n5444 = n5443 ^ n5427 ;
  assign n5445 = ~n1051 & ~n5444 ;
  assign n5446 = n5445 ^ n5427 ;
  assign n8747 = n5429 & n5446 ;
  assign n5458 = ~x419 & ~x420 ;
  assign n5459 = x415 & x416 ;
  assign n1055 = x416 ^ x415 ;
  assign n5460 = n5459 ^ n1055 ;
  assign n5461 = n5460 ^ x418 ;
  assign n5462 = n5460 ^ x417 ;
  assign n5463 = ~n5461 & ~n5462 ;
  assign n5464 = n5463 ^ n5460 ;
  assign n1054 = x420 ^ x419 ;
  assign n5465 = n5458 ^ n1054 ;
  assign n5466 = n5465 ^ n5459 ;
  assign n5467 = n5461 ^ n5459 ;
  assign n5468 = n5467 ^ n5462 ;
  assign n5469 = ~n5466 & n5468 ;
  assign n5470 = n5469 ^ n5460 ;
  assign n5471 = n5464 & n5470 ;
  assign n5472 = n5471 ^ n5460 ;
  assign n5473 = n5472 ^ n5459 ;
  assign n5474 = ~n5458 & n5473 ;
  assign n5476 = x417 & x418 ;
  assign n5480 = ~n5459 & n5465 ;
  assign n5481 = n5476 & n5480 ;
  assign n5482 = n5481 ^ n5476 ;
  assign n8746 = ~n5474 & ~n5482 ;
  assign n8748 = n8747 ^ n8746 ;
  assign n5479 = ~n5465 & n5476 ;
  assign n5483 = n5482 ^ n5479 ;
  assign n1056 = x418 ^ x417 ;
  assign n1057 = n1056 ^ n1055 ;
  assign n5475 = ~x416 & n1057 ;
  assign n5477 = n5458 & ~n5476 ;
  assign n5478 = n5475 & n5477 ;
  assign n5484 = n5483 ^ n5478 ;
  assign n5485 = n5476 ^ n1056 ;
  assign n5486 = n5465 & ~n5485 ;
  assign n5494 = x416 & n5486 ;
  assign n5495 = ~n5458 & n5494 ;
  assign n5496 = n5495 ^ n5458 ;
  assign n5487 = n5486 ^ n5479 ;
  assign n5488 = n5487 ^ n5458 ;
  assign n5497 = n5496 ^ n5488 ;
  assign n5498 = ~x415 & n5497 ;
  assign n5499 = ~n5484 & ~n5498 ;
  assign n5500 = ~n5474 & n5499 ;
  assign n5430 = ~x421 & n5429 ;
  assign n5433 = n5432 ^ x422 ;
  assign n5436 = n5435 ^ x422 ;
  assign n5437 = n5433 & n5436 ;
  assign n5438 = n5437 ^ x422 ;
  assign n5439 = n5430 & n5438 ;
  assign n5440 = n5439 ^ x421 ;
  assign n5453 = ~x422 & n5422 ;
  assign n5454 = ~n5432 & n5453 ;
  assign n5455 = n5454 ^ n5432 ;
  assign n5447 = n5446 ^ n5432 ;
  assign n5456 = n5455 ^ n5447 ;
  assign n5457 = n5440 & n5456 ;
  assign n5501 = n5500 ^ n5457 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1053 = n1052 ^ n1049 ;
  assign n1058 = n1057 ^ n1054 ;
  assign n5503 = n1053 & n1058 ;
  assign n8743 = n5503 ^ n5500 ;
  assign n8744 = ~n5501 & n8743 ;
  assign n8745 = n8744 ^ n5503 ;
  assign n8749 = n8748 ^ n8745 ;
  assign n8723 = ~x427 & ~x428 ;
  assign n5514 = ~x429 & ~x430 ;
  assign n1061 = x430 ^ x429 ;
  assign n5515 = n5514 ^ n1061 ;
  assign n8724 = x432 & ~n5515 ;
  assign n8725 = ~x431 & ~x432 ;
  assign n8726 = ~n5514 & ~n8725 ;
  assign n1060 = x432 ^ x431 ;
  assign n8727 = n8725 ^ n1060 ;
  assign n8728 = n5515 & n8727 ;
  assign n8729 = ~n8726 & n8728 ;
  assign n8730 = x427 & x428 ;
  assign n8731 = ~n8729 & n8730 ;
  assign n8732 = n8731 ^ x431 ;
  assign n8733 = n8724 & n8732 ;
  assign n8734 = n8733 ^ n8731 ;
  assign n8735 = n8728 ^ n8726 ;
  assign n8736 = n8735 ^ n8729 ;
  assign n8737 = ~n8734 & n8736 ;
  assign n8740 = n8723 & n8737 ;
  assign n8738 = n8737 ^ n8734 ;
  assign n8741 = n8740 ^ n8738 ;
  assign n5509 = ~x435 & ~x436 ;
  assign n8698 = ~x437 & ~x438 ;
  assign n8701 = ~n5509 & ~n8698 ;
  assign n1066 = x436 ^ x435 ;
  assign n5510 = n5509 ^ n1066 ;
  assign n8706 = n8701 ^ n5510 ;
  assign n1065 = x438 ^ x437 ;
  assign n8699 = n8698 ^ n1065 ;
  assign n8700 = n8699 ^ n5510 ;
  assign n8704 = n8700 ^ x433 ;
  assign n8707 = n8706 ^ n8704 ;
  assign n8708 = n8707 ^ x434 ;
  assign n8709 = n8708 ^ n8706 ;
  assign n8712 = n5510 ^ x434 ;
  assign n8713 = n8712 ^ n8706 ;
  assign n8714 = ~n8709 & n8713 ;
  assign n8715 = n8714 ^ n8699 ;
  assign n8716 = n8714 ^ x434 ;
  assign n8717 = n8716 ^ n5510 ;
  assign n8718 = ~n8700 & ~n8717 ;
  assign n8719 = ~n8709 & n8718 ;
  assign n8720 = n8715 & n8719 ;
  assign n8721 = n8720 ^ n8718 ;
  assign n8722 = n8721 ^ n8716 ;
  assign n8742 = n8741 ^ n8722 ;
  assign n8750 = n8749 ^ n8742 ;
  assign n5527 = x437 ^ x434 ;
  assign n5530 = n5509 ^ x437 ;
  assign n5531 = ~n5527 & n5530 ;
  assign n5528 = n5527 ^ n5509 ;
  assign n5529 = x433 & ~n5528 ;
  assign n5532 = n5531 ^ n5529 ;
  assign n5518 = x431 ^ x428 ;
  assign n5521 = n5514 ^ x431 ;
  assign n5522 = ~n5518 & n5521 ;
  assign n5519 = n5518 ^ n5514 ;
  assign n5520 = x427 & n5519 ;
  assign n5523 = n5522 ^ n5520 ;
  assign n1062 = x428 ^ x427 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n5513 = n1063 ^ x431 ;
  assign n5516 = n5515 ^ x432 ;
  assign n5517 = n5513 & n5516 ;
  assign n5524 = n5523 ^ n5517 ;
  assign n5525 = n5524 ^ x433 ;
  assign n1067 = x434 ^ x433 ;
  assign n1068 = n1067 ^ n1066 ;
  assign n5508 = n1068 ^ x437 ;
  assign n5511 = n5510 ^ x438 ;
  assign n5512 = n5508 & n5511 ;
  assign n5526 = n5525 ^ n5512 ;
  assign n5533 = n5532 ^ n5526 ;
  assign n1064 = n1063 ^ n1060 ;
  assign n1069 = n1068 ^ n1065 ;
  assign n5502 = n1064 & n1069 ;
  assign n8751 = n5524 ^ n5502 ;
  assign n8752 = n5533 & ~n8751 ;
  assign n8753 = n8752 ^ n5524 ;
  assign n8761 = n5533 ^ n5502 ;
  assign n1059 = n1058 ^ n1053 ;
  assign n1070 = n1069 ^ n1064 ;
  assign n5504 = n1059 & n1070 ;
  assign n8759 = n5504 ^ n5502 ;
  assign n8762 = n8761 ^ n8759 ;
  assign n8769 = n8762 ^ n5503 ;
  assign n8757 = n8769 ^ n5502 ;
  assign n8758 = n8757 ^ n5501 ;
  assign n8770 = n8759 ^ n8758 ;
  assign n8775 = n8770 ^ n5502 ;
  assign n8779 = ~n5533 & n8775 ;
  assign n8772 = n8762 ^ n8758 ;
  assign n8771 = n8770 ^ n5503 ;
  assign n8773 = n8772 ^ n8771 ;
  assign n8774 = n8769 & ~n8773 ;
  assign n8780 = n8779 ^ n8774 ;
  assign n8781 = n8780 ^ n8772 ;
  assign n8782 = n8779 ^ n8770 ;
  assign n8783 = n8782 ^ n8772 ;
  assign n8784 = ~n8781 & n8783 ;
  assign n8785 = n8758 & n8784 ;
  assign n8786 = n8785 ^ n8779 ;
  assign n8787 = n8786 ^ n5533 ;
  assign n8754 = n5503 ^ n5501 ;
  assign n8798 = n8787 ^ n8754 ;
  assign n8799 = n8798 ^ n5502 ;
  assign n8800 = n8799 ^ n8754 ;
  assign n12041 = n8722 & n8741 ;
  assign n12042 = n8800 & ~n12041 ;
  assign n12043 = ~n8753 & n12042 ;
  assign n12044 = n12043 ^ n12041 ;
  assign n8801 = n8800 ^ n8753 ;
  assign n12045 = n12044 ^ n8801 ;
  assign n12046 = n12045 ^ n8749 ;
  assign n12047 = n12046 ^ n12044 ;
  assign n12048 = ~n8750 & ~n12047 ;
  assign n12049 = n12048 ^ n12045 ;
  assign n1088 = x460 ^ x459 ;
  assign n5536 = x461 & x462 ;
  assign n5537 = n5536 ^ x460 ;
  assign n5538 = n1088 & ~n5537 ;
  assign n5539 = n5538 ^ x459 ;
  assign n1089 = x462 ^ x461 ;
  assign n5540 = n5536 ^ n1089 ;
  assign n5541 = x458 & n5540 ;
  assign n5542 = x459 & x460 ;
  assign n5543 = n5536 & n5542 ;
  assign n5544 = ~n5541 & ~n5543 ;
  assign n5545 = n5539 & n5544 ;
  assign n5546 = n5545 ^ n5539 ;
  assign n5563 = x457 & x458 ;
  assign n5564 = n5542 & n5563 ;
  assign n5577 = ~x462 & n5564 ;
  assign n1090 = x458 ^ x457 ;
  assign n5551 = n5543 ^ n5537 ;
  assign n5552 = n5551 ^ n5538 ;
  assign n5567 = n5552 ^ n5539 ;
  assign n5568 = n5567 ^ n5542 ;
  assign n5569 = n5568 ^ n5539 ;
  assign n5572 = x458 & n5569 ;
  assign n5573 = n5572 ^ n5539 ;
  assign n5574 = ~n1090 & n5573 ;
  assign n5575 = n5574 ^ n5539 ;
  assign n5576 = n5540 & n5575 ;
  assign n5579 = n5577 ^ n5576 ;
  assign n8814 = ~n5546 & ~n5579 ;
  assign n1079 = x444 ^ x443 ;
  assign n1078 = x442 ^ x441 ;
  assign n1080 = n1079 ^ n1078 ;
  assign n1077 = x440 ^ x439 ;
  assign n1081 = n1080 ^ n1077 ;
  assign n1074 = x450 ^ x449 ;
  assign n1073 = x448 ^ x447 ;
  assign n1075 = n1074 ^ n1073 ;
  assign n1072 = x446 ^ x445 ;
  assign n1076 = n1075 ^ n1072 ;
  assign n1082 = n1081 ^ n1076 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1092 = n1091 ^ n1088 ;
  assign n1085 = x452 ^ x451 ;
  assign n1084 = x456 ^ x455 ;
  assign n1086 = n1085 ^ n1084 ;
  assign n1083 = x454 ^ x453 ;
  assign n1087 = n1086 ^ n1083 ;
  assign n1093 = n1092 ^ n1087 ;
  assign n5718 = n1082 & n1093 ;
  assign n5587 = x453 & x454 ;
  assign n5608 = x451 & x452 ;
  assign n5609 = n5587 & n5608 ;
  assign n5610 = x455 & n5609 ;
  assign n5581 = x455 & x456 ;
  assign n5585 = n5581 ^ n1084 ;
  assign n5586 = x452 & n5585 ;
  assign n5593 = n5585 ^ x451 ;
  assign n5594 = n5593 ^ x452 ;
  assign n5595 = ~n5586 & n5594 ;
  assign n5588 = n5581 & n5587 ;
  assign n5582 = n5581 ^ x454 ;
  assign n5596 = n5588 ^ n5582 ;
  assign n5583 = n1083 & ~n5582 ;
  assign n5597 = n5596 ^ n5583 ;
  assign n5598 = n5597 ^ x452 ;
  assign n5599 = n5598 ^ n5587 ;
  assign n5600 = n5599 ^ n5597 ;
  assign n5603 = ~n1085 & ~n5600 ;
  assign n5604 = n5603 ^ n5597 ;
  assign n5605 = ~n5595 & ~n5604 ;
  assign n5606 = n5605 ^ n5597 ;
  assign n5584 = n5583 ^ x453 ;
  assign n5589 = ~n5586 & ~n5588 ;
  assign n5590 = n5584 & n5589 ;
  assign n5591 = n5590 ^ n5584 ;
  assign n5592 = ~x451 & n5591 ;
  assign n5607 = n5606 ^ n5592 ;
  assign n5611 = n5610 ^ n5607 ;
  assign n5622 = ~x456 & n5609 ;
  assign n5612 = n5597 ^ n5584 ;
  assign n5613 = n5612 ^ n5587 ;
  assign n5614 = n5613 ^ n5584 ;
  assign n5617 = x452 & n5614 ;
  assign n5618 = n5617 ^ n5584 ;
  assign n5619 = ~n1085 & n5618 ;
  assign n5620 = n5619 ^ n5584 ;
  assign n5621 = n5585 & n5620 ;
  assign n5624 = n5622 ^ n5621 ;
  assign n5625 = n5611 & ~n5624 ;
  assign n5565 = x461 & n5564 ;
  assign n5548 = n5540 ^ x457 ;
  assign n5549 = n5548 ^ x458 ;
  assign n5550 = ~n5541 & n5549 ;
  assign n5553 = n5552 ^ x458 ;
  assign n5554 = n5553 ^ n5542 ;
  assign n5555 = n5554 ^ n5552 ;
  assign n5558 = ~n1090 & ~n5555 ;
  assign n5559 = n5558 ^ n5552 ;
  assign n5560 = ~n5550 & ~n5559 ;
  assign n5561 = n5560 ^ n5552 ;
  assign n5547 = ~x457 & n5546 ;
  assign n5562 = n5561 ^ n5547 ;
  assign n5566 = n5565 ^ n5562 ;
  assign n5580 = n5566 & ~n5579 ;
  assign n5626 = n5625 ^ n5580 ;
  assign n8810 = n5718 ^ n5626 ;
  assign n5719 = n1076 & n1081 ;
  assign n5672 = x441 ^ x440 ;
  assign n5673 = ~n1078 & ~n5672 ;
  assign n5674 = x444 ^ x439 ;
  assign n5677 = ~x442 & ~n5674 ;
  assign n5678 = n5677 ^ x439 ;
  assign n5679 = n5673 & n5678 ;
  assign n5680 = ~x443 & n5679 ;
  assign n5708 = x443 ^ x442 ;
  assign n5712 = ~n1079 & ~n5708 ;
  assign n5710 = n1080 & ~n5672 ;
  assign n5681 = ~x441 & ~x442 ;
  assign n5693 = x443 & x444 ;
  assign n5695 = n5681 & ~n5693 ;
  assign n5694 = n5693 ^ n1079 ;
  assign n5696 = n5695 ^ n5694 ;
  assign n5697 = n5696 ^ x443 ;
  assign n5689 = n5681 ^ n1078 ;
  assign n5690 = n5689 ^ x444 ;
  assign n5691 = n5690 ^ n5681 ;
  assign n5692 = n5691 ^ n5689 ;
  assign n5698 = n5697 ^ n5692 ;
  assign n8836 = n5693 ^ n5689 ;
  assign n8837 = n8836 ^ n1079 ;
  assign n5700 = n8837 ^ x439 ;
  assign n5701 = ~n5698 & n5700 ;
  assign n5702 = n5694 ^ x440 ;
  assign n5703 = ~n5701 & n5702 ;
  assign n5686 = n1079 & ~n5692 ;
  assign n5687 = n5686 & n5691 ;
  assign n5688 = n5690 ^ n5687 ;
  assign n5704 = n5703 ^ n5688 ;
  assign n5705 = x440 & ~n5704 ;
  assign n5706 = n5705 ^ n5703 ;
  assign n5711 = n5710 ^ n5706 ;
  assign n5713 = n5712 ^ n5711 ;
  assign n5714 = ~x439 & n5713 ;
  assign n5715 = n5714 ^ n5706 ;
  assign n5716 = ~n5680 & ~n5715 ;
  assign n5627 = x447 ^ x446 ;
  assign n5628 = ~n1073 & ~n5627 ;
  assign n5629 = x450 ^ x445 ;
  assign n5632 = ~x448 & ~n5629 ;
  assign n5633 = n5632 ^ x445 ;
  assign n5634 = n5628 & n5633 ;
  assign n5635 = ~x449 & n5634 ;
  assign n5662 = x449 ^ x448 ;
  assign n5667 = ~n1074 & ~n5662 ;
  assign n5665 = n1075 & ~n5627 ;
  assign n5648 = x449 & x450 ;
  assign n5650 = n5648 ^ n1074 ;
  assign n5636 = ~x447 & ~x448 ;
  assign n5649 = n5636 & ~n5648 ;
  assign n5651 = n5650 ^ n5649 ;
  assign n5652 = n5651 ^ x449 ;
  assign n5644 = n5636 ^ n1073 ;
  assign n5645 = n5644 ^ x450 ;
  assign n5646 = n5645 ^ n5636 ;
  assign n5647 = n5646 ^ n5644 ;
  assign n5653 = n5652 ^ n5647 ;
  assign n8824 = n5648 ^ n5644 ;
  assign n8825 = n8824 ^ n1074 ;
  assign n5655 = n8825 ^ x445 ;
  assign n5656 = ~n5653 & n5655 ;
  assign n5657 = n5650 ^ x446 ;
  assign n5658 = ~n5656 & n5657 ;
  assign n5641 = n1074 & ~n5647 ;
  assign n5642 = n5641 & n5646 ;
  assign n5643 = n5645 ^ n5642 ;
  assign n5659 = n5658 ^ n5643 ;
  assign n5660 = x446 & ~n5659 ;
  assign n5661 = n5660 ^ n5658 ;
  assign n5666 = n5665 ^ n5661 ;
  assign n5668 = n5667 ^ n5666 ;
  assign n5669 = ~x445 & n5668 ;
  assign n5670 = n5669 ^ n5661 ;
  assign n5671 = ~n5635 & ~n5670 ;
  assign n5717 = n5716 ^ n5671 ;
  assign n8808 = n5719 ^ n5717 ;
  assign n8811 = n8808 ^ n5626 ;
  assign n8812 = ~n8810 & n8811 ;
  assign n5720 = n1087 & n1092 ;
  assign n8809 = ~n5720 & n8808 ;
  assign n8813 = n8812 ^ n8809 ;
  assign n8815 = n8814 ^ n8813 ;
  assign n8819 = ~n5591 & ~n5624 ;
  assign n12059 = n8819 ^ n8814 ;
  assign n12060 = n8815 & n12059 ;
  assign n12061 = n12060 ^ n8819 ;
  assign n8840 = ~x440 & n5694 ;
  assign n8841 = n8840 ^ n5694 ;
  assign n8842 = n5695 ^ n1078 ;
  assign n8843 = n8841 & ~n8842 ;
  assign n8844 = n8843 ^ n8836 ;
  assign n8845 = n8840 ^ n1079 ;
  assign n8846 = n8845 ^ n8843 ;
  assign n8847 = ~n8844 & ~n8846 ;
  assign n8848 = n8847 ^ n5689 ;
  assign n8849 = x439 & n8848 ;
  assign n8850 = n5706 & n8849 ;
  assign n8851 = n8850 ^ n8848 ;
  assign n8852 = n8851 ^ n5644 ;
  assign n8828 = ~x446 & n5650 ;
  assign n8829 = n8828 ^ n5650 ;
  assign n8830 = n5649 ^ n1073 ;
  assign n8831 = n8829 & ~n8830 ;
  assign n8832 = n8831 ^ n8824 ;
  assign n8833 = n8828 ^ n1074 ;
  assign n8834 = n8833 ^ n8831 ;
  assign n8835 = ~n8832 & ~n8834 ;
  assign n8853 = n8852 ^ n8835 ;
  assign n8854 = n8853 ^ n8851 ;
  assign n8855 = x445 & n5661 ;
  assign n8856 = n8854 & n8855 ;
  assign n8857 = n8856 ^ n8853 ;
  assign n8821 = n5719 ^ n5716 ;
  assign n8822 = ~n5717 & n8821 ;
  assign n8823 = n8822 ^ n5719 ;
  assign n8858 = n8857 ^ n8823 ;
  assign n8816 = n5720 ^ n5625 ;
  assign n8817 = ~n5626 & n8816 ;
  assign n8818 = n8817 ^ n5720 ;
  assign n8820 = n8819 ^ n8818 ;
  assign n8859 = n8858 ^ n8820 ;
  assign n8860 = n8859 ^ n8815 ;
  assign n12062 = n8860 ^ n8818 ;
  assign n12063 = n8860 ^ n8858 ;
  assign n12064 = ~n12062 & ~n12063 ;
  assign n12065 = n12064 ^ n8860 ;
  assign n12066 = n12061 & n12065 ;
  assign n12067 = n8858 & ~n8860 ;
  assign n12068 = ~n12061 & n12067 ;
  assign n12070 = n8851 ^ n8823 ;
  assign n12071 = n8857 & ~n12070 ;
  assign n12072 = n12071 ^ n8851 ;
  assign n12645 = ~n12068 & n12072 ;
  assign n12646 = ~n12066 & n12645 ;
  assign n12647 = n12646 ^ n12066 ;
  assign n12649 = n12647 ^ n12044 ;
  assign n12050 = n8747 ^ n8745 ;
  assign n12051 = n8748 & ~n12050 ;
  assign n12052 = n12051 ^ n8747 ;
  assign n12648 = n12647 ^ n12052 ;
  assign n12650 = n12649 ^ n12648 ;
  assign n12651 = ~n12049 & ~n12650 ;
  assign n12652 = n12651 ^ n12649 ;
  assign n1071 = n1070 ^ n1059 ;
  assign n1094 = n1093 ^ n1082 ;
  assign n5420 = n1071 & n1094 ;
  assign n5535 = n8758 ^ n5420 ;
  assign n8802 = n8801 ^ n8750 ;
  assign n5721 = n5720 ^ n5719 ;
  assign n5722 = n5721 ^ n5718 ;
  assign n5723 = n5722 ^ n5717 ;
  assign n5724 = n5723 ^ n5626 ;
  assign n8803 = n8802 ^ n5724 ;
  assign n8804 = n8803 ^ n8758 ;
  assign n8805 = n8804 ^ n8802 ;
  assign n8806 = ~n5535 & n8805 ;
  assign n8807 = n8806 ^ n8803 ;
  assign n12053 = n12052 ^ n12049 ;
  assign n12055 = n12053 ^ n8802 ;
  assign n12054 = n12053 ^ n8860 ;
  assign n12056 = n12055 ^ n12054 ;
  assign n12057 = ~n8807 & ~n12056 ;
  assign n12058 = n12057 ^ n12055 ;
  assign n12069 = n12068 ^ n12066 ;
  assign n12073 = n12072 ^ n12069 ;
  assign n12653 = n12073 ^ n12053 ;
  assign n12654 = ~n12058 & n12653 ;
  assign n12655 = n12654 ^ n12053 ;
  assign n12902 = n12655 ^ n12647 ;
  assign n12903 = ~n12652 & ~n12902 ;
  assign n12904 = n12903 ^ n12647 ;
  assign n12908 = n12907 ^ n12904 ;
  assign n12674 = n12673 ^ n12670 ;
  assign n12656 = n12655 ^ n12652 ;
  assign n12675 = n12674 ^ n12656 ;
  assign n12074 = n12073 ^ n12058 ;
  assign n6031 = n6030 ^ n5891 ;
  assign n5725 = n5724 ^ n5535 ;
  assign n6032 = n6031 ^ n5725 ;
  assign n8861 = n8860 ^ n8807 ;
  assign n8862 = n8861 ^ n5725 ;
  assign n1048 = n1047 ^ n1024 ;
  assign n1095 = n1094 ^ n1071 ;
  assign n5417 = n1048 & n1095 ;
  assign n8863 = n8862 ^ n5417 ;
  assign n8864 = n8863 ^ n8861 ;
  assign n8865 = ~n6032 & n8864 ;
  assign n8866 = n8865 ^ n8862 ;
  assign n8971 = n8970 ^ n8917 ;
  assign n12038 = n8971 ^ n8861 ;
  assign n12039 = ~n8866 & n12038 ;
  assign n12040 = n12039 ^ n8861 ;
  assign n12075 = n12074 ^ n12040 ;
  assign n12115 = n12114 ^ n12099 ;
  assign n12642 = n12115 ^ n12040 ;
  assign n12643 = ~n12075 & n12642 ;
  assign n12644 = n12643 ^ n12115 ;
  assign n12909 = n12674 ^ n12644 ;
  assign n12910 = n12675 & n12909 ;
  assign n12911 = n12910 ^ n12674 ;
  assign n13149 = n12911 ^ n12907 ;
  assign n13150 = ~n12908 & n13149 ;
  assign n13151 = n13150 ^ n12911 ;
  assign n8972 = n8971 ^ n8866 ;
  assign n1096 = n1095 ^ n1048 ;
  assign n1185 = x284 ^ x283 ;
  assign n1184 = x286 ^ x285 ;
  assign n1186 = n1185 ^ n1184 ;
  assign n1183 = x288 ^ x287 ;
  assign n1187 = n1186 ^ n1183 ;
  assign n1180 = x276 ^ x275 ;
  assign n1179 = x274 ^ x273 ;
  assign n1181 = n1180 ^ n1179 ;
  assign n1178 = x272 ^ x271 ;
  assign n1182 = n1181 ^ n1178 ;
  assign n1188 = n1187 ^ n1182 ;
  assign n1174 = x278 ^ x277 ;
  assign n1173 = x282 ^ x281 ;
  assign n1175 = n1174 ^ n1173 ;
  assign n1172 = x280 ^ x279 ;
  assign n1176 = n1175 ^ n1172 ;
  assign n1169 = x290 ^ x289 ;
  assign n1168 = x292 ^ x291 ;
  assign n1170 = n1169 ^ n1168 ;
  assign n1167 = x294 ^ x293 ;
  assign n1171 = n1170 ^ n1167 ;
  assign n1177 = n1176 ^ n1171 ;
  assign n1189 = n1188 ^ n1177 ;
  assign n1163 = x306 ^ x305 ;
  assign n1161 = x304 ^ x303 ;
  assign n1160 = x302 ^ x301 ;
  assign n1162 = n1161 ^ n1160 ;
  assign n1164 = n1163 ^ n1162 ;
  assign n6062 = x299 ^ x297 ;
  assign n6074 = n6062 ^ x298 ;
  assign n6075 = n6074 ^ x300 ;
  assign n1155 = x296 ^ x295 ;
  assign n1159 = n6075 ^ n1155 ;
  assign n1165 = n1164 ^ n1159 ;
  assign n1152 = x318 ^ x317 ;
  assign n1150 = x316 ^ x315 ;
  assign n1149 = x314 ^ x313 ;
  assign n1151 = n1150 ^ n1149 ;
  assign n1153 = n1152 ^ n1151 ;
  assign n1146 = x312 ^ x311 ;
  assign n1145 = x310 ^ x309 ;
  assign n1147 = n1146 ^ n1145 ;
  assign n1144 = x308 ^ x307 ;
  assign n1148 = n1147 ^ n1144 ;
  assign n1154 = n1153 ^ n1148 ;
  assign n1166 = n1165 ^ n1154 ;
  assign n1190 = n1189 ^ n1166 ;
  assign n1138 = x356 ^ x355 ;
  assign n1137 = x358 ^ x357 ;
  assign n1139 = n1138 ^ n1137 ;
  assign n1136 = x360 ^ x359 ;
  assign n1140 = n1139 ^ n1136 ;
  assign n1133 = x362 ^ x361 ;
  assign n1132 = x364 ^ x363 ;
  assign n1134 = n1133 ^ n1132 ;
  assign n1131 = x366 ^ x365 ;
  assign n1135 = n1134 ^ n1131 ;
  assign n1141 = n1140 ^ n1135 ;
  assign n1128 = x348 ^ x347 ;
  assign n1126 = x346 ^ x345 ;
  assign n1125 = x344 ^ x343 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1129 = n1128 ^ n1127 ;
  assign n1123 = x354 ^ x353 ;
  assign n1121 = x352 ^ x351 ;
  assign n1120 = x350 ^ x349 ;
  assign n1122 = n1121 ^ n1120 ;
  assign n1124 = n1123 ^ n1122 ;
  assign n1130 = n1129 ^ n1124 ;
  assign n1142 = n1141 ^ n1130 ;
  assign n1116 = x336 ^ x335 ;
  assign n1114 = x334 ^ x333 ;
  assign n1113 = x332 ^ x331 ;
  assign n1115 = n1114 ^ n1113 ;
  assign n1117 = n1116 ^ n1115 ;
  assign n1111 = x340 ^ x339 ;
  assign n1109 = x342 ^ x341 ;
  assign n1108 = x338 ^ x337 ;
  assign n1110 = n1109 ^ n1108 ;
  assign n1112 = n1111 ^ n1110 ;
  assign n1118 = n1117 ^ n1112 ;
  assign n1104 = x320 ^ x319 ;
  assign n1103 = x322 ^ x321 ;
  assign n1105 = n1104 ^ n1103 ;
  assign n1102 = x324 ^ x323 ;
  assign n1106 = n1105 ^ n1102 ;
  assign n1100 = x330 ^ x329 ;
  assign n1098 = x328 ^ x327 ;
  assign n1097 = x326 ^ x325 ;
  assign n1099 = n1098 ^ n1097 ;
  assign n1101 = n1100 ^ n1099 ;
  assign n1107 = n1106 ^ n1101 ;
  assign n1119 = n1118 ^ n1107 ;
  assign n1143 = n1142 ^ n1119 ;
  assign n1191 = n1190 ^ n1143 ;
  assign n5418 = n1096 & n1191 ;
  assign n5419 = n5418 ^ n5417 ;
  assign n6033 = n6032 ^ n5419 ;
  assign n6367 = ~x291 & ~x292 ;
  assign n6365 = ~x293 & ~x294 ;
  assign n6376 = n6367 ^ n6365 ;
  assign n6375 = n6365 & n6367 ;
  assign n6377 = n6376 ^ n6375 ;
  assign n6366 = n6365 ^ n1167 ;
  assign n6368 = n6367 ^ n1168 ;
  assign n6370 = n6366 & n6368 ;
  assign n6378 = n6377 ^ n6370 ;
  assign n6386 = n6365 ^ n1169 ;
  assign n6387 = n6386 ^ n6367 ;
  assign n6388 = ~n6375 & ~n6387 ;
  assign n6389 = ~n6378 & ~n6388 ;
  assign n6369 = n6368 ^ n6366 ;
  assign n6371 = n6370 ^ n6369 ;
  assign n6372 = x289 & x290 ;
  assign n6373 = n6371 & n6372 ;
  assign n6374 = n6373 ^ n6370 ;
  assign n6379 = n6377 ^ n1169 ;
  assign n6380 = ~n6378 & n6379 ;
  assign n6381 = ~n6374 & n6380 ;
  assign n6382 = n6381 ^ n6373 ;
  assign n6383 = n6371 & ~n6382 ;
  assign n6384 = n6383 ^ n6382 ;
  assign n6385 = n6384 ^ n6372 ;
  assign n6390 = n6389 ^ n6385 ;
  assign n6341 = ~x285 & ~x286 ;
  assign n6339 = ~x287 & ~x288 ;
  assign n6350 = n6341 ^ n6339 ;
  assign n6349 = n6339 & n6341 ;
  assign n6351 = n6350 ^ n6349 ;
  assign n6340 = n6339 ^ n1183 ;
  assign n6342 = n6341 ^ n1184 ;
  assign n6344 = n6340 & n6342 ;
  assign n6352 = n6351 ^ n6344 ;
  assign n6360 = n6339 ^ n1185 ;
  assign n6361 = n6360 ^ n6341 ;
  assign n6362 = ~n6349 & ~n6361 ;
  assign n6363 = ~n6352 & ~n6362 ;
  assign n6343 = n6342 ^ n6340 ;
  assign n6345 = n6344 ^ n6343 ;
  assign n6346 = x283 & x284 ;
  assign n6347 = n6345 & n6346 ;
  assign n6348 = n6347 ^ n1185 ;
  assign n6353 = n6344 ^ n1185 ;
  assign n6354 = ~n6352 & n6353 ;
  assign n6355 = n6348 & n6354 ;
  assign n6356 = n6355 ^ n6347 ;
  assign n6357 = n6345 & ~n6356 ;
  assign n6358 = n6357 ^ n6356 ;
  assign n6359 = n6358 ^ n6346 ;
  assign n6364 = n6363 ^ n6359 ;
  assign n6391 = n6390 ^ n6364 ;
  assign n6333 = n1187 ^ n1171 ;
  assign n6336 = n6333 ^ n1182 ;
  assign n6337 = ~n1176 & n6336 ;
  assign n6334 = n1182 ^ n1171 ;
  assign n6335 = ~n6333 & ~n6334 ;
  assign n6338 = n6337 ^ n6335 ;
  assign n6392 = n6391 ^ n6338 ;
  assign n6284 = x276 ^ x272 ;
  assign n6283 = x276 ^ x274 ;
  assign n6285 = n6284 ^ n6283 ;
  assign n6286 = n6285 ^ x276 ;
  assign n6288 = x272 & n6286 ;
  assign n6289 = n6288 ^ x276 ;
  assign n6317 = x273 ^ x272 ;
  assign n6294 = n6317 ^ n1178 ;
  assign n6295 = n6285 ^ n1178 ;
  assign n6296 = n6295 ^ n6284 ;
  assign n6297 = n6296 ^ x276 ;
  assign n6298 = ~n6294 & n6297 ;
  assign n6301 = n6298 ^ x274 ;
  assign n6302 = ~n6289 & ~n6301 ;
  assign n6305 = ~x275 & n6302 ;
  assign n6315 = n6284 ^ n1179 ;
  assign n6292 = x276 ^ x273 ;
  assign n6318 = ~n6292 & ~n6317 ;
  assign n6321 = n6318 ^ x274 ;
  assign n6322 = n6321 ^ n6284 ;
  assign n6316 = x275 ^ x274 ;
  assign n6323 = n6322 ^ n6316 ;
  assign n6324 = n6318 & n6323 ;
  assign n6325 = n6324 ^ n6316 ;
  assign n6326 = ~n6315 & n6325 ;
  assign n6327 = n6326 ^ n6321 ;
  assign n6306 = ~x275 & ~x276 ;
  assign n6307 = n6306 ^ n1180 ;
  assign n6308 = n6307 ^ x274 ;
  assign n6309 = x272 & ~n6306 ;
  assign n6312 = n6309 ^ n6307 ;
  assign n6313 = n6308 & n6312 ;
  assign n6310 = n6309 ^ n6308 ;
  assign n6311 = x273 & n6310 ;
  assign n6314 = n6313 ^ n6311 ;
  assign n6328 = n6327 ^ n6314 ;
  assign n6329 = ~x271 & n6328 ;
  assign n6330 = n6329 ^ n6327 ;
  assign n6331 = ~n6305 & ~n6330 ;
  assign n6252 = ~x281 & ~x282 ;
  assign n6253 = n6252 ^ n1173 ;
  assign n6245 = ~x279 & ~x280 ;
  assign n6254 = n6245 ^ n1172 ;
  assign n6255 = ~n6253 & ~n6254 ;
  assign n6246 = x281 ^ x278 ;
  assign n6249 = n1173 & n6246 ;
  assign n6250 = n6249 ^ x281 ;
  assign n6251 = n6245 & ~n6250 ;
  assign n6256 = n6255 ^ n6251 ;
  assign n6257 = ~x277 & n6256 ;
  assign n6261 = x277 & x278 ;
  assign n6266 = n6261 ^ n1174 ;
  assign n6267 = n6266 ^ x280 ;
  assign n6268 = n6266 ^ x279 ;
  assign n6269 = ~n6267 & ~n6268 ;
  assign n6270 = n6269 ^ n6266 ;
  assign n6271 = n6261 ^ n6253 ;
  assign n6272 = n6267 ^ n6261 ;
  assign n6273 = n6272 ^ n6268 ;
  assign n6274 = ~n6271 & n6273 ;
  assign n6275 = n6274 ^ n6266 ;
  assign n6276 = n6270 & n6275 ;
  assign n6277 = n6276 ^ n6266 ;
  assign n6278 = n6277 ^ n6261 ;
  assign n6279 = ~n6252 & n6278 ;
  assign n6262 = n6253 & ~n6254 ;
  assign n6263 = ~n6261 & n6262 ;
  assign n6264 = n6263 ^ n6254 ;
  assign n6265 = n6264 ^ n6255 ;
  assign n6280 = n6279 ^ n6265 ;
  assign n6258 = ~x278 & n1176 ;
  assign n6259 = n6252 & n6254 ;
  assign n6260 = n6258 & n6259 ;
  assign n6281 = n6280 ^ n6260 ;
  assign n6282 = ~n6257 & n6281 ;
  assign n6332 = n6331 ^ n6282 ;
  assign n6393 = n6392 ^ n6332 ;
  assign n6187 = x312 ^ x308 ;
  assign n6186 = x312 ^ x310 ;
  assign n6188 = n6187 ^ n6186 ;
  assign n6189 = n6188 ^ x312 ;
  assign n6191 = x308 & n6189 ;
  assign n6192 = n6191 ^ x312 ;
  assign n6195 = x312 ^ x309 ;
  assign n6196 = n6195 ^ n6187 ;
  assign n6197 = n6196 ^ n1144 ;
  assign n6198 = n6188 ^ n1144 ;
  assign n6199 = n6198 ^ n6187 ;
  assign n6200 = n6199 ^ x312 ;
  assign n6201 = ~n6197 & n6200 ;
  assign n6204 = n6201 ^ x310 ;
  assign n6205 = ~n6192 & ~n6204 ;
  assign n6208 = ~x311 & n6205 ;
  assign n6220 = x311 ^ x308 ;
  assign n6221 = n6220 ^ x310 ;
  assign n6222 = n6221 ^ x312 ;
  assign n6218 = x311 ^ x309 ;
  assign n6223 = n6222 ^ n6218 ;
  assign n6229 = ~n6186 & ~n6188 ;
  assign n6233 = n6229 ^ x309 ;
  assign n6234 = n6233 ^ n6218 ;
  assign n6235 = n6229 & n6234 ;
  assign n6236 = n6235 ^ n6218 ;
  assign n6237 = ~n6223 & n6236 ;
  assign n6238 = n6237 ^ n6233 ;
  assign n6209 = ~x311 & ~x312 ;
  assign n6210 = n6209 ^ n1146 ;
  assign n6211 = n6210 ^ x310 ;
  assign n6212 = x308 & ~n6209 ;
  assign n6215 = n6212 ^ n6210 ;
  assign n6216 = n6211 & n6215 ;
  assign n6213 = n6212 ^ n6211 ;
  assign n6214 = x309 & n6213 ;
  assign n6217 = n6216 ^ n6214 ;
  assign n6239 = n6238 ^ n6217 ;
  assign n6240 = ~x307 & n6239 ;
  assign n6241 = n6240 ^ n6238 ;
  assign n6242 = ~n6208 & ~n6241 ;
  assign n6139 = x315 & x316 ;
  assign n6140 = n6139 ^ x314 ;
  assign n6143 = n1150 ^ x313 ;
  assign n6144 = ~x318 & n6143 ;
  assign n6145 = n6144 ^ x313 ;
  assign n6146 = ~n6139 & n6145 ;
  assign n6147 = n6146 ^ x313 ;
  assign n6148 = ~n6140 & n6147 ;
  assign n6149 = ~x317 & n6148 ;
  assign n6150 = x317 & x318 ;
  assign n6151 = n6150 ^ n1152 ;
  assign n6156 = n6139 & n6150 ;
  assign n6152 = n6150 ^ x316 ;
  assign n6157 = n6156 ^ n6152 ;
  assign n6153 = n1150 & ~n6152 ;
  assign n6158 = n6157 ^ n6153 ;
  assign n6154 = n6153 ^ x315 ;
  assign n6155 = n6154 ^ n6139 ;
  assign n6159 = n6158 ^ n6155 ;
  assign n6160 = n6159 ^ n6154 ;
  assign n6163 = x314 & n6160 ;
  assign n6164 = n6163 ^ n6154 ;
  assign n6165 = ~n1149 & n6164 ;
  assign n6166 = n6165 ^ n6154 ;
  assign n6167 = n6151 & n6166 ;
  assign n6168 = x313 & x314 ;
  assign n6169 = ~x318 & n6139 ;
  assign n6170 = n6168 & n6169 ;
  assign n6171 = ~n6167 & ~n6170 ;
  assign n6172 = ~x313 & n6171 ;
  assign n6173 = x314 & n6151 ;
  assign n6181 = ~n6158 & ~n6173 ;
  assign n6174 = n6154 & ~n6156 ;
  assign n6175 = ~n6173 & n6174 ;
  assign n6176 = n6175 ^ n6154 ;
  assign n6182 = n6181 ^ n6176 ;
  assign n6183 = n6172 & n6182 ;
  assign n6184 = n6183 ^ n6171 ;
  assign n6185 = ~n6149 & n6184 ;
  assign n6243 = n6242 ^ n6185 ;
  assign n6045 = x299 & x300 ;
  assign n6048 = ~x297 & ~x298 ;
  assign n1157 = x298 ^ x297 ;
  assign n6056 = n6048 ^ n1157 ;
  assign n6130 = ~n6045 & n6056 ;
  assign n6064 = x299 ^ x296 ;
  assign n6065 = n6064 ^ x298 ;
  assign n6066 = n6065 ^ x300 ;
  assign n6067 = n6066 ^ n6062 ;
  assign n6068 = n6067 ^ x300 ;
  assign n6069 = n6068 ^ x299 ;
  assign n6070 = n6069 ^ n6062 ;
  assign n6076 = n6075 ^ n6062 ;
  assign n6077 = ~n6070 & ~n6076 ;
  assign n6078 = ~x299 & n6077 ;
  assign n6081 = n6078 ^ n6077 ;
  assign n6079 = n6078 ^ n6062 ;
  assign n6080 = n6067 & n6079 ;
  assign n6082 = n6081 ^ n6080 ;
  assign n6083 = n6082 ^ x299 ;
  assign n6132 = x295 & n6083 ;
  assign n6131 = n6083 ^ x295 ;
  assign n6133 = n6132 ^ n6131 ;
  assign n6134 = n6130 & ~n6133 ;
  assign n6091 = x305 ^ x304 ;
  assign n6095 = ~n1163 & ~n6091 ;
  assign n6090 = x303 ^ x302 ;
  assign n6092 = n6091 ^ x303 ;
  assign n6093 = n6092 ^ x306 ;
  assign n6094 = ~n6090 & n6093 ;
  assign n6096 = n6095 ^ n6094 ;
  assign n6097 = ~x301 & n6096 ;
  assign n6098 = ~n1161 & ~n6090 ;
  assign n6099 = x306 ^ x301 ;
  assign n6102 = ~x304 & ~n6099 ;
  assign n6103 = n6102 ^ x301 ;
  assign n6104 = n6098 & n6103 ;
  assign n6105 = ~x305 & n6104 ;
  assign n6106 = ~x303 & ~x304 ;
  assign n6109 = n6106 ^ n1161 ;
  assign n6110 = x301 & x302 ;
  assign n6111 = x306 & n6110 ;
  assign n6112 = ~n6109 & n6111 ;
  assign n6113 = n6112 ^ n6110 ;
  assign n6107 = ~x305 & ~x306 ;
  assign n6108 = ~n6106 & ~n6107 ;
  assign n6114 = n6113 ^ n6108 ;
  assign n6115 = n6107 ^ n1163 ;
  assign n6120 = n6109 & n6115 ;
  assign n6121 = n6120 ^ n6108 ;
  assign n6122 = n6114 & n6121 ;
  assign n6123 = n6122 ^ n6113 ;
  assign n6124 = ~n1160 & n6123 ;
  assign n6125 = n6122 & n6124 ;
  assign n6126 = n6125 ^ n6123 ;
  assign n6127 = ~n6105 & ~n6126 ;
  assign n6128 = ~n6097 & n6127 ;
  assign n6129 = n6128 ^ n6083 ;
  assign n6135 = n6134 ^ n6129 ;
  assign n6057 = n6056 ^ n6045 ;
  assign n1156 = x300 ^ x299 ;
  assign n6046 = n6045 ^ n1156 ;
  assign n6047 = n6046 ^ x296 ;
  assign n6049 = n6048 ^ n6047 ;
  assign n6058 = n6049 ^ n6045 ;
  assign n6051 = ~n6046 & n6048 ;
  assign n6050 = n6048 ^ n6046 ;
  assign n6052 = n6051 ^ n6050 ;
  assign n6053 = ~n6049 & ~n6052 ;
  assign n6059 = n6058 ^ n6053 ;
  assign n6060 = ~n6057 & n6059 ;
  assign n6061 = n6060 ^ n6056 ;
  assign n6087 = ~x295 & ~n6082 ;
  assign n6088 = n6087 ^ x299 ;
  assign n6089 = ~n6061 & ~n6088 ;
  assign n6136 = n6135 ^ n6089 ;
  assign n6054 = n6051 ^ x295 ;
  assign n6055 = ~n6053 & ~n6054 ;
  assign n6137 = n6136 ^ n6055 ;
  assign n6042 = n1159 & n1164 ;
  assign n6040 = n1148 & n1153 ;
  assign n8652 = n6042 ^ n6040 ;
  assign n6037 = n1159 ^ n1154 ;
  assign n6038 = n1165 & ~n6037 ;
  assign n6039 = n6038 ^ n1164 ;
  assign n8653 = n8652 ^ n6039 ;
  assign n6044 = n8653 ^ n6042 ;
  assign n6138 = n6137 ^ n6044 ;
  assign n6244 = n6243 ^ n6138 ;
  assign n6394 = n6393 ^ n6244 ;
  assign n6035 = n1166 & n1189 ;
  assign n8473 = n6394 ^ n6035 ;
  assign n6034 = n1143 & n1190 ;
  assign n8474 = n8473 ^ n6034 ;
  assign n6657 = x329 ^ x328 ;
  assign n6661 = ~n1100 & ~n6657 ;
  assign n6656 = x327 ^ x326 ;
  assign n6658 = n6657 ^ x327 ;
  assign n6659 = n6658 ^ x330 ;
  assign n6660 = ~n6656 & n6659 ;
  assign n6662 = n6661 ^ n6660 ;
  assign n6663 = ~x325 & n6662 ;
  assign n6664 = ~n1098 & ~n6656 ;
  assign n6665 = x330 ^ x325 ;
  assign n6668 = ~x328 & ~n6665 ;
  assign n6669 = n6668 ^ x325 ;
  assign n6670 = n6664 & n6669 ;
  assign n6671 = ~x329 & n6670 ;
  assign n6672 = ~x327 & ~x328 ;
  assign n6675 = n6672 ^ n1098 ;
  assign n6676 = x325 & x326 ;
  assign n6677 = x330 & n6676 ;
  assign n6678 = ~n6675 & n6677 ;
  assign n6679 = n6678 ^ n6676 ;
  assign n6673 = ~x329 & ~x330 ;
  assign n6674 = ~n6672 & ~n6673 ;
  assign n6680 = n6679 ^ n6674 ;
  assign n6681 = n6673 ^ n1100 ;
  assign n6686 = n6675 & n6681 ;
  assign n6687 = n6686 ^ n6674 ;
  assign n6688 = n6680 & n6687 ;
  assign n6689 = n6688 ^ n6679 ;
  assign n6690 = ~n1097 & n6689 ;
  assign n6691 = n6688 & n6690 ;
  assign n6692 = n6691 ^ n6689 ;
  assign n6693 = ~n6671 & ~n6692 ;
  assign n6694 = ~n6663 & n6693 ;
  assign n6655 = n1101 & n1106 ;
  assign n6695 = n6694 ^ n6655 ;
  assign n6617 = x323 ^ x322 ;
  assign n6621 = ~n1102 & ~n6617 ;
  assign n6616 = x321 ^ x320 ;
  assign n6618 = n6617 ^ x321 ;
  assign n6619 = n6618 ^ x324 ;
  assign n6620 = ~n6616 & n6619 ;
  assign n6622 = n6621 ^ n6620 ;
  assign n6623 = ~x319 & n6622 ;
  assign n6624 = ~n1103 & ~n6616 ;
  assign n6625 = x324 ^ x319 ;
  assign n6628 = ~x322 & ~n6625 ;
  assign n6629 = n6628 ^ x319 ;
  assign n6630 = n6624 & n6629 ;
  assign n6631 = ~x323 & n6630 ;
  assign n6632 = ~x321 & ~x322 ;
  assign n6635 = n6632 ^ n1103 ;
  assign n6636 = x319 & x320 ;
  assign n6637 = x324 & n6636 ;
  assign n6638 = ~n6635 & n6637 ;
  assign n6639 = n6638 ^ n6636 ;
  assign n6633 = ~x323 & ~x324 ;
  assign n6634 = ~n6632 & ~n6633 ;
  assign n6640 = n6639 ^ n6634 ;
  assign n6641 = n6633 ^ n1102 ;
  assign n6646 = n6635 & n6641 ;
  assign n6647 = n6646 ^ n6634 ;
  assign n6648 = n6640 & n6647 ;
  assign n6649 = n6648 ^ n6639 ;
  assign n6650 = ~n1104 & n6649 ;
  assign n6651 = n6648 & n6650 ;
  assign n6652 = n6651 ^ n6649 ;
  assign n6653 = ~n6631 & ~n6652 ;
  assign n6654 = ~n6623 & n6653 ;
  assign n6696 = n6695 ^ n6654 ;
  assign n6613 = n1112 & n1117 ;
  assign n6593 = x339 & x340 ;
  assign n6595 = n6593 ^ n1111 ;
  assign n6592 = x341 & x342 ;
  assign n6596 = n6592 ^ n1109 ;
  assign n6597 = n6595 & n6596 ;
  assign n6606 = n6597 ^ x338 ;
  assign n6594 = n6593 ^ n6592 ;
  assign n6598 = n6597 ^ n6593 ;
  assign n6599 = n6598 ^ n1108 ;
  assign n6600 = ~n6594 & ~n6599 ;
  assign n6601 = n6600 ^ n6597 ;
  assign n6602 = n1111 ^ n1109 ;
  assign n6603 = n6602 ^ n6594 ;
  assign n6604 = n6603 ^ n6600 ;
  assign n6605 = ~n6601 & ~n6604 ;
  assign n6607 = n6606 ^ n6605 ;
  assign n6611 = n1108 & ~n6607 ;
  assign n6609 = n6600 ^ x337 ;
  assign n6612 = n6611 ^ n6609 ;
  assign n6614 = n6613 ^ n6612 ;
  assign n6572 = x335 & x336 ;
  assign n6574 = n6572 ^ n1116 ;
  assign n6571 = x333 & x334 ;
  assign n6575 = n6571 ^ n1114 ;
  assign n6576 = n6574 & n6575 ;
  assign n6585 = n6576 ^ x332 ;
  assign n6573 = n6572 ^ n6571 ;
  assign n6577 = n6576 ^ n6572 ;
  assign n6578 = n6577 ^ n1113 ;
  assign n6579 = ~n6573 & ~n6578 ;
  assign n6580 = n6579 ^ n6576 ;
  assign n6581 = n1116 ^ n1114 ;
  assign n6582 = n6581 ^ n6573 ;
  assign n6583 = n6582 ^ n6579 ;
  assign n6584 = ~n6580 & ~n6583 ;
  assign n6586 = n6585 ^ n6584 ;
  assign n6590 = n1113 & ~n6586 ;
  assign n6588 = n6579 ^ x331 ;
  assign n6591 = n6590 ^ n6588 ;
  assign n6615 = n6614 ^ n6591 ;
  assign n6697 = n6696 ^ n6615 ;
  assign n6521 = x345 & x346 ;
  assign n6522 = n6521 ^ x344 ;
  assign n6525 = n1126 ^ x343 ;
  assign n6526 = ~x348 & n6525 ;
  assign n6527 = n6526 ^ x343 ;
  assign n6528 = ~n6521 & n6527 ;
  assign n6529 = n6528 ^ x343 ;
  assign n6530 = ~n6522 & n6529 ;
  assign n6531 = ~x347 & n6530 ;
  assign n6532 = x347 & x348 ;
  assign n6533 = n6532 ^ n1128 ;
  assign n6538 = n6521 & n6532 ;
  assign n6534 = n6532 ^ x346 ;
  assign n6539 = n6538 ^ n6534 ;
  assign n6535 = n1126 & ~n6534 ;
  assign n6540 = n6539 ^ n6535 ;
  assign n6536 = n6535 ^ x345 ;
  assign n6537 = n6536 ^ n6521 ;
  assign n6541 = n6540 ^ n6537 ;
  assign n6542 = n6541 ^ n6536 ;
  assign n6545 = x344 & n6542 ;
  assign n6546 = n6545 ^ n6536 ;
  assign n6547 = ~n1125 & n6546 ;
  assign n6548 = n6547 ^ n6536 ;
  assign n6549 = n6533 & n6548 ;
  assign n6550 = x343 & x344 ;
  assign n6551 = ~x348 & n6521 ;
  assign n6552 = n6550 & n6551 ;
  assign n6553 = ~n6549 & ~n6552 ;
  assign n6554 = ~x343 & n6553 ;
  assign n6555 = x344 & n6533 ;
  assign n6563 = ~n6540 & ~n6555 ;
  assign n6556 = n6536 & ~n6538 ;
  assign n6557 = ~n6555 & n6556 ;
  assign n6558 = n6557 ^ n6536 ;
  assign n6564 = n6563 ^ n6558 ;
  assign n6565 = n6554 & n6564 ;
  assign n6566 = n6565 ^ n6553 ;
  assign n6567 = ~n6531 & n6566 ;
  assign n6519 = n1124 & n1129 ;
  assign n6482 = ~x349 & ~n1121 ;
  assign n6484 = ~x351 & ~x352 ;
  assign n6485 = n6484 ^ n1121 ;
  assign n6504 = n6485 ^ x350 ;
  assign n6505 = n6484 ^ n1120 ;
  assign n6506 = ~x353 & ~n6505 ;
  assign n6507 = n1121 ^ x354 ;
  assign n6508 = n6507 ^ n1120 ;
  assign n6509 = n6506 & n6508 ;
  assign n6510 = n6504 & n6509 ;
  assign n6489 = x353 & x354 ;
  assign n6490 = n6489 ^ n1123 ;
  assign n6491 = ~n6484 & n6490 ;
  assign n6483 = x349 & x350 ;
  assign n6486 = x354 & ~n6485 ;
  assign n6487 = n6483 & n6486 ;
  assign n6488 = n6487 ^ n6483 ;
  assign n6492 = n6491 ^ n6488 ;
  assign n6497 = n6485 & ~n6489 ;
  assign n6498 = n6497 ^ n6488 ;
  assign n6499 = n6492 & ~n6498 ;
  assign n6501 = ~n1120 & n6491 ;
  assign n6502 = n6499 & n6501 ;
  assign n6500 = n6499 ^ n6488 ;
  assign n6503 = n6502 ^ n6500 ;
  assign n6511 = n6510 ^ n6503 ;
  assign n6512 = x353 ^ x350 ;
  assign n6513 = ~n1123 & n6512 ;
  assign n6514 = n6513 ^ x350 ;
  assign n6515 = n6514 ^ x351 ;
  assign n6516 = ~n6511 & ~n6515 ;
  assign n6517 = n6482 & n6516 ;
  assign n6518 = n6517 ^ n6511 ;
  assign n6520 = n6519 ^ n6518 ;
  assign n6568 = n6567 ^ n6520 ;
  assign n6479 = n1130 & n1141 ;
  assign n6478 = n1135 & n1140 ;
  assign n6480 = n6479 ^ n6478 ;
  assign n6439 = x359 ^ x358 ;
  assign n6443 = ~n1136 & ~n6439 ;
  assign n6438 = x357 ^ x356 ;
  assign n6440 = n6439 ^ x357 ;
  assign n6441 = n6440 ^ x360 ;
  assign n6442 = ~n6438 & n6441 ;
  assign n6444 = n6443 ^ n6442 ;
  assign n6445 = ~x355 & n6444 ;
  assign n6446 = ~n1137 & ~n6438 ;
  assign n6447 = x360 ^ x355 ;
  assign n6450 = ~x358 & ~n6447 ;
  assign n6451 = n6450 ^ x355 ;
  assign n6452 = n6446 & n6451 ;
  assign n6453 = ~x359 & n6452 ;
  assign n6454 = ~x357 & ~x358 ;
  assign n6457 = n6454 ^ n1137 ;
  assign n6458 = x355 & x356 ;
  assign n6459 = x360 & n6458 ;
  assign n6460 = ~n6457 & n6459 ;
  assign n6461 = n6460 ^ n6458 ;
  assign n6455 = ~x359 & ~x360 ;
  assign n6456 = ~n6454 & ~n6455 ;
  assign n6462 = n6461 ^ n6456 ;
  assign n6463 = n6455 ^ n1136 ;
  assign n6468 = n6457 & n6463 ;
  assign n6469 = n6468 ^ n6456 ;
  assign n6470 = n6462 & n6469 ;
  assign n6471 = n6470 ^ n6461 ;
  assign n6472 = ~n1138 & n6471 ;
  assign n6473 = n6470 & n6472 ;
  assign n6474 = n6473 ^ n6471 ;
  assign n6475 = ~n6453 & ~n6474 ;
  assign n6476 = ~n6445 & n6475 ;
  assign n6400 = x365 ^ x364 ;
  assign n6404 = ~n1131 & ~n6400 ;
  assign n6399 = x363 ^ x362 ;
  assign n6401 = n6400 ^ x363 ;
  assign n6402 = n6401 ^ x366 ;
  assign n6403 = ~n6399 & n6402 ;
  assign n6405 = n6404 ^ n6403 ;
  assign n6406 = ~x361 & n6405 ;
  assign n6407 = ~n1132 & ~n6399 ;
  assign n6408 = x366 ^ x361 ;
  assign n6411 = ~x364 & ~n6408 ;
  assign n6412 = n6411 ^ x361 ;
  assign n6413 = n6407 & n6412 ;
  assign n6414 = ~x365 & n6413 ;
  assign n6415 = ~x363 & ~x364 ;
  assign n6418 = n6415 ^ n1132 ;
  assign n6419 = x361 & x362 ;
  assign n6420 = x366 & n6419 ;
  assign n6421 = ~n6418 & n6420 ;
  assign n6422 = n6421 ^ n6419 ;
  assign n6416 = ~x365 & ~x366 ;
  assign n6417 = ~n6415 & ~n6416 ;
  assign n6423 = n6422 ^ n6417 ;
  assign n6424 = n6416 ^ n1131 ;
  assign n6429 = n6418 & n6424 ;
  assign n6430 = n6429 ^ n6417 ;
  assign n6431 = n6423 & n6430 ;
  assign n6432 = n6431 ^ n6422 ;
  assign n6433 = ~n1133 & n6432 ;
  assign n6434 = n6431 & n6433 ;
  assign n6435 = n6434 ^ n6432 ;
  assign n6436 = ~n6414 & ~n6435 ;
  assign n6437 = ~n6406 & n6436 ;
  assign n6477 = n6476 ^ n6437 ;
  assign n6481 = n6480 ^ n6477 ;
  assign n6569 = n6568 ^ n6481 ;
  assign n6397 = n1119 & n1142 ;
  assign n6396 = n1107 & n1118 ;
  assign n6398 = n6397 ^ n6396 ;
  assign n6570 = n6569 ^ n6398 ;
  assign n6698 = n6697 ^ n6570 ;
  assign n6699 = n8474 ^ n6698 ;
  assign n8689 = n6699 ^ n5418 ;
  assign n8696 = n6033 & ~n8689 ;
  assign n8697 = n8696 ^ n6699 ;
  assign n8973 = n8972 ^ n8697 ;
  assign n8676 = n6211 ^ x309 ;
  assign n8677 = n6215 & n8676 ;
  assign n8678 = n8677 ^ n1145 ;
  assign n8679 = ~x310 & ~n8678 ;
  assign n8680 = ~n8677 & n8679 ;
  assign n8681 = n8680 ^ n8678 ;
  assign n8682 = x307 & n6238 ;
  assign n8683 = n8681 & n8682 ;
  assign n8684 = n8683 ^ n8681 ;
  assign n8673 = n6185 ^ n6040 ;
  assign n8674 = n6243 & n8673 ;
  assign n8675 = n8674 ^ n6185 ;
  assign n8685 = n8684 ^ n8675 ;
  assign n8665 = n6061 & ~n6132 ;
  assign n8659 = n6115 ^ n6109 ;
  assign n8660 = x302 & n6108 ;
  assign n8661 = n8660 ^ n6109 ;
  assign n8662 = n8659 & ~n8661 ;
  assign n8663 = n8662 ^ n6109 ;
  assign n8664 = ~n6126 & n8663 ;
  assign n8666 = n8665 ^ n8664 ;
  assign n8667 = n6128 ^ n6042 ;
  assign n8668 = ~n6137 & n8667 ;
  assign n8669 = n8668 ^ n6128 ;
  assign n11988 = n8669 ^ n8665 ;
  assign n11989 = n8666 & ~n11988 ;
  assign n11990 = n11989 ^ n8665 ;
  assign n8658 = n6171 & ~n6176 ;
  assign n12000 = n11990 ^ n8658 ;
  assign n8670 = n8669 ^ n8666 ;
  assign n11995 = n11990 ^ n8670 ;
  assign n12002 = n12000 ^ n11995 ;
  assign n8650 = n6137 ^ n6042 ;
  assign n8656 = ~n8650 & n8653 ;
  assign n8651 = n8650 ^ n6040 ;
  assign n8654 = n8653 ^ n8651 ;
  assign n8655 = n6243 & ~n8654 ;
  assign n8657 = n8656 ^ n8655 ;
  assign n8672 = n12002 ^ n8657 ;
  assign n8686 = n8685 ^ n8672 ;
  assign n8638 = x271 & n6327 ;
  assign n8613 = n1176 & n1182 ;
  assign n8629 = n8613 ^ n6282 ;
  assign n8630 = n6332 & n8629 ;
  assign n8631 = n8630 ^ n6282 ;
  assign n8632 = n8631 ^ n1179 ;
  assign n8627 = n6308 ^ x273 ;
  assign n8628 = n6312 & n8627 ;
  assign n8633 = n8632 ^ n8628 ;
  assign n8634 = n8633 ^ n8631 ;
  assign n8635 = ~x274 & ~n8628 ;
  assign n8636 = ~n8634 & n8635 ;
  assign n8637 = n8636 ^ n8633 ;
  assign n8639 = n8637 ^ n8631 ;
  assign n8640 = n8638 & n8639 ;
  assign n8641 = n8640 ^ n8637 ;
  assign n8625 = n6383 ^ n6357 ;
  assign n8615 = n1171 & n1187 ;
  assign n8622 = n8615 ^ n6364 ;
  assign n8623 = n6391 & ~n8622 ;
  assign n8624 = n8623 ^ n6390 ;
  assign n8626 = n8625 ^ n8624 ;
  assign n8642 = n8641 ^ n8626 ;
  assign n8614 = n8613 ^ n6332 ;
  assign n8617 = n8613 ^ n6338 ;
  assign n8620 = n8614 & ~n8617 ;
  assign n8616 = n8615 ^ n8614 ;
  assign n8618 = n8617 ^ n8616 ;
  assign n8619 = n6391 & ~n8618 ;
  assign n8621 = n8620 ^ n8619 ;
  assign n8643 = n8642 ^ n8621 ;
  assign n8612 = n6264 & ~n6279 ;
  assign n8644 = n8643 ^ n8612 ;
  assign n8645 = n8644 ^ n6393 ;
  assign n8646 = n8645 ^ n6035 ;
  assign n8647 = n8646 ^ n8644 ;
  assign n8648 = n6394 & ~n8647 ;
  assign n8649 = n8648 ^ n8645 ;
  assign n8687 = n8686 ^ n8649 ;
  assign n8594 = n6424 ^ n6418 ;
  assign n8595 = x362 & n6417 ;
  assign n8596 = n8595 ^ n6418 ;
  assign n8597 = n8594 & ~n8596 ;
  assign n8598 = n8597 ^ n6418 ;
  assign n8599 = ~n6435 & ~n8598 ;
  assign n8600 = n8599 ^ n6435 ;
  assign n8588 = n6463 ^ n6457 ;
  assign n8589 = x356 & n6456 ;
  assign n8590 = n8589 ^ n6457 ;
  assign n8591 = n8588 & ~n8590 ;
  assign n8592 = n8591 ^ n6457 ;
  assign n8593 = ~n6474 & n8592 ;
  assign n8601 = n8600 ^ n8593 ;
  assign n8585 = n6478 ^ n6437 ;
  assign n8586 = ~n6477 & n8585 ;
  assign n8587 = n8586 ^ n6478 ;
  assign n8602 = n8601 ^ n8587 ;
  assign n8582 = n6568 ^ n6479 ;
  assign n8583 = ~n6481 & ~n8582 ;
  assign n8584 = n8583 ^ n6568 ;
  assign n8603 = n8602 ^ n8584 ;
  assign n8578 = n6567 ^ n6518 ;
  assign n8579 = n6520 & ~n8578 ;
  assign n8580 = n8579 ^ n6567 ;
  assign n8575 = ~n6485 & n6514 ;
  assign n8576 = ~n6503 & n8575 ;
  assign n8572 = n6553 & ~n6558 ;
  assign n8573 = n8572 ^ n6503 ;
  assign n8577 = n8576 ^ n8573 ;
  assign n8581 = n8580 ^ n8577 ;
  assign n8604 = n8603 ^ n8581 ;
  assign n8563 = n6593 ^ x338 ;
  assign n8542 = n6598 ^ n6594 ;
  assign n8548 = n8563 ^ n8542 ;
  assign n8552 = n1108 & n8548 ;
  assign n8546 = n6593 & ~n6597 ;
  assign n8553 = n8552 ^ n8546 ;
  assign n8539 = n6593 ^ x337 ;
  assign n8540 = n8539 ^ n6598 ;
  assign n8544 = n8540 ^ n6594 ;
  assign n8554 = n8553 ^ n8544 ;
  assign n8555 = n8552 ^ n8542 ;
  assign n8556 = n8555 ^ n8544 ;
  assign n8557 = n8554 & n8556 ;
  assign n8558 = ~n6594 & n8557 ;
  assign n8559 = n8558 ^ n8552 ;
  assign n8560 = n8559 ^ n1108 ;
  assign n8566 = n8560 ^ n6593 ;
  assign n8567 = n8566 ^ n8563 ;
  assign n8531 = n6572 ^ x332 ;
  assign n8510 = n6577 ^ n6573 ;
  assign n8516 = n8531 ^ n8510 ;
  assign n8520 = n1113 & n8516 ;
  assign n8514 = n6572 & ~n6576 ;
  assign n8521 = n8520 ^ n8514 ;
  assign n8507 = n6572 ^ x331 ;
  assign n8508 = n8507 ^ n6577 ;
  assign n8512 = n8508 ^ n6573 ;
  assign n8522 = n8521 ^ n8512 ;
  assign n8523 = n8520 ^ n8510 ;
  assign n8524 = n8523 ^ n8512 ;
  assign n8525 = n8522 & n8524 ;
  assign n8526 = ~n6573 & n8525 ;
  assign n8527 = n8526 ^ n8520 ;
  assign n8528 = n8527 ^ n1113 ;
  assign n8534 = n8528 ^ n6572 ;
  assign n8535 = n8534 ^ n8531 ;
  assign n8568 = n8567 ^ n8535 ;
  assign n8501 = n6612 ^ n6591 ;
  assign n8502 = n6614 & n8501 ;
  assign n8503 = n8502 ^ n6591 ;
  assign n8569 = n8568 ^ n8503 ;
  assign n8492 = n6641 ^ n6635 ;
  assign n8493 = x320 & n6634 ;
  assign n8494 = n8493 ^ n6635 ;
  assign n8495 = n8492 & ~n8494 ;
  assign n8496 = n8495 ^ n6635 ;
  assign n8497 = ~n6652 & ~n8496 ;
  assign n8498 = n8497 ^ n6652 ;
  assign n8486 = n6681 ^ n6675 ;
  assign n8487 = x326 & n6674 ;
  assign n8488 = n8487 ^ n6675 ;
  assign n8489 = n8486 & ~n8488 ;
  assign n8490 = n8489 ^ n6675 ;
  assign n8491 = ~n6692 & n8490 ;
  assign n8499 = n8498 ^ n8491 ;
  assign n8483 = n6655 ^ n6654 ;
  assign n8484 = n6695 & n8483 ;
  assign n8485 = n8484 ^ n6655 ;
  assign n8500 = n8499 ^ n8485 ;
  assign n8570 = n8569 ^ n8500 ;
  assign n8480 = n6615 ^ n6396 ;
  assign n8481 = n6697 & n8480 ;
  assign n8482 = n8481 ^ n6615 ;
  assign n8571 = n8570 ^ n8482 ;
  assign n8605 = n8604 ^ n8571 ;
  assign n8475 = n6569 ^ n6397 ;
  assign n8476 = n6697 ^ n6397 ;
  assign n8477 = n8476 ^ n6396 ;
  assign n8478 = ~n8475 & ~n8477 ;
  assign n8479 = n8478 ^ n6569 ;
  assign n8606 = n8605 ^ n8479 ;
  assign n8607 = n8606 ^ n6698 ;
  assign n8608 = n8607 ^ n6034 ;
  assign n8609 = n8608 ^ n8606 ;
  assign n8610 = ~n8474 & ~n8609 ;
  assign n8611 = n8610 ^ n8607 ;
  assign n8688 = n8687 ^ n8611 ;
  assign n12117 = n8697 ^ n8688 ;
  assign n12118 = n8973 & ~n12117 ;
  assign n12119 = n12118 ^ n8688 ;
  assign n12116 = n12115 ^ n12075 ;
  assign n12120 = n12119 ^ n12116 ;
  assign n12676 = n12675 ^ n12644 ;
  assign n12677 = n12676 ^ n12119 ;
  assign n11991 = ~n8675 & n8684 ;
  assign n11992 = n11991 ^ n8685 ;
  assign n11997 = ~n8670 & ~n11992 ;
  assign n11998 = n11997 ^ n11990 ;
  assign n12006 = n11992 ^ n8670 ;
  assign n12007 = n12006 ^ n11990 ;
  assign n11993 = n11992 ^ n11990 ;
  assign n12003 = n12002 ^ n11993 ;
  assign n12004 = n12003 ^ n11990 ;
  assign n12020 = n8658 ^ n8657 ;
  assign n12005 = n12004 & n12020 ;
  assign n12008 = n12007 ^ n12005 ;
  assign n12009 = n11998 & n12008 ;
  assign n12010 = n12009 ^ n11990 ;
  assign n12013 = ~n8672 & n11991 ;
  assign n12014 = ~n12010 & n12013 ;
  assign n12015 = n12014 ^ n12010 ;
  assign n12016 = n8670 & ~n12015 ;
  assign n12017 = n8684 ^ n8670 ;
  assign n12021 = n12017 ^ n8675 ;
  assign n12022 = n12021 ^ n8657 ;
  assign n12023 = n12020 & ~n12022 ;
  assign n12028 = n8657 & n12023 ;
  assign n12029 = n12028 ^ n12017 ;
  assign n12030 = ~n8685 & n12029 ;
  assign n12024 = n12017 ^ n11990 ;
  assign n12025 = n12024 ^ n12023 ;
  assign n12031 = n12030 ^ n12025 ;
  assign n12032 = n12031 ^ n11990 ;
  assign n12033 = n8657 & ~n12032 ;
  assign n12034 = n12016 & n12033 ;
  assign n12035 = n12034 ^ n12031 ;
  assign n11971 = n8631 ^ n8621 ;
  assign n11972 = ~n8641 & n11971 ;
  assign n11973 = n11972 ^ n8631 ;
  assign n11979 = n8626 & ~n8644 ;
  assign n11980 = n11973 & n11979 ;
  assign n11974 = n8626 ^ n8612 ;
  assign n11976 = n8643 & ~n11974 ;
  assign n11977 = n11976 ^ n8612 ;
  assign n11978 = ~n11973 & n11977 ;
  assign n11981 = n11980 ^ n11978 ;
  assign n11968 = n8624 ^ n6357 ;
  assign n11969 = n8625 & n11968 ;
  assign n11970 = n11969 ^ n6383 ;
  assign n11982 = n11981 ^ n11970 ;
  assign n11984 = n11982 ^ n8644 ;
  assign n11983 = n11982 ^ n8686 ;
  assign n11985 = n11984 ^ n11983 ;
  assign n11986 = ~n8649 & n11985 ;
  assign n11987 = n11986 ^ n11984 ;
  assign n12036 = n12035 ^ n11987 ;
  assign n11961 = n8584 ^ n8581 ;
  assign n11962 = ~n8603 & n11961 ;
  assign n11963 = n11962 ^ n8581 ;
  assign n11957 = n8580 ^ n8572 ;
  assign n11958 = ~n8577 & ~n11957 ;
  assign n11959 = n11958 ^ n8572 ;
  assign n11954 = n8600 ^ n8587 ;
  assign n11955 = ~n8601 & n11954 ;
  assign n11956 = n11955 ^ n8600 ;
  assign n11960 = n11959 ^ n11956 ;
  assign n11964 = n11963 ^ n11960 ;
  assign n11950 = n8567 ^ n8503 ;
  assign n11951 = n8568 & ~n11950 ;
  assign n11952 = n11951 ^ n8567 ;
  assign n11947 = n8569 ^ n8482 ;
  assign n11948 = n8570 & ~n11947 ;
  assign n11942 = n8498 ^ n8485 ;
  assign n11943 = ~n8499 & n11942 ;
  assign n11944 = n11943 ^ n8498 ;
  assign n11945 = n11944 ^ n8569 ;
  assign n11949 = n11948 ^ n11945 ;
  assign n11953 = n11952 ^ n11949 ;
  assign n11965 = n11964 ^ n11953 ;
  assign n11939 = n8571 ^ n8479 ;
  assign n11940 = ~n8605 & n11939 ;
  assign n11941 = n11940 ^ n8604 ;
  assign n11966 = n11965 ^ n11941 ;
  assign n11936 = n8687 ^ n8606 ;
  assign n11937 = ~n8611 & ~n11936 ;
  assign n11938 = n11937 ^ n8606 ;
  assign n11967 = n11966 ^ n11938 ;
  assign n12037 = n12036 ^ n11967 ;
  assign n12678 = n12677 ^ n12037 ;
  assign n12679 = n12678 ^ n12676 ;
  assign n12680 = ~n12120 & n12679 ;
  assign n12681 = n12680 ^ n12677 ;
  assign n12696 = n11956 & ~n11959 ;
  assign n12697 = ~n11941 & n12696 ;
  assign n12703 = n12697 ^ n11960 ;
  assign n12701 = n12696 ^ n11960 ;
  assign n12702 = n11941 & n12701 ;
  assign n12704 = n12703 ^ n12702 ;
  assign n12705 = n12704 ^ n11941 ;
  assign n12693 = n11952 ^ n11944 ;
  assign n12694 = ~n11949 & n12693 ;
  assign n12695 = n12694 ^ n11944 ;
  assign n12725 = ~n11953 & ~n11963 ;
  assign n12726 = n12695 & n12725 ;
  assign n12727 = ~n12705 & n12726 ;
  assign n12698 = n12697 ^ n12695 ;
  assign n12699 = ~n11953 & ~n12698 ;
  assign n12712 = ~n11963 & n12699 ;
  assign n12713 = ~n12705 & n12712 ;
  assign n12714 = n12713 ^ n12705 ;
  assign n12700 = n12699 ^ n11953 ;
  assign n12706 = n12705 ^ n12700 ;
  assign n12715 = n12714 ^ n12706 ;
  assign n12716 = ~n12695 & n12715 ;
  assign n12717 = n12702 ^ n11963 ;
  assign n12718 = n12702 ^ n11953 ;
  assign n12719 = n12705 & n12718 ;
  assign n12720 = n12717 & n12719 ;
  assign n12721 = n12720 ^ n12702 ;
  assign n12723 = ~n12716 & ~n12721 ;
  assign n12728 = n12727 ^ n12723 ;
  assign n12722 = n12721 ^ n12716 ;
  assign n12724 = n12723 ^ n12722 ;
  assign n12729 = n12728 ^ n12724 ;
  assign n12688 = n12035 ^ n11982 ;
  assign n12689 = n11987 & n12688 ;
  assign n12690 = n12689 ^ n11982 ;
  assign n12691 = n12690 ^ n12015 ;
  assign n12685 = n11970 & ~n11981 ;
  assign n12686 = n12685 ^ n11978 ;
  assign n12682 = n12036 ^ n11938 ;
  assign n12683 = ~n11967 & n12682 ;
  assign n12684 = n12683 ^ n12036 ;
  assign n12687 = n12686 ^ n12684 ;
  assign n12692 = n12691 ^ n12687 ;
  assign n12730 = n12729 ^ n12692 ;
  assign n12913 = n12730 ^ n12676 ;
  assign n12914 = ~n12681 & ~n12913 ;
  assign n12915 = n12914 ^ n12676 ;
  assign n13156 = n13151 ^ n12915 ;
  assign n13152 = n12915 & n13151 ;
  assign n13153 = n12907 & n12911 ;
  assign n13154 = n12904 & n13153 ;
  assign n13155 = n13152 & ~n13154 ;
  assign n13157 = n13156 ^ n13155 ;
  assign n12916 = n12015 & ~n12726 ;
  assign n12917 = ~n12684 & ~n12690 ;
  assign n12918 = n12916 & n12917 ;
  assign n12919 = n12686 & ~n12918 ;
  assign n12920 = ~n12724 & n12919 ;
  assign n12921 = n12690 ^ n12684 ;
  assign n12922 = ~n12691 & n12921 ;
  assign n12923 = n12922 ^ n12690 ;
  assign n12924 = n12920 & ~n12923 ;
  assign n12925 = n12924 ^ n12919 ;
  assign n12929 = n12723 ^ n12015 ;
  assign n12930 = n12929 ^ n12690 ;
  assign n12933 = n12684 & n12930 ;
  assign n12934 = n12933 ^ n12723 ;
  assign n12935 = n12929 ^ n12727 ;
  assign n12936 = n12933 ^ n12930 ;
  assign n12937 = n12935 & n12936 ;
  assign n12938 = n12937 ^ n12929 ;
  assign n12939 = n12934 & ~n12938 ;
  assign n12940 = n12939 ^ n12723 ;
  assign n12941 = n12925 & ~n12940 ;
  assign n12944 = ~n12684 & ~n12728 ;
  assign n12942 = ~n12686 & ~n12723 ;
  assign n12945 = n12944 ^ n12942 ;
  assign n12946 = n12945 ^ n12684 ;
  assign n12947 = ~n12690 & ~n12946 ;
  assign n12950 = n12724 & n12944 ;
  assign n12951 = n12947 & n12950 ;
  assign n12943 = ~n12684 & n12942 ;
  assign n12948 = n12947 ^ n12943 ;
  assign n12952 = n12951 ^ n12948 ;
  assign n12953 = n12952 ^ n12943 ;
  assign n12954 = n12953 ^ n12952 ;
  assign n12955 = n12954 ^ n12727 ;
  assign n12956 = n12955 ^ n12954 ;
  assign n12957 = n12954 ^ n12686 ;
  assign n12958 = n12957 ^ n12954 ;
  assign n12959 = n12956 & ~n12958 ;
  assign n12960 = n12959 ^ n12954 ;
  assign n12961 = n12690 & n12960 ;
  assign n12962 = n12961 ^ n12953 ;
  assign n12963 = ~n12015 & n12962 ;
  assign n12964 = n12963 ^ n12952 ;
  assign n12965 = n12690 & ~n12724 ;
  assign n12966 = n12942 & n12965 ;
  assign n12969 = n12966 ^ n12015 ;
  assign n12970 = n12969 ^ n12966 ;
  assign n12967 = n12966 ^ n12724 ;
  assign n12971 = n12966 ^ n12684 ;
  assign n12972 = n12971 ^ n12966 ;
  assign n12975 = ~n12967 & n12972 ;
  assign n12976 = ~n12970 & n12975 ;
  assign n12977 = n12976 ^ n12970 ;
  assign n12978 = n12977 ^ n12969 ;
  assign n12979 = ~n12964 & ~n12978 ;
  assign n12980 = ~n12941 & n12979 ;
  assign n13158 = n12721 ^ n12692 ;
  assign n13159 = n12716 ^ n12692 ;
  assign n13160 = ~n13158 & n13159 ;
  assign n13161 = n13160 ^ n12721 ;
  assign n13162 = n12015 & n12952 ;
  assign n13163 = ~n13161 & n13162 ;
  assign n13164 = n13163 ^ n13161 ;
  assign n13165 = ~n12941 & ~n13164 ;
  assign n12912 = n12911 ^ n12908 ;
  assign n13166 = n13165 ^ n12912 ;
  assign n13167 = n13166 ^ n13151 ;
  assign n13168 = n13167 ^ n13154 ;
  assign n13169 = ~n12980 & n13168 ;
  assign n13170 = n13157 & n13169 ;
  assign n13171 = n13164 ^ n13154 ;
  assign n13172 = n13171 ^ n13164 ;
  assign n13173 = n13164 ^ n13152 ;
  assign n13174 = n12979 & n13173 ;
  assign n13175 = n13174 ^ n13164 ;
  assign n13176 = ~n13172 & ~n13175 ;
  assign n13177 = n13176 ^ n13164 ;
  assign n13178 = ~n12941 & ~n13177 ;
  assign n13179 = ~n13170 & ~n13178 ;
  assign n13301 = n12558 & ~n12881 ;
  assign n13302 = n12837 & n13299 ;
  assign n13303 = n13301 & n13302 ;
  assign n13304 = n13179 & ~n13303 ;
  assign n13305 = ~n13300 & n13304 ;
  assign n13306 = n13305 ^ n13179 ;
  assign n12838 = n12837 ^ n12835 ;
  assign n13138 = n12837 ^ n12832 ;
  assign n13139 = ~n12838 & ~n13138 ;
  assign n13140 = n13139 ^ n12832 ;
  assign n12839 = n12838 ^ n12832 ;
  assign n12895 = n12894 ^ n12839 ;
  assign n13135 = n12839 ^ n12829 ;
  assign n13136 = n12895 & n13135 ;
  assign n13137 = n13136 ^ n12894 ;
  assign n13141 = n13140 ^ n13137 ;
  assign n12731 = n12730 ^ n12681 ;
  assign n12641 = n12640 ^ n12571 ;
  assign n12732 = n12731 ^ n12641 ;
  assign n12896 = n12895 ^ n12829 ;
  assign n12897 = n12896 ^ n12641 ;
  assign n12898 = n12897 ^ n12896 ;
  assign n11933 = n11932 ^ n11850 ;
  assign n8469 = n8468 ^ n8148 ;
  assign n11934 = n11933 ^ n8469 ;
  assign n8974 = n8973 ^ n8688 ;
  assign n7940 = n7939 ^ n7396 ;
  assign n6700 = n6699 ^ n6033 ;
  assign n7941 = n7940 ^ n6700 ;
  assign n1192 = n1191 ^ n1096 ;
  assign n1383 = n1382 ^ n1287 ;
  assign n4128 = n1192 & n1383 ;
  assign n8470 = n7940 ^ n4128 ;
  assign n8471 = n7941 & n8470 ;
  assign n8472 = n8471 ^ n7940 ;
  assign n8975 = n8974 ^ n8472 ;
  assign n11758 = n8472 ^ n8469 ;
  assign n11759 = n8975 & n11758 ;
  assign n11935 = n11934 ^ n11759 ;
  assign n12121 = n12120 ^ n12037 ;
  assign n12536 = n12121 ^ n11933 ;
  assign n12537 = n11935 & n12536 ;
  assign n12538 = n12537 ^ n12121 ;
  assign n12899 = n12898 ^ n12538 ;
  assign n12900 = n12732 & n12899 ;
  assign n12901 = n12900 ^ n12897 ;
  assign n12981 = n12980 ^ n12915 ;
  assign n12982 = n12981 ^ n12912 ;
  assign n13146 = n12982 ^ n12896 ;
  assign n13147 = ~n12901 & ~n13146 ;
  assign n13148 = n13147 ^ n12896 ;
  assign n13307 = n13148 ^ n13140 ;
  assign n13308 = n13307 ^ n13137 ;
  assign n13309 = n13308 ^ n13140 ;
  assign n13310 = ~n13141 & n13309 ;
  assign n13311 = n13310 ^ n13308 ;
  assign n13312 = n13311 ^ n13179 ;
  assign n13313 = n13312 ^ n13311 ;
  assign n13316 = n13311 ^ n13137 ;
  assign n13317 = n13316 ^ n13311 ;
  assign n13318 = n13310 & n13317 ;
  assign n13319 = n13313 & n13318 ;
  assign n13320 = n13319 ^ n13313 ;
  assign n13321 = n13320 ^ n13312 ;
  assign n13322 = n13144 & n13321 ;
  assign n13323 = n13322 ^ n12886 ;
  assign n13324 = n13323 ^ n13322 ;
  assign n13325 = n13322 ^ n12852 ;
  assign n13326 = n13325 ^ n13322 ;
  assign n13327 = ~n13324 & n13326 ;
  assign n13328 = n13327 ^ n13322 ;
  assign n13329 = n13306 & ~n13328 ;
  assign n13330 = n13329 ^ n13322 ;
  assign n13331 = n13148 ^ n13137 ;
  assign n13332 = n13331 ^ n13148 ;
  assign n13333 = ~n13179 & n13332 ;
  assign n13334 = n13333 ^ n13148 ;
  assign n13335 = n13179 ^ n13141 ;
  assign n13336 = n13335 ^ n13144 ;
  assign n13337 = n13334 & ~n13336 ;
  assign n13338 = n13337 ^ n13179 ;
  assign n13339 = ~n13144 & ~n13338 ;
  assign n13340 = ~n13330 & ~n13339 ;
  assign n13261 = n12980 & ~n13154 ;
  assign n13262 = ~n13152 & n13261 ;
  assign n13263 = ~n13164 & n13262 ;
  assign n13264 = n13263 ^ n13261 ;
  assign n13265 = n13264 ^ n13154 ;
  assign n13266 = ~n13165 & n13170 ;
  assign n13267 = ~n13265 & n13266 ;
  assign n13268 = n13267 ^ n13265 ;
  assign n13341 = n13340 ^ n13268 ;
  assign n4306 = ~x969 & ~x970 ;
  assign n1506 = x970 ^ x969 ;
  assign n4307 = n4306 ^ n1506 ;
  assign n4312 = ~x971 & ~x972 ;
  assign n1507 = x972 ^ x971 ;
  assign n4313 = n4312 ^ n1507 ;
  assign n4314 = n4307 & n4313 ;
  assign n4308 = x967 & x968 ;
  assign n4309 = ~n4307 & n4308 ;
  assign n4310 = x972 & n4309 ;
  assign n4311 = n4310 ^ n4308 ;
  assign n4315 = n4314 ^ n4311 ;
  assign n4320 = ~n4306 & ~n4312 ;
  assign n4321 = n4320 ^ n4311 ;
  assign n4322 = ~n4315 & n4321 ;
  assign n1509 = x968 ^ x967 ;
  assign n4323 = n4322 ^ n4311 ;
  assign n4324 = ~n1509 & n4323 ;
  assign n4325 = n4322 & n4324 ;
  assign n4326 = n4325 ^ n4323 ;
  assign n9692 = n4313 ^ n4307 ;
  assign n9693 = n9692 ^ n4314 ;
  assign n9694 = ~n4309 & n9693 ;
  assign n9695 = ~n4326 & n9694 ;
  assign n4336 = x975 & x976 ;
  assign n4346 = x973 & x974 ;
  assign n4347 = n4336 & n4346 ;
  assign n4348 = ~x978 & n4347 ;
  assign n4329 = x977 & x978 ;
  assign n1512 = x978 ^ x977 ;
  assign n4330 = n4329 ^ n1512 ;
  assign n1511 = x974 ^ x973 ;
  assign n4337 = n4329 & n4336 ;
  assign n4331 = n4329 ^ x976 ;
  assign n4338 = n4337 ^ n4331 ;
  assign n1514 = x976 ^ x975 ;
  assign n4332 = n1514 & ~n4331 ;
  assign n4339 = n4338 ^ n4332 ;
  assign n4340 = n4339 ^ n4336 ;
  assign n4341 = x974 & n4340 ;
  assign n4333 = n4332 ^ x975 ;
  assign n4342 = n4341 ^ n4333 ;
  assign n4343 = ~n1511 & n4342 ;
  assign n4344 = n4343 ^ n4333 ;
  assign n4345 = n4330 & n4344 ;
  assign n4350 = n4348 ^ n4345 ;
  assign n4351 = x974 & n4330 ;
  assign n4352 = n4333 & ~n4337 ;
  assign n4353 = ~n4351 & n4352 ;
  assign n4354 = n4353 ^ n4333 ;
  assign n9696 = ~n4350 & ~n4354 ;
  assign n12433 = ~n9695 & ~n9696 ;
  assign n9697 = n9696 ^ n9695 ;
  assign n4374 = ~x983 & ~x984 ;
  assign n1501 = x984 ^ x983 ;
  assign n4375 = n4374 ^ n1501 ;
  assign n4378 = n4375 ^ x982 ;
  assign n4376 = x981 & x982 ;
  assign n4377 = ~n4375 & n4376 ;
  assign n4434 = n4378 ^ n4377 ;
  assign n1502 = x982 ^ x981 ;
  assign n4379 = n1502 & n4378 ;
  assign n4435 = n4434 ^ n4379 ;
  assign n4436 = ~x980 & n4435 ;
  assign n4380 = n4379 ^ x981 ;
  assign n4428 = n4380 ^ n4374 ;
  assign n4427 = ~n4374 & n4380 ;
  assign n4429 = n4428 ^ n4427 ;
  assign n1503 = n1502 ^ n1501 ;
  assign n1500 = x980 ^ x979 ;
  assign n1504 = n1503 ^ n1500 ;
  assign n4430 = n4429 ^ n1504 ;
  assign n4431 = n1504 ^ x979 ;
  assign n4432 = ~n4430 & n4431 ;
  assign n4388 = x987 & x988 ;
  assign n4406 = n4388 ^ x986 ;
  assign n1496 = x988 ^ x987 ;
  assign n4409 = n1496 ^ x985 ;
  assign n4410 = ~x990 & n4409 ;
  assign n4411 = n4410 ^ x985 ;
  assign n4412 = ~n4388 & n4411 ;
  assign n4413 = n4412 ^ x985 ;
  assign n4414 = ~n4406 & n4413 ;
  assign n4423 = x989 & n4414 ;
  assign n4386 = ~x989 & ~x990 ;
  assign n1495 = x990 ^ x989 ;
  assign n4387 = n4386 ^ n1495 ;
  assign n4390 = n4387 ^ x988 ;
  assign n4392 = n1496 & n4390 ;
  assign n4397 = n4392 ^ x987 ;
  assign n4389 = ~n4387 & n4388 ;
  assign n4394 = x986 & ~n4386 ;
  assign n4417 = ~n4389 & ~n4394 ;
  assign n4418 = n4397 & n4417 ;
  assign n4419 = n4418 ^ n4397 ;
  assign n4415 = x990 & n4414 ;
  assign n4398 = n4397 ^ n4386 ;
  assign n4399 = n4398 ^ x986 ;
  assign n4400 = n4399 ^ n4397 ;
  assign n4391 = n4390 ^ n4389 ;
  assign n4393 = n4392 ^ n4391 ;
  assign n4401 = x986 & ~n4393 ;
  assign n4402 = n4401 ^ n4397 ;
  assign n4403 = n4400 & n4402 ;
  assign n4404 = n4403 ^ n4397 ;
  assign n4405 = x985 & n4404 ;
  assign n4416 = n4415 ^ n4405 ;
  assign n4420 = n4419 ^ n4416 ;
  assign n4421 = n4416 ^ n4414 ;
  assign n4422 = ~n4420 & ~n4421 ;
  assign n4424 = n4423 ^ n4422 ;
  assign n4395 = ~x985 & ~n4394 ;
  assign n4396 = n4393 & n4395 ;
  assign n4425 = n4424 ^ n4396 ;
  assign n4381 = ~n4377 & n4380 ;
  assign n4382 = x980 & n4381 ;
  assign n4383 = ~n4374 & n4382 ;
  assign n4384 = n4383 ^ n4381 ;
  assign n4385 = n4384 ^ n4380 ;
  assign n4426 = n4425 ^ n4385 ;
  assign n4433 = n4432 ^ n4426 ;
  assign n4437 = n4436 ^ n4433 ;
  assign n4368 = x977 & n4347 ;
  assign n4356 = n4330 ^ x973 ;
  assign n4357 = n4356 ^ x974 ;
  assign n4358 = ~n4351 & n4357 ;
  assign n4359 = n4340 ^ x974 ;
  assign n4360 = n4359 ^ n4339 ;
  assign n4363 = ~n1511 & ~n4360 ;
  assign n4364 = n4363 ^ n4339 ;
  assign n4365 = ~n4358 & ~n4364 ;
  assign n4366 = n4365 ^ n4339 ;
  assign n4355 = ~x973 & n4354 ;
  assign n4367 = n4366 ^ n4355 ;
  assign n4369 = n4368 ^ n4367 ;
  assign n4370 = ~n4350 & n4369 ;
  assign n4291 = x971 ^ x970 ;
  assign n4295 = ~n1507 & ~n4291 ;
  assign n1508 = n1507 ^ n1506 ;
  assign n4290 = x969 ^ x968 ;
  assign n4294 = n1508 & ~n4290 ;
  assign n4296 = n4295 ^ n4294 ;
  assign n4297 = ~x967 & n4296 ;
  assign n4298 = ~n1506 & ~n4290 ;
  assign n4299 = x972 ^ x967 ;
  assign n4302 = ~x970 & ~n4299 ;
  assign n4303 = n4302 ^ x967 ;
  assign n4304 = n4298 & n4303 ;
  assign n4305 = ~x971 & n4304 ;
  assign n4327 = ~n4305 & ~n4326 ;
  assign n4328 = ~n4297 & n4327 ;
  assign n4371 = n4370 ^ n4328 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1515 = n1514 ^ n1513 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1516 = n1515 ^ n1510 ;
  assign n1497 = x986 ^ x985 ;
  assign n1498 = n1497 ^ n1496 ;
  assign n1499 = n1498 ^ n1495 ;
  assign n1505 = n1504 ^ n1499 ;
  assign n4284 = n1510 ^ n1505 ;
  assign n4285 = ~n1516 & n4284 ;
  assign n4286 = n4285 ^ n1505 ;
  assign n4287 = n1499 & ~n4286 ;
  assign n4288 = ~n4285 & n4287 ;
  assign n4289 = n4288 ^ n4286 ;
  assign n4372 = n4371 ^ n4289 ;
  assign n4281 = n1499 & n1504 ;
  assign n4282 = n1510 & n1515 ;
  assign n4283 = n4281 & n4282 ;
  assign n4373 = n4372 ^ n4283 ;
  assign n9680 = n4373 ^ n4281 ;
  assign n9681 = n4437 & n9680 ;
  assign n9682 = n9681 ^ n4281 ;
  assign n9683 = n4289 ^ n4282 ;
  assign n9686 = ~n4371 & ~n9683 ;
  assign n9687 = n9686 ^ n4282 ;
  assign n9688 = ~n9682 & ~n9687 ;
  assign n11477 = n9697 ^ n9688 ;
  assign n9689 = n4328 ^ n4282 ;
  assign n9690 = n4371 & n9689 ;
  assign n9691 = n9690 ^ n4328 ;
  assign n11478 = n11477 ^ n9691 ;
  assign n11473 = n9691 ^ n9688 ;
  assign n11474 = n9695 ^ n9688 ;
  assign n11475 = ~n11473 & ~n11474 ;
  assign n11480 = n11475 ^ n9688 ;
  assign n11481 = n9691 & n11480 ;
  assign n9712 = ~n4416 & ~n4419 ;
  assign n9707 = x979 & n4427 ;
  assign n9702 = n4429 ^ n4377 ;
  assign n9703 = x979 & ~n4435 ;
  assign n9704 = ~n9702 & n9703 ;
  assign n9708 = n9707 ^ n9704 ;
  assign n9709 = ~x980 & n9708 ;
  assign n9710 = n9709 ^ n9704 ;
  assign n9711 = ~n4385 & ~n9710 ;
  assign n9713 = n9712 ^ n9711 ;
  assign n9699 = n4425 ^ n4281 ;
  assign n9700 = ~n4437 & n9699 ;
  assign n9701 = n9700 ^ n4425 ;
  assign n9714 = n9713 ^ n9701 ;
  assign n9698 = n9697 ^ n9691 ;
  assign n9715 = n9714 ^ n9698 ;
  assign n9716 = n9715 ^ n9688 ;
  assign n11479 = n9716 ^ n9696 ;
  assign n11482 = n11481 ^ n11479 ;
  assign n11483 = ~n11478 & ~n11482 ;
  assign n11469 = n9712 ^ n9701 ;
  assign n11470 = n9713 & ~n11469 ;
  assign n11471 = n11470 ^ n9712 ;
  assign n11468 = n9714 ^ n9695 ;
  assign n11472 = n11471 ^ n11468 ;
  assign n11476 = n11475 ^ n11472 ;
  assign n11484 = n11483 ^ n11476 ;
  assign n12443 = n9714 & n11478 ;
  assign n12444 = n11475 ^ n9695 ;
  assign n12445 = n11471 & ~n12444 ;
  assign n12446 = n12443 & n12445 ;
  assign n4184 = x965 ^ x962 ;
  assign n4185 = n4184 ^ x964 ;
  assign n4186 = n4185 ^ x966 ;
  assign n4182 = x965 ^ x963 ;
  assign n4187 = n4186 ^ n4182 ;
  assign n4159 = x966 ^ x964 ;
  assign n4160 = x966 ^ x962 ;
  assign n4161 = n4160 ^ n4159 ;
  assign n4193 = ~n4159 & ~n4161 ;
  assign n4197 = n4193 ^ x963 ;
  assign n4198 = n4197 ^ n4182 ;
  assign n4199 = n4193 & n4198 ;
  assign n4200 = n4199 ^ n4182 ;
  assign n4201 = ~n4187 & n4200 ;
  assign n4202 = n4201 ^ n4197 ;
  assign n9591 = x961 & n4202 ;
  assign n4203 = x965 & x966 ;
  assign n1489 = x966 ^ x965 ;
  assign n4204 = n4203 ^ n1489 ;
  assign n4205 = x962 & n4204 ;
  assign n4209 = n4205 ^ n4203 ;
  assign n4206 = n4203 ^ x964 ;
  assign n9594 = n4206 ^ x963 ;
  assign n9595 = ~n4209 & ~n9594 ;
  assign n1490 = x964 ^ x963 ;
  assign n9596 = n9595 ^ n1490 ;
  assign n9597 = ~n9591 & ~n9596 ;
  assign n4243 = x959 ^ x956 ;
  assign n4244 = n4243 ^ x958 ;
  assign n4245 = n4244 ^ x960 ;
  assign n4241 = x959 ^ x957 ;
  assign n4246 = n4245 ^ n4241 ;
  assign n4218 = x960 ^ x958 ;
  assign n4219 = x960 ^ x956 ;
  assign n4220 = n4219 ^ n4218 ;
  assign n4252 = ~n4218 & ~n4220 ;
  assign n4256 = n4252 ^ x957 ;
  assign n4257 = n4256 ^ n4241 ;
  assign n4258 = n4252 & n4257 ;
  assign n4259 = n4258 ^ n4241 ;
  assign n4260 = ~n4246 & n4259 ;
  assign n4261 = n4260 ^ n4256 ;
  assign n9580 = x955 & n4261 ;
  assign n4262 = x959 & x960 ;
  assign n4265 = n4262 ^ x958 ;
  assign n1484 = x960 ^ x959 ;
  assign n4263 = n4262 ^ n1484 ;
  assign n4264 = x956 & n4263 ;
  assign n4266 = n4265 ^ n4264 ;
  assign n9581 = n4265 ^ x957 ;
  assign n9584 = ~n4266 & ~n9581 ;
  assign n9585 = n9584 ^ n4265 ;
  assign n9586 = ~n9580 & n9585 ;
  assign n9587 = n9586 ^ n9580 ;
  assign n9588 = ~x958 & ~n4262 ;
  assign n9589 = ~n9587 & n9588 ;
  assign n9590 = n9589 ^ n9586 ;
  assign n9592 = n9591 ^ n9590 ;
  assign n9600 = n9597 ^ n9592 ;
  assign n9598 = ~x963 & ~n9595 ;
  assign n9599 = n9597 & n9598 ;
  assign n9601 = n9600 ^ n9599 ;
  assign n4221 = n4220 ^ x960 ;
  assign n4223 = x956 & n4221 ;
  assign n4224 = n4223 ^ x960 ;
  assign n4227 = x960 ^ x957 ;
  assign n4228 = n4227 ^ n4219 ;
  assign n1483 = x956 ^ x955 ;
  assign n4229 = n4228 ^ n1483 ;
  assign n4230 = n4220 ^ n1483 ;
  assign n4231 = n4230 ^ n4219 ;
  assign n4232 = n4231 ^ x960 ;
  assign n4233 = ~n4229 & n4232 ;
  assign n4236 = n4233 ^ x958 ;
  assign n4237 = ~n4224 & ~n4236 ;
  assign n4240 = ~x959 & n4237 ;
  assign n4268 = n4264 ^ n4262 ;
  assign n4269 = ~n4265 & ~n4268 ;
  assign n4267 = x957 & ~n4266 ;
  assign n4270 = n4269 ^ n4267 ;
  assign n4271 = n4270 ^ n4261 ;
  assign n4274 = x955 & n4271 ;
  assign n4275 = n4274 ^ n4270 ;
  assign n4276 = ~n4240 & ~n4275 ;
  assign n4162 = n4161 ^ x966 ;
  assign n4164 = x962 & n4162 ;
  assign n4165 = n4164 ^ x966 ;
  assign n4168 = x966 ^ x963 ;
  assign n4169 = n4168 ^ n4160 ;
  assign n1488 = x962 ^ x961 ;
  assign n4170 = n4169 ^ n1488 ;
  assign n4171 = n4161 ^ n1488 ;
  assign n4172 = n4171 ^ n4160 ;
  assign n4173 = n4172 ^ x966 ;
  assign n4174 = ~n4170 & n4173 ;
  assign n4177 = n4174 ^ x964 ;
  assign n4178 = ~n4165 & ~n4177 ;
  assign n4181 = ~x965 & n4178 ;
  assign n4210 = ~n4206 & ~n4209 ;
  assign n4207 = n4206 ^ n4205 ;
  assign n4208 = x963 & ~n4207 ;
  assign n4211 = n4210 ^ n4208 ;
  assign n4212 = n4211 ^ n4202 ;
  assign n4215 = x961 & n4212 ;
  assign n4216 = n4215 ^ n4211 ;
  assign n4217 = ~n4181 & ~n4216 ;
  assign n4277 = n4276 ^ n4217 ;
  assign n1485 = x958 ^ x957 ;
  assign n1486 = n1485 ^ n1484 ;
  assign n1487 = n1486 ^ n1483 ;
  assign n1491 = n1490 ^ n1489 ;
  assign n1492 = n1491 ^ n1488 ;
  assign n4150 = n1487 & n1492 ;
  assign n9602 = n4217 ^ n4150 ;
  assign n9603 = ~n4277 & n9602 ;
  assign n9604 = n9603 ^ n4150 ;
  assign n11490 = n9604 ^ n9590 ;
  assign n11491 = n9601 & ~n11490 ;
  assign n11492 = n11491 ^ n9604 ;
  assign n9605 = n9604 ^ n9601 ;
  assign n1493 = n1492 ^ n1487 ;
  assign n1480 = x954 ^ x953 ;
  assign n1478 = x952 ^ x951 ;
  assign n1477 = x950 ^ x949 ;
  assign n1479 = n1478 ^ n1477 ;
  assign n1481 = n1480 ^ n1479 ;
  assign n1475 = x948 ^ x947 ;
  assign n1473 = x946 ^ x945 ;
  assign n1472 = x944 ^ x943 ;
  assign n1474 = n1473 ^ n1472 ;
  assign n1476 = n1475 ^ n1474 ;
  assign n1482 = n1481 ^ n1476 ;
  assign n4153 = n1487 ^ n1482 ;
  assign n4154 = ~n1493 & n4153 ;
  assign n4155 = n4154 ^ n1482 ;
  assign n4156 = n1481 & ~n4155 ;
  assign n4157 = ~n4154 & n4156 ;
  assign n4158 = n4157 ^ n4155 ;
  assign n9572 = n4158 ^ n4150 ;
  assign n9573 = ~n4277 & ~n9572 ;
  assign n9574 = n9573 ^ n4150 ;
  assign n4147 = n1475 ^ n1473 ;
  assign n4148 = n1474 & n4147 ;
  assign n4144 = ~x945 & ~x946 ;
  assign n4142 = x947 & ~n1475 ;
  assign n4141 = x943 & ~n1472 ;
  assign n4143 = n4142 ^ n4141 ;
  assign n4145 = n4144 ^ n4143 ;
  assign n4138 = ~x951 & ~x952 ;
  assign n4136 = x953 & ~n1480 ;
  assign n4135 = x949 & ~n1477 ;
  assign n4137 = n4136 ^ n4135 ;
  assign n4139 = n4138 ^ n4137 ;
  assign n4133 = n1480 ^ n1478 ;
  assign n4134 = n1479 & n4133 ;
  assign n4140 = n4139 ^ n4134 ;
  assign n4146 = n4145 ^ n4140 ;
  assign n4149 = n4148 ^ n4146 ;
  assign n4278 = n4277 ^ n4158 ;
  assign n4151 = n1476 & n1481 ;
  assign n4152 = n4150 & n4151 ;
  assign n4279 = n4278 ^ n4152 ;
  assign n9575 = n4279 ^ n4151 ;
  assign n9577 = n4149 & n9575 ;
  assign n9578 = n9577 ^ n4279 ;
  assign n9579 = ~n9574 & ~n9578 ;
  assign n12434 = n9605 ^ n9579 ;
  assign n9606 = n4151 ^ n4140 ;
  assign n9607 = ~n4149 & ~n9606 ;
  assign n9608 = n9607 ^ n4151 ;
  assign n12435 = n9608 ^ n9579 ;
  assign n12436 = ~n12434 & n12435 ;
  assign n12437 = n12436 ^ n9579 ;
  assign n12438 = ~n11492 & ~n12437 ;
  assign n9609 = n4144 ^ n1473 ;
  assign n9610 = n9609 ^ n4142 ;
  assign n9611 = n4142 ^ n1475 ;
  assign n9612 = ~n4144 & n9611 ;
  assign n9617 = x944 & n9612 ;
  assign n9618 = n9617 ^ n9609 ;
  assign n9619 = ~n9610 & n9618 ;
  assign n9620 = n9619 ^ n4142 ;
  assign n9624 = ~n4142 & n9609 ;
  assign n9621 = x948 & n4141 ;
  assign n9622 = ~n9609 & n9621 ;
  assign n9623 = n9622 ^ n4141 ;
  assign n9625 = n9624 ^ n9623 ;
  assign n9626 = n9624 ^ n9612 ;
  assign n9627 = ~n9625 & n9626 ;
  assign n9635 = ~n1472 & n9627 ;
  assign n9636 = ~n9624 & n9635 ;
  assign n9637 = n9636 ^ n9624 ;
  assign n9628 = n9627 ^ n9623 ;
  assign n9629 = n9628 ^ n9624 ;
  assign n9638 = n9637 ^ n9629 ;
  assign n9639 = ~n9620 & ~n9638 ;
  assign n9640 = n4138 ^ n1478 ;
  assign n9641 = n9640 ^ n4136 ;
  assign n9642 = n4136 ^ n1480 ;
  assign n9643 = ~n4138 & n9642 ;
  assign n9648 = x950 & n9643 ;
  assign n9649 = n9648 ^ n9640 ;
  assign n9650 = ~n9641 & n9649 ;
  assign n9651 = n9650 ^ n4136 ;
  assign n9655 = ~n4136 & n9640 ;
  assign n9652 = x954 & n4135 ;
  assign n9653 = ~n9640 & n9652 ;
  assign n9654 = n9653 ^ n4135 ;
  assign n9656 = n9655 ^ n9654 ;
  assign n9657 = n9655 ^ n9643 ;
  assign n9658 = ~n9656 & n9657 ;
  assign n9666 = ~n1477 & n9658 ;
  assign n9667 = ~n9655 & n9666 ;
  assign n9668 = n9667 ^ n9655 ;
  assign n9659 = n9658 ^ n9654 ;
  assign n9660 = n9659 ^ n9655 ;
  assign n9669 = n9668 ^ n9660 ;
  assign n9670 = ~n9651 & ~n9669 ;
  assign n11496 = n9639 & n9670 ;
  assign n9671 = n9670 ^ n9639 ;
  assign n11497 = n11496 ^ n9671 ;
  assign n11504 = ~n9608 & n11496 ;
  assign n9672 = n9671 ^ n9608 ;
  assign n9673 = n9672 ^ n9605 ;
  assign n9674 = n9673 ^ n9579 ;
  assign n11493 = n9674 ^ n9605 ;
  assign n11500 = ~n9579 & n11497 ;
  assign n11501 = n11500 ^ n9674 ;
  assign n11502 = n11493 & n11501 ;
  assign n11503 = n11502 ^ n11492 ;
  assign n11505 = n11504 ^ n11503 ;
  assign n12439 = n11497 & ~n11505 ;
  assign n12440 = ~n12438 & n12439 ;
  assign n12441 = n12440 ^ n12438 ;
  assign n12442 = n12441 ^ n11471 ;
  assign n12447 = n12446 ^ n12442 ;
  assign n12448 = n12447 ^ n12441 ;
  assign n12449 = n11484 & ~n12448 ;
  assign n12452 = n12433 & n12449 ;
  assign n12450 = n12449 ^ n12447 ;
  assign n12453 = n12452 ^ n12450 ;
  assign n1494 = n1493 ^ n1482 ;
  assign n1517 = n1516 ^ n1505 ;
  assign n4439 = n1494 & n1517 ;
  assign n4438 = n4437 ^ n4373 ;
  assign n4440 = n4439 ^ n4438 ;
  assign n9675 = n9674 ^ n4439 ;
  assign n4280 = n4279 ^ n4149 ;
  assign n9676 = n9675 ^ n4280 ;
  assign n9677 = n9676 ^ n9674 ;
  assign n9678 = ~n4440 & n9677 ;
  assign n9679 = n9678 ^ n9675 ;
  assign n11486 = n11484 ^ n9674 ;
  assign n11485 = n11484 ^ n9716 ;
  assign n11487 = n11486 ^ n11485 ;
  assign n11488 = ~n9679 & ~n11487 ;
  assign n11489 = n11488 ^ n11486 ;
  assign n12454 = n11505 ^ n11484 ;
  assign n12455 = ~n11489 & ~n12454 ;
  assign n12456 = n12455 ^ n11484 ;
  assign n13035 = n12456 ^ n12441 ;
  assign n13036 = n12453 & ~n13035 ;
  assign n13037 = n13036 ^ n12441 ;
  assign n1463 = x62 ^ x61 ;
  assign n4620 = ~x63 & ~x64 ;
  assign n4618 = x65 & x66 ;
  assign n4626 = n4620 ^ n4618 ;
  assign n1464 = x64 ^ x63 ;
  assign n4623 = n1464 & n4618 ;
  assign n4627 = n4626 ^ n4623 ;
  assign n4631 = n4627 ^ x62 ;
  assign n4621 = n4620 ^ n1464 ;
  assign n1466 = x66 ^ x65 ;
  assign n4619 = n4618 ^ n1466 ;
  assign n4628 = n4621 ^ n4619 ;
  assign n4622 = n4619 & ~n4621 ;
  assign n4629 = n4628 ^ n4622 ;
  assign n4632 = n4631 ^ n4629 ;
  assign n4633 = n1463 & ~n4632 ;
  assign n4634 = n4633 ^ x61 ;
  assign n4630 = ~n4627 & ~n4629 ;
  assign n4636 = n4634 ^ n4630 ;
  assign n4635 = ~n4630 & ~n4634 ;
  assign n4637 = n4636 ^ n4635 ;
  assign n4624 = n4623 ^ n4622 ;
  assign n4625 = n1463 & n4624 ;
  assign n4638 = n4637 ^ n4625 ;
  assign n4639 = n4638 ^ n4635 ;
  assign n4582 = ~x57 & ~x58 ;
  assign n4581 = ~x59 & ~x60 ;
  assign n1461 = x60 ^ x59 ;
  assign n4585 = n4581 ^ n1461 ;
  assign n4586 = ~n4582 & ~n4585 ;
  assign n1459 = x58 ^ x57 ;
  assign n4583 = n4582 ^ n1459 ;
  assign n4584 = ~n4581 & ~n4583 ;
  assign n4588 = n4586 ^ n4584 ;
  assign n4587 = ~n4584 & ~n4586 ;
  assign n4589 = n4588 ^ n4587 ;
  assign n4590 = ~x55 & n4589 ;
  assign n4591 = n4583 ^ n4581 ;
  assign n4592 = n4591 ^ n4584 ;
  assign n4593 = n4592 ^ x56 ;
  assign n4594 = n4585 ^ n4582 ;
  assign n4595 = n4594 ^ n4586 ;
  assign n4596 = n4595 ^ x56 ;
  assign n4597 = n4593 & n4596 ;
  assign n4598 = n4597 ^ x56 ;
  assign n4599 = n4590 & n4598 ;
  assign n4600 = n4599 ^ x55 ;
  assign n4613 = ~x56 & n4582 ;
  assign n4614 = ~n4592 & n4613 ;
  assign n4615 = n4614 ^ n4592 ;
  assign n1458 = x56 ^ x55 ;
  assign n4601 = n4592 ^ n4589 ;
  assign n4602 = x56 & n4595 ;
  assign n4603 = ~n4601 & n4602 ;
  assign n4604 = n4603 ^ n4587 ;
  assign n4605 = ~n1458 & ~n4604 ;
  assign n4606 = n4605 ^ n4587 ;
  assign n4607 = n4606 ^ n4592 ;
  assign n4616 = n4615 ^ n4607 ;
  assign n4617 = n4600 & n4616 ;
  assign n4640 = n4639 ^ n4617 ;
  assign n1460 = n1459 ^ n1458 ;
  assign n1462 = n1461 ^ n1460 ;
  assign n1465 = n1464 ^ n1463 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n4580 = n1462 & n1467 ;
  assign n9530 = n4639 ^ n4580 ;
  assign n9531 = n4640 & n9530 ;
  assign n9532 = n9531 ^ n4639 ;
  assign n1450 = x72 ^ x71 ;
  assign n1448 = x70 ^ x69 ;
  assign n1447 = x68 ^ x67 ;
  assign n1449 = n1448 ^ n1447 ;
  assign n1451 = n1450 ^ n1449 ;
  assign n1455 = x78 ^ x77 ;
  assign n1453 = x76 ^ x75 ;
  assign n1452 = x74 ^ x73 ;
  assign n1454 = n1453 ^ n1452 ;
  assign n1456 = n1455 ^ n1454 ;
  assign n9517 = n1451 & n1456 ;
  assign n4687 = x77 ^ x76 ;
  assign n4691 = ~n1455 & ~n4687 ;
  assign n4686 = x75 ^ x74 ;
  assign n4688 = n4687 ^ x75 ;
  assign n4689 = n4688 ^ x78 ;
  assign n4690 = ~n4686 & n4689 ;
  assign n4692 = n4691 ^ n4690 ;
  assign n4693 = ~x73 & n4692 ;
  assign n4694 = ~n1453 & ~n4686 ;
  assign n4695 = x78 ^ x73 ;
  assign n4698 = ~x76 & ~n4695 ;
  assign n4699 = n4698 ^ x73 ;
  assign n4700 = n4694 & n4699 ;
  assign n4701 = ~x77 & n4700 ;
  assign n4702 = ~x75 & ~x76 ;
  assign n4705 = n4702 ^ n1453 ;
  assign n4706 = x73 & x74 ;
  assign n4707 = x78 & n4706 ;
  assign n4708 = ~n4705 & n4707 ;
  assign n4709 = n4708 ^ n4706 ;
  assign n4703 = ~x77 & ~x78 ;
  assign n4704 = ~n4702 & ~n4703 ;
  assign n4710 = n4709 ^ n4704 ;
  assign n4711 = n4703 ^ n1455 ;
  assign n4716 = n4705 & n4711 ;
  assign n4717 = n4716 ^ n4704 ;
  assign n4718 = n4710 & n4717 ;
  assign n4719 = n4718 ^ n4709 ;
  assign n4720 = ~n1452 & n4719 ;
  assign n4721 = n4718 & n4720 ;
  assign n4722 = n4721 ^ n4719 ;
  assign n4723 = ~n4701 & ~n4722 ;
  assign n4724 = ~n4693 & n4723 ;
  assign n4648 = x71 ^ x70 ;
  assign n4652 = ~n1450 & ~n4648 ;
  assign n4647 = x69 ^ x68 ;
  assign n4649 = n4648 ^ x69 ;
  assign n4650 = n4649 ^ x72 ;
  assign n4651 = ~n4647 & n4650 ;
  assign n4653 = n4652 ^ n4651 ;
  assign n4654 = ~x67 & n4653 ;
  assign n4655 = ~n1448 & ~n4647 ;
  assign n4656 = x72 ^ x67 ;
  assign n4659 = ~x70 & ~n4656 ;
  assign n4660 = n4659 ^ x67 ;
  assign n4661 = n4655 & n4660 ;
  assign n4662 = ~x71 & n4661 ;
  assign n4663 = ~x69 & ~x70 ;
  assign n4666 = n4663 ^ n1448 ;
  assign n4667 = x67 & x68 ;
  assign n4668 = x72 & n4667 ;
  assign n4669 = ~n4666 & n4668 ;
  assign n4670 = n4669 ^ n4667 ;
  assign n4664 = ~x71 & ~x72 ;
  assign n4665 = ~n4663 & ~n4664 ;
  assign n4671 = n4670 ^ n4665 ;
  assign n4672 = n4664 ^ n1450 ;
  assign n4677 = n4666 & n4672 ;
  assign n4678 = n4677 ^ n4665 ;
  assign n4679 = n4671 & n4678 ;
  assign n4680 = n4679 ^ n4670 ;
  assign n4681 = ~n1447 & n4680 ;
  assign n4682 = n4679 & n4681 ;
  assign n4683 = n4682 ^ n4680 ;
  assign n4684 = ~n4662 & ~n4683 ;
  assign n4685 = ~n4654 & n4684 ;
  assign n4725 = n4724 ^ n4685 ;
  assign n9518 = n9517 ^ n4725 ;
  assign n1457 = n1456 ^ n1451 ;
  assign n1468 = n1467 ^ n1462 ;
  assign n4644 = n1468 ^ n1451 ;
  assign n4645 = ~n1457 & n4644 ;
  assign n4641 = n4640 ^ n4580 ;
  assign n4642 = n4641 ^ n1468 ;
  assign n4646 = n4645 ^ n4642 ;
  assign n4726 = n4725 ^ n4646 ;
  assign n9516 = n4726 ^ n4580 ;
  assign n9519 = n9518 ^ n9516 ;
  assign n9520 = ~n4640 & ~n9519 ;
  assign n9521 = n9520 ^ n4580 ;
  assign n9522 = n9518 ^ n4646 ;
  assign n9523 = n9520 ^ n9519 ;
  assign n9524 = ~n9522 & ~n9523 ;
  assign n9525 = n9524 ^ n4646 ;
  assign n9526 = n9525 ^ n9522 ;
  assign n9527 = n9521 & n9526 ;
  assign n9528 = n9527 ^ n9524 ;
  assign n9529 = n9528 ^ n9518 ;
  assign n11551 = n9532 ^ n9529 ;
  assign n9533 = n4618 & ~n4621 ;
  assign n9534 = n4638 & n9533 ;
  assign n9535 = n9534 ^ n4638 ;
  assign n11562 = n9535 ^ n9532 ;
  assign n9536 = n4589 & n4606 ;
  assign n9537 = n9536 ^ n9535 ;
  assign n11555 = n9537 ^ n9529 ;
  assign n11556 = n11555 ^ n9532 ;
  assign n11563 = n11562 ^ n11556 ;
  assign n11553 = ~n11551 & ~n11563 ;
  assign n11554 = n11553 ^ n9536 ;
  assign n9553 = n9517 ^ n4724 ;
  assign n9554 = n4725 & n9553 ;
  assign n9555 = n9554 ^ n4724 ;
  assign n9545 = n4711 ^ n4705 ;
  assign n9546 = x74 & n4704 ;
  assign n9547 = n9546 ^ n4705 ;
  assign n9548 = n9545 & ~n9547 ;
  assign n9549 = n9548 ^ n4705 ;
  assign n9550 = ~n4722 & ~n9549 ;
  assign n9551 = n9550 ^ n4722 ;
  assign n9539 = n4672 ^ n4666 ;
  assign n9540 = x68 & n4665 ;
  assign n9541 = n9540 ^ n4666 ;
  assign n9542 = n9539 & ~n9541 ;
  assign n9543 = n9542 ^ n4666 ;
  assign n9544 = ~n4683 & n9543 ;
  assign n9552 = n9551 ^ n9544 ;
  assign n9556 = n9555 ^ n9552 ;
  assign n11557 = n9556 ^ n9535 ;
  assign n9538 = n9537 ^ n9532 ;
  assign n11559 = n11557 ^ n9538 ;
  assign n11560 = n9535 ^ n9529 ;
  assign n11561 = n11560 ^ n11557 ;
  assign n11564 = n11561 & n11563 ;
  assign n11565 = ~n11559 & n11564 ;
  assign n11566 = n11565 ^ n9535 ;
  assign n11567 = n11566 ^ n11556 ;
  assign n11568 = n11557 & ~n11567 ;
  assign n11569 = n11556 & n11568 ;
  assign n11570 = n11569 ^ n9535 ;
  assign n12397 = n11554 & n11570 ;
  assign n9557 = n9556 ^ n9538 ;
  assign n9558 = n9557 ^ n9529 ;
  assign n11575 = ~n9556 & n9558 ;
  assign n11576 = n11575 ^ n11570 ;
  assign n11577 = ~n11554 & n11576 ;
  assign n11578 = n11577 ^ n11570 ;
  assign n11579 = n9555 ^ n9551 ;
  assign n11580 = ~n9552 & n11579 ;
  assign n11581 = n11580 ^ n9551 ;
  assign n12396 = ~n11578 & ~n11581 ;
  assign n12398 = n12397 ^ n12396 ;
  assign n4496 = ~x39 & ~x40 ;
  assign n1425 = x40 ^ x39 ;
  assign n9490 = n4496 ^ n1425 ;
  assign n4492 = x37 & x38 ;
  assign n9491 = x42 & n4492 ;
  assign n9492 = ~n9490 & n9491 ;
  assign n9493 = n9492 ^ n4492 ;
  assign n4494 = ~x41 & ~x42 ;
  assign n9488 = ~n4494 & ~n4496 ;
  assign n9494 = n9493 ^ n9488 ;
  assign n1427 = x42 ^ x41 ;
  assign n9495 = n4494 ^ n1427 ;
  assign n9500 = n9490 & n9495 ;
  assign n9501 = n9500 ^ n9488 ;
  assign n9502 = n9494 & n9501 ;
  assign n9504 = n9502 ^ n9493 ;
  assign n1424 = x38 ^ x37 ;
  assign n9489 = ~n1424 & n9488 ;
  assign n9503 = n9489 & n9502 ;
  assign n9505 = n9504 ^ n9503 ;
  assign n9506 = n9495 ^ n9490 ;
  assign n9507 = x38 & n9488 ;
  assign n9508 = n9507 ^ n9490 ;
  assign n9509 = n9506 & ~n9508 ;
  assign n9510 = n9509 ^ n9490 ;
  assign n9511 = ~n9505 & ~n9510 ;
  assign n9512 = n9511 ^ n9505 ;
  assign n4447 = x35 & x36 ;
  assign n4450 = ~x33 & ~x34 ;
  assign n1431 = x34 ^ x33 ;
  assign n4458 = n4450 ^ n1431 ;
  assign n4502 = ~n4447 & n4458 ;
  assign n4466 = x35 ^ x32 ;
  assign n4467 = n4466 ^ x34 ;
  assign n4468 = n4467 ^ x36 ;
  assign n4464 = x35 ^ x33 ;
  assign n4469 = n4468 ^ n4464 ;
  assign n4470 = n4469 ^ x36 ;
  assign n4471 = n4470 ^ x35 ;
  assign n4472 = n4471 ^ n4464 ;
  assign n4476 = n4464 ^ x34 ;
  assign n4477 = n4476 ^ x36 ;
  assign n4478 = n4477 ^ n4464 ;
  assign n4479 = ~n4472 & ~n4478 ;
  assign n4480 = ~x35 & n4479 ;
  assign n4483 = n4480 ^ n4479 ;
  assign n4481 = n4480 ^ n4464 ;
  assign n4482 = n4469 & n4481 ;
  assign n4484 = n4483 ^ n4482 ;
  assign n4485 = n4484 ^ x35 ;
  assign n4504 = x31 & n4485 ;
  assign n4503 = n4485 ^ x31 ;
  assign n4505 = n4504 ^ n4503 ;
  assign n4506 = n4502 & ~n4505 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n4498 = n1427 ^ n1425 ;
  assign n4499 = ~n1426 & n4498 ;
  assign n4493 = n4492 ^ n1425 ;
  assign n4495 = n4494 ^ n4493 ;
  assign n4497 = n4496 ^ n4495 ;
  assign n4500 = n4499 ^ n4497 ;
  assign n4501 = n4500 ^ n4485 ;
  assign n4507 = n4506 ^ n4501 ;
  assign n4459 = n4458 ^ n4447 ;
  assign n1430 = x36 ^ x35 ;
  assign n4448 = n4447 ^ n1430 ;
  assign n4449 = n4448 ^ x32 ;
  assign n4451 = n4450 ^ n4449 ;
  assign n4460 = n4451 ^ n4447 ;
  assign n4453 = ~n4448 & n4450 ;
  assign n4452 = n4450 ^ n4448 ;
  assign n4454 = n4453 ^ n4452 ;
  assign n4455 = ~n4451 & ~n4454 ;
  assign n4461 = n4460 ^ n4455 ;
  assign n4462 = ~n4459 & n4461 ;
  assign n4463 = n4462 ^ n4458 ;
  assign n4489 = ~x31 & ~n4484 ;
  assign n4490 = n4489 ^ x35 ;
  assign n4491 = ~n4463 & ~n4490 ;
  assign n4508 = n4507 ^ n4491 ;
  assign n4456 = n4453 ^ x31 ;
  assign n4457 = ~n4455 & ~n4456 ;
  assign n4509 = n4508 ^ n4457 ;
  assign n9482 = n4463 & ~n4504 ;
  assign n1428 = n1427 ^ n1426 ;
  assign n1429 = x32 ^ x31 ;
  assign n1433 = n4477 ^ n1429 ;
  assign n4517 = n1428 & n1433 ;
  assign n9483 = n9482 ^ n4517 ;
  assign n9484 = n9483 ^ n4500 ;
  assign n9485 = n9484 ^ n9482 ;
  assign n9486 = n4509 & n9485 ;
  assign n9487 = n9486 ^ n9483 ;
  assign n9513 = n9512 ^ n9487 ;
  assign n4570 = x51 & x52 ;
  assign n4569 = x53 & x54 ;
  assign n4571 = n4570 ^ n4569 ;
  assign n1438 = x54 ^ x53 ;
  assign n4572 = n4569 ^ n1438 ;
  assign n1436 = x52 ^ x51 ;
  assign n4573 = n4570 ^ n1436 ;
  assign n4574 = n4572 & n4573 ;
  assign n4575 = n4574 ^ n4570 ;
  assign n4576 = ~n4571 & ~n4575 ;
  assign n4522 = n1438 ^ x50 ;
  assign n4523 = n4522 ^ n1436 ;
  assign n1443 = x48 ^ x47 ;
  assign n4525 = x47 ^ x46 ;
  assign n4529 = ~n1443 & ~n4525 ;
  assign n4524 = x45 ^ x44 ;
  assign n4526 = n4525 ^ x45 ;
  assign n4527 = n4526 ^ x48 ;
  assign n4528 = ~n4524 & n4527 ;
  assign n4530 = n4529 ^ n4528 ;
  assign n4531 = ~x43 & n4530 ;
  assign n1441 = x46 ^ x45 ;
  assign n4532 = ~n1441 & ~n4524 ;
  assign n4533 = x48 ^ x43 ;
  assign n4536 = ~x46 & ~n4533 ;
  assign n4537 = n4536 ^ x43 ;
  assign n4538 = n4532 & n4537 ;
  assign n4539 = ~x47 & n4538 ;
  assign n4540 = ~x45 & ~x46 ;
  assign n4543 = n4540 ^ n1441 ;
  assign n4544 = x43 & x44 ;
  assign n4545 = x48 & n4544 ;
  assign n4546 = ~n4543 & n4545 ;
  assign n4547 = n4546 ^ n4544 ;
  assign n4541 = ~x47 & ~x48 ;
  assign n4542 = ~n4540 & ~n4541 ;
  assign n4548 = n4547 ^ n4542 ;
  assign n4549 = n4541 ^ n1443 ;
  assign n4554 = n4543 & n4549 ;
  assign n4555 = n4554 ^ n4542 ;
  assign n4556 = n4548 & n4555 ;
  assign n1440 = x44 ^ x43 ;
  assign n4557 = n4556 ^ n4547 ;
  assign n4558 = ~n1440 & n4557 ;
  assign n4559 = n4556 & n4558 ;
  assign n4560 = n4559 ^ n4557 ;
  assign n4561 = ~n4539 & ~n4560 ;
  assign n4562 = ~n4531 & n4561 ;
  assign n4563 = n4562 ^ x49 ;
  assign n4564 = n4563 ^ n1438 ;
  assign n4565 = n4564 ^ n1436 ;
  assign n4566 = n4565 ^ n4562 ;
  assign n4567 = ~n4523 & n4566 ;
  assign n4568 = n4567 ^ n4563 ;
  assign n4577 = n4576 ^ n4568 ;
  assign n1435 = x50 ^ x49 ;
  assign n1437 = n1436 ^ n1435 ;
  assign n1439 = n1438 ^ n1437 ;
  assign n1442 = n1441 ^ n1440 ;
  assign n1444 = n1443 ^ n1442 ;
  assign n9447 = n1439 & n1444 ;
  assign n9477 = n9447 ^ n4562 ;
  assign n9478 = ~n4577 & n9477 ;
  assign n9479 = n9478 ^ n4562 ;
  assign n9465 = n4574 ^ x50 ;
  assign n9466 = n4571 ^ x49 ;
  assign n9467 = n9466 ^ n4574 ;
  assign n9468 = n9465 & ~n9467 ;
  assign n9471 = n9468 ^ n4574 ;
  assign n9469 = n9468 ^ n4575 ;
  assign n9470 = ~n4571 & n9469 ;
  assign n9472 = n9471 ^ n9470 ;
  assign n9473 = x49 & n9470 ;
  assign n9474 = ~n9472 & n9473 ;
  assign n9475 = n9474 ^ n9472 ;
  assign n9459 = n4549 ^ n4543 ;
  assign n9460 = x44 & n4542 ;
  assign n9461 = n9460 ^ n4543 ;
  assign n9462 = n9459 & ~n9461 ;
  assign n9463 = n9462 ^ n4543 ;
  assign n9464 = ~n4560 & n9463 ;
  assign n9476 = n9475 ^ n9464 ;
  assign n9480 = n9479 ^ n9476 ;
  assign n4510 = n1444 ^ n1433 ;
  assign n4511 = n4510 ^ n1428 ;
  assign n1445 = n1444 ^ n1439 ;
  assign n4512 = ~n1445 & ~n4510 ;
  assign n4513 = n4511 & n4512 ;
  assign n4514 = n4513 ^ n1428 ;
  assign n4518 = n4517 ^ n4512 ;
  assign n4515 = n1445 ^ n1433 ;
  assign n4516 = ~n4514 & n4515 ;
  assign n4519 = n4518 ^ n4516 ;
  assign n4520 = ~n4514 & n4519 ;
  assign n4521 = n4520 ^ n4509 ;
  assign n9448 = n9447 ^ n4521 ;
  assign n9450 = ~n4577 & n9448 ;
  assign n9451 = n9450 ^ n4521 ;
  assign n9456 = n4509 & n4519 ;
  assign n9457 = n9456 ^ n4517 ;
  assign n9458 = ~n9451 & ~n9457 ;
  assign n9481 = n9480 ^ n9458 ;
  assign n9514 = n9513 ^ n9481 ;
  assign n9559 = n9558 ^ n9514 ;
  assign n1434 = n1433 ^ n1428 ;
  assign n1446 = n1445 ^ n1434 ;
  assign n1469 = n1468 ^ n1457 ;
  assign n4579 = n1446 & n1469 ;
  assign n4727 = n4726 ^ n4579 ;
  assign n4578 = n4577 ^ n4521 ;
  assign n9444 = n4726 ^ n4578 ;
  assign n9445 = n4727 & ~n9444 ;
  assign n9446 = n9445 ^ n4726 ;
  assign n11547 = n9558 ^ n9446 ;
  assign n11548 = ~n9559 & ~n11547 ;
  assign n11549 = n11548 ^ n9558 ;
  assign n11536 = n9512 ^ n9482 ;
  assign n11537 = ~n9487 & ~n11536 ;
  assign n11538 = n11537 ^ n9482 ;
  assign n11539 = n9479 ^ n9475 ;
  assign n11540 = ~n9476 & n11539 ;
  assign n11541 = n11540 ^ n9475 ;
  assign n11543 = n9513 ^ n9480 ;
  assign n11544 = ~n9481 & n11543 ;
  assign n11545 = n11544 ^ n9480 ;
  assign n12402 = n11541 & ~n11545 ;
  assign n12403 = ~n11538 & n12402 ;
  assign n11542 = n11541 ^ n11538 ;
  assign n12404 = n12403 ^ n11542 ;
  assign n12399 = n11545 ^ n11538 ;
  assign n12400 = n11542 & n12399 ;
  assign n12405 = n12404 ^ n12400 ;
  assign n12406 = n11549 & n12405 ;
  assign n12401 = n12400 ^ n11542 ;
  assign n11582 = n11581 ^ n11578 ;
  assign n12409 = n12400 ^ n11545 ;
  assign n12407 = n12405 ^ n11549 ;
  assign n12408 = n12407 ^ n12406 ;
  assign n12411 = n12409 ^ n12408 ;
  assign n12410 = n12408 & n12409 ;
  assign n12412 = n12411 ^ n12410 ;
  assign n12413 = ~n11582 & n12412 ;
  assign n12414 = ~n12398 & n12413 ;
  assign n12415 = ~n12401 & n12414 ;
  assign n12416 = n12415 ^ n12413 ;
  assign n12423 = n12403 & n12416 ;
  assign n12417 = n12410 ^ n12397 ;
  assign n12418 = n11582 & n12417 ;
  assign n12419 = ~n12416 & ~n12418 ;
  assign n12424 = n12423 ^ n12419 ;
  assign n12425 = ~n12406 & ~n12424 ;
  assign n12426 = n12425 ^ n12419 ;
  assign n12427 = n12398 & ~n12426 ;
  assign n12428 = n12427 ^ n12419 ;
  assign n9560 = n9559 ^ n9446 ;
  assign n1413 = x999 ^ x998 ;
  assign n4951 = x998 ^ x997 ;
  assign n4952 = ~n1413 & n4951 ;
  assign n4953 = n4952 ^ x997 ;
  assign n1408 = x2 ^ x1 ;
  assign n1409 = n1408 ^ x0 ;
  assign n1410 = x5 ^ x4 ;
  assign n1411 = n1410 ^ x3 ;
  assign n4941 = n1409 & n1411 ;
  assign n9262 = n4953 ^ n4941 ;
  assign n1412 = n1411 ^ n1409 ;
  assign n1414 = n1413 ^ x997 ;
  assign n1415 = n1414 ^ x6 ;
  assign n4939 = n1412 & n1415 ;
  assign n9263 = n9262 ^ n4939 ;
  assign n4943 = x1 ^ x0 ;
  assign n4944 = ~n1408 & n4943 ;
  assign n4945 = n4944 ^ x0 ;
  assign n4946 = n4945 ^ x3 ;
  assign n4947 = n4946 ^ x4 ;
  assign n4948 = n4947 ^ n4945 ;
  assign n4949 = ~n1410 & n4948 ;
  assign n4950 = n4949 ^ n4946 ;
  assign n9264 = n9263 ^ n4950 ;
  assign n9265 = n9264 ^ n4953 ;
  assign n4938 = x6 & n1414 ;
  assign n9269 = n9265 ^ n4938 ;
  assign n9275 = n9269 ^ n4953 ;
  assign n1416 = n1415 ^ n1412 ;
  assign n1420 = x996 ^ x995 ;
  assign n1418 = x994 ^ x993 ;
  assign n1417 = x992 ^ x991 ;
  assign n1419 = n1418 ^ n1417 ;
  assign n1421 = n1420 ^ n1419 ;
  assign n4937 = n1416 & n1421 ;
  assign n4956 = n9275 ^ n4937 ;
  assign n4899 = x995 ^ x994 ;
  assign n4903 = ~n1420 & ~n4899 ;
  assign n4898 = x993 ^ x992 ;
  assign n4900 = n4899 ^ x993 ;
  assign n4901 = n4900 ^ x996 ;
  assign n4902 = ~n4898 & n4901 ;
  assign n4904 = n4903 ^ n4902 ;
  assign n4905 = ~x991 & n4904 ;
  assign n4906 = ~n1418 & ~n4898 ;
  assign n4907 = x996 ^ x991 ;
  assign n4910 = ~x994 & ~n4907 ;
  assign n4911 = n4910 ^ x991 ;
  assign n4912 = n4906 & n4911 ;
  assign n4913 = ~x995 & n4912 ;
  assign n4914 = ~x993 & ~x994 ;
  assign n4917 = n4914 ^ n1418 ;
  assign n4918 = x991 & x992 ;
  assign n4919 = x996 & n4918 ;
  assign n4920 = ~n4917 & n4919 ;
  assign n4921 = n4920 ^ n4918 ;
  assign n4915 = ~x995 & ~x996 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4922 = n4921 ^ n4916 ;
  assign n4923 = n4915 ^ n1420 ;
  assign n4928 = n4917 & n4923 ;
  assign n4929 = n4928 ^ n4916 ;
  assign n4930 = n4922 & n4929 ;
  assign n4931 = n4930 ^ n4921 ;
  assign n4932 = ~n1417 & n4931 ;
  assign n4933 = n4930 & n4932 ;
  assign n4934 = n4933 ^ n4931 ;
  assign n4935 = ~n4913 & ~n4934 ;
  assign n4936 = ~n4905 & n4935 ;
  assign n4957 = n4956 ^ n4936 ;
  assign n4847 = x11 & x12 ;
  assign n1399 = x12 ^ x11 ;
  assign n4849 = n4847 ^ n1399 ;
  assign n4850 = x8 & n4849 ;
  assign n4848 = n4847 ^ x10 ;
  assign n4853 = n4850 ^ n4848 ;
  assign n4854 = x9 & ~n4853 ;
  assign n4851 = n4850 ^ n4847 ;
  assign n4852 = ~n4848 & ~n4851 ;
  assign n4855 = n4854 ^ n4852 ;
  assign n4856 = ~x7 & n4855 ;
  assign n1397 = x10 ^ x9 ;
  assign n4857 = x7 & n1397 ;
  assign n4858 = ~x11 & ~n4857 ;
  assign n4859 = ~x9 & ~x10 ;
  assign n4860 = n4859 ^ n1397 ;
  assign n4861 = n4860 ^ x8 ;
  assign n4862 = x12 ^ x7 ;
  assign n4865 = n4860 & ~n4862 ;
  assign n4866 = n4865 ^ x7 ;
  assign n4867 = n4861 & n4866 ;
  assign n4868 = n4858 & n4867 ;
  assign n4873 = n4849 & ~n4859 ;
  assign n1396 = x8 ^ x7 ;
  assign n4869 = n1396 ^ x12 ;
  assign n4870 = x9 & n4869 ;
  assign n4874 = n4873 ^ n4870 ;
  assign n4875 = ~x8 & ~n4874 ;
  assign n4876 = n4875 ^ n4870 ;
  assign n4877 = x7 & ~n4876 ;
  assign n4884 = ~n4847 & n4860 ;
  assign n4878 = n4857 ^ n4850 ;
  assign n4879 = n4878 ^ n4877 ;
  assign n4885 = n4884 ^ n4879 ;
  assign n4886 = n4877 & n4885 ;
  assign n4887 = n4886 ^ n4879 ;
  assign n4888 = n4887 ^ n4877 ;
  assign n4889 = n4877 ^ n4857 ;
  assign n4890 = ~n4886 & ~n4889 ;
  assign n4891 = ~n4888 & n4890 ;
  assign n4892 = n4891 ^ n4887 ;
  assign n4893 = ~n4868 & n4892 ;
  assign n4894 = ~n4856 & n4893 ;
  assign n1403 = x16 ^ x15 ;
  assign n4807 = x15 ^ x14 ;
  assign n4808 = ~n1403 & ~n4807 ;
  assign n4809 = x18 ^ x13 ;
  assign n4812 = ~x16 & ~n4809 ;
  assign n4813 = n4812 ^ x13 ;
  assign n4814 = n4808 & n4813 ;
  assign n4815 = ~x17 & n4814 ;
  assign n1402 = x18 ^ x17 ;
  assign n4838 = x17 ^ x16 ;
  assign n4842 = ~n1402 & ~n4838 ;
  assign n1404 = n1403 ^ n1402 ;
  assign n4840 = n1404 & ~n4807 ;
  assign n4817 = x15 & x16 ;
  assign n4823 = n4817 ^ n1403 ;
  assign n4824 = ~x17 & ~x18 ;
  assign n4825 = n4824 ^ n1402 ;
  assign n4826 = n4823 & ~n4825 ;
  assign n4827 = n4824 ^ x14 ;
  assign n4828 = ~n4826 & ~n4827 ;
  assign n4816 = n1403 ^ x17 ;
  assign n4818 = n4817 ^ x18 ;
  assign n4819 = n4818 ^ n1403 ;
  assign n4820 = ~n4817 & n4819 ;
  assign n4821 = ~n4816 & n4820 ;
  assign n4822 = n4821 ^ n4818 ;
  assign n4829 = n4824 ^ n4822 ;
  assign n4830 = n4829 ^ n4817 ;
  assign n4831 = n4830 ^ n4822 ;
  assign n4832 = n4831 ^ x13 ;
  assign n4833 = n4828 & n4832 ;
  assign n4834 = n4833 ^ n4829 ;
  assign n4835 = ~x14 & ~n4834 ;
  assign n4836 = n4835 ^ n4822 ;
  assign n4841 = n4840 ^ n4836 ;
  assign n4843 = n4842 ^ n4841 ;
  assign n4844 = ~x13 & n4843 ;
  assign n4845 = n4844 ^ n4836 ;
  assign n4846 = ~n4815 & ~n4845 ;
  assign n4895 = n4894 ^ n4846 ;
  assign n1388 = x24 ^ x23 ;
  assign n4779 = x23 ^ x22 ;
  assign n4783 = ~n1388 & ~n4779 ;
  assign n4778 = x21 ^ x20 ;
  assign n4780 = n4779 ^ x21 ;
  assign n4781 = n4780 ^ x24 ;
  assign n4782 = ~n4778 & n4781 ;
  assign n4784 = n4783 ^ n4782 ;
  assign n4785 = ~x19 & n4784 ;
  assign n4786 = ~x21 & ~x22 ;
  assign n4787 = ~x23 & ~x24 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4789 = n4788 ^ x20 ;
  assign n1386 = x22 ^ x21 ;
  assign n4790 = n4786 ^ n1386 ;
  assign n4791 = n4787 ^ n1388 ;
  assign n4792 = n4790 & n4791 ;
  assign n4793 = n4792 ^ x20 ;
  assign n4794 = n4789 & ~n4793 ;
  assign n4795 = n4794 ^ x20 ;
  assign n4796 = x19 & ~n4795 ;
  assign n4797 = n4796 ^ x19 ;
  assign n4798 = n4797 ^ x23 ;
  assign n4799 = x24 ^ x22 ;
  assign n4800 = ~n1386 & ~n4778 ;
  assign n4801 = ~n4799 & n4800 ;
  assign n4802 = ~n4798 & ~n4801 ;
  assign n4803 = n4802 ^ x23 ;
  assign n4804 = ~n4785 & n4803 ;
  assign n1392 = x28 ^ x27 ;
  assign n4735 = x27 ^ x26 ;
  assign n4736 = ~n1392 & ~n4735 ;
  assign n4737 = x30 ^ x25 ;
  assign n4740 = ~x28 & ~n4737 ;
  assign n4741 = n4740 ^ x25 ;
  assign n4742 = n4736 & n4741 ;
  assign n4743 = ~x29 & n4742 ;
  assign n4757 = ~x29 & ~x30 ;
  assign n4760 = n4757 ^ x29 ;
  assign n4761 = n4760 ^ x30 ;
  assign n4750 = x27 & x28 ;
  assign n4756 = n4750 ^ n1392 ;
  assign n4759 = ~n4756 & ~n4761 ;
  assign n4762 = n4761 ^ n4759 ;
  assign n4763 = n4757 ^ x26 ;
  assign n4764 = n4762 & ~n4763 ;
  assign n4749 = n1392 ^ x29 ;
  assign n4751 = n4750 ^ x30 ;
  assign n4752 = n4751 ^ n1392 ;
  assign n4753 = ~n4750 & n4752 ;
  assign n4754 = ~n4749 & n4753 ;
  assign n4755 = n4754 ^ n4751 ;
  assign n4765 = n4757 ^ n4755 ;
  assign n4766 = n4765 ^ n4750 ;
  assign n4767 = n4766 ^ n4755 ;
  assign n4768 = n4767 ^ x25 ;
  assign n4769 = n4764 & n4768 ;
  assign n4770 = n4769 ^ n4765 ;
  assign n4771 = ~x26 & ~n4770 ;
  assign n4772 = n4771 ^ n4755 ;
  assign n1391 = x30 ^ x29 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n4748 = n1393 & ~n4735 ;
  assign n4773 = n4772 ^ n4748 ;
  assign n4744 = x29 ^ x28 ;
  assign n4745 = ~n1391 & ~n4744 ;
  assign n4774 = n4773 ^ n4745 ;
  assign n4775 = ~x25 & n4774 ;
  assign n4776 = n4775 ^ n4772 ;
  assign n4777 = ~n4743 & ~n4776 ;
  assign n4805 = n4804 ^ n4777 ;
  assign n1385 = x20 ^ x19 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1390 = x26 ^ x25 ;
  assign n1394 = n1393 ^ n1390 ;
  assign n4734 = n1389 & n1394 ;
  assign n4806 = n4805 ^ n4734 ;
  assign n4896 = n4895 ^ n4806 ;
  assign n1401 = x14 ^ x13 ;
  assign n1405 = n1404 ^ n1401 ;
  assign n1398 = n1397 ^ n1396 ;
  assign n1400 = n1399 ^ n1398 ;
  assign n1406 = n1405 ^ n1400 ;
  assign n1395 = n1394 ^ n1389 ;
  assign n1407 = n1406 ^ n1395 ;
  assign n1422 = n1421 ^ n1416 ;
  assign n4732 = n1407 & n1422 ;
  assign n4729 = n1400 ^ n1395 ;
  assign n4730 = n1406 & ~n4729 ;
  assign n4731 = n4730 ^ n1405 ;
  assign n4733 = n4732 ^ n4731 ;
  assign n4897 = n4896 ^ n4733 ;
  assign n4958 = n4957 ^ n4897 ;
  assign n4728 = n4727 ^ n4578 ;
  assign n4959 = n4958 ^ n4728 ;
  assign n1423 = n1422 ^ n1407 ;
  assign n1470 = n1469 ^ n1446 ;
  assign n9440 = n1423 & n1470 ;
  assign n9441 = n9440 ^ n4958 ;
  assign n9442 = ~n4959 & n9441 ;
  assign n9443 = n9442 ^ n4958 ;
  assign n9561 = n9560 ^ n9443 ;
  assign n9383 = n1400 & n1405 ;
  assign n9432 = n9383 ^ n4846 ;
  assign n9433 = n4895 & n9432 ;
  assign n9434 = n9433 ^ n4846 ;
  assign n9419 = x13 & n4836 ;
  assign n9421 = x14 & ~n4824 ;
  assign n9420 = n9419 ^ n4817 ;
  assign n9422 = n9421 ^ n9420 ;
  assign n9423 = n4826 ^ n4825 ;
  assign n9426 = ~n4817 & n9423 ;
  assign n9427 = n9426 ^ n4825 ;
  assign n9428 = n9422 & n9427 ;
  assign n9429 = n9428 ^ n4817 ;
  assign n9430 = ~n9419 & ~n9429 ;
  assign n9412 = n4860 ^ n4847 ;
  assign n9413 = n4850 & ~n4859 ;
  assign n9414 = n9413 ^ n4860 ;
  assign n9415 = ~n9412 & ~n9414 ;
  assign n9416 = n9415 ^ n4860 ;
  assign n9417 = n4892 & ~n9416 ;
  assign n9418 = n9417 ^ n4892 ;
  assign n9431 = n9430 ^ n9418 ;
  assign n9435 = n9434 ^ n9431 ;
  assign n9398 = x25 & n4772 ;
  assign n9400 = x26 & ~n4757 ;
  assign n9399 = n9398 ^ n4750 ;
  assign n9401 = n9400 ^ n9399 ;
  assign n9405 = ~n4750 & ~n4759 ;
  assign n9406 = n9405 ^ n4761 ;
  assign n9407 = n9401 & n9406 ;
  assign n9408 = n9407 ^ n4750 ;
  assign n9409 = ~n9398 & ~n9408 ;
  assign n9392 = n4791 ^ n4790 ;
  assign n9393 = x20 & n4788 ;
  assign n9394 = n9393 ^ n4790 ;
  assign n9395 = n9392 & ~n9394 ;
  assign n9396 = n9395 ^ n4790 ;
  assign n9397 = ~n4797 & n9396 ;
  assign n9410 = n9409 ^ n9397 ;
  assign n9389 = n4777 ^ n4734 ;
  assign n9390 = n4805 & n9389 ;
  assign n9391 = n9390 ^ n4777 ;
  assign n9411 = n9410 ^ n9391 ;
  assign n9436 = n9435 ^ n9411 ;
  assign n9387 = n4731 & n4806 ;
  assign n9384 = n9383 ^ n4806 ;
  assign n9385 = n9384 ^ n4731 ;
  assign n9386 = n4895 & n9385 ;
  assign n9388 = n9387 ^ n9386 ;
  assign n9437 = n9436 ^ n9388 ;
  assign n9374 = n4923 ^ n4917 ;
  assign n9375 = x992 & n4916 ;
  assign n9376 = n9375 ^ n4917 ;
  assign n9377 = n9374 & ~n9376 ;
  assign n9378 = n9377 ^ n4917 ;
  assign n9379 = ~n4934 & ~n9378 ;
  assign n9380 = n9379 ^ n4934 ;
  assign n9371 = n4945 ^ n4941 ;
  assign n9372 = n4950 & n9371 ;
  assign n9373 = n9372 ^ n4945 ;
  assign n9381 = n9380 ^ n9373 ;
  assign n9355 = n4953 ^ n4938 ;
  assign n9360 = n9355 ^ n4941 ;
  assign n9351 = n9265 ^ n4950 ;
  assign n9352 = n9351 ^ n9264 ;
  assign n9349 = n9265 ^ n4939 ;
  assign n9350 = n9349 ^ n9264 ;
  assign n9353 = n9352 ^ n9350 ;
  assign n9317 = n9269 ^ n4939 ;
  assign n9318 = n9355 ^ n9317 ;
  assign n9300 = ~n9269 & n9355 ;
  assign n9301 = n9300 ^ n9262 ;
  assign n9302 = n9318 ^ n9301 ;
  assign n9303 = n9302 ^ n9264 ;
  assign n9305 = n9360 ^ n9264 ;
  assign n9306 = n9303 & ~n9305 ;
  assign n9329 = n9360 ^ n9269 ;
  assign n9319 = n9318 ^ n4938 ;
  assign n9307 = n9319 ^ n4941 ;
  assign n9308 = n9329 ^ n9307 ;
  assign n9311 = n9308 & ~n9353 ;
  assign n9312 = n9306 & n9311 ;
  assign n9313 = n9312 ^ n9300 ;
  assign n9346 = n9353 ^ n9313 ;
  assign n9347 = n9346 ^ n4938 ;
  assign n9348 = n9347 ^ n4941 ;
  assign n9354 = n9353 ^ n9348 ;
  assign n9365 = n9360 ^ n9354 ;
  assign n9366 = n9365 ^ n4937 ;
  assign n9367 = n9366 ^ n4936 ;
  assign n9368 = n9367 ^ n9365 ;
  assign n9369 = n4956 & n9368 ;
  assign n9370 = n9369 ^ n9366 ;
  assign n9382 = n9381 ^ n9370 ;
  assign n9438 = n9437 ^ n9382 ;
  assign n9259 = n4957 ^ n4732 ;
  assign n9260 = ~n4897 & n9259 ;
  assign n9261 = n9260 ^ n4957 ;
  assign n9439 = n9438 ^ n9261 ;
  assign n11533 = n9443 ^ n9439 ;
  assign n11534 = ~n9561 & n11533 ;
  assign n11526 = n9435 ^ n9388 ;
  assign n11527 = n9436 & n11526 ;
  assign n11528 = n11527 ^ n9435 ;
  assign n11523 = n9373 & n9380 ;
  assign n11520 = n9381 ^ n9365 ;
  assign n11521 = ~n9370 & n11520 ;
  assign n11522 = n11521 ^ n9381 ;
  assign n11524 = n11523 ^ n11522 ;
  assign n11516 = n9409 ^ n9391 ;
  assign n11517 = n9410 & ~n11516 ;
  assign n11518 = n11517 ^ n9409 ;
  assign n11513 = n9434 ^ n9418 ;
  assign n11514 = ~n9431 & ~n11513 ;
  assign n11515 = n11514 ^ n9434 ;
  assign n11519 = n11518 ^ n11515 ;
  assign n11525 = n11524 ^ n11519 ;
  assign n11529 = n11528 ^ n11525 ;
  assign n11510 = n9382 ^ n9261 ;
  assign n11511 = n9438 & n11510 ;
  assign n11512 = n11511 ^ n9382 ;
  assign n11530 = n11529 ^ n11512 ;
  assign n11531 = n11530 ^ n9443 ;
  assign n11535 = n11534 ^ n11531 ;
  assign n12361 = ~n11522 & ~n11523 ;
  assign n12363 = n12361 ^ n11524 ;
  assign n12364 = ~n11512 & n12363 ;
  assign n12362 = n11518 & n12361 ;
  assign n12365 = n12364 ^ n12362 ;
  assign n12366 = ~n11515 & ~n11530 ;
  assign n12367 = n12366 ^ n12364 ;
  assign n12368 = n12365 & n12367 ;
  assign n12369 = n12368 ^ n12364 ;
  assign n12370 = ~n11528 & n12369 ;
  assign n12386 = ~n11512 & ~n11515 ;
  assign n12387 = n12362 & n12386 ;
  assign n12388 = n12387 ^ n12362 ;
  assign n12371 = n12364 ^ n11518 ;
  assign n12372 = n12371 ^ n11528 ;
  assign n12373 = n12371 ^ n11515 ;
  assign n12374 = ~n12372 & ~n12373 ;
  assign n12375 = n12374 ^ n12371 ;
  assign n12376 = ~n12361 & ~n12375 ;
  assign n12377 = n12364 & n12376 ;
  assign n12378 = ~n12374 & n12377 ;
  assign n12379 = n12378 ^ n12376 ;
  assign n12380 = n12379 ^ n12362 ;
  assign n12389 = n12388 ^ n12380 ;
  assign n12390 = ~n12370 & ~n12389 ;
  assign n12391 = n12390 ^ n11530 ;
  assign n11546 = n11545 ^ n11542 ;
  assign n11550 = n11549 ^ n11546 ;
  assign n11583 = n11582 ^ n11550 ;
  assign n12392 = n12391 ^ n11583 ;
  assign n12393 = n12392 ^ n12390 ;
  assign n12394 = ~n11535 & ~n12393 ;
  assign n12395 = n12394 ^ n12391 ;
  assign n12429 = n12428 ^ n12395 ;
  assign n13038 = n13037 ^ n12429 ;
  assign n12457 = n12456 ^ n12453 ;
  assign n11584 = n11583 ^ n11535 ;
  assign n9717 = n9716 ^ n9679 ;
  assign n4441 = n4440 ^ n4280 ;
  assign n9563 = n9440 ^ n4441 ;
  assign n9564 = n9563 ^ n4959 ;
  assign n1518 = n1517 ^ n1494 ;
  assign n4132 = n1518 ^ n1423 ;
  assign n4442 = n4441 ^ n1470 ;
  assign n4443 = n4442 ^ n1518 ;
  assign n4444 = n4443 ^ n4441 ;
  assign n4445 = ~n4132 & n4444 ;
  assign n4446 = n4445 ^ n4442 ;
  assign n9565 = n9564 ^ n4446 ;
  assign n9566 = n9564 ^ n9440 ;
  assign n9567 = n9565 & n9566 ;
  assign n9568 = n9567 ^ n9563 ;
  assign n9569 = n4441 & ~n9568 ;
  assign n9570 = ~n9567 & n9569 ;
  assign n9571 = n9570 ^ n9568 ;
  assign n9718 = n9717 ^ n9571 ;
  assign n9562 = n9561 ^ n9439 ;
  assign n11507 = n9571 ^ n9562 ;
  assign n11508 = ~n9718 & n11507 ;
  assign n11509 = n11508 ^ n9562 ;
  assign n11585 = n11584 ^ n11509 ;
  assign n11506 = n11505 ^ n11489 ;
  assign n12430 = n11509 ^ n11506 ;
  assign n12431 = n11585 & ~n12430 ;
  assign n12432 = n12431 ^ n11509 ;
  assign n12458 = n12457 ^ n12432 ;
  assign n13033 = n12432 ^ n12429 ;
  assign n13034 = n12458 & ~n13033 ;
  assign n13039 = n13038 ^ n13034 ;
  assign n13030 = n12428 ^ n12390 ;
  assign n13031 = n12395 & ~n13030 ;
  assign n13028 = n12428 ^ n12379 ;
  assign n13019 = ~n12397 & ~n12410 ;
  assign n13013 = n12403 ^ n11582 ;
  assign n13014 = n13013 ^ n12416 ;
  assign n13020 = n13019 ^ n13014 ;
  assign n13021 = n11582 & ~n13020 ;
  assign n13022 = n13021 ^ n13014 ;
  assign n13023 = n13022 ^ n12403 ;
  assign n13024 = n12416 ^ n12403 ;
  assign n13025 = ~n13021 & n13024 ;
  assign n13026 = ~n13023 & n13025 ;
  assign n13027 = n13026 ^ n13022 ;
  assign n13029 = n13028 ^ n13027 ;
  assign n13032 = n13031 ^ n13029 ;
  assign n13201 = n13037 ^ n13032 ;
  assign n13202 = ~n13039 & ~n13201 ;
  assign n13203 = n13202 ^ n13037 ;
  assign n13204 = n13203 ^ n13032 ;
  assign n13205 = n13204 ^ n13203 ;
  assign n13206 = ~n12379 & n13027 ;
  assign n13207 = ~n13205 & n13206 ;
  assign n13208 = n13207 ^ n13204 ;
  assign n13249 = ~n13203 & ~n13208 ;
  assign n1602 = x920 ^ x919 ;
  assign n5092 = ~x923 & ~x924 ;
  assign n5093 = ~x921 & ~x922 ;
  assign n1601 = x922 ^ x921 ;
  assign n5094 = n5093 ^ n1601 ;
  assign n5096 = ~n5092 & ~n5094 ;
  assign n1604 = x924 ^ x923 ;
  assign n5098 = n5092 ^ n1604 ;
  assign n5109 = ~n5093 & ~n5098 ;
  assign n5110 = ~n5096 & ~n5109 ;
  assign n5111 = n1602 & ~n5110 ;
  assign n5095 = n5094 ^ n5092 ;
  assign n5097 = n5096 ^ n5095 ;
  assign n5102 = n5097 ^ x920 ;
  assign n5099 = n5098 ^ x922 ;
  assign n5100 = ~n1601 & n5099 ;
  assign n5103 = n5102 ^ n5100 ;
  assign n5104 = n1602 & n5103 ;
  assign n5105 = n5104 ^ x919 ;
  assign n5101 = n5097 & ~n5100 ;
  assign n5107 = n5105 ^ n5101 ;
  assign n5106 = ~n5101 & ~n5105 ;
  assign n5108 = n5107 ^ n5106 ;
  assign n5112 = n5111 ^ n5108 ;
  assign n9245 = n5109 ^ n5096 ;
  assign n9246 = n9245 ^ n5110 ;
  assign n9247 = n5112 & n9246 ;
  assign n5126 = x925 & x926 ;
  assign n5122 = ~x927 & ~x928 ;
  assign n1607 = x928 ^ x927 ;
  assign n5127 = n5122 ^ n1607 ;
  assign n5128 = x930 & ~n5127 ;
  assign n5129 = n5126 & n5128 ;
  assign n5130 = n5129 ^ n5126 ;
  assign n5123 = ~x929 & ~x930 ;
  assign n5124 = ~n5122 & ~n5123 ;
  assign n5131 = n5130 ^ n5124 ;
  assign n1609 = x930 ^ x929 ;
  assign n5132 = n5123 ^ n1609 ;
  assign n5137 = n5127 & n5132 ;
  assign n5138 = n5137 ^ n5124 ;
  assign n5139 = n5131 & n5138 ;
  assign n5141 = n5139 ^ n5130 ;
  assign n1606 = x926 ^ x925 ;
  assign n5125 = ~n1606 & n5124 ;
  assign n5140 = n5125 & n5139 ;
  assign n5142 = n5141 ^ n5140 ;
  assign n9238 = n5132 ^ n5127 ;
  assign n9239 = x926 & n5124 ;
  assign n9240 = n9239 ^ n5127 ;
  assign n9241 = n9238 & ~n9240 ;
  assign n9242 = n9241 ^ n5127 ;
  assign n9243 = ~n5142 & ~n9242 ;
  assign n9244 = n9243 ^ n5142 ;
  assign n9248 = n9247 ^ n9244 ;
  assign n5197 = x939 & x940 ;
  assign n5196 = x941 & x942 ;
  assign n5198 = n5197 ^ n5196 ;
  assign n1598 = x942 ^ x941 ;
  assign n5199 = n5196 ^ n1598 ;
  assign n1595 = x940 ^ x939 ;
  assign n5200 = n5197 ^ n1595 ;
  assign n5201 = n5199 & n5200 ;
  assign n5202 = n5201 ^ n5197 ;
  assign n5203 = ~n5198 & ~n5202 ;
  assign n1596 = x938 ^ x937 ;
  assign n5192 = n1595 ^ x937 ;
  assign n5193 = n5192 ^ n1598 ;
  assign n5194 = n1596 & n5193 ;
  assign n5195 = n5194 ^ x937 ;
  assign n5204 = n5203 ^ n5195 ;
  assign n5156 = ~x933 & ~x934 ;
  assign n5155 = ~x935 & ~x936 ;
  assign n1593 = x936 ^ x935 ;
  assign n5159 = n5155 ^ n1593 ;
  assign n5160 = ~n5156 & ~n5159 ;
  assign n1591 = x934 ^ x933 ;
  assign n5157 = n5156 ^ n1591 ;
  assign n5158 = ~n5155 & ~n5157 ;
  assign n5162 = n5160 ^ n5158 ;
  assign n5161 = ~n5158 & ~n5160 ;
  assign n5163 = n5162 ^ n5161 ;
  assign n5164 = ~x931 & n5163 ;
  assign n5165 = n5159 ^ n5156 ;
  assign n5166 = n5165 ^ n5160 ;
  assign n5167 = n5166 ^ x932 ;
  assign n5168 = n5157 ^ n5155 ;
  assign n5169 = n5168 ^ n5158 ;
  assign n5170 = n5169 ^ x932 ;
  assign n5171 = n5167 & n5170 ;
  assign n5172 = n5171 ^ x932 ;
  assign n5173 = n5164 & n5172 ;
  assign n5174 = n5173 ^ x931 ;
  assign n5187 = ~x932 & n5156 ;
  assign n5188 = ~n5169 & n5187 ;
  assign n5189 = n5188 ^ n5169 ;
  assign n1590 = x932 ^ x931 ;
  assign n5175 = n5169 ^ n5163 ;
  assign n5176 = x932 & n5166 ;
  assign n5177 = ~n5175 & n5176 ;
  assign n5178 = n5177 ^ n5161 ;
  assign n5179 = ~n1590 & ~n5178 ;
  assign n5180 = n5179 ^ n5161 ;
  assign n5181 = n5180 ^ n5169 ;
  assign n5190 = n5189 ^ n5181 ;
  assign n5191 = n5174 & n5190 ;
  assign n5205 = n5204 ^ n5191 ;
  assign n1592 = n1591 ^ n1590 ;
  assign n1594 = n1593 ^ n1592 ;
  assign n1597 = n1596 ^ n1595 ;
  assign n1599 = n1598 ^ n1597 ;
  assign n5088 = n1594 & n1599 ;
  assign n9234 = n5204 ^ n5088 ;
  assign n9235 = n5205 & ~n9234 ;
  assign n9236 = n9235 ^ n5088 ;
  assign n9221 = n5198 ^ x937 ;
  assign n9222 = n9221 ^ n5201 ;
  assign n9223 = n5201 ^ x938 ;
  assign n9224 = ~n9222 & n9223 ;
  assign n9225 = n9224 ^ n5202 ;
  assign n9226 = ~n5198 & n9225 ;
  assign n9227 = ~n5197 & n9226 ;
  assign n9228 = n9224 ^ n5201 ;
  assign n9229 = n9228 ^ n9226 ;
  assign n9230 = n9229 ^ x937 ;
  assign n9231 = n9227 & n9230 ;
  assign n9232 = n9231 ^ n9229 ;
  assign n9220 = n5163 & n5180 ;
  assign n9233 = n9232 ^ n9220 ;
  assign n9237 = n9236 ^ n9233 ;
  assign n9249 = n9248 ^ n9237 ;
  assign n5115 = x929 ^ x928 ;
  assign n5119 = ~n1609 & ~n5115 ;
  assign n5114 = x927 ^ x926 ;
  assign n5116 = n5115 ^ x927 ;
  assign n5117 = n5116 ^ x930 ;
  assign n5118 = ~n5114 & n5117 ;
  assign n5120 = n5119 ^ n5118 ;
  assign n5121 = ~x925 & n5120 ;
  assign n5143 = ~n1607 & ~n5114 ;
  assign n5144 = x930 ^ x925 ;
  assign n5147 = ~x928 & ~n5144 ;
  assign n5148 = n5147 ^ x925 ;
  assign n5149 = n5143 & n5148 ;
  assign n5150 = ~x929 & n5149 ;
  assign n5151 = ~n5142 & ~n5150 ;
  assign n5152 = ~n5121 & n5151 ;
  assign n5113 = n5112 ^ n5106 ;
  assign n5153 = n5152 ^ n5113 ;
  assign n1603 = n1602 ^ n1601 ;
  assign n1605 = n1604 ^ n1603 ;
  assign n1608 = n1607 ^ n1606 ;
  assign n1610 = n1609 ^ n1608 ;
  assign n5090 = n1605 & n1610 ;
  assign n9217 = n5152 ^ n5090 ;
  assign n9218 = n5153 & n9217 ;
  assign n9219 = n9218 ^ n5152 ;
  assign n9250 = n9249 ^ n9219 ;
  assign n9210 = n5205 ^ n5088 ;
  assign n1600 = n1599 ^ n1594 ;
  assign n1611 = n1610 ^ n1605 ;
  assign n5087 = n1600 & n1611 ;
  assign n9212 = n5090 ^ n5087 ;
  assign n9215 = ~n9210 & n9212 ;
  assign n9211 = n9210 ^ n5090 ;
  assign n9213 = n9212 ^ n9211 ;
  assign n9214 = n5153 & ~n9213 ;
  assign n9216 = n9215 ^ n9214 ;
  assign n11623 = n9216 & n9250 ;
  assign n11624 = n9236 ^ n9232 ;
  assign n11625 = n9233 & n11624 ;
  assign n11630 = n11625 ^ n9233 ;
  assign n11628 = ~n9220 & n9232 ;
  assign n11629 = n9236 & n11628 ;
  assign n11631 = n11630 ^ n11629 ;
  assign n11632 = n9244 & ~n11631 ;
  assign n11626 = n11625 ^ n9236 ;
  assign n11633 = n11632 ^ n11626 ;
  assign n11634 = ~n9247 & n11633 ;
  assign n11627 = n9244 & n11626 ;
  assign n11635 = n11634 ^ n11627 ;
  assign n11636 = n11635 ^ n11629 ;
  assign n11637 = ~n11623 & n11636 ;
  assign n11642 = ~n9219 & n11637 ;
  assign n11643 = n11642 ^ n9216 ;
  assign n11644 = n9250 & n11643 ;
  assign n11645 = n11644 ^ n11637 ;
  assign n11646 = n11645 ^ n11623 ;
  assign n11647 = n9249 ^ n9247 ;
  assign n11648 = n11647 ^ n11632 ;
  assign n11653 = ~n11632 & ~n11648 ;
  assign n11649 = n11648 ^ n11626 ;
  assign n11654 = n11653 ^ n11649 ;
  assign n11655 = ~n9219 & n11654 ;
  assign n11656 = n11655 ^ n11649 ;
  assign n11657 = n9249 & n11656 ;
  assign n11658 = n11657 ^ n11649 ;
  assign n11659 = ~n11646 & ~n11658 ;
  assign n11660 = n11659 ^ n11623 ;
  assign n12514 = n9236 & n9244 ;
  assign n12508 = n11660 ^ n11628 ;
  assign n12509 = n12508 ^ n11645 ;
  assign n12515 = n12514 ^ n12509 ;
  assign n12516 = n11660 & n12515 ;
  assign n12517 = n12516 ^ n12509 ;
  assign n12518 = n12517 ^ n11628 ;
  assign n12519 = n12517 ^ n11660 ;
  assign n12520 = ~n12516 & ~n12519 ;
  assign n12521 = n12518 & n12520 ;
  assign n12522 = n12521 ^ n12517 ;
  assign n5000 = x899 & x900 ;
  assign n4999 = x897 & x898 ;
  assign n5001 = n5000 ^ n4999 ;
  assign n1570 = x900 ^ x899 ;
  assign n5002 = n5000 ^ n1570 ;
  assign n1568 = x898 ^ x897 ;
  assign n5003 = n4999 ^ n1568 ;
  assign n5004 = n5002 & n5003 ;
  assign n5005 = n5004 ^ n5000 ;
  assign n5006 = ~n5001 & ~n5005 ;
  assign n4969 = n1568 ^ x896 ;
  assign n4970 = n4969 ^ n1570 ;
  assign n1573 = x902 ^ x901 ;
  assign n4971 = ~x903 & ~x904 ;
  assign n1572 = x904 ^ x903 ;
  assign n4972 = n4971 ^ n1572 ;
  assign n4973 = x905 & x906 ;
  assign n1575 = x906 ^ x905 ;
  assign n4974 = n4973 ^ n1575 ;
  assign n4976 = ~n4972 & n4974 ;
  assign n4988 = ~n4971 & n4973 ;
  assign n4989 = ~n4976 & ~n4988 ;
  assign n4990 = n1573 & ~n4989 ;
  assign n4975 = n4974 ^ n4972 ;
  assign n4977 = n4976 ^ n4975 ;
  assign n4981 = n4977 ^ x902 ;
  assign n4978 = n4973 ^ x904 ;
  assign n4979 = ~n1572 & ~n4978 ;
  assign n4982 = n4981 ^ n4979 ;
  assign n4983 = n1573 & ~n4982 ;
  assign n4984 = n4983 ^ x901 ;
  assign n4980 = ~n4977 & ~n4979 ;
  assign n4986 = n4984 ^ n4980 ;
  assign n4985 = ~n4980 & ~n4984 ;
  assign n4987 = n4986 ^ n4985 ;
  assign n4991 = n4990 ^ n4987 ;
  assign n4992 = n4991 ^ n4985 ;
  assign n4993 = n4992 ^ x895 ;
  assign n4994 = n4993 ^ n1568 ;
  assign n4995 = n4994 ^ n1570 ;
  assign n4996 = n4995 ^ n4992 ;
  assign n4997 = ~n4970 & n4996 ;
  assign n4998 = n4997 ^ n4993 ;
  assign n5007 = n5006 ^ n4998 ;
  assign n1567 = x896 ^ x895 ;
  assign n1569 = n1568 ^ n1567 ;
  assign n1571 = n1570 ^ n1569 ;
  assign n1574 = n1573 ^ n1572 ;
  assign n1576 = n1575 ^ n1574 ;
  assign n4967 = n1571 & n1576 ;
  assign n9167 = n4992 ^ n4967 ;
  assign n9168 = ~n5007 & n9167 ;
  assign n9169 = n9168 ^ n4992 ;
  assign n5022 = ~x915 & ~x916 ;
  assign n1586 = x916 ^ x915 ;
  assign n5031 = n5022 ^ n1586 ;
  assign n5029 = ~x917 & ~x918 ;
  assign n1584 = x918 ^ x917 ;
  assign n5030 = n5029 ^ n1584 ;
  assign n5032 = n5031 ^ n5030 ;
  assign n5033 = ~n5022 & ~n5029 ;
  assign n5038 = x914 & n5033 ;
  assign n5039 = n5038 ^ n5030 ;
  assign n5040 = n5032 & n5039 ;
  assign n5041 = n5040 ^ n5031 ;
  assign n5067 = x913 & x914 ;
  assign n5068 = x918 & ~n5031 ;
  assign n5069 = n5067 & n5068 ;
  assign n5070 = n5069 ^ n5067 ;
  assign n5071 = n5070 ^ n5033 ;
  assign n5076 = n5030 & n5031 ;
  assign n5077 = n5076 ^ n5070 ;
  assign n5078 = n5071 & ~n5077 ;
  assign n1583 = x914 ^ x913 ;
  assign n5079 = n5078 ^ n5070 ;
  assign n5080 = ~n1583 & n5079 ;
  assign n5081 = n5078 & n5080 ;
  assign n5082 = n5081 ^ n5079 ;
  assign n9170 = n5041 & ~n5082 ;
  assign n5023 = x917 ^ x914 ;
  assign n5026 = n1584 & n5023 ;
  assign n5027 = n5026 ^ x917 ;
  assign n5028 = n5022 & ~n5027 ;
  assign n5042 = n5041 ^ n5028 ;
  assign n5043 = ~x913 & ~n5042 ;
  assign n5045 = x918 ^ x914 ;
  assign n5044 = x918 ^ x916 ;
  assign n5046 = n5045 ^ n5044 ;
  assign n5047 = n5046 ^ x918 ;
  assign n5049 = x914 & n5047 ;
  assign n5050 = n5049 ^ x918 ;
  assign n5053 = x918 ^ x915 ;
  assign n5054 = n5053 ^ n5045 ;
  assign n5055 = n5054 ^ n1583 ;
  assign n5056 = n5046 ^ n1583 ;
  assign n5057 = n5056 ^ n5045 ;
  assign n5058 = n5057 ^ x918 ;
  assign n5059 = ~n5055 & n5058 ;
  assign n5062 = n5059 ^ x916 ;
  assign n5063 = ~n5050 & ~n5062 ;
  assign n5066 = ~x917 & n5063 ;
  assign n5083 = ~n5066 & ~n5082 ;
  assign n5084 = ~n5043 & n5083 ;
  assign n1579 = x908 ^ x907 ;
  assign n1578 = x912 ^ x911 ;
  assign n5017 = n1578 ^ x908 ;
  assign n1581 = x910 ^ x909 ;
  assign n5018 = n5017 ^ n1581 ;
  assign n5019 = n1579 & ~n5018 ;
  assign n5020 = n5019 ^ x907 ;
  assign n5010 = x911 & x912 ;
  assign n5009 = x909 & x910 ;
  assign n5011 = n5010 ^ n5009 ;
  assign n5012 = n5009 ^ n1581 ;
  assign n5013 = n5010 ^ n1578 ;
  assign n5014 = n5012 & n5013 ;
  assign n5015 = n5014 ^ n5009 ;
  assign n5016 = ~n5011 & ~n5015 ;
  assign n5021 = n5020 ^ n5016 ;
  assign n5085 = n5084 ^ n5021 ;
  assign n1580 = n1579 ^ n1578 ;
  assign n1582 = n1581 ^ n1580 ;
  assign n1585 = n1584 ^ n1583 ;
  assign n1587 = n1586 ^ n1585 ;
  assign n4965 = n1582 & n1587 ;
  assign n9188 = n5021 ^ n4965 ;
  assign n9189 = ~n5085 & ~n9188 ;
  assign n9190 = n9189 ^ n5021 ;
  assign n9191 = n5014 ^ x908 ;
  assign n9192 = n5011 ^ x907 ;
  assign n9193 = n9192 ^ n5014 ;
  assign n9194 = n9191 & ~n9193 ;
  assign n9197 = n9194 ^ n5014 ;
  assign n9195 = n9194 ^ n5015 ;
  assign n9196 = ~n5011 & n9195 ;
  assign n9198 = n9197 ^ n9196 ;
  assign n9199 = x907 & n9196 ;
  assign n9200 = ~n9198 & n9199 ;
  assign n9201 = n9200 ^ n9198 ;
  assign n11602 = n9190 & ~n9201 ;
  assign n11603 = n9170 & n11602 ;
  assign n9171 = n5004 ^ x896 ;
  assign n9172 = n5001 ^ x895 ;
  assign n9173 = n9172 ^ n5004 ;
  assign n9174 = n9171 & ~n9173 ;
  assign n9177 = n9174 ^ n5004 ;
  assign n9175 = n9174 ^ n5005 ;
  assign n9176 = ~n5001 & n9175 ;
  assign n9178 = n9177 ^ n9176 ;
  assign n9179 = x895 & n9176 ;
  assign n9180 = ~n9178 & n9179 ;
  assign n9181 = n9180 ^ n9178 ;
  assign n9182 = n4988 ^ n4976 ;
  assign n9183 = n9182 ^ n4989 ;
  assign n9184 = n4991 & n9183 ;
  assign n11605 = ~n9181 & n9184 ;
  assign n12499 = ~n11603 & n11605 ;
  assign n12500 = ~n9169 & n12499 ;
  assign n12501 = n12500 ^ n11603 ;
  assign n9202 = n9201 ^ n9190 ;
  assign n11612 = n11602 ^ n9202 ;
  assign n11613 = ~n9170 & n11612 ;
  assign n9185 = n9184 ^ n9181 ;
  assign n9186 = n9185 ^ n9170 ;
  assign n9187 = n9186 ^ n9169 ;
  assign n9203 = n9202 ^ n9187 ;
  assign n11614 = n11603 ^ n9203 ;
  assign n11615 = n11614 ^ n11605 ;
  assign n11616 = n11615 ^ n9169 ;
  assign n11617 = n11616 ^ n11613 ;
  assign n11596 = n9202 ^ n9170 ;
  assign n11597 = n9185 & ~n11596 ;
  assign n11618 = n11617 ^ n11597 ;
  assign n9143 = n5085 ^ n4965 ;
  assign n1577 = n1576 ^ n1571 ;
  assign n1588 = n1587 ^ n1582 ;
  assign n4964 = n1577 & n1588 ;
  assign n9146 = n9143 ^ n4964 ;
  assign n9147 = n9146 ^ n4967 ;
  assign n9148 = n9147 ^ n5007 ;
  assign n9149 = n9148 ^ n4967 ;
  assign n9150 = n9149 ^ n9143 ;
  assign n9157 = ~n5007 & ~n9150 ;
  assign n9144 = n9143 ^ n5007 ;
  assign n9152 = n9148 ^ n9144 ;
  assign n9158 = n9157 ^ n9152 ;
  assign n9160 = n9157 ^ n5007 ;
  assign n9161 = n5085 & ~n9160 ;
  assign n9162 = n9161 ^ n4965 ;
  assign n9163 = n9162 ^ n5085 ;
  assign n9164 = ~n9158 & ~n9163 ;
  assign n9165 = n9164 ^ n9161 ;
  assign n9166 = n9165 ^ n9143 ;
  assign n11604 = n11603 ^ n9169 ;
  assign n11606 = n11605 ^ n9169 ;
  assign n11607 = n11604 & n11606 ;
  assign n11608 = n11607 ^ n9169 ;
  assign n11609 = ~n9166 & ~n11608 ;
  assign n11610 = n11609 ^ n9169 ;
  assign n11611 = ~n9203 & ~n11610 ;
  assign n11619 = n11618 ^ n11611 ;
  assign n11598 = n9169 & n11597 ;
  assign n11599 = ~n9166 & n11598 ;
  assign n11620 = n11619 ^ n11599 ;
  assign n12504 = n12500 ^ n11620 ;
  assign n12505 = ~n11613 & n12504 ;
  assign n12506 = ~n12501 & n12505 ;
  assign n9204 = n9203 ^ n9166 ;
  assign n11621 = n11620 ^ n9204 ;
  assign n1589 = n1588 ^ n1577 ;
  assign n1612 = n1611 ^ n1600 ;
  assign n5207 = n1589 & n1612 ;
  assign n5089 = n5088 ^ n5087 ;
  assign n5091 = n5090 ^ n5089 ;
  assign n5154 = n5153 ^ n5091 ;
  assign n5206 = n5205 ^ n5154 ;
  assign n5208 = n5207 ^ n5206 ;
  assign n9207 = n9148 ^ n5206 ;
  assign n9208 = ~n5208 & ~n9207 ;
  assign n9205 = n9204 ^ n5206 ;
  assign n9209 = n9208 ^ n9205 ;
  assign n9251 = n9250 ^ n9216 ;
  assign n11594 = n9251 ^ n9204 ;
  assign n11595 = ~n9209 & n11594 ;
  assign n11622 = n11621 ^ n11595 ;
  assign n12496 = n11660 ^ n11620 ;
  assign n12497 = ~n11622 & n12496 ;
  assign n12498 = n12497 ^ n11660 ;
  assign n12502 = n12501 ^ n12498 ;
  assign n12507 = n12506 ^ n12502 ;
  assign n12523 = n12522 ^ n12507 ;
  assign n1549 = x856 ^ x855 ;
  assign n5228 = ~x857 & ~x858 ;
  assign n1551 = x858 ^ x857 ;
  assign n5232 = n5228 ^ n1551 ;
  assign n5233 = n5232 ^ x856 ;
  assign n5234 = n1549 & n5233 ;
  assign n5235 = n5234 ^ x855 ;
  assign n5237 = ~x855 & ~x856 ;
  assign n5238 = n5232 & n5237 ;
  assign n5236 = n5234 ^ n5233 ;
  assign n5239 = n5238 ^ n5236 ;
  assign n5240 = n5235 & ~n5239 ;
  assign n5242 = x854 & ~n5228 ;
  assign n5243 = n5240 & n5242 ;
  assign n5244 = n5243 ^ n5239 ;
  assign n5246 = n5237 ^ n1549 ;
  assign n5249 = ~n5244 & n5246 ;
  assign n5245 = n5244 ^ n5238 ;
  assign n5247 = n5246 ^ n5245 ;
  assign n5248 = ~x854 & ~n5247 ;
  assign n5250 = n5249 ^ n5248 ;
  assign n1548 = x854 ^ x853 ;
  assign n1550 = n1549 ^ n1548 ;
  assign n1552 = n1551 ^ n1550 ;
  assign n5229 = n5228 ^ n1552 ;
  assign n5230 = n5228 ^ x853 ;
  assign n5231 = ~n5229 & n5230 ;
  assign n5251 = n5250 ^ n5231 ;
  assign n5213 = x849 & x850 ;
  assign n5211 = x851 & x852 ;
  assign n5216 = n5213 ^ n5211 ;
  assign n1546 = x852 ^ x851 ;
  assign n5212 = n5211 ^ n1546 ;
  assign n1544 = x850 ^ x849 ;
  assign n5214 = n5213 ^ n1544 ;
  assign n5218 = n5212 & n5214 ;
  assign n5219 = n5218 ^ n5211 ;
  assign n5220 = ~n5216 & n5219 ;
  assign n5215 = n5214 ^ n5212 ;
  assign n5227 = n5220 ^ n5215 ;
  assign n5252 = n5251 ^ n5227 ;
  assign n1543 = x848 ^ x847 ;
  assign n5217 = n5216 ^ x848 ;
  assign n5221 = ~n5217 & n5220 ;
  assign n5222 = n5221 ^ n5217 ;
  assign n5223 = n5222 ^ n5215 ;
  assign n5224 = ~n1543 & n5223 ;
  assign n5253 = n5252 ^ n5224 ;
  assign n5226 = n5221 & n5224 ;
  assign n5254 = n5253 ^ n5226 ;
  assign n1562 = x864 ^ x863 ;
  assign n5299 = x863 ^ x862 ;
  assign n5303 = ~n1562 & ~n5299 ;
  assign n5298 = x861 ^ x860 ;
  assign n5300 = n5299 ^ x861 ;
  assign n5301 = n5300 ^ x864 ;
  assign n5302 = ~n5298 & n5301 ;
  assign n5304 = n5303 ^ n5302 ;
  assign n5305 = ~x859 & n5304 ;
  assign n1560 = x862 ^ x861 ;
  assign n5306 = ~n1560 & ~n5298 ;
  assign n5307 = x864 ^ x859 ;
  assign n5310 = ~x862 & ~n5307 ;
  assign n5311 = n5310 ^ x859 ;
  assign n5312 = n5306 & n5311 ;
  assign n5313 = ~x863 & n5312 ;
  assign n5314 = ~x861 & ~x862 ;
  assign n5317 = n5314 ^ n1560 ;
  assign n5318 = x859 & x860 ;
  assign n5319 = x864 & n5318 ;
  assign n5320 = ~n5317 & n5319 ;
  assign n5321 = n5320 ^ n5318 ;
  assign n5315 = ~x863 & ~x864 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5322 = n5321 ^ n5316 ;
  assign n5323 = n5315 ^ n1562 ;
  assign n5328 = n5317 & n5323 ;
  assign n5329 = n5328 ^ n5316 ;
  assign n5330 = n5322 & n5329 ;
  assign n1559 = x860 ^ x859 ;
  assign n5331 = n5330 ^ n5321 ;
  assign n5332 = ~n1559 & n5331 ;
  assign n5333 = n5330 & n5332 ;
  assign n5334 = n5333 ^ n5331 ;
  assign n5335 = ~n5313 & ~n5334 ;
  assign n5336 = ~n5305 & n5335 ;
  assign n1557 = x870 ^ x869 ;
  assign n5260 = x869 ^ x868 ;
  assign n5264 = ~n1557 & ~n5260 ;
  assign n5259 = x867 ^ x866 ;
  assign n5261 = n5260 ^ x867 ;
  assign n5262 = n5261 ^ x870 ;
  assign n5263 = ~n5259 & n5262 ;
  assign n5265 = n5264 ^ n5263 ;
  assign n5266 = ~x865 & n5265 ;
  assign n1555 = x868 ^ x867 ;
  assign n5267 = ~n1555 & ~n5259 ;
  assign n5268 = x870 ^ x865 ;
  assign n5271 = ~x868 & ~n5268 ;
  assign n5272 = n5271 ^ x865 ;
  assign n5273 = n5267 & n5272 ;
  assign n5274 = ~x869 & n5273 ;
  assign n5275 = ~x867 & ~x868 ;
  assign n5278 = n5275 ^ n1555 ;
  assign n5279 = x865 & x866 ;
  assign n5280 = x870 & n5279 ;
  assign n5281 = ~n5278 & n5280 ;
  assign n5282 = n5281 ^ n5279 ;
  assign n5276 = ~x869 & ~x870 ;
  assign n5277 = ~n5275 & ~n5276 ;
  assign n5283 = n5282 ^ n5277 ;
  assign n5284 = n5276 ^ n1557 ;
  assign n5289 = n5278 & n5284 ;
  assign n5290 = n5289 ^ n5277 ;
  assign n5291 = n5283 & n5290 ;
  assign n1554 = x866 ^ x865 ;
  assign n5292 = n5291 ^ n5282 ;
  assign n5293 = ~n1554 & n5292 ;
  assign n5294 = n5291 & n5293 ;
  assign n5295 = n5294 ^ n5292 ;
  assign n5296 = ~n5274 & ~n5295 ;
  assign n5297 = ~n5266 & n5296 ;
  assign n5337 = n5336 ^ n5297 ;
  assign n1556 = n1555 ^ n1554 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1561 = n1560 ^ n1559 ;
  assign n1563 = n1562 ^ n1561 ;
  assign n5257 = n1558 & n1563 ;
  assign n1545 = n1544 ^ n1543 ;
  assign n1547 = n1546 ^ n1545 ;
  assign n1553 = n1552 ^ n1547 ;
  assign n1564 = n1563 ^ n1558 ;
  assign n5256 = n1553 & n1564 ;
  assign n5258 = n5257 ^ n5256 ;
  assign n5338 = n5337 ^ n5258 ;
  assign n5210 = n1547 & n1552 ;
  assign n5255 = n5254 ^ n5210 ;
  assign n8977 = n5256 ^ n5255 ;
  assign n8978 = n5338 & n8977 ;
  assign n8979 = n8978 ^ n5256 ;
  assign n8980 = n8979 ^ n5251 ;
  assign n8981 = n8980 ^ n5210 ;
  assign n8982 = n8981 ^ n8979 ;
  assign n8983 = n5254 & n8982 ;
  assign n8984 = n8983 ^ n8980 ;
  assign n8999 = n5297 ^ n5257 ;
  assign n9000 = n5337 & n8999 ;
  assign n9001 = n9000 ^ n5297 ;
  assign n8991 = n5323 ^ n5317 ;
  assign n8992 = x860 & n5316 ;
  assign n8993 = n8992 ^ n5317 ;
  assign n8994 = n8991 & ~n8993 ;
  assign n8995 = n8994 ^ n5317 ;
  assign n8996 = ~n5334 & ~n8995 ;
  assign n8997 = n8996 ^ n5334 ;
  assign n8985 = n5284 ^ n5278 ;
  assign n8986 = x866 & n5277 ;
  assign n8987 = n8986 ^ n5278 ;
  assign n8988 = n8985 & ~n8987 ;
  assign n8989 = n8988 ^ n5278 ;
  assign n8990 = ~n5295 & n8989 ;
  assign n8998 = n8997 ^ n8990 ;
  assign n9002 = n9001 ^ n8998 ;
  assign n11671 = n9002 ^ n8979 ;
  assign n11672 = ~n8984 & ~n11671 ;
  assign n11673 = n11672 ^ n9002 ;
  assign n9019 = x853 & x854 ;
  assign n9020 = ~x858 & ~n5246 ;
  assign n9021 = n9019 & n9020 ;
  assign n9024 = n5238 ^ n5235 ;
  assign n9025 = n9024 ^ n5246 ;
  assign n9026 = n9025 ^ n5235 ;
  assign n9027 = x854 & n9026 ;
  assign n9028 = n9027 ^ n5235 ;
  assign n9029 = ~n1548 & n9028 ;
  assign n9030 = n9029 ^ n5235 ;
  assign n9031 = ~n5228 & n9030 ;
  assign n9032 = ~n9021 & ~n9031 ;
  assign n9033 = ~n5244 & n9032 ;
  assign n9009 = n5218 ^ n5213 ;
  assign n9004 = n5218 ^ x848 ;
  assign n9005 = n5218 ^ n5216 ;
  assign n9006 = n9005 ^ x847 ;
  assign n9007 = n9004 & ~n9006 ;
  assign n9010 = n9009 ^ n9007 ;
  assign n9011 = ~n5216 & n9010 ;
  assign n9014 = x847 & n9011 ;
  assign n9015 = n9007 ^ n5218 ;
  assign n9016 = n9014 & n9015 ;
  assign n9008 = n9007 ^ n9004 ;
  assign n9012 = n9011 ^ n9008 ;
  assign n9013 = n9012 ^ n5213 ;
  assign n9017 = n9016 ^ n9013 ;
  assign n9003 = n5217 ^ n5211 ;
  assign n9018 = n9017 ^ n9003 ;
  assign n9034 = n9033 ^ n9018 ;
  assign n9035 = n9034 ^ n9002 ;
  assign n11684 = n11673 ^ n9035 ;
  assign n11685 = n11684 ^ n8984 ;
  assign n11681 = n9001 ^ n8997 ;
  assign n11682 = ~n8998 & n11681 ;
  assign n11683 = n11682 ^ n8997 ;
  assign n11686 = n11685 ^ n11683 ;
  assign n11666 = n9018 ^ n9002 ;
  assign n11676 = n9002 & ~n11673 ;
  assign n11677 = ~n11666 & n11676 ;
  assign n11678 = n11677 ^ n11666 ;
  assign n11679 = n11678 ^ n8984 ;
  assign n11680 = n9034 & n11679 ;
  assign n11687 = n11686 ^ n11680 ;
  assign n12471 = n9018 & ~n9033 ;
  assign n12465 = n11687 ^ n11673 ;
  assign n12466 = n12465 ^ n11683 ;
  assign n12472 = n12471 ^ n12466 ;
  assign n12473 = n11687 & ~n12472 ;
  assign n12474 = n12473 ^ n12466 ;
  assign n12475 = n12474 ^ n11673 ;
  assign n12476 = n12474 ^ n11687 ;
  assign n12478 = n12475 & n12476 ;
  assign n12479 = n12478 ^ n12474 ;
  assign n9113 = ~x871 & ~x872 ;
  assign n5349 = ~x873 & ~x874 ;
  assign n1532 = x874 ^ x873 ;
  assign n5378 = n5349 ^ n1532 ;
  assign n9114 = x876 & ~n5378 ;
  assign n9115 = ~x875 & ~x876 ;
  assign n9116 = ~n5349 & ~n9115 ;
  assign n1534 = x876 ^ x875 ;
  assign n9117 = n9115 ^ n1534 ;
  assign n9118 = n5378 & n9117 ;
  assign n9119 = ~n9116 & n9118 ;
  assign n9120 = x871 & x872 ;
  assign n9121 = ~n9119 & n9120 ;
  assign n9122 = n9121 ^ x875 ;
  assign n9123 = n9114 & n9122 ;
  assign n9124 = n9123 ^ n9121 ;
  assign n9125 = n9118 ^ n9116 ;
  assign n9126 = n9125 ^ n9119 ;
  assign n9127 = ~n9124 & n9126 ;
  assign n9130 = n9113 & n9127 ;
  assign n9128 = n9127 ^ n9124 ;
  assign n9131 = n9130 ^ n9128 ;
  assign n5357 = x879 & x880 ;
  assign n5355 = x881 & x882 ;
  assign n5360 = n5357 ^ n5355 ;
  assign n1539 = x882 ^ x881 ;
  assign n5356 = n5355 ^ n1539 ;
  assign n1537 = x880 ^ x879 ;
  assign n5358 = n5357 ^ n1537 ;
  assign n5361 = n5356 & n5358 ;
  assign n9093 = n5361 ^ x878 ;
  assign n9096 = n5355 ^ x877 ;
  assign n9097 = n9096 ^ n5360 ;
  assign n9095 = n5355 ^ x878 ;
  assign n9098 = n9097 ^ n9095 ;
  assign n9099 = n9093 & n9098 ;
  assign n5362 = n5361 ^ n5355 ;
  assign n9100 = n9099 ^ n5362 ;
  assign n9101 = ~n5360 & n9100 ;
  assign n9104 = x877 & n9101 ;
  assign n9105 = n9099 ^ n5361 ;
  assign n9106 = n9104 & n9105 ;
  assign n9102 = n9101 ^ n9093 ;
  assign n9103 = n9102 ^ n9099 ;
  assign n9107 = n9106 ^ n9103 ;
  assign n9110 = n9107 ^ n5355 ;
  assign n9112 = n9110 ^ n9095 ;
  assign n9132 = n9131 ^ n9112 ;
  assign n5396 = x893 & x894 ;
  assign n1528 = x894 ^ x893 ;
  assign n5398 = n5396 ^ n1528 ;
  assign n5395 = x891 & x892 ;
  assign n1526 = x892 ^ x891 ;
  assign n5399 = n5395 ^ n1526 ;
  assign n5400 = n5398 & n5399 ;
  assign n9081 = n5400 ^ x890 ;
  assign n5397 = n5396 ^ n5395 ;
  assign n9082 = n5397 ^ x889 ;
  assign n9083 = n9082 ^ n5400 ;
  assign n9084 = n9081 & ~n9083 ;
  assign n9087 = n9084 ^ n5400 ;
  assign n5401 = n5400 ^ n5396 ;
  assign n9085 = n9084 ^ n5401 ;
  assign n9086 = ~n5397 & n9085 ;
  assign n9088 = n9087 ^ n9086 ;
  assign n9089 = x889 & n9086 ;
  assign n9090 = ~n9088 & n9089 ;
  assign n9091 = n9090 ^ n9088 ;
  assign n5385 = ~x885 & ~x886 ;
  assign n9056 = ~x887 & ~x888 ;
  assign n9059 = ~n5385 & ~n9056 ;
  assign n1522 = x886 ^ x885 ;
  assign n5406 = n5385 ^ n1522 ;
  assign n9064 = n9059 ^ n5406 ;
  assign n1520 = x888 ^ x887 ;
  assign n9057 = n9056 ^ n1520 ;
  assign n9058 = n9057 ^ n5406 ;
  assign n9062 = n9058 ^ x883 ;
  assign n9065 = n9064 ^ n9062 ;
  assign n9066 = n9065 ^ x884 ;
  assign n9067 = n9066 ^ n9064 ;
  assign n9070 = n5406 ^ x884 ;
  assign n9071 = n9070 ^ n9064 ;
  assign n9072 = ~n9067 & n9071 ;
  assign n9073 = n9072 ^ n9057 ;
  assign n9074 = n9072 ^ x884 ;
  assign n9075 = n9074 ^ n5406 ;
  assign n9076 = ~n9058 & ~n9075 ;
  assign n9077 = ~n9067 & n9076 ;
  assign n9078 = n9073 & n9077 ;
  assign n9079 = n9078 ^ n9076 ;
  assign n9080 = n9079 ^ n9074 ;
  assign n9092 = n9091 ^ n9080 ;
  assign n9133 = n9132 ^ n9092 ;
  assign n1521 = x884 ^ x883 ;
  assign n1523 = n1522 ^ n1521 ;
  assign n5405 = n1523 ^ x887 ;
  assign n5407 = n5406 ^ x888 ;
  assign n5408 = n5405 & n5407 ;
  assign n5402 = ~n5397 & ~n5401 ;
  assign n1525 = x890 ^ x889 ;
  assign n5391 = n1528 ^ x890 ;
  assign n5392 = n5391 ^ n1526 ;
  assign n5393 = n1525 & ~n5392 ;
  assign n5394 = n5393 ^ x889 ;
  assign n5403 = n5402 ^ n5394 ;
  assign n5383 = x887 ^ x884 ;
  assign n5386 = n5385 ^ x887 ;
  assign n5389 = ~n5383 & n5386 ;
  assign n5387 = n5386 ^ x884 ;
  assign n5388 = x883 & n5387 ;
  assign n5390 = n5389 ^ n5388 ;
  assign n5404 = n5403 ^ n5390 ;
  assign n5409 = n5408 ^ n5404 ;
  assign n1524 = n1523 ^ n1520 ;
  assign n1527 = n1526 ^ n1525 ;
  assign n1529 = n1528 ^ n1527 ;
  assign n5344 = n1524 & n1529 ;
  assign n9053 = n5403 ^ n5344 ;
  assign n9054 = n5409 & ~n9053 ;
  assign n9055 = n9054 ^ n5403 ;
  assign n9134 = n9133 ^ n9055 ;
  assign n5379 = n5378 ^ x876 ;
  assign n1531 = x872 ^ x871 ;
  assign n1533 = n1532 ^ n1531 ;
  assign n5380 = n1533 ^ x875 ;
  assign n5381 = n5379 & n5380 ;
  assign n5363 = ~n5360 & n5362 ;
  assign n5365 = n5360 ^ x878 ;
  assign n5359 = n5358 ^ n5356 ;
  assign n5364 = n5363 ^ n5359 ;
  assign n5366 = n5365 ^ n5364 ;
  assign n5367 = n5366 ^ n5363 ;
  assign n5368 = n5367 ^ n5364 ;
  assign n5370 = n5363 & n5368 ;
  assign n1536 = x878 ^ x877 ;
  assign n5371 = n5370 ^ n5367 ;
  assign n5372 = ~n1536 & n5371 ;
  assign n5375 = n5370 & n5372 ;
  assign n5373 = n5372 ^ n5364 ;
  assign n5376 = n5375 ^ n5373 ;
  assign n5347 = x875 ^ x872 ;
  assign n5350 = n5349 ^ x875 ;
  assign n5353 = ~n5347 & n5350 ;
  assign n5351 = n5350 ^ x872 ;
  assign n5352 = x871 & n5351 ;
  assign n5354 = n5353 ^ n5352 ;
  assign n5377 = n5376 ^ n5354 ;
  assign n5382 = n5381 ^ n5377 ;
  assign n9045 = n5382 ^ n5344 ;
  assign n1535 = n1534 ^ n1533 ;
  assign n1538 = n1537 ^ n1536 ;
  assign n1540 = n1539 ^ n1538 ;
  assign n9046 = n1535 & n1540 ;
  assign n1541 = n1540 ^ n1535 ;
  assign n1530 = n1529 ^ n1524 ;
  assign n5340 = n1535 ^ n1530 ;
  assign n5341 = n1541 & ~n5340 ;
  assign n5342 = n5341 ^ n1540 ;
  assign n9047 = n9046 ^ n5342 ;
  assign n9048 = ~n9045 & n9047 ;
  assign n9042 = n5409 ^ n5344 ;
  assign n9043 = n5382 ^ n5342 ;
  assign n9044 = n9042 & ~n9043 ;
  assign n9049 = n9048 ^ n9044 ;
  assign n9050 = n9046 ^ n5376 ;
  assign n9051 = ~n5382 & n9050 ;
  assign n9052 = n9051 ^ n5376 ;
  assign n11713 = n9112 ^ n9052 ;
  assign n11692 = ~n9055 & n9091 ;
  assign n11693 = n9080 & n11692 ;
  assign n11690 = n9055 & ~n9091 ;
  assign n11691 = ~n9080 & n11690 ;
  assign n11694 = n11693 ^ n11691 ;
  assign n11722 = ~n9131 & n11694 ;
  assign n11717 = n11693 ^ n9052 ;
  assign n11723 = n11722 ^ n11717 ;
  assign n11724 = ~n11713 & ~n11723 ;
  assign n11710 = n9112 & n11693 ;
  assign n11695 = n11694 ^ n9092 ;
  assign n11696 = n11695 ^ n9055 ;
  assign n11708 = ~n9112 & ~n11696 ;
  assign n11709 = ~n9052 & n11708 ;
  assign n11711 = n11710 ^ n11709 ;
  assign n11714 = n11711 ^ n11693 ;
  assign n11725 = n11724 ^ n11714 ;
  assign n11726 = n11725 ^ n11693 ;
  assign n11712 = n11711 ^ n9131 ;
  assign n11727 = n11726 ^ n11712 ;
  assign n11728 = n9131 & n11725 ;
  assign n11729 = n11728 ^ n11712 ;
  assign n11730 = n11691 ^ n9131 ;
  assign n11733 = ~n11729 & n11730 ;
  assign n11734 = ~n11727 & n11733 ;
  assign n11735 = n11734 ^ n11728 ;
  assign n11736 = n11735 ^ n11711 ;
  assign n11737 = ~n9052 & ~n11736 ;
  assign n11702 = n9112 & ~n11691 ;
  assign n11703 = n11702 ^ n11696 ;
  assign n11704 = ~n9132 & n11703 ;
  assign n11699 = n11696 ^ n11693 ;
  assign n11705 = n11704 ^ n11699 ;
  assign n11738 = n11737 ^ n11705 ;
  assign n11739 = ~n9049 & ~n11738 ;
  assign n11740 = n11739 ^ n11705 ;
  assign n11741 = ~n9134 & ~n11740 ;
  assign n12480 = n11709 ^ n9112 ;
  assign n12481 = n12480 ^ n11691 ;
  assign n11746 = n9049 & n9052 ;
  assign n11747 = n11746 ^ n11736 ;
  assign n11748 = ~n11705 & ~n11747 ;
  assign n12482 = n11748 ^ n9112 ;
  assign n12483 = n12482 ^ n11691 ;
  assign n12488 = n9131 & ~n12483 ;
  assign n12489 = n12481 & n12488 ;
  assign n12490 = n12489 ^ n11748 ;
  assign n12491 = n12490 ^ n11709 ;
  assign n12492 = ~n11691 & ~n12491 ;
  assign n12493 = ~n11709 & n12492 ;
  assign n12494 = ~n11741 & n12493 ;
  assign n12991 = n12479 & ~n12494 ;
  assign n12495 = n12494 ^ n12479 ;
  assign n12994 = n12991 ^ n12495 ;
  assign n12995 = n12523 & ~n12994 ;
  assign n11661 = n11660 ^ n11622 ;
  assign n9135 = n9134 ^ n9052 ;
  assign n9136 = n9135 ^ n9049 ;
  assign n5410 = n5409 ^ n5382 ;
  assign n1542 = n1541 ^ n1530 ;
  assign n1565 = n1564 ^ n1553 ;
  assign n5343 = n1542 & n1565 ;
  assign n5345 = n5344 ^ n5343 ;
  assign n5346 = n5345 ^ n5342 ;
  assign n5411 = n5410 ^ n5346 ;
  assign n5339 = n5338 ^ n5255 ;
  assign n9039 = n5343 ^ n5339 ;
  assign n9040 = ~n5411 & n9039 ;
  assign n9036 = n9035 ^ n8984 ;
  assign n9037 = n9036 ^ n5343 ;
  assign n9041 = n9040 ^ n9037 ;
  assign n9137 = n9136 ^ n9041 ;
  assign n11662 = n11661 ^ n9137 ;
  assign n5412 = n5411 ^ n5339 ;
  assign n5209 = n9148 ^ n5208 ;
  assign n5413 = n5412 ^ n5209 ;
  assign n1566 = n1565 ^ n1542 ;
  assign n1613 = n1612 ^ n1589 ;
  assign n4962 = n1566 & n1613 ;
  assign n9140 = n5209 ^ n4962 ;
  assign n9141 = n5413 & ~n9140 ;
  assign n9138 = n9137 ^ n5209 ;
  assign n9142 = n9141 ^ n9138 ;
  assign n9252 = n9251 ^ n9209 ;
  assign n11592 = n9252 ^ n9137 ;
  assign n11593 = n9142 & n11592 ;
  assign n11663 = n11662 ^ n11593 ;
  assign n11749 = ~n11741 & ~n11748 ;
  assign n11688 = n11687 ^ n9036 ;
  assign n11664 = n9136 ^ n9036 ;
  assign n11665 = n9041 & ~n11664 ;
  assign n11689 = n11688 ^ n11665 ;
  assign n11750 = n11749 ^ n11689 ;
  assign n12525 = n11750 ^ n11661 ;
  assign n12526 = n11663 & ~n12525 ;
  assign n12527 = n12526 ^ n11750 ;
  assign n12528 = n11749 ^ n11687 ;
  assign n12529 = n11689 & ~n12528 ;
  assign n12530 = n12529 ^ n11687 ;
  assign n12990 = ~n12527 & n12530 ;
  assign n12531 = n12530 ^ n12527 ;
  assign n12996 = n12990 ^ n12531 ;
  assign n12997 = n12995 & n12996 ;
  assign n12999 = ~n12523 & ~n12996 ;
  assign n13188 = n12994 & n12999 ;
  assign n13003 = ~n12990 & n12991 ;
  assign n13004 = n13003 ^ n12994 ;
  assign n13005 = ~n12999 & n13004 ;
  assign n13006 = n13005 ^ n12994 ;
  assign n13189 = n13188 ^ n13006 ;
  assign n12987 = n12522 ^ n12498 ;
  assign n12988 = n12507 & n12987 ;
  assign n12989 = n12988 ^ n12522 ;
  assign n13190 = n13189 ^ n12989 ;
  assign n13191 = n13190 ^ n13189 ;
  assign n12992 = ~n12523 & ~n12991 ;
  assign n12993 = n12990 & n12992 ;
  assign n13192 = n13189 ^ n12993 ;
  assign n13193 = n13192 ^ n13189 ;
  assign n13195 = n13189 ^ n13188 ;
  assign n13196 = ~n13193 & ~n13195 ;
  assign n13197 = ~n13191 & n13196 ;
  assign n13198 = n13197 ^ n13191 ;
  assign n13199 = n13198 ^ n13190 ;
  assign n13200 = ~n12997 & ~n13199 ;
  assign n13209 = n13208 ^ n13200 ;
  assign n13040 = n13039 ^ n13032 ;
  assign n12459 = n12458 ^ n12429 ;
  assign n13041 = n13040 ^ n12459 ;
  assign n1471 = n1470 ^ n1423 ;
  assign n1519 = n1518 ^ n1471 ;
  assign n1614 = n1613 ^ n1566 ;
  assign n4961 = n1519 & n1614 ;
  assign n4963 = n4962 ^ n4961 ;
  assign n5414 = n5413 ^ n4963 ;
  assign n4960 = n4959 ^ n4446 ;
  assign n9256 = n4961 ^ n4960 ;
  assign n9257 = n5414 & n9256 ;
  assign n9253 = n9252 ^ n9142 ;
  assign n9254 = n9253 ^ n4961 ;
  assign n9258 = n9257 ^ n9254 ;
  assign n11586 = n11585 ^ n11506 ;
  assign n11588 = n11586 ^ n9253 ;
  assign n9719 = n9718 ^ n9562 ;
  assign n11587 = n11586 ^ n9719 ;
  assign n11589 = n11588 ^ n11587 ;
  assign n11590 = ~n9258 & n11589 ;
  assign n11591 = n11590 ^ n11588 ;
  assign n12461 = n12459 ^ n11586 ;
  assign n11751 = n11750 ^ n11663 ;
  assign n12460 = n12459 ^ n11751 ;
  assign n12462 = n12461 ^ n12460 ;
  assign n12463 = ~n11591 & n12462 ;
  assign n12464 = n12463 ^ n12461 ;
  assign n12524 = n12523 ^ n12495 ;
  assign n12532 = n12531 ^ n12524 ;
  assign n13009 = n12532 ^ n12459 ;
  assign n13010 = ~n12464 & n13009 ;
  assign n13042 = n13041 ^ n13010 ;
  assign n12998 = n12997 ^ n12993 ;
  assign n13007 = ~n12998 & ~n13006 ;
  assign n13008 = n13007 ^ n12989 ;
  assign n13185 = n13040 ^ n13008 ;
  assign n13186 = n13042 & ~n13185 ;
  assign n13187 = n13186 ^ n13040 ;
  assign n13210 = n13209 ^ n13187 ;
  assign n13043 = n13042 ^ n13008 ;
  assign n12533 = n12532 ^ n12464 ;
  assign n11752 = n11751 ^ n11591 ;
  assign n12534 = n12533 ^ n11752 ;
  assign n5415 = n5414 ^ n4960 ;
  assign n1615 = n1614 ^ n1519 ;
  assign n4130 = ~n1383 & n1615 ;
  assign n9725 = n4130 ^ n4128 ;
  assign n4127 = ~n1192 & n1615 ;
  assign n9726 = n9725 ^ n4127 ;
  assign n9727 = n5415 & n9726 ;
  assign n9721 = n5415 ^ n4130 ;
  assign n9722 = n9721 ^ n4127 ;
  assign n9723 = n7941 & n9722 ;
  assign n9720 = n9719 ^ n9258 ;
  assign n9724 = n9723 ^ n9720 ;
  assign n9728 = n9727 ^ n9724 ;
  assign n11753 = n11752 ^ n9720 ;
  assign n11754 = n11753 ^ n11752 ;
  assign n8976 = n8975 ^ n8469 ;
  assign n11755 = n11754 ^ n8976 ;
  assign n11756 = n9728 & ~n11755 ;
  assign n11757 = n11756 ^ n11753 ;
  assign n12122 = n12121 ^ n11935 ;
  assign n12359 = n12122 ^ n11752 ;
  assign n12360 = ~n11757 & ~n12359 ;
  assign n12535 = n12534 ^ n12360 ;
  assign n12733 = n12732 ^ n12538 ;
  assign n12984 = n12733 ^ n12533 ;
  assign n12985 = n12535 & ~n12984 ;
  assign n12986 = n12985 ^ n12733 ;
  assign n13044 = n13043 ^ n12986 ;
  assign n12983 = n12982 ^ n12901 ;
  assign n13182 = n12986 ^ n12983 ;
  assign n13183 = n13044 & ~n13182 ;
  assign n13184 = n13183 ^ n12983 ;
  assign n13211 = n13210 ^ n13184 ;
  assign n13180 = n13179 ^ n13148 ;
  assign n13145 = n13144 ^ n13141 ;
  assign n13181 = n13180 ^ n13145 ;
  assign n13250 = n13184 ^ n13181 ;
  assign n13251 = ~n13211 & ~n13250 ;
  assign n13252 = n13251 ^ n13184 ;
  assign n13253 = n13252 ^ n13208 ;
  assign n13254 = n13253 ^ n13187 ;
  assign n13255 = n13254 ^ n13252 ;
  assign n13256 = n13209 & ~n13255 ;
  assign n13257 = n13256 ^ n13253 ;
  assign n13258 = n13257 ^ n13252 ;
  assign n13259 = n13249 & ~n13258 ;
  assign n13260 = n13259 ^ n13257 ;
  assign n13342 = n13341 ^ n13260 ;
  assign n1921 = x690 ^ x689 ;
  assign n1920 = x688 ^ x687 ;
  assign n1922 = n1921 ^ n1920 ;
  assign n1919 = x686 ^ x685 ;
  assign n1923 = n1922 ^ n1919 ;
  assign n1917 = x682 ^ x681 ;
  assign n1915 = x684 ^ x683 ;
  assign n1914 = x680 ^ x679 ;
  assign n1916 = n1915 ^ n1914 ;
  assign n1918 = n1917 ^ n1916 ;
  assign n1924 = n1923 ^ n1918 ;
  assign n1910 = x694 ^ x693 ;
  assign n1909 = x696 ^ x695 ;
  assign n1911 = n1910 ^ n1909 ;
  assign n1908 = x692 ^ x691 ;
  assign n1912 = n1911 ^ n1908 ;
  assign n1905 = x702 ^ x701 ;
  assign n1904 = x700 ^ x699 ;
  assign n1906 = n1905 ^ n1904 ;
  assign n1903 = x698 ^ x697 ;
  assign n1907 = n1906 ^ n1903 ;
  assign n1913 = n1912 ^ n1907 ;
  assign n2054 = n1923 ^ n1913 ;
  assign n2055 = n1924 & n2054 ;
  assign n2043 = x681 & x682 ;
  assign n2042 = x683 & x684 ;
  assign n2044 = n2043 ^ n2042 ;
  assign n2045 = n2043 ^ n1917 ;
  assign n2046 = n2042 ^ n1915 ;
  assign n2047 = n2045 & n2046 ;
  assign n2048 = n2047 ^ n2043 ;
  assign n2049 = ~n2044 & ~n2048 ;
  assign n2038 = n1917 ^ x680 ;
  assign n2039 = n2038 ^ n1915 ;
  assign n2040 = n1914 & ~n2039 ;
  assign n2041 = n2040 ^ x679 ;
  assign n2050 = n2049 ^ n2041 ;
  assign n2014 = x689 & x690 ;
  assign n2015 = n2014 ^ n1921 ;
  assign n2016 = ~x687 & ~x688 ;
  assign n2020 = ~n2014 & n2016 ;
  assign n2017 = n2016 ^ n1920 ;
  assign n2018 = n2014 & ~n2017 ;
  assign n2021 = n2020 ^ n2018 ;
  assign n2019 = n2014 ^ x688 ;
  assign n2022 = n2021 ^ n2019 ;
  assign n2023 = n2022 ^ x687 ;
  assign n2034 = n2015 & ~n2023 ;
  assign n2033 = n2023 ^ n2015 ;
  assign n2035 = n2034 ^ n2033 ;
  assign n2036 = ~x686 & n2035 ;
  assign n2029 = n2020 ^ n1923 ;
  assign n2030 = n1923 ^ x685 ;
  assign n2031 = ~n2029 & n2030 ;
  assign n2024 = ~n2018 & ~n2023 ;
  assign n2025 = x686 & n2024 ;
  assign n2026 = n2015 & n2025 ;
  assign n2027 = n2026 ^ n2024 ;
  assign n2028 = n2027 ^ n2023 ;
  assign n2032 = n2031 ^ n2028 ;
  assign n2037 = n2036 ^ n2032 ;
  assign n2051 = n2050 ^ n2037 ;
  assign n2052 = n2051 ^ n1923 ;
  assign n2056 = n2055 ^ n2052 ;
  assign n2106 = x691 & ~x692 ;
  assign n2107 = x696 ^ x693 ;
  assign n2108 = x695 ^ x694 ;
  assign n2109 = n2108 ^ x696 ;
  assign n2110 = n2107 & ~n2109 ;
  assign n2111 = n2110 ^ x696 ;
  assign n2112 = n2106 & ~n2111 ;
  assign n2114 = n2112 ^ n2106 ;
  assign n2115 = ~x694 & ~x695 ;
  assign n2116 = n2114 & n2115 ;
  assign n2113 = n2112 ^ x691 ;
  assign n2117 = n2116 ^ n2113 ;
  assign n2118 = x695 ^ x693 ;
  assign n2119 = ~n1910 & n2118 ;
  assign n2120 = n2119 ^ n1909 ;
  assign n2121 = n2120 ^ n1910 ;
  assign n2126 = x696 & ~n2119 ;
  assign n2127 = n2121 & n2126 ;
  assign n2128 = n2127 ^ n2121 ;
  assign n2129 = n2128 ^ n1910 ;
  assign n2130 = x692 & ~n2129 ;
  assign n2131 = n2117 & ~n2130 ;
  assign n2133 = x693 ^ x692 ;
  assign n2136 = n1911 & ~n2133 ;
  assign n2132 = ~n1909 & ~n2108 ;
  assign n2137 = n2136 ^ n2132 ;
  assign n2138 = ~x691 & n2137 ;
  assign n2139 = ~n2131 & ~n2138 ;
  assign n2140 = ~n1910 & ~n2133 ;
  assign n2141 = x696 ^ x691 ;
  assign n2144 = ~x694 & ~n2141 ;
  assign n2145 = n2144 ^ x691 ;
  assign n2146 = n2140 & n2145 ;
  assign n2147 = ~x695 & n2146 ;
  assign n2148 = n2139 & ~n2147 ;
  assign n2070 = x701 ^ x698 ;
  assign n2071 = n2070 ^ x700 ;
  assign n2072 = n2071 ^ x702 ;
  assign n2068 = x701 ^ x699 ;
  assign n2073 = n2072 ^ n2068 ;
  assign n2074 = n2073 ^ x702 ;
  assign n2075 = n2074 ^ x701 ;
  assign n2076 = n2075 ^ n2068 ;
  assign n2082 = n2068 ^ n1906 ;
  assign n2083 = ~n2076 & ~n2082 ;
  assign n2084 = ~x701 & n2083 ;
  assign n2087 = n2084 ^ n2083 ;
  assign n2085 = n2084 ^ n2068 ;
  assign n2086 = n2073 & n2085 ;
  assign n2088 = n2087 ^ n2086 ;
  assign n2089 = n2088 ^ x701 ;
  assign n2149 = n2148 ^ n2089 ;
  assign n2058 = ~x699 & ~x700 ;
  assign n2092 = n2058 ^ n1904 ;
  assign n2060 = ~x701 & ~x702 ;
  assign n2091 = n2060 ^ n1905 ;
  assign n2095 = n2092 ^ n2091 ;
  assign n2059 = n2058 ^ x698 ;
  assign n2061 = n2060 ^ n2059 ;
  assign n2096 = n2092 ^ n2061 ;
  assign n2063 = n2060 ^ n2058 ;
  assign n2062 = n2058 & n2060 ;
  assign n2064 = n2063 ^ n2062 ;
  assign n2065 = n2061 & n2064 ;
  assign n2097 = n2096 ^ n2065 ;
  assign n2098 = n2095 & n2097 ;
  assign n2099 = n2098 ^ n2091 ;
  assign n2103 = ~x697 & ~n2088 ;
  assign n2104 = n2103 ^ x701 ;
  assign n2105 = ~n2099 & ~n2104 ;
  assign n2150 = n2149 ^ n2105 ;
  assign n2090 = ~x697 & ~n2089 ;
  assign n2093 = n2091 & n2092 ;
  assign n2094 = n2090 & n2093 ;
  assign n2151 = n2150 ^ n2094 ;
  assign n2066 = n2062 ^ x697 ;
  assign n2067 = ~n2065 & ~n2066 ;
  assign n2152 = n2151 ^ n2067 ;
  assign n2057 = n1907 & n1912 ;
  assign n2153 = n2152 ^ n2057 ;
  assign n10984 = n2153 ^ n2051 ;
  assign n10985 = ~n2056 & n10984 ;
  assign n10986 = n10985 ^ n2051 ;
  assign n10959 = x694 ^ x692 ;
  assign n10964 = n2133 & n10959 ;
  assign n10965 = n10964 ^ x692 ;
  assign n10975 = n1910 ^ x692 ;
  assign n10971 = n2108 ^ x693 ;
  assign n10972 = n10971 ^ x692 ;
  assign n10973 = ~n1909 & n10972 ;
  assign n10976 = n10975 ^ n10973 ;
  assign n10977 = n10965 & n10976 ;
  assign n10980 = ~n2131 & ~n10977 ;
  assign n10956 = n2089 ^ x697 ;
  assign n10957 = n10956 ^ n2090 ;
  assign n10958 = n2099 & n10957 ;
  assign n10981 = n10980 ^ n10958 ;
  assign n10953 = n2148 ^ n2057 ;
  assign n10954 = ~n2152 & n10953 ;
  assign n10955 = n10954 ^ n2148 ;
  assign n10982 = n10981 ^ n10955 ;
  assign n10940 = n2047 ^ x680 ;
  assign n10941 = n2044 ^ x679 ;
  assign n10942 = n10941 ^ n2047 ;
  assign n10943 = n10940 & ~n10942 ;
  assign n10946 = n10943 ^ n2047 ;
  assign n10944 = n10943 ^ n2048 ;
  assign n10945 = ~n2044 & n10944 ;
  assign n10947 = n10946 ^ n10945 ;
  assign n10948 = x679 & n10945 ;
  assign n10949 = ~n10947 & n10948 ;
  assign n10950 = n10949 ^ n10947 ;
  assign n10934 = ~n2021 & ~n2035 ;
  assign n10935 = n10934 ^ n2034 ;
  assign n10936 = x686 & n10935 ;
  assign n10937 = n10936 ^ n2034 ;
  assign n10938 = x685 & n10937 ;
  assign n10939 = n2028 & ~n10938 ;
  assign n10951 = n10950 ^ n10939 ;
  assign n10931 = n2037 & ~n2050 ;
  assign n10952 = n10951 ^ n10931 ;
  assign n10983 = n10982 ^ n10952 ;
  assign n10987 = n10986 ^ n10983 ;
  assign n2284 = x677 ^ x673 ;
  assign n2285 = n2284 ^ x678 ;
  assign n1944 = x674 ^ x673 ;
  assign n1943 = x676 ^ x675 ;
  assign n1945 = n1944 ^ n1943 ;
  assign n2286 = n2285 ^ n1945 ;
  assign n1942 = x678 ^ x677 ;
  assign n2272 = x675 & x676 ;
  assign n2292 = ~x678 & ~n2272 ;
  assign n2293 = ~n1942 & n2292 ;
  assign n2294 = n2293 ^ n1942 ;
  assign n2295 = n2294 ^ n1945 ;
  assign n2296 = n2286 & ~n2295 ;
  assign n2269 = ~x677 & ~x678 ;
  assign n2270 = n2269 ^ n1942 ;
  assign n2273 = ~n2270 & n2272 ;
  assign n2271 = n2270 ^ x676 ;
  assign n2275 = n1943 & n2271 ;
  assign n2278 = n2275 ^ x675 ;
  assign n2279 = ~n2273 & n2278 ;
  assign n2280 = x674 & n2279 ;
  assign n2281 = ~n2269 & n2280 ;
  assign n2282 = n2281 ^ n2279 ;
  assign n2283 = n2282 ^ n2278 ;
  assign n2297 = n2296 ^ n2283 ;
  assign n2274 = n2273 ^ n2271 ;
  assign n2276 = n2275 ^ n2274 ;
  assign n2277 = ~x674 & n2276 ;
  assign n2298 = n2297 ^ n2277 ;
  assign n2211 = x672 ^ x668 ;
  assign n2210 = x672 ^ x670 ;
  assign n2212 = n2211 ^ n2210 ;
  assign n2213 = n2212 ^ x672 ;
  assign n2215 = x668 & n2213 ;
  assign n2216 = n2215 ^ x672 ;
  assign n2219 = x672 ^ x669 ;
  assign n2220 = n2219 ^ n2211 ;
  assign n1937 = x668 ^ x667 ;
  assign n2221 = n2220 ^ n1937 ;
  assign n2222 = n2212 ^ n1937 ;
  assign n2223 = n2222 ^ n2211 ;
  assign n2224 = n2223 ^ x672 ;
  assign n2225 = ~n2221 & n2224 ;
  assign n2228 = n2225 ^ x670 ;
  assign n2229 = ~n2216 & ~n2228 ;
  assign n2232 = ~x671 & n2229 ;
  assign n2254 = x671 & x672 ;
  assign n2257 = n2254 ^ x670 ;
  assign n1939 = x672 ^ x671 ;
  assign n2255 = n2254 ^ n1939 ;
  assign n2256 = x668 & n2255 ;
  assign n2260 = n2256 ^ n2254 ;
  assign n2261 = ~n2257 & ~n2260 ;
  assign n2258 = n2257 ^ n2256 ;
  assign n2259 = x669 & ~n2258 ;
  assign n2262 = n2261 ^ n2259 ;
  assign n2235 = x671 ^ x668 ;
  assign n2236 = n2235 ^ x670 ;
  assign n2237 = n2236 ^ x672 ;
  assign n2233 = x671 ^ x669 ;
  assign n2238 = n2237 ^ n2233 ;
  assign n2244 = ~n2210 & ~n2212 ;
  assign n2248 = n2244 ^ x669 ;
  assign n2249 = n2248 ^ n2233 ;
  assign n2250 = n2244 & n2249 ;
  assign n2251 = n2250 ^ n2233 ;
  assign n2252 = ~n2238 & n2251 ;
  assign n2253 = n2252 ^ n2248 ;
  assign n2263 = n2262 ^ n2253 ;
  assign n2266 = x667 & n2263 ;
  assign n2267 = n2266 ^ n2262 ;
  assign n2268 = ~n2232 & ~n2267 ;
  assign n2299 = n2298 ^ n2268 ;
  assign n2200 = x659 & x660 ;
  assign n2199 = x657 & x658 ;
  assign n2201 = n2200 ^ n2199 ;
  assign n1934 = x660 ^ x659 ;
  assign n2202 = n2200 ^ n1934 ;
  assign n1932 = x658 ^ x657 ;
  assign n2203 = n2199 ^ n1932 ;
  assign n2204 = n2202 & n2203 ;
  assign n2205 = n2204 ^ n2200 ;
  assign n2206 = ~n2201 & ~n2205 ;
  assign n1931 = x656 ^ x655 ;
  assign n2195 = n1934 ^ x656 ;
  assign n2196 = n2195 ^ n1932 ;
  assign n2197 = n1931 & ~n2196 ;
  assign n2198 = n2197 ^ x655 ;
  assign n2207 = n2206 ^ n2198 ;
  assign n2164 = ~x663 & ~x664 ;
  assign n1927 = x664 ^ x663 ;
  assign n2171 = n2164 ^ n1927 ;
  assign n2163 = x665 & x666 ;
  assign n1929 = x666 ^ x665 ;
  assign n2168 = n2163 ^ n1929 ;
  assign n2176 = n2171 ^ n2168 ;
  assign n2172 = n2168 & ~n2171 ;
  assign n2177 = n2176 ^ n2172 ;
  assign n2178 = ~x662 & n2177 ;
  assign n2166 = n2163 & ~n2164 ;
  assign n2174 = n2172 ^ n2166 ;
  assign n2173 = ~n2166 & ~n2172 ;
  assign n2175 = n2174 ^ n2173 ;
  assign n2179 = n2178 ^ n2175 ;
  assign n2165 = n2164 ^ n2163 ;
  assign n2167 = n2166 ^ n2165 ;
  assign n2169 = n2168 ^ x662 ;
  assign n2170 = n2167 & n2169 ;
  assign n2180 = n2179 ^ n2170 ;
  assign n2181 = ~x661 & ~n2180 ;
  assign n2192 = n2164 & n2178 ;
  assign n1926 = x662 ^ x661 ;
  assign n2182 = n2175 ^ n2167 ;
  assign n2183 = x662 & ~n2177 ;
  assign n2184 = n2182 & n2183 ;
  assign n2185 = n2184 ^ n2173 ;
  assign n2186 = ~n1926 & ~n2185 ;
  assign n2187 = n2186 ^ n2173 ;
  assign n2193 = n2192 ^ n2187 ;
  assign n2194 = ~n2181 & n2193 ;
  assign n2208 = n2207 ^ n2194 ;
  assign n1928 = n1927 ^ n1926 ;
  assign n1930 = n1929 ^ n1928 ;
  assign n1933 = n1932 ^ n1931 ;
  assign n1935 = n1934 ^ n1933 ;
  assign n2159 = n1930 & n1935 ;
  assign n1946 = n1945 ^ n1942 ;
  assign n1938 = x670 ^ x669 ;
  assign n1940 = n1939 ^ n1938 ;
  assign n1941 = n1940 ^ n1937 ;
  assign n1947 = n1946 ^ n1941 ;
  assign n1936 = n1935 ^ n1930 ;
  assign n2156 = n1941 ^ n1936 ;
  assign n2157 = n1947 & ~n2156 ;
  assign n2158 = n2157 ^ n1946 ;
  assign n2160 = n2159 ^ n2158 ;
  assign n2209 = n2208 ^ n2160 ;
  assign n2300 = n2299 ^ n2209 ;
  assign n2154 = n2153 ^ n2056 ;
  assign n2301 = n2300 ^ n2154 ;
  assign n1925 = n1924 ^ n1913 ;
  assign n1948 = n1947 ^ n1936 ;
  assign n2012 = n1925 & n1948 ;
  assign n10928 = n2154 ^ n2012 ;
  assign n10929 = n2301 & n10928 ;
  assign n10930 = n10929 ^ n2154 ;
  assign n10988 = n10987 ^ n10930 ;
  assign n10921 = x667 & n2253 ;
  assign n10888 = n2257 ^ x669 ;
  assign n10889 = ~n2260 & ~n10888 ;
  assign n10890 = n10889 ^ n1938 ;
  assign n10918 = ~x670 & ~n10889 ;
  assign n10919 = ~n10890 & n10918 ;
  assign n10891 = x673 & ~n2283 ;
  assign n10894 = x677 ^ x674 ;
  assign n10895 = n10894 ^ x676 ;
  assign n10896 = n10895 ^ x678 ;
  assign n10892 = x677 ^ x675 ;
  assign n10897 = n10896 ^ n10892 ;
  assign n10898 = n10897 ^ x678 ;
  assign n10899 = n10898 ^ x677 ;
  assign n10900 = n10899 ^ n10892 ;
  assign n10903 = x678 ^ x676 ;
  assign n10904 = ~n10900 & ~n10903 ;
  assign n10908 = n10904 ^ x675 ;
  assign n10909 = n10908 ^ n10892 ;
  assign n10910 = n10904 & n10909 ;
  assign n10911 = n10910 ^ n10892 ;
  assign n10912 = ~n10897 & n10911 ;
  assign n10913 = n10912 ^ n10908 ;
  assign n10914 = n10891 & n10913 ;
  assign n10915 = n10914 ^ n2283 ;
  assign n10916 = n10915 ^ n10890 ;
  assign n10920 = n10919 ^ n10916 ;
  assign n10922 = n10920 ^ n10915 ;
  assign n10923 = n10921 & n10922 ;
  assign n10924 = n10923 ^ n10920 ;
  assign n2155 = n1941 & n1946 ;
  assign n10885 = n2298 ^ n2155 ;
  assign n10886 = ~n2299 & ~n10885 ;
  assign n10887 = n10886 ^ n2298 ;
  assign n10925 = n10924 ^ n10887 ;
  assign n10883 = n2158 & n2209 ;
  assign n10881 = n2209 ^ n2155 ;
  assign n10882 = ~n2299 & ~n10881 ;
  assign n10884 = n10883 ^ n10882 ;
  assign n10926 = n10925 ^ n10884 ;
  assign n10869 = n2204 ^ x656 ;
  assign n10870 = n2201 ^ x655 ;
  assign n10871 = n10870 ^ n2204 ;
  assign n10872 = n10869 & ~n10871 ;
  assign n10875 = n10872 ^ n2204 ;
  assign n10873 = n10872 ^ n2205 ;
  assign n10874 = ~n2201 & n10873 ;
  assign n10876 = n10875 ^ n10874 ;
  assign n10877 = x655 & n10874 ;
  assign n10878 = ~n10876 & n10877 ;
  assign n10879 = n10878 ^ n10876 ;
  assign n10867 = n2175 & n2187 ;
  assign n10864 = n2207 ^ n2159 ;
  assign n10865 = ~n2208 & ~n10864 ;
  assign n10866 = n10865 ^ n2207 ;
  assign n10868 = n10867 ^ n10866 ;
  assign n10880 = n10879 ^ n10868 ;
  assign n10927 = n10926 ^ n10880 ;
  assign n10989 = n10988 ^ n10927 ;
  assign n1952 = x736 ^ x735 ;
  assign n1951 = x734 ^ x733 ;
  assign n1953 = n1952 ^ n1951 ;
  assign n2329 = n1953 ^ x737 ;
  assign n2310 = ~x735 & ~x736 ;
  assign n2330 = n2310 ^ n1952 ;
  assign n2331 = n2330 ^ x738 ;
  assign n2332 = n2329 & n2331 ;
  assign n1956 = x730 ^ x729 ;
  assign n1957 = x732 ^ x731 ;
  assign n2318 = x731 ^ x728 ;
  assign n2319 = n2318 ^ n1956 ;
  assign n2320 = n1957 & n2319 ;
  assign n2321 = n2320 ^ x731 ;
  assign n10804 = n2321 ^ x730 ;
  assign n10803 = n2321 ^ x728 ;
  assign n10805 = n10804 ^ n10803 ;
  assign n2326 = ~n1956 & n10805 ;
  assign n1958 = n1957 ^ n1956 ;
  assign n1955 = x728 ^ x727 ;
  assign n1959 = n1958 ^ n1955 ;
  assign n2316 = x727 & ~n1959 ;
  assign n2317 = n2316 ^ x728 ;
  assign n2322 = n2321 ^ n2317 ;
  assign n2327 = n2326 ^ n2322 ;
  assign n2308 = x737 ^ x734 ;
  assign n2311 = n2310 ^ x737 ;
  assign n2314 = ~n2308 & n2311 ;
  assign n2312 = n2311 ^ x734 ;
  assign n2313 = x733 & n2312 ;
  assign n2315 = n2314 ^ n2313 ;
  assign n2328 = n2327 ^ n2315 ;
  assign n2333 = n2332 ^ n2328 ;
  assign n1950 = x738 ^ x737 ;
  assign n1954 = n1953 ^ n1950 ;
  assign n2306 = n1954 & n1959 ;
  assign n10857 = n2327 ^ n2306 ;
  assign n10858 = n2333 & n10857 ;
  assign n10859 = n10858 ^ n2306 ;
  assign n10828 = ~x737 & ~x738 ;
  assign n10835 = n10828 ^ n1950 ;
  assign n10836 = n10835 ^ n2330 ;
  assign n10829 = ~n2310 & ~n10828 ;
  assign n10843 = x734 & n10829 ;
  assign n10844 = n10843 ^ n10835 ;
  assign n10845 = n10836 & n10844 ;
  assign n10846 = n10845 ^ n2330 ;
  assign n10847 = n10846 ^ n10836 ;
  assign n10830 = x733 & x734 ;
  assign n10831 = x738 & ~n2330 ;
  assign n10832 = n10830 & n10831 ;
  assign n10833 = n10832 ^ n10830 ;
  assign n10834 = n10833 ^ n10829 ;
  assign n10837 = n10836 ^ n10829 ;
  assign n10838 = ~n10834 & n10837 ;
  assign n10848 = n10847 ^ n10838 ;
  assign n10849 = n10848 ^ n10846 ;
  assign n10850 = ~n10835 & ~n10838 ;
  assign n10851 = ~n10849 & n10850 ;
  assign n10852 = n10851 ^ n10848 ;
  assign n10854 = ~n1951 & ~n10833 ;
  assign n10855 = ~n10852 & n10854 ;
  assign n10853 = n10852 ^ n10846 ;
  assign n10856 = n10855 ^ n10853 ;
  assign n10860 = n10859 ^ n10856 ;
  assign n1964 = x750 ^ x749 ;
  assign n2358 = ~x747 & ~x748 ;
  assign n1962 = x748 ^ x747 ;
  assign n2359 = n2358 ^ n1962 ;
  assign n2360 = x745 & x746 ;
  assign n2361 = ~n2359 & n2360 ;
  assign n2435 = ~n1964 & n2361 ;
  assign n2335 = ~x749 & ~x750 ;
  assign n1961 = x746 ^ x745 ;
  assign n2365 = n2335 ^ n1961 ;
  assign n2339 = n2335 ^ n1964 ;
  assign n2372 = n2339 & n2358 ;
  assign n2366 = n2359 ^ x746 ;
  assign n2373 = n2372 ^ n2366 ;
  assign n2374 = ~n2365 & n2373 ;
  assign n2431 = n2374 ^ n2359 ;
  assign n2375 = n2374 ^ n2366 ;
  assign n2429 = ~n2335 & n2375 ;
  assign n2432 = ~x745 & n2429 ;
  assign n2433 = n2431 & n2432 ;
  assign n2377 = ~x741 & ~x742 ;
  assign n1967 = x742 ^ x741 ;
  assign n2411 = n2377 ^ n1967 ;
  assign n2379 = ~x743 & ~x744 ;
  assign n1968 = x744 ^ x743 ;
  assign n2387 = n2379 ^ n1968 ;
  assign n2414 = n2411 ^ n2387 ;
  assign n2378 = n2377 ^ x740 ;
  assign n2380 = n2379 ^ n2378 ;
  assign n2415 = n2387 ^ n2380 ;
  assign n2382 = n2379 ^ n2377 ;
  assign n2381 = n2377 & n2379 ;
  assign n2383 = n2382 ^ n2381 ;
  assign n2384 = n2380 & n2383 ;
  assign n2416 = n2415 ^ n2384 ;
  assign n2417 = n2414 & n2416 ;
  assign n2418 = n2417 ^ n2411 ;
  assign n2390 = x743 ^ x740 ;
  assign n2391 = n2390 ^ x742 ;
  assign n2392 = n2391 ^ x744 ;
  assign n2388 = x743 ^ x741 ;
  assign n2393 = n2392 ^ n2388 ;
  assign n2394 = n2393 ^ x744 ;
  assign n2395 = n2394 ^ x743 ;
  assign n2396 = n2395 ^ n2388 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n2402 = n2388 ^ n1969 ;
  assign n2403 = ~n2396 & ~n2402 ;
  assign n2404 = ~x743 & n2403 ;
  assign n2407 = n2404 ^ n2403 ;
  assign n2405 = n2404 ^ n2388 ;
  assign n2406 = n2393 & n2405 ;
  assign n2408 = n2407 ^ n2406 ;
  assign n2422 = ~x739 & ~n2408 ;
  assign n2423 = n2422 ^ x743 ;
  assign n2424 = ~n2418 & ~n2423 ;
  assign n2409 = n2408 ^ x743 ;
  assign n2425 = n2424 ^ n2409 ;
  assign n2410 = ~x739 & ~n2409 ;
  assign n2412 = n2410 & n2411 ;
  assign n2413 = n2387 & n2412 ;
  assign n2426 = n2425 ^ n2413 ;
  assign n2385 = n2381 ^ x739 ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2427 = n2426 ^ n2386 ;
  assign n2356 = ~n2339 & ~n2359 ;
  assign n2370 = n2366 ^ n2358 ;
  assign n2340 = n2370 ^ n2339 ;
  assign n2345 = n1961 & ~n2340 ;
  assign n2342 = n1961 ^ x747 ;
  assign n2343 = n2342 ^ n2340 ;
  assign n2346 = n2345 ^ n2343 ;
  assign n2347 = n2339 ^ n1961 ;
  assign n2348 = n2347 ^ n2340 ;
  assign n2349 = n2348 ^ n2343 ;
  assign n2350 = ~n2346 & n2349 ;
  assign n2351 = ~n1962 & n2350 ;
  assign n2352 = n2351 ^ n2345 ;
  assign n2353 = n2352 ^ x745 ;
  assign n2354 = ~n2335 & n2353 ;
  assign n2357 = n2356 ^ n2354 ;
  assign n2362 = ~x750 & n2361 ;
  assign n2363 = ~n2357 & n2362 ;
  assign n2364 = n2363 ^ n2357 ;
  assign n2376 = n2375 ^ n2364 ;
  assign n2428 = n2427 ^ n2376 ;
  assign n2430 = n2429 ^ n2428 ;
  assign n2434 = n2433 ^ n2430 ;
  assign n2436 = n2435 ^ n2434 ;
  assign n1963 = n1962 ^ n1961 ;
  assign n1965 = n1964 ^ n1963 ;
  assign n1966 = x740 ^ x739 ;
  assign n1970 = n1969 ^ n1966 ;
  assign n2304 = n1965 & n1970 ;
  assign n10821 = n2436 ^ n2304 ;
  assign n1960 = n1959 ^ n1954 ;
  assign n1971 = n1970 ^ n1965 ;
  assign n2303 = n1960 & n1971 ;
  assign n10823 = n2306 ^ n2303 ;
  assign n10826 = n10821 & n10823 ;
  assign n10822 = n10821 ^ n2306 ;
  assign n10824 = n10823 ^ n10822 ;
  assign n10825 = ~n2333 & n10824 ;
  assign n10827 = n10826 ^ n10825 ;
  assign n10861 = n10860 ^ n10827 ;
  assign n10815 = n2409 ^ x739 ;
  assign n10816 = n10815 ^ n2410 ;
  assign n10817 = n2418 & n10816 ;
  assign n10818 = n10817 ^ n2364 ;
  assign n10812 = n2427 ^ n2304 ;
  assign n10813 = n2436 & ~n10812 ;
  assign n10814 = n10813 ^ n2427 ;
  assign n10819 = n10818 ^ n10814 ;
  assign n10802 = n2321 ^ n2316 ;
  assign n10808 = n1956 & n10805 ;
  assign n10809 = n10808 ^ n10804 ;
  assign n10810 = n10802 & ~n10809 ;
  assign n10811 = n10810 ^ n2316 ;
  assign n10820 = n10819 ^ n10811 ;
  assign n10862 = n10861 ^ n10820 ;
  assign n1972 = n1971 ^ n1960 ;
  assign n1992 = x708 ^ x707 ;
  assign n1990 = x704 ^ x703 ;
  assign n1989 = x706 ^ x705 ;
  assign n1991 = n1990 ^ n1989 ;
  assign n1993 = n1992 ^ n1991 ;
  assign n1987 = x714 ^ x713 ;
  assign n1985 = x710 ^ x709 ;
  assign n1984 = x712 ^ x711 ;
  assign n1986 = n1985 ^ n1984 ;
  assign n1988 = n1987 ^ n1986 ;
  assign n1994 = n1993 ^ n1988 ;
  assign n1980 = x724 ^ x723 ;
  assign n1979 = x722 ^ x721 ;
  assign n1981 = n1980 ^ n1979 ;
  assign n1978 = x726 ^ x725 ;
  assign n1982 = n1981 ^ n1978 ;
  assign n1975 = x716 ^ x715 ;
  assign n1974 = x718 ^ x717 ;
  assign n1976 = n1975 ^ n1974 ;
  assign n1973 = x720 ^ x719 ;
  assign n1977 = n1976 ^ n1973 ;
  assign n1983 = n1982 ^ n1977 ;
  assign n1995 = n1994 ^ n1983 ;
  assign n2484 = n1972 & n1995 ;
  assign n2480 = ~x705 & ~x706 ;
  assign n2477 = x707 & ~n1992 ;
  assign n2476 = x703 & ~n1990 ;
  assign n2478 = n2477 ^ n2476 ;
  assign n2474 = n1992 ^ n1990 ;
  assign n2475 = n1991 & ~n2474 ;
  assign n2479 = n2478 ^ n2475 ;
  assign n2481 = n2480 ^ n2479 ;
  assign n2472 = ~x711 & ~x712 ;
  assign n2469 = x713 & ~n1987 ;
  assign n2468 = x709 & ~n1985 ;
  assign n2470 = n2469 ^ n2468 ;
  assign n2466 = n1987 ^ n1985 ;
  assign n2467 = n1986 & ~n2466 ;
  assign n2471 = n2470 ^ n2467 ;
  assign n2473 = n2472 ^ n2471 ;
  assign n2482 = n2481 ^ n2473 ;
  assign n2459 = x715 & x716 ;
  assign n2460 = n2459 ^ n1973 ;
  assign n2458 = ~x719 & ~x720 ;
  assign n2461 = n2460 ^ n2458 ;
  assign n2457 = ~x717 & ~x718 ;
  assign n2462 = n2461 ^ n2457 ;
  assign n2452 = x721 & x722 ;
  assign n2453 = n2452 ^ n1978 ;
  assign n2451 = ~x725 & ~x726 ;
  assign n2454 = n2453 ^ n2451 ;
  assign n2450 = ~x723 & ~x724 ;
  assign n2455 = n2454 ^ n2450 ;
  assign n2448 = n1979 ^ n1978 ;
  assign n2449 = n1981 & ~n2448 ;
  assign n2456 = n2455 ^ n2449 ;
  assign n2463 = n2462 ^ n2456 ;
  assign n2446 = n1974 ^ n1973 ;
  assign n2447 = n1976 & n2446 ;
  assign n2464 = n2463 ^ n2447 ;
  assign n2443 = n1977 & n1982 ;
  assign n2441 = n1988 & n1993 ;
  assign n2438 = n1988 ^ n1983 ;
  assign n2439 = n1994 & ~n2438 ;
  assign n2440 = n2439 ^ n1993 ;
  assign n2442 = n2441 ^ n2440 ;
  assign n2444 = n2443 ^ n2442 ;
  assign n2445 = n2444 ^ n2441 ;
  assign n2465 = n2464 ^ n2445 ;
  assign n2483 = n2482 ^ n2465 ;
  assign n2485 = n2484 ^ n2483 ;
  assign n2305 = n2304 ^ n2303 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2334 = n2333 ^ n2307 ;
  assign n2437 = n2436 ^ n2334 ;
  assign n10799 = n2484 ^ n2437 ;
  assign n10800 = n2485 & ~n10799 ;
  assign n10772 = n2480 ^ n1989 ;
  assign n10773 = x708 & n2476 ;
  assign n10774 = ~n10772 & n10773 ;
  assign n10775 = n10774 ^ n2476 ;
  assign n10769 = n2477 ^ n1992 ;
  assign n10770 = ~n2480 & n10769 ;
  assign n10776 = n10775 ^ n10770 ;
  assign n10781 = ~n2477 & n10772 ;
  assign n10782 = n10781 ^ n10770 ;
  assign n10783 = n10776 & n10782 ;
  assign n10785 = n10783 ^ n10775 ;
  assign n10771 = ~n1990 & n10770 ;
  assign n10784 = n10771 & n10783 ;
  assign n10786 = n10785 ^ n10784 ;
  assign n10787 = n10772 ^ n2477 ;
  assign n10788 = x704 & n10770 ;
  assign n10789 = n10788 ^ n2477 ;
  assign n10790 = ~n10787 & n10789 ;
  assign n10791 = n10790 ^ n2477 ;
  assign n10792 = ~n10786 & n10791 ;
  assign n10793 = n10792 ^ n10786 ;
  assign n10734 = n2472 ^ n1984 ;
  assign n10735 = n10734 ^ n2469 ;
  assign n10736 = n2469 ^ n1987 ;
  assign n10737 = ~n2472 & n10736 ;
  assign n10742 = x710 & n10737 ;
  assign n10743 = n10742 ^ n10734 ;
  assign n10744 = ~n10735 & n10743 ;
  assign n10745 = n10744 ^ n2469 ;
  assign n10746 = x714 & n2468 ;
  assign n10747 = ~n10734 & n10746 ;
  assign n10748 = n10747 ^ n2468 ;
  assign n10749 = n10748 ^ n10737 ;
  assign n10754 = ~n2469 & n10734 ;
  assign n10755 = n10754 ^ n10748 ;
  assign n10756 = n10749 & ~n10755 ;
  assign n10764 = n10737 & n10756 ;
  assign n10765 = ~n1985 & n10764 ;
  assign n10766 = n10765 ^ n1985 ;
  assign n10757 = n10756 ^ n10748 ;
  assign n10758 = n10757 ^ n1985 ;
  assign n10767 = n10766 ^ n10758 ;
  assign n10768 = ~n10745 & ~n10767 ;
  assign n10794 = n10793 ^ n10768 ;
  assign n10731 = n2473 ^ n2441 ;
  assign n10732 = n2482 & ~n10731 ;
  assign n10733 = n10732 ^ n2473 ;
  assign n10795 = n10794 ^ n10733 ;
  assign n10705 = n2450 ^ n1980 ;
  assign n10706 = x726 & n2452 ;
  assign n10707 = ~n10705 & n10706 ;
  assign n10708 = n10707 ^ n2452 ;
  assign n10703 = ~n2450 & ~n2451 ;
  assign n10709 = n10708 ^ n10703 ;
  assign n10710 = n2451 ^ n1978 ;
  assign n10715 = n10705 & n10710 ;
  assign n10716 = n10715 ^ n10703 ;
  assign n10717 = n10709 & n10716 ;
  assign n10719 = n10717 ^ n10708 ;
  assign n10704 = ~n1979 & n10703 ;
  assign n10718 = n10704 & n10717 ;
  assign n10720 = n10719 ^ n10718 ;
  assign n10721 = n10710 ^ n10705 ;
  assign n10722 = x722 & n10703 ;
  assign n10723 = n10722 ^ n10705 ;
  assign n10724 = n10721 & ~n10723 ;
  assign n10725 = n10724 ^ n10705 ;
  assign n10726 = ~n10720 & ~n10725 ;
  assign n10727 = n10726 ^ n10720 ;
  assign n10669 = n2458 ^ n1973 ;
  assign n10668 = n2457 ^ n1974 ;
  assign n10670 = n10669 ^ n10668 ;
  assign n10671 = ~n2457 & ~n2458 ;
  assign n10676 = x716 & n10671 ;
  assign n10677 = n10676 ^ n10668 ;
  assign n10678 = n10670 & n10677 ;
  assign n10679 = n10678 ^ n10669 ;
  assign n10680 = x720 & n2459 ;
  assign n10681 = ~n10668 & n10680 ;
  assign n10682 = n10681 ^ n2459 ;
  assign n10683 = n10682 ^ n10671 ;
  assign n10688 = n10668 & n10669 ;
  assign n10689 = n10688 ^ n10682 ;
  assign n10690 = n10683 & ~n10689 ;
  assign n10698 = ~n1975 & n10690 ;
  assign n10699 = n10671 & n10698 ;
  assign n10700 = n10699 ^ n10671 ;
  assign n10691 = n10690 ^ n10682 ;
  assign n10692 = n10691 ^ n10671 ;
  assign n10701 = n10700 ^ n10692 ;
  assign n10702 = n10679 & ~n10701 ;
  assign n10728 = n10727 ^ n10702 ;
  assign n10665 = n2456 ^ n2443 ;
  assign n10666 = n2464 & n10665 ;
  assign n10667 = n10666 ^ n2456 ;
  assign n10729 = n10728 ^ n10667 ;
  assign n10658 = n2464 ^ n2443 ;
  assign n10662 = n2443 ^ n2441 ;
  assign n10663 = n10658 & ~n10662 ;
  assign n10657 = n2482 ^ n2464 ;
  assign n10659 = n10658 ^ n2441 ;
  assign n10660 = n10659 ^ n2440 ;
  assign n10661 = n10657 & n10660 ;
  assign n10664 = n10663 ^ n10661 ;
  assign n10730 = n10729 ^ n10664 ;
  assign n10796 = n10795 ^ n10730 ;
  assign n10797 = n10796 ^ n2484 ;
  assign n10801 = n10800 ^ n10797 ;
  assign n10863 = n10862 ^ n10801 ;
  assign n10990 = n10989 ^ n10863 ;
  assign n2486 = n2485 ^ n2437 ;
  assign n1949 = n1948 ^ n1925 ;
  assign n1996 = n1995 ^ n1972 ;
  assign n2011 = n1949 & n1996 ;
  assign n10652 = n2486 ^ n2011 ;
  assign n10653 = n2301 ^ n2012 ;
  assign n10654 = n10653 ^ n2011 ;
  assign n10655 = ~n10652 & ~n10654 ;
  assign n10656 = n10655 ^ n2486 ;
  assign n10991 = n10990 ^ n10656 ;
  assign n2585 = x771 & x772 ;
  assign n2584 = x773 & x774 ;
  assign n2586 = n2585 ^ n2584 ;
  assign n1869 = x774 ^ x773 ;
  assign n2587 = n2584 ^ n1869 ;
  assign n1867 = x772 ^ x771 ;
  assign n2588 = n2585 ^ n1867 ;
  assign n2589 = n2587 & n2588 ;
  assign n2590 = n2589 ^ n2584 ;
  assign n2591 = ~n2586 & ~n2590 ;
  assign n2563 = n1867 ^ x770 ;
  assign n2564 = n2563 ^ n1869 ;
  assign n1872 = x766 ^ x765 ;
  assign n2572 = n1872 ^ x767 ;
  assign n1871 = x764 ^ x763 ;
  assign n2573 = n2572 ^ n1871 ;
  assign n2574 = n1872 ^ x768 ;
  assign n2566 = ~x765 & ~x766 ;
  assign n2575 = n2574 ^ n2566 ;
  assign n2576 = n2573 & n2575 ;
  assign n2565 = x767 ^ x764 ;
  assign n2569 = n2566 ^ n2565 ;
  assign n2570 = x763 & n2569 ;
  assign n2567 = n2566 ^ x767 ;
  assign n2568 = ~n2565 & n2567 ;
  assign n2571 = n2570 ^ n2568 ;
  assign n2577 = n2576 ^ n2571 ;
  assign n2578 = n2577 ^ x769 ;
  assign n2579 = n2578 ^ n1867 ;
  assign n2580 = n2579 ^ n1869 ;
  assign n2581 = n2580 ^ n2577 ;
  assign n2582 = ~n2564 & n2581 ;
  assign n2583 = n2582 ^ n2578 ;
  assign n2592 = n2591 ^ n2583 ;
  assign n1866 = x770 ^ x769 ;
  assign n1868 = n1867 ^ n1866 ;
  assign n1870 = n1869 ^ n1868 ;
  assign n1874 = x768 ^ x767 ;
  assign n1873 = n1872 ^ n1871 ;
  assign n1875 = n1874 ^ n1873 ;
  assign n10580 = n1870 & n1875 ;
  assign n10643 = n10580 ^ n2577 ;
  assign n10644 = n2592 & ~n10643 ;
  assign n10645 = n10644 ^ n2577 ;
  assign n10598 = n2589 ^ x770 ;
  assign n10599 = n2586 ^ x769 ;
  assign n10600 = n10599 ^ n2589 ;
  assign n10601 = n10598 & ~n10600 ;
  assign n10602 = n10601 ^ n2590 ;
  assign n10603 = ~n2586 & n10602 ;
  assign n10604 = x769 & n10603 ;
  assign n10605 = n10601 ^ n2589 ;
  assign n10606 = n10605 ^ n10603 ;
  assign n10641 = n10604 & ~n10606 ;
  assign n10636 = n2572 ^ x768 ;
  assign n10609 = n1874 & n2574 ;
  assign n10610 = n10609 ^ x767 ;
  assign n10611 = ~n2566 & n10610 ;
  assign n10612 = n10611 ^ x764 ;
  assign n10613 = ~n1871 & n10612 ;
  assign n10637 = n10636 ^ n10613 ;
  assign n10621 = ~n2572 & ~n10636 ;
  assign n10622 = n10621 ^ n10613 ;
  assign n10631 = n10613 ^ x768 ;
  assign n10624 = n10637 ^ x767 ;
  assign n10623 = n10637 ^ x766 ;
  assign n10625 = n10624 ^ n10623 ;
  assign n10619 = n10637 ^ x768 ;
  assign n10626 = n10623 ^ n10619 ;
  assign n10627 = n10637 ^ n10626 ;
  assign n10628 = n10627 ^ n10613 ;
  assign n10629 = ~n10625 & ~n10628 ;
  assign n10632 = n10631 ^ n10629 ;
  assign n10633 = ~n10622 & ~n10632 ;
  assign n10638 = n10637 ^ n10633 ;
  assign n10639 = n10638 ^ n10606 ;
  assign n10642 = n10641 ^ n10639 ;
  assign n10646 = n10645 ^ n10642 ;
  assign n2511 = ~x755 & ~x756 ;
  assign n1858 = x756 ^ x755 ;
  assign n2514 = n2511 ^ n1858 ;
  assign n2512 = ~x753 & ~x754 ;
  assign n1856 = x754 ^ x753 ;
  assign n2515 = n2512 ^ n1856 ;
  assign n2516 = n2514 & n2515 ;
  assign n2513 = ~n2511 & ~n2512 ;
  assign n2518 = n2516 ^ n2513 ;
  assign n2517 = ~n2513 & n2516 ;
  assign n2519 = n2518 ^ n2517 ;
  assign n2520 = ~x752 & n2519 ;
  assign n2522 = n2520 ^ x751 ;
  assign n2521 = x751 & ~n2520 ;
  assign n2523 = n2522 ^ n2521 ;
  assign n2524 = n2523 ^ n2519 ;
  assign n2525 = n2515 ^ n2514 ;
  assign n2526 = n2525 ^ n2516 ;
  assign n2527 = ~n2524 & n2526 ;
  assign n2537 = x751 & x752 ;
  assign n2542 = x756 & ~n2515 ;
  assign n2543 = n2542 ^ n2517 ;
  assign n2544 = n2537 & ~n2543 ;
  assign n10596 = n2527 & ~n2544 ;
  assign n1860 = x758 ^ x757 ;
  assign n2490 = x761 & x762 ;
  assign n1863 = x762 ^ x761 ;
  assign n2491 = n2490 ^ n1863 ;
  assign n2492 = x759 & x760 ;
  assign n1861 = x760 ^ x759 ;
  assign n2493 = n2492 ^ n1861 ;
  assign n2494 = n2491 & n2493 ;
  assign n2500 = n2494 ^ n2490 ;
  assign n10585 = n2500 ^ n2492 ;
  assign n10586 = n10585 ^ x758 ;
  assign n10587 = n1860 & n10586 ;
  assign n10591 = n10587 ^ x757 ;
  assign n2496 = n2492 ^ n2490 ;
  assign n10588 = n2490 ^ x757 ;
  assign n10589 = n10588 ^ n10587 ;
  assign n10590 = ~n2496 & n10589 ;
  assign n10592 = n10591 ^ n10590 ;
  assign n10593 = n2494 & n10590 ;
  assign n10594 = ~n10592 & n10593 ;
  assign n10595 = n10594 ^ n10592 ;
  assign n10597 = n10596 ^ n10595 ;
  assign n10647 = n10646 ^ n10597 ;
  assign n1855 = x752 ^ x751 ;
  assign n1857 = n1856 ^ n1855 ;
  assign n1859 = n1858 ^ n1857 ;
  assign n1862 = n1861 ^ n1860 ;
  assign n1864 = n1863 ^ n1862 ;
  assign n2561 = n1859 & n1864 ;
  assign n2501 = n2500 ^ n1860 ;
  assign n2502 = ~n2496 & ~n2501 ;
  assign n2495 = n1863 ^ n1861 ;
  assign n2497 = n2496 ^ n2495 ;
  assign n2498 = n2497 ^ x758 ;
  assign n2499 = n2498 ^ n2494 ;
  assign n2503 = n2502 ^ n2499 ;
  assign n2504 = n2503 ^ n2498 ;
  assign n2506 = n2494 ^ x758 ;
  assign n2507 = n2506 ^ n2498 ;
  assign n2508 = n2504 & ~n2507 ;
  assign n2509 = n2508 ^ n2498 ;
  assign n2558 = n1860 & n2509 ;
  assign n2555 = n2502 ^ x757 ;
  assign n2529 = x755 ^ x752 ;
  assign n2532 = ~n1858 & n2529 ;
  assign n2533 = n2532 ^ x752 ;
  assign n2534 = n2512 & ~n2533 ;
  assign n2535 = n2534 ^ n2527 ;
  assign n2536 = ~n2521 & ~n2535 ;
  assign n2545 = n1856 ^ x751 ;
  assign n2546 = n2512 ^ n1855 ;
  assign n2547 = ~x755 & ~n2546 ;
  assign n2548 = n1856 ^ x756 ;
  assign n2549 = n2548 ^ n1855 ;
  assign n2550 = n2547 & n2549 ;
  assign n2551 = n2545 & n2550 ;
  assign n2552 = n2551 ^ n2544 ;
  assign n2553 = ~n2536 & ~n2552 ;
  assign n2556 = n2555 ^ n2553 ;
  assign n2559 = n2558 ^ n2556 ;
  assign n2560 = n2559 ^ n1875 ;
  assign n2562 = n2561 ^ n2560 ;
  assign n2593 = n2592 ^ n2562 ;
  assign n1876 = n1875 ^ n1870 ;
  assign n1865 = n1864 ^ n1859 ;
  assign n2488 = n1870 ^ n1865 ;
  assign n2489 = n1876 & ~n2488 ;
  assign n2594 = n2593 ^ n2489 ;
  assign n10577 = n2594 ^ n2559 ;
  assign n10581 = n10580 ^ n2592 ;
  assign n10582 = n10581 ^ n2594 ;
  assign n10583 = ~n10577 & ~n10582 ;
  assign n10579 = ~n2553 & n2559 ;
  assign n10584 = n10583 ^ n10579 ;
  assign n10648 = n10647 ^ n10584 ;
  assign n2724 = x779 & x780 ;
  assign n2723 = x777 & x778 ;
  assign n2725 = n2724 ^ n2723 ;
  assign n1892 = x780 ^ x779 ;
  assign n2726 = n2724 ^ n1892 ;
  assign n1890 = x778 ^ x777 ;
  assign n2727 = n2723 ^ n1890 ;
  assign n2728 = n2726 & n2727 ;
  assign n2729 = n2728 ^ n2724 ;
  assign n2730 = ~n2725 & ~n2729 ;
  assign n2676 = n1892 ^ x776 ;
  assign n2677 = n2676 ^ n1890 ;
  assign n1897 = x786 ^ x785 ;
  assign n2679 = x785 ^ x784 ;
  assign n2683 = ~n1897 & ~n2679 ;
  assign n2678 = x783 ^ x782 ;
  assign n2680 = n2679 ^ x783 ;
  assign n2681 = n2680 ^ x786 ;
  assign n2682 = ~n2678 & n2681 ;
  assign n2684 = n2683 ^ n2682 ;
  assign n2685 = ~x781 & n2684 ;
  assign n1895 = x784 ^ x783 ;
  assign n2686 = ~n1895 & ~n2678 ;
  assign n2687 = x786 ^ x781 ;
  assign n2690 = ~x784 & ~n2687 ;
  assign n2691 = n2690 ^ x781 ;
  assign n2692 = n2686 & n2691 ;
  assign n2693 = ~x785 & n2692 ;
  assign n2694 = ~x783 & ~x784 ;
  assign n2697 = n2694 ^ n1895 ;
  assign n2698 = x781 & x782 ;
  assign n2699 = x786 & n2698 ;
  assign n2700 = ~n2697 & n2699 ;
  assign n2701 = n2700 ^ n2698 ;
  assign n2695 = ~x785 & ~x786 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2702 = n2701 ^ n2696 ;
  assign n2703 = n2695 ^ n1897 ;
  assign n2708 = n2697 & n2703 ;
  assign n2709 = n2708 ^ n2696 ;
  assign n2710 = n2702 & n2709 ;
  assign n1894 = x782 ^ x781 ;
  assign n2711 = n2710 ^ n2701 ;
  assign n2712 = ~n1894 & n2711 ;
  assign n2713 = n2710 & n2712 ;
  assign n2714 = n2713 ^ n2711 ;
  assign n2715 = ~n2693 & ~n2714 ;
  assign n2716 = ~n2685 & n2715 ;
  assign n2717 = n2716 ^ x775 ;
  assign n2718 = n2717 ^ n1892 ;
  assign n2719 = n2718 ^ n1890 ;
  assign n2720 = n2719 ^ n2716 ;
  assign n2721 = ~n2677 & n2720 ;
  assign n2722 = n2721 ^ n2717 ;
  assign n2731 = n2730 ^ n2722 ;
  assign n1889 = x776 ^ x775 ;
  assign n1891 = n1890 ^ n1889 ;
  assign n1893 = n1892 ^ n1891 ;
  assign n10555 = n2731 ^ n1893 ;
  assign n1896 = n1895 ^ n1894 ;
  assign n1898 = n1897 ^ n1896 ;
  assign n1899 = n1898 ^ n1893 ;
  assign n1881 = x792 ^ x791 ;
  assign n1879 = x790 ^ x789 ;
  assign n1878 = x788 ^ x787 ;
  assign n1880 = n1879 ^ n1878 ;
  assign n1882 = n1881 ^ n1880 ;
  assign n1886 = x798 ^ x797 ;
  assign n1884 = x796 ^ x795 ;
  assign n1883 = x794 ^ x793 ;
  assign n1885 = n1884 ^ n1883 ;
  assign n1887 = n1886 ^ n1885 ;
  assign n1888 = n1887 ^ n1882 ;
  assign n1900 = n1899 ^ n1888 ;
  assign n2738 = ~n1882 & n1900 ;
  assign n2636 = x791 ^ x790 ;
  assign n2640 = ~n1881 & ~n2636 ;
  assign n2635 = x789 ^ x788 ;
  assign n2637 = n2636 ^ x789 ;
  assign n2638 = n2637 ^ x792 ;
  assign n2639 = ~n2635 & n2638 ;
  assign n2641 = n2640 ^ n2639 ;
  assign n2642 = ~x787 & n2641 ;
  assign n2643 = ~n1879 & ~n2635 ;
  assign n2644 = x792 ^ x787 ;
  assign n2647 = ~x790 & ~n2644 ;
  assign n2648 = n2647 ^ x787 ;
  assign n2649 = n2643 & n2648 ;
  assign n2650 = ~x791 & n2649 ;
  assign n2651 = ~x789 & ~x790 ;
  assign n2654 = n2651 ^ n1879 ;
  assign n2655 = x787 & x788 ;
  assign n2656 = x792 & n2655 ;
  assign n2657 = ~n2654 & n2656 ;
  assign n2658 = n2657 ^ n2655 ;
  assign n2652 = ~x791 & ~x792 ;
  assign n2653 = ~n2651 & ~n2652 ;
  assign n2659 = n2658 ^ n2653 ;
  assign n2660 = n2652 ^ n1881 ;
  assign n2665 = n2654 & n2660 ;
  assign n2666 = n2665 ^ n2653 ;
  assign n2667 = n2659 & n2666 ;
  assign n2668 = n2667 ^ n2658 ;
  assign n2669 = ~n1878 & n2668 ;
  assign n2670 = n2667 & n2669 ;
  assign n2671 = n2670 ^ n2668 ;
  assign n2672 = ~n2650 & ~n2671 ;
  assign n2673 = ~n2642 & n2672 ;
  assign n2597 = x797 ^ x796 ;
  assign n2601 = ~n1886 & ~n2597 ;
  assign n2596 = x795 ^ x794 ;
  assign n2598 = n2597 ^ x795 ;
  assign n2599 = n2598 ^ x798 ;
  assign n2600 = ~n2596 & n2599 ;
  assign n2602 = n2601 ^ n2600 ;
  assign n2603 = ~x793 & n2602 ;
  assign n2604 = ~n1884 & ~n2596 ;
  assign n2605 = x798 ^ x793 ;
  assign n2608 = ~x796 & ~n2605 ;
  assign n2609 = n2608 ^ x793 ;
  assign n2610 = n2604 & n2609 ;
  assign n2611 = ~x797 & n2610 ;
  assign n2612 = ~x795 & ~x796 ;
  assign n2615 = n2612 ^ n1884 ;
  assign n2616 = x793 & x794 ;
  assign n2617 = x798 & n2616 ;
  assign n2618 = ~n2615 & n2617 ;
  assign n2619 = n2618 ^ n2616 ;
  assign n2613 = ~x797 & ~x798 ;
  assign n2614 = ~n2612 & ~n2613 ;
  assign n2620 = n2619 ^ n2614 ;
  assign n2621 = n2613 ^ n1886 ;
  assign n2626 = n2615 & n2621 ;
  assign n2627 = n2626 ^ n2614 ;
  assign n2628 = n2620 & n2627 ;
  assign n2629 = n2628 ^ n2619 ;
  assign n2630 = ~n1883 & n2629 ;
  assign n2631 = n2628 & n2630 ;
  assign n2632 = n2631 ^ n2629 ;
  assign n2633 = ~n2611 & ~n2632 ;
  assign n2634 = ~n2603 & n2633 ;
  assign n2674 = n2673 ^ n2634 ;
  assign n10556 = n2738 ^ n2674 ;
  assign n2736 = n1893 & n1898 ;
  assign n10561 = n2731 & ~n2736 ;
  assign n10562 = n10561 ^ n2738 ;
  assign n10563 = ~n10556 & ~n10562 ;
  assign n10564 = n10563 ^ n2674 ;
  assign n2734 = ~n1887 & ~n1899 ;
  assign n2595 = n1882 & n1887 ;
  assign n2735 = n2734 ^ n2595 ;
  assign n10568 = ~n2674 & n2735 ;
  assign n10569 = n10568 ^ n2595 ;
  assign n10570 = n10564 & ~n10569 ;
  assign n10571 = ~n1899 & n10570 ;
  assign n10572 = n10555 & n10571 ;
  assign n10573 = n10572 ^ n10570 ;
  assign n10551 = n2736 ^ n2716 ;
  assign n10552 = ~n2731 & n10551 ;
  assign n10553 = n10552 ^ n2716 ;
  assign n10546 = n2673 ^ n2595 ;
  assign n10547 = n2674 & n10546 ;
  assign n10548 = n10547 ^ n2673 ;
  assign n10538 = n2660 ^ n2654 ;
  assign n10539 = x788 & n2653 ;
  assign n10540 = n10539 ^ n2654 ;
  assign n10541 = n10538 & ~n10540 ;
  assign n10542 = n10541 ^ n2654 ;
  assign n10543 = ~n2671 & ~n10542 ;
  assign n10544 = n10543 ^ n2671 ;
  assign n10532 = n2621 ^ n2615 ;
  assign n10533 = x794 & n2614 ;
  assign n10534 = n10533 ^ n2615 ;
  assign n10535 = n10532 & ~n10534 ;
  assign n10536 = n10535 ^ n2615 ;
  assign n10537 = ~n2632 & n10536 ;
  assign n10545 = n10544 ^ n10537 ;
  assign n10549 = n10548 ^ n10545 ;
  assign n10524 = n2703 ^ n2697 ;
  assign n10525 = x782 & n2696 ;
  assign n10526 = n10525 ^ n2697 ;
  assign n10527 = n10524 & ~n10526 ;
  assign n10528 = n10527 ^ n2697 ;
  assign n10529 = ~n2714 & ~n10528 ;
  assign n10530 = n10529 ^ n2714 ;
  assign n10513 = n2728 ^ x776 ;
  assign n10514 = n2725 ^ x775 ;
  assign n10515 = n10514 ^ n2728 ;
  assign n10516 = n10513 & ~n10515 ;
  assign n10519 = n10516 ^ n2728 ;
  assign n10517 = n10516 ^ n2729 ;
  assign n10518 = ~n2725 & n10517 ;
  assign n10520 = n10519 ^ n10518 ;
  assign n10521 = x775 & n10518 ;
  assign n10522 = ~n10520 & n10521 ;
  assign n10523 = n10522 ^ n10520 ;
  assign n10531 = n10530 ^ n10523 ;
  assign n10550 = n10549 ^ n10531 ;
  assign n10554 = n10553 ^ n10550 ;
  assign n10574 = n10573 ^ n10554 ;
  assign n1877 = n1876 ^ n1865 ;
  assign n2733 = n1877 & n1900 ;
  assign n10575 = n10574 ^ n2733 ;
  assign n2737 = n2736 ^ n2735 ;
  assign n2739 = n2738 ^ n2737 ;
  assign n2740 = n2739 ^ n2733 ;
  assign n2675 = n2674 ^ n2595 ;
  assign n2732 = n2731 ^ n2675 ;
  assign n2741 = n2740 ^ n2732 ;
  assign n10511 = n2733 ^ n2594 ;
  assign n10512 = n2741 & ~n10511 ;
  assign n10576 = n10575 ^ n10512 ;
  assign n10649 = n10648 ^ n10576 ;
  assign n2994 = x825 & x826 ;
  assign n2995 = n2994 ^ x824 ;
  assign n1837 = x826 ^ x825 ;
  assign n2998 = n1837 ^ x823 ;
  assign n2999 = ~x828 & n2998 ;
  assign n3000 = n2999 ^ x823 ;
  assign n3001 = ~n2994 & n3000 ;
  assign n3002 = n3001 ^ x823 ;
  assign n3003 = ~n2995 & n3002 ;
  assign n3004 = ~x827 & n3003 ;
  assign n3005 = ~x823 & ~n3004 ;
  assign n3006 = x827 & x828 ;
  assign n1839 = x828 ^ x827 ;
  assign n3007 = n3006 ^ n1839 ;
  assign n3008 = x824 & n3007 ;
  assign n3010 = n3006 ^ x826 ;
  assign n3009 = n2994 & n3006 ;
  assign n3016 = n3010 ^ n3009 ;
  assign n3011 = n1837 & ~n3010 ;
  assign n3017 = n3016 ^ n3011 ;
  assign n3022 = ~n3008 & ~n3017 ;
  assign n3012 = n3011 ^ x825 ;
  assign n3013 = ~n3009 & n3012 ;
  assign n3014 = ~n3008 & n3013 ;
  assign n3015 = n3014 ^ n3012 ;
  assign n3023 = n3022 ^ n3015 ;
  assign n3024 = n3005 & n3023 ;
  assign n3025 = n3024 ^ n3004 ;
  assign n1836 = x824 ^ x823 ;
  assign n3028 = n3017 ^ n3012 ;
  assign n3029 = n3028 ^ n2994 ;
  assign n3030 = n3029 ^ n3012 ;
  assign n3031 = x824 & n3030 ;
  assign n3032 = n3031 ^ n3012 ;
  assign n3033 = ~n1836 & n3032 ;
  assign n3034 = n3033 ^ n3012 ;
  assign n3035 = n3007 & n3034 ;
  assign n3036 = x823 & x824 ;
  assign n3037 = ~x828 & n2994 ;
  assign n3038 = n3036 & n3037 ;
  assign n3039 = ~n3035 & ~n3038 ;
  assign n3040 = ~n3025 & n3039 ;
  assign n1833 = x830 ^ x829 ;
  assign n1832 = x832 ^ x831 ;
  assign n1834 = n1833 ^ n1832 ;
  assign n1831 = x834 ^ x833 ;
  assign n1835 = n1834 ^ n1831 ;
  assign n1838 = n1837 ^ n1836 ;
  assign n1840 = n1839 ^ n1838 ;
  assign n2993 = n1835 & n1840 ;
  assign n3041 = n3040 ^ n2993 ;
  assign n2959 = ~x833 & ~x834 ;
  assign n2960 = ~x831 & ~x832 ;
  assign n2963 = n2959 ^ n1831 ;
  assign n2966 = n2960 & n2963 ;
  assign n2982 = n2966 ^ x829 ;
  assign n2983 = n2959 ^ n1834 ;
  assign n2984 = n2983 ^ n2966 ;
  assign n2985 = n2982 & n2984 ;
  assign n2988 = ~n2966 & n2985 ;
  assign n2970 = n1833 & ~n2959 ;
  assign n2964 = n2963 ^ x832 ;
  assign n2965 = n1832 & n2964 ;
  assign n2973 = n2965 ^ x831 ;
  assign n2978 = n2970 & n2973 ;
  assign n2974 = x829 & x830 ;
  assign n2967 = n2966 ^ n2964 ;
  assign n2968 = n2967 ^ n2965 ;
  assign n2961 = n2960 ^ n1832 ;
  assign n2962 = n2959 & n2961 ;
  assign n2969 = n2968 ^ n2962 ;
  assign n2975 = ~n2966 & ~n2969 ;
  assign n2976 = n2974 & n2975 ;
  assign n2979 = n2978 ^ n2976 ;
  assign n2989 = n2988 ^ n2979 ;
  assign n2990 = ~n2959 & n2989 ;
  assign n2991 = n2990 ^ n2985 ;
  assign n2971 = ~x830 & ~n2970 ;
  assign n2972 = n2969 & n2971 ;
  assign n2992 = n2991 ^ n2972 ;
  assign n3042 = n3041 ^ n2992 ;
  assign n1841 = n1840 ^ n1835 ;
  assign n1850 = x840 ^ x839 ;
  assign n1848 = x836 ^ x835 ;
  assign n1847 = x838 ^ x837 ;
  assign n1849 = n1848 ^ n1847 ;
  assign n1851 = n1850 ^ n1849 ;
  assign n1845 = x846 ^ x845 ;
  assign n1843 = x842 ^ x841 ;
  assign n1842 = x844 ^ x843 ;
  assign n1844 = n1843 ^ n1842 ;
  assign n1846 = n1845 ^ n1844 ;
  assign n1852 = n1851 ^ n1846 ;
  assign n2956 = n1841 & n1852 ;
  assign n2955 = n1846 & n1851 ;
  assign n2957 = n2956 ^ n2955 ;
  assign n2952 = ~x837 & ~x838 ;
  assign n2949 = x839 & ~n1850 ;
  assign n2948 = x835 & ~n1848 ;
  assign n2950 = n2949 ^ n2948 ;
  assign n2946 = n1850 ^ n1848 ;
  assign n2947 = n1849 & ~n2946 ;
  assign n2951 = n2950 ^ n2947 ;
  assign n2953 = n2952 ^ n2951 ;
  assign n2944 = ~x843 & ~x844 ;
  assign n2941 = x845 & ~n1845 ;
  assign n2940 = x841 & ~n1843 ;
  assign n2942 = n2941 ^ n2940 ;
  assign n2938 = n1845 ^ n1843 ;
  assign n2939 = n1844 & ~n2938 ;
  assign n2943 = n2942 ^ n2939 ;
  assign n2945 = n2944 ^ n2943 ;
  assign n2954 = n2953 ^ n2945 ;
  assign n2958 = n2957 ^ n2954 ;
  assign n3043 = n3042 ^ n2958 ;
  assign n1826 = x818 ^ x817 ;
  assign n1825 = x822 ^ x821 ;
  assign n1827 = n1826 ^ n1825 ;
  assign n1824 = x820 ^ x819 ;
  assign n1828 = n1827 ^ n1824 ;
  assign n1821 = x812 ^ x811 ;
  assign n1820 = x816 ^ x815 ;
  assign n1822 = n1821 ^ n1820 ;
  assign n1819 = x814 ^ x813 ;
  assign n1823 = n1822 ^ n1819 ;
  assign n1829 = n1828 ^ n1823 ;
  assign n1815 = x802 ^ x801 ;
  assign n1814 = x800 ^ x799 ;
  assign n1816 = n1815 ^ n1814 ;
  assign n1813 = x804 ^ x803 ;
  assign n1817 = n1816 ^ n1813 ;
  assign n1810 = x806 ^ x805 ;
  assign n1809 = x808 ^ x807 ;
  assign n1811 = n1810 ^ n1809 ;
  assign n1808 = x810 ^ x809 ;
  assign n1812 = n1811 ^ n1808 ;
  assign n1818 = n1817 ^ n1812 ;
  assign n1830 = n1829 ^ n1818 ;
  assign n1853 = n1852 ^ n1841 ;
  assign n2937 = n1830 & n1853 ;
  assign n3044 = n3043 ^ n2937 ;
  assign n2896 = x809 ^ x808 ;
  assign n2900 = ~n1808 & ~n2896 ;
  assign n2895 = x807 ^ x806 ;
  assign n2897 = n2896 ^ x807 ;
  assign n2898 = n2897 ^ x810 ;
  assign n2899 = ~n2895 & n2898 ;
  assign n2901 = n2900 ^ n2899 ;
  assign n2902 = ~x805 & n2901 ;
  assign n2903 = ~n1809 & ~n2895 ;
  assign n2904 = x810 ^ x805 ;
  assign n2907 = ~x808 & ~n2904 ;
  assign n2908 = n2907 ^ x805 ;
  assign n2909 = n2903 & n2908 ;
  assign n2910 = ~x809 & n2909 ;
  assign n2911 = ~x807 & ~x808 ;
  assign n2914 = n2911 ^ n1809 ;
  assign n2915 = x805 & x806 ;
  assign n2916 = x810 & n2915 ;
  assign n2917 = ~n2914 & n2916 ;
  assign n2918 = n2917 ^ n2915 ;
  assign n2912 = ~x809 & ~x810 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2919 = n2918 ^ n2913 ;
  assign n2920 = n2912 ^ n1808 ;
  assign n2925 = n2914 & n2920 ;
  assign n2926 = n2925 ^ n2913 ;
  assign n2927 = n2919 & n2926 ;
  assign n2928 = n2927 ^ n2918 ;
  assign n2929 = ~n1810 & n2928 ;
  assign n2930 = n2927 & n2929 ;
  assign n2931 = n2930 ^ n2928 ;
  assign n2932 = ~n2910 & ~n2931 ;
  assign n2933 = ~n2902 & n2932 ;
  assign n2885 = n1815 ^ n1813 ;
  assign n2876 = x803 & x804 ;
  assign n2875 = x801 & x802 ;
  assign n2877 = n2876 ^ n2875 ;
  assign n2886 = n2885 ^ n2877 ;
  assign n2887 = n2886 ^ x800 ;
  assign n2893 = n1814 & n2887 ;
  assign n2879 = n2876 ^ n1813 ;
  assign n2880 = n2875 ^ n1815 ;
  assign n2881 = n2879 & n2880 ;
  assign n2878 = n2875 ^ n1814 ;
  assign n2882 = n2881 ^ n2878 ;
  assign n2883 = ~n2877 & ~n2882 ;
  assign n2884 = n2883 ^ x799 ;
  assign n2894 = n2893 ^ n2884 ;
  assign n2934 = n2933 ^ n2894 ;
  assign n2873 = n1818 & n1829 ;
  assign n2871 = n1812 & n1817 ;
  assign n2870 = n1823 & n1828 ;
  assign n2872 = n2871 ^ n2870 ;
  assign n2874 = n2873 ^ n2872 ;
  assign n2935 = n2934 ^ n2874 ;
  assign n2808 = ~x813 & ~x814 ;
  assign n2820 = x815 ^ x812 ;
  assign n2823 = n1820 & n2820 ;
  assign n2824 = n2823 ^ x815 ;
  assign n2825 = n2808 & ~n2824 ;
  assign n2809 = n2808 ^ n1819 ;
  assign n2806 = ~x815 & ~x816 ;
  assign n2807 = n2806 ^ n1820 ;
  assign n2810 = n2809 ^ n2807 ;
  assign n2811 = ~n2806 & ~n2808 ;
  assign n2816 = x812 & n2811 ;
  assign n2817 = n2816 ^ n2807 ;
  assign n2818 = n2810 & n2817 ;
  assign n2819 = n2818 ^ n2809 ;
  assign n2826 = n2825 ^ n2819 ;
  assign n2827 = ~x811 & ~n2826 ;
  assign n2829 = x816 ^ x812 ;
  assign n2828 = x816 ^ x814 ;
  assign n2830 = n2829 ^ n2828 ;
  assign n2831 = n2830 ^ x816 ;
  assign n2833 = x812 & n2831 ;
  assign n2834 = n2833 ^ x816 ;
  assign n2837 = x816 ^ x813 ;
  assign n2838 = n2837 ^ n2829 ;
  assign n2839 = n2838 ^ n1821 ;
  assign n2840 = n2830 ^ n1821 ;
  assign n2841 = n2840 ^ n2829 ;
  assign n2842 = n2841 ^ x816 ;
  assign n2843 = ~n2839 & n2842 ;
  assign n2846 = n2843 ^ x814 ;
  assign n2847 = ~n2834 & ~n2846 ;
  assign n2850 = ~x815 & n2847 ;
  assign n2851 = x811 & x812 ;
  assign n2852 = x816 & ~n2809 ;
  assign n2853 = n2851 & n2852 ;
  assign n2854 = n2853 ^ n2851 ;
  assign n2855 = n2854 ^ n2811 ;
  assign n2860 = n2807 & n2809 ;
  assign n2861 = n2860 ^ n2854 ;
  assign n2862 = n2855 & ~n2861 ;
  assign n2863 = n2862 ^ n2854 ;
  assign n2864 = ~n1821 & n2863 ;
  assign n2865 = n2862 & n2864 ;
  assign n2866 = n2865 ^ n2863 ;
  assign n2867 = ~n2850 & ~n2866 ;
  assign n2868 = ~n2827 & n2867 ;
  assign n2745 = ~x819 & ~x820 ;
  assign n2757 = x821 ^ x818 ;
  assign n2760 = n1825 & n2757 ;
  assign n2761 = n2760 ^ x821 ;
  assign n2762 = n2745 & ~n2761 ;
  assign n2746 = n2745 ^ n1824 ;
  assign n2743 = ~x821 & ~x822 ;
  assign n2744 = n2743 ^ n1825 ;
  assign n2747 = n2746 ^ n2744 ;
  assign n2748 = ~n2743 & ~n2745 ;
  assign n2753 = x818 & n2748 ;
  assign n2754 = n2753 ^ n2744 ;
  assign n2755 = n2747 & n2754 ;
  assign n2756 = n2755 ^ n2746 ;
  assign n2763 = n2762 ^ n2756 ;
  assign n2764 = ~x817 & ~n2763 ;
  assign n2766 = x822 ^ x818 ;
  assign n2765 = x822 ^ x820 ;
  assign n2767 = n2766 ^ n2765 ;
  assign n2768 = n2767 ^ x822 ;
  assign n2770 = x818 & n2768 ;
  assign n2771 = n2770 ^ x822 ;
  assign n2774 = x822 ^ x819 ;
  assign n2775 = n2774 ^ n2766 ;
  assign n2776 = n2775 ^ n1826 ;
  assign n2777 = n2767 ^ n1826 ;
  assign n2778 = n2777 ^ n2766 ;
  assign n2779 = n2778 ^ x822 ;
  assign n2780 = ~n2776 & n2779 ;
  assign n2783 = n2780 ^ x820 ;
  assign n2784 = ~n2771 & ~n2783 ;
  assign n2787 = ~x821 & n2784 ;
  assign n2788 = x817 & x818 ;
  assign n2789 = x822 & ~n2746 ;
  assign n2790 = n2788 & n2789 ;
  assign n2791 = n2790 ^ n2788 ;
  assign n2792 = n2791 ^ n2748 ;
  assign n2797 = n2744 & n2746 ;
  assign n2798 = n2797 ^ n2791 ;
  assign n2799 = n2792 & ~n2798 ;
  assign n2800 = n2799 ^ n2791 ;
  assign n2801 = ~n1826 & n2800 ;
  assign n2802 = n2799 & n2801 ;
  assign n2803 = n2802 ^ n2800 ;
  assign n2804 = ~n2787 & ~n2803 ;
  assign n2805 = ~n2764 & n2804 ;
  assign n2869 = n2868 ^ n2805 ;
  assign n2936 = n2935 ^ n2869 ;
  assign n3045 = n3044 ^ n2936 ;
  assign n2742 = n2741 ^ n2594 ;
  assign n3046 = n3045 ^ n2742 ;
  assign n1854 = n1853 ^ n1830 ;
  assign n1901 = n1900 ^ n1877 ;
  assign n2003 = n1854 & n1901 ;
  assign n10508 = n3045 ^ n2003 ;
  assign n10509 = ~n3046 & n10508 ;
  assign n10510 = n10509 ^ n3045 ;
  assign n10650 = n10649 ^ n10510 ;
  assign n10490 = n2756 & ~n2803 ;
  assign n10489 = n2819 & ~n2866 ;
  assign n10491 = n10490 ^ n10489 ;
  assign n10486 = n2870 ^ n2805 ;
  assign n10487 = ~n2869 & n10486 ;
  assign n10488 = n10487 ^ n2870 ;
  assign n10492 = n10491 ^ n10488 ;
  assign n10460 = n2876 ^ x800 ;
  assign n10450 = n2876 ^ x799 ;
  assign n10455 = n10450 ^ n2877 ;
  assign n10461 = n10460 ^ n10455 ;
  assign n10452 = n2881 ^ n2876 ;
  assign n10453 = n10452 ^ n10450 ;
  assign n10462 = n10461 ^ n10453 ;
  assign n10463 = n10462 ^ n2877 ;
  assign n10465 = n10461 & n10463 ;
  assign n10459 = ~x799 & n2876 ;
  assign n10466 = n10465 ^ n10459 ;
  assign n10457 = n10453 ^ n2877 ;
  assign n10467 = n10466 ^ n10457 ;
  assign n10468 = n10465 ^ n10455 ;
  assign n10469 = n10468 ^ n10457 ;
  assign n10470 = n10467 & n10469 ;
  assign n10471 = ~n2877 & n10470 ;
  assign n10472 = n10471 ^ n10465 ;
  assign n10473 = n10472 ^ n10463 ;
  assign n10476 = n10473 ^ n2876 ;
  assign n10477 = n10476 ^ n10460 ;
  assign n11343 = n10492 ^ n10477 ;
  assign n10478 = n2920 ^ n2914 ;
  assign n10479 = x806 & n2913 ;
  assign n10480 = n10479 ^ n2914 ;
  assign n10481 = n10478 & ~n10480 ;
  assign n10482 = n10481 ^ n2914 ;
  assign n10483 = ~n2931 & ~n10482 ;
  assign n10484 = n10483 ^ n2931 ;
  assign n11344 = n11343 ^ n10484 ;
  assign n10502 = ~n2894 & n2933 ;
  assign n10496 = n2873 ^ n2871 ;
  assign n10503 = n2936 & n10496 ;
  assign n10504 = n10502 & n10503 ;
  assign n10494 = n2870 ^ n2869 ;
  assign n10495 = ~n2936 & ~n10494 ;
  assign n10497 = n10496 ^ n10495 ;
  assign n10498 = n10496 ^ n2894 ;
  assign n10499 = n2934 & n10498 ;
  assign n10500 = ~n10497 & n10499 ;
  assign n10501 = n10500 ^ n10495 ;
  assign n10505 = n10504 ^ n10501 ;
  assign n11346 = n11344 ^ n10505 ;
  assign n10445 = n3043 ^ n2936 ;
  assign n10446 = ~n3044 & n10445 ;
  assign n10439 = ~n2968 & ~n2979 ;
  assign n10438 = ~n3015 & n3039 ;
  assign n10440 = n10439 ^ n10438 ;
  assign n10435 = n2993 ^ n2992 ;
  assign n10436 = n3041 & ~n10435 ;
  assign n10437 = n10436 ^ n2993 ;
  assign n10441 = n10440 ^ n10437 ;
  assign n10401 = n2952 ^ n1847 ;
  assign n10402 = n10401 ^ n2949 ;
  assign n10403 = n2949 ^ n1850 ;
  assign n10404 = ~n2952 & n10403 ;
  assign n10409 = x836 & n10404 ;
  assign n10410 = n10409 ^ n10401 ;
  assign n10411 = ~n10402 & n10410 ;
  assign n10412 = n10411 ^ n2949 ;
  assign n10416 = ~n2949 & n10401 ;
  assign n10413 = x840 & n2948 ;
  assign n10414 = ~n10401 & n10413 ;
  assign n10415 = n10414 ^ n2948 ;
  assign n10417 = n10416 ^ n10415 ;
  assign n10418 = n10416 ^ n10404 ;
  assign n10419 = ~n10417 & n10418 ;
  assign n10427 = ~n1848 & n10419 ;
  assign n10428 = ~n10416 & n10427 ;
  assign n10429 = n10428 ^ n10416 ;
  assign n10420 = n10419 ^ n10415 ;
  assign n10421 = n10420 ^ n10416 ;
  assign n10430 = n10429 ^ n10421 ;
  assign n10431 = ~n10412 & ~n10430 ;
  assign n10370 = n2944 ^ n1842 ;
  assign n10371 = n10370 ^ n2941 ;
  assign n10372 = n2941 ^ n1845 ;
  assign n10373 = ~n2944 & n10372 ;
  assign n10378 = x842 & n10373 ;
  assign n10379 = n10378 ^ n10370 ;
  assign n10380 = ~n10371 & n10379 ;
  assign n10381 = n10380 ^ n2941 ;
  assign n10385 = ~n2941 & n10370 ;
  assign n10382 = x846 & n2940 ;
  assign n10383 = ~n10370 & n10382 ;
  assign n10384 = n10383 ^ n2940 ;
  assign n10386 = n10385 ^ n10384 ;
  assign n10387 = n10385 ^ n10373 ;
  assign n10388 = ~n10386 & n10387 ;
  assign n10396 = ~n1843 & n10388 ;
  assign n10397 = ~n10385 & n10396 ;
  assign n10398 = n10397 ^ n10385 ;
  assign n10389 = n10388 ^ n10384 ;
  assign n10390 = n10389 ^ n10385 ;
  assign n10399 = n10398 ^ n10390 ;
  assign n10400 = ~n10381 & ~n10399 ;
  assign n10432 = n10431 ^ n10400 ;
  assign n10367 = n2955 ^ n2945 ;
  assign n10368 = ~n2954 & ~n10367 ;
  assign n10369 = n10368 ^ n2955 ;
  assign n10433 = n10432 ^ n10369 ;
  assign n10364 = n3042 ^ n2956 ;
  assign n10365 = ~n2958 & ~n10364 ;
  assign n10366 = n10365 ^ n3042 ;
  assign n10434 = n10433 ^ n10366 ;
  assign n10442 = n10441 ^ n10434 ;
  assign n10443 = n10442 ^ n3043 ;
  assign n10447 = n10446 ^ n10443 ;
  assign n10507 = n11346 ^ n10447 ;
  assign n10651 = n10650 ^ n10507 ;
  assign n10992 = n10991 ^ n10651 ;
  assign n2487 = n10654 ^ n2486 ;
  assign n1902 = n1901 ^ n1854 ;
  assign n1997 = n1996 ^ n1949 ;
  assign n2001 = ~n1902 & ~n1997 ;
  assign n1998 = n1997 ^ n1902 ;
  assign n2002 = n2001 ^ n1998 ;
  assign n10355 = n2487 ^ n2002 ;
  assign n10360 = n2002 & ~n2003 ;
  assign n10361 = n10360 ^ n3046 ;
  assign n10362 = n10355 & ~n10361 ;
  assign n10363 = n10362 ^ n2487 ;
  assign n10993 = n10992 ^ n10363 ;
  assign n1753 = x472 ^ x471 ;
  assign n1752 = x474 ^ x473 ;
  assign n1754 = n1753 ^ n1752 ;
  assign n1751 = x470 ^ x469 ;
  assign n1755 = n1754 ^ n1751 ;
  assign n1749 = x466 ^ x465 ;
  assign n1747 = x468 ^ x467 ;
  assign n1746 = x464 ^ x463 ;
  assign n1748 = n1747 ^ n1746 ;
  assign n1750 = n1749 ^ n1748 ;
  assign n1756 = n1755 ^ n1750 ;
  assign n1743 = x480 ^ x479 ;
  assign n1741 = x476 ^ x475 ;
  assign n1740 = x478 ^ x477 ;
  assign n1742 = n1741 ^ n1740 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1738 = x486 ^ x485 ;
  assign n1736 = x484 ^ x483 ;
  assign n1735 = x482 ^ x481 ;
  assign n1737 = n1736 ^ n1735 ;
  assign n1739 = n1738 ^ n1737 ;
  assign n1745 = n1744 ^ n1739 ;
  assign n1757 = n1756 ^ n1745 ;
  assign n1731 = x488 ^ x487 ;
  assign n1729 = x490 ^ x489 ;
  assign n1728 = x492 ^ x491 ;
  assign n1730 = n1729 ^ n1728 ;
  assign n1732 = n1731 ^ n1730 ;
  assign n1726 = x498 ^ x497 ;
  assign n1724 = x496 ^ x495 ;
  assign n1723 = x494 ^ x493 ;
  assign n1725 = n1724 ^ n1723 ;
  assign n1727 = n1726 ^ n1725 ;
  assign n1733 = n1732 ^ n1727 ;
  assign n1720 = x504 ^ x503 ;
  assign n1718 = x502 ^ x501 ;
  assign n1717 = x500 ^ x499 ;
  assign n1719 = n1718 ^ n1717 ;
  assign n1721 = n1720 ^ n1719 ;
  assign n1715 = x510 ^ x509 ;
  assign n1713 = x506 ^ x505 ;
  assign n1712 = x508 ^ x507 ;
  assign n1714 = n1713 ^ n1712 ;
  assign n1716 = n1715 ^ n1714 ;
  assign n1722 = n1721 ^ n1716 ;
  assign n1734 = n1733 ^ n1722 ;
  assign n1758 = n1757 ^ n1734 ;
  assign n1800 = x546 ^ x545 ;
  assign n1799 = x544 ^ x543 ;
  assign n1801 = n1800 ^ n1799 ;
  assign n1798 = x542 ^ x541 ;
  assign n1802 = n1801 ^ n1798 ;
  assign n1796 = x540 ^ x539 ;
  assign n1794 = x536 ^ x535 ;
  assign n1793 = x538 ^ x537 ;
  assign n1795 = n1794 ^ n1793 ;
  assign n1797 = n1796 ^ n1795 ;
  assign n1803 = n1802 ^ n1797 ;
  assign n1790 = x548 ^ x547 ;
  assign n1788 = x552 ^ x551 ;
  assign n1787 = x550 ^ x549 ;
  assign n1789 = n1788 ^ n1787 ;
  assign n1791 = n1790 ^ n1789 ;
  assign n1785 = x558 ^ x557 ;
  assign n1783 = x556 ^ x555 ;
  assign n1782 = x554 ^ x553 ;
  assign n1784 = n1783 ^ n1782 ;
  assign n1786 = n1785 ^ n1784 ;
  assign n1792 = n1791 ^ n1786 ;
  assign n1804 = n1803 ^ n1792 ;
  assign n1778 = x534 ^ x533 ;
  assign n1776 = x532 ^ x531 ;
  assign n1775 = x530 ^ x529 ;
  assign n1777 = n1776 ^ n1775 ;
  assign n1779 = n1778 ^ n1777 ;
  assign n1773 = x528 ^ x527 ;
  assign n1771 = x526 ^ x525 ;
  assign n1770 = x524 ^ x523 ;
  assign n1772 = n1771 ^ n1770 ;
  assign n1774 = n1773 ^ n1772 ;
  assign n1780 = n1779 ^ n1774 ;
  assign n1767 = x516 ^ x515 ;
  assign n1765 = x512 ^ x511 ;
  assign n1764 = x514 ^ x513 ;
  assign n1766 = n1765 ^ n1764 ;
  assign n1768 = n1767 ^ n1766 ;
  assign n1762 = x522 ^ x521 ;
  assign n1760 = x520 ^ x519 ;
  assign n1759 = x518 ^ x517 ;
  assign n1761 = n1760 ^ n1759 ;
  assign n1763 = n1762 ^ n1761 ;
  assign n1769 = n1768 ^ n1763 ;
  assign n1781 = n1780 ^ n1769 ;
  assign n1805 = n1804 ^ n1781 ;
  assign n3673 = n1758 & n1805 ;
  assign n3671 = n1734 & n1757 ;
  assign n9747 = n3673 ^ n3671 ;
  assign n3776 = x501 & x502 ;
  assign n3778 = n3776 ^ n1718 ;
  assign n3775 = x503 & x504 ;
  assign n3779 = n3775 ^ n1720 ;
  assign n3780 = n3778 & n3779 ;
  assign n3789 = n3780 ^ x500 ;
  assign n3777 = n3776 ^ n3775 ;
  assign n3781 = n3780 ^ n3776 ;
  assign n3782 = n3781 ^ n1717 ;
  assign n3783 = ~n3777 & ~n3782 ;
  assign n3784 = n3783 ^ n3780 ;
  assign n3785 = n3777 ^ n1718 ;
  assign n3786 = n3785 ^ n1720 ;
  assign n3787 = n3786 ^ n3783 ;
  assign n3788 = ~n3784 & ~n3787 ;
  assign n3790 = n3789 ^ n3788 ;
  assign n3794 = n1717 & ~n3790 ;
  assign n3792 = n3783 ^ x499 ;
  assign n3795 = n3794 ^ n3792 ;
  assign n3733 = x509 & x510 ;
  assign n3741 = n3733 ^ n1715 ;
  assign n3742 = ~x508 & ~n3741 ;
  assign n3734 = x508 & n3733 ;
  assign n3740 = n3734 ^ n1715 ;
  assign n3743 = n3742 ^ n3740 ;
  assign n3744 = n3743 ^ x508 ;
  assign n3748 = n3742 ^ x507 ;
  assign n3747 = ~x507 & n3742 ;
  assign n3749 = n3748 ^ n3747 ;
  assign n3752 = n3744 & ~n3749 ;
  assign n3753 = ~x506 & n3752 ;
  assign n3754 = n3753 ^ x506 ;
  assign n3736 = n3734 ^ x507 ;
  assign n3735 = ~x507 & ~n3734 ;
  assign n3737 = n3736 ^ n3735 ;
  assign n3738 = n3737 ^ x506 ;
  assign n3755 = n3754 ^ n3738 ;
  assign n3756 = ~x505 & ~n3755 ;
  assign n3757 = x505 & x506 ;
  assign n3772 = n3747 & ~n3757 ;
  assign n3758 = n3737 & n3757 ;
  assign n3759 = n3758 ^ n3744 ;
  assign n3762 = n1713 & ~n3735 ;
  assign n3763 = n3762 ^ n3749 ;
  assign n3764 = ~n3758 & ~n3763 ;
  assign n3765 = n3764 ^ n3749 ;
  assign n3766 = ~n3759 & ~n3765 ;
  assign n3767 = n3766 ^ n3758 ;
  assign n3773 = n3772 ^ n3767 ;
  assign n3774 = ~n3756 & ~n3773 ;
  assign n3796 = n3795 ^ n3774 ;
  assign n3730 = n1716 & n1721 ;
  assign n10121 = n3796 ^ n3730 ;
  assign n3727 = n1727 ^ n1722 ;
  assign n3728 = n1733 & ~n3727 ;
  assign n3729 = n3728 ^ n1732 ;
  assign n10123 = n10121 ^ n3729 ;
  assign n3675 = ~x489 & ~x490 ;
  assign n3676 = x491 & x492 ;
  assign n3677 = n3675 & ~n3676 ;
  assign n3678 = n3675 ^ n1729 ;
  assign n3679 = n3676 ^ n1728 ;
  assign n3680 = n3678 & ~n3679 ;
  assign n3681 = ~n3677 & ~n3680 ;
  assign n3684 = n3676 & ~n3678 ;
  assign n3682 = n3680 ^ n3677 ;
  assign n3683 = n3682 ^ n3681 ;
  assign n3685 = n3684 ^ n3683 ;
  assign n3686 = n3685 ^ x488 ;
  assign n3687 = ~n1731 & n3686 ;
  assign n3688 = n3687 ^ n3685 ;
  assign n3723 = n3687 & ~n3688 ;
  assign n3724 = n3681 & n3723 ;
  assign n3725 = n3724 ^ ~n3688 ;
  assign n3715 = x488 & ~n3684 ;
  assign n3716 = n3715 ^ n1730 ;
  assign n3717 = ~n1731 & n3716 ;
  assign n3718 = n3717 ^ n1730 ;
  assign n3719 = n3681 & n3718 ;
  assign n3689 = x497 & x498 ;
  assign n3690 = n3689 ^ n1726 ;
  assign n3692 = x495 & x496 ;
  assign n3693 = n3692 ^ n1724 ;
  assign n3697 = n3690 & n3693 ;
  assign n3698 = n3697 ^ n1723 ;
  assign n3700 = n3692 ^ n3689 ;
  assign n3696 = ~n3689 & ~n3692 ;
  assign n3701 = n3700 ^ n3696 ;
  assign n3702 = x493 & x494 ;
  assign n3703 = n3701 & n3702 ;
  assign n3704 = n3703 ^ n3696 ;
  assign n3705 = n3703 ^ n3697 ;
  assign n3706 = ~n3704 & n3705 ;
  assign n3707 = ~n3698 & n3706 ;
  assign n3708 = n3707 ^ n3703 ;
  assign n3710 = n3708 ^ x493 ;
  assign n3709 = n3701 & ~n3708 ;
  assign n3711 = n3710 ^ n3709 ;
  assign n3699 = n3696 & ~n3698 ;
  assign n3712 = n3711 ^ n3699 ;
  assign n3691 = n3690 ^ x494 ;
  assign n3694 = n3693 ^ n3691 ;
  assign n3695 = n1723 & n3694 ;
  assign n3713 = n3712 ^ n3695 ;
  assign n3720 = n3719 ^ n3713 ;
  assign n3726 = n3725 ^ n3720 ;
  assign n10124 = n10123 ^ n3726 ;
  assign n3891 = ~x473 & ~x474 ;
  assign n3892 = n3891 ^ n1752 ;
  assign n3895 = n3892 ^ x472 ;
  assign n3897 = n1753 & n3895 ;
  assign n3893 = x471 & x472 ;
  assign n3894 = ~n3892 & n3893 ;
  assign n3896 = n3895 ^ n3894 ;
  assign n3898 = n3897 ^ n3896 ;
  assign n3899 = x469 & ~n3898 ;
  assign n3900 = n3897 ^ x471 ;
  assign n3902 = ~n3891 & n3900 ;
  assign n3901 = n3900 ^ n3891 ;
  assign n3903 = n3902 ^ n3901 ;
  assign n3904 = n3903 ^ n3894 ;
  assign n3905 = n3899 & ~n3904 ;
  assign n3906 = n3905 ^ n3902 ;
  assign n3907 = x469 & ~x470 ;
  assign n3908 = n3906 & n3907 ;
  assign n3909 = n3908 ^ n3905 ;
  assign n3910 = ~x470 & n3903 ;
  assign n3911 = n3910 ^ x469 ;
  assign n3912 = x470 & ~n3891 ;
  assign n3921 = n3898 & ~n3912 ;
  assign n3913 = ~n3894 & n3900 ;
  assign n3914 = ~n3912 & n3913 ;
  assign n3915 = n3914 ^ n3900 ;
  assign n3916 = n3915 ^ n3910 ;
  assign n3922 = n3921 ^ n3916 ;
  assign n3923 = ~n3911 & ~n3922 ;
  assign n3924 = n3923 ^ x469 ;
  assign n3925 = ~n3909 & n3924 ;
  assign n3871 = x467 & x468 ;
  assign n3873 = n3871 ^ n1747 ;
  assign n3870 = x465 & x466 ;
  assign n3874 = n3870 ^ n1749 ;
  assign n3875 = n3873 & n3874 ;
  assign n3884 = n3875 ^ x464 ;
  assign n3872 = n3871 ^ n3870 ;
  assign n3876 = n3875 ^ n3871 ;
  assign n3877 = n3876 ^ n1746 ;
  assign n3878 = ~n3872 & ~n3877 ;
  assign n3879 = n3878 ^ n3875 ;
  assign n3880 = n1749 ^ n1747 ;
  assign n3881 = n3880 ^ n3872 ;
  assign n3882 = n3881 ^ n3878 ;
  assign n3883 = ~n3879 & ~n3882 ;
  assign n3885 = n3884 ^ n3883 ;
  assign n3889 = n1746 & ~n3885 ;
  assign n3887 = n3878 ^ x463 ;
  assign n3890 = n3889 ^ n3887 ;
  assign n3926 = n3925 ^ n3890 ;
  assign n3865 = n1750 & n1755 ;
  assign n9985 = n3926 ^ n3865 ;
  assign n3867 = n1739 & n1744 ;
  assign n9987 = n9985 ^ n3867 ;
  assign n3864 = n1745 & n1756 ;
  assign n9988 = n9987 ^ n3864 ;
  assign n3799 = x477 & x478 ;
  assign n3798 = x479 & x480 ;
  assign n3800 = n3799 ^ n3798 ;
  assign n3804 = n3798 ^ n1743 ;
  assign n3805 = n3799 ^ n1740 ;
  assign n3806 = n3804 & n3805 ;
  assign n3808 = n3806 ^ n3798 ;
  assign n3809 = n3808 ^ n1741 ;
  assign n3810 = ~n3800 & ~n3809 ;
  assign n3801 = n3800 ^ n1743 ;
  assign n3802 = n3801 ^ n1740 ;
  assign n3803 = n3802 ^ x476 ;
  assign n3807 = n3806 ^ n3803 ;
  assign n3811 = n3810 ^ n3807 ;
  assign n3812 = n3811 ^ n3803 ;
  assign n3814 = n3806 ^ x476 ;
  assign n3815 = n3814 ^ n3803 ;
  assign n3816 = n3812 & ~n3815 ;
  assign n3817 = n3816 ^ n3803 ;
  assign n3862 = n1741 & n3817 ;
  assign n3859 = n3810 ^ x475 ;
  assign n3820 = x485 ^ x484 ;
  assign n3824 = ~n1738 & ~n3820 ;
  assign n3819 = x483 ^ x482 ;
  assign n3821 = n3820 ^ x483 ;
  assign n3822 = n3821 ^ x486 ;
  assign n3823 = ~n3819 & n3822 ;
  assign n3825 = n3824 ^ n3823 ;
  assign n3826 = ~x481 & n3825 ;
  assign n3827 = ~n1736 & ~n3819 ;
  assign n3828 = x486 ^ x481 ;
  assign n3831 = ~x484 & ~n3828 ;
  assign n3832 = n3831 ^ x481 ;
  assign n3833 = n3827 & n3832 ;
  assign n3834 = ~x485 & n3833 ;
  assign n3835 = ~x483 & ~x484 ;
  assign n3838 = n3835 ^ n1736 ;
  assign n3839 = x481 & x482 ;
  assign n3840 = x486 & n3839 ;
  assign n3841 = ~n3838 & n3840 ;
  assign n3842 = n3841 ^ n3839 ;
  assign n3836 = ~x485 & ~x486 ;
  assign n3837 = ~n3835 & ~n3836 ;
  assign n3843 = n3842 ^ n3837 ;
  assign n3844 = n3836 ^ n1738 ;
  assign n3849 = n3838 & n3844 ;
  assign n3850 = n3849 ^ n3837 ;
  assign n3851 = n3843 & n3850 ;
  assign n3852 = n3851 ^ n3842 ;
  assign n3853 = ~n1735 & n3852 ;
  assign n3854 = n3851 & n3853 ;
  assign n3855 = n3854 ^ n3852 ;
  assign n3856 = ~n3834 & ~n3855 ;
  assign n3857 = ~n3826 & n3856 ;
  assign n3860 = n3859 ^ n3857 ;
  assign n3863 = n3862 ^ n3860 ;
  assign n9989 = n9988 ^ n3863 ;
  assign n3928 = n10124 ^ n9989 ;
  assign n9748 = n9747 ^ n3928 ;
  assign n3670 = n1781 & n1804 ;
  assign n9749 = n9748 ^ n3670 ;
  assign n4006 = x533 & x534 ;
  assign n4005 = x531 & x532 ;
  assign n4007 = n4006 ^ n4005 ;
  assign n4008 = n4005 ^ n1776 ;
  assign n4009 = n4006 ^ n1778 ;
  assign n4010 = n4008 & n4009 ;
  assign n4011 = n4010 ^ n4005 ;
  assign n4012 = ~n4007 & ~n4011 ;
  assign n3984 = n1776 ^ x530 ;
  assign n3985 = n3984 ^ n1778 ;
  assign n3991 = x527 & x528 ;
  assign n3990 = x525 & x526 ;
  assign n3992 = n3991 ^ n3990 ;
  assign n3993 = n3991 ^ n1773 ;
  assign n3994 = n3990 ^ n1771 ;
  assign n3995 = n3993 & n3994 ;
  assign n3996 = n3995 ^ n3991 ;
  assign n3997 = ~n3992 & ~n3996 ;
  assign n3986 = n1773 ^ x524 ;
  assign n3987 = n3986 ^ n1771 ;
  assign n3988 = n1770 & ~n3987 ;
  assign n3989 = n3988 ^ x523 ;
  assign n3998 = n3997 ^ n3989 ;
  assign n3999 = n3998 ^ x529 ;
  assign n4000 = n3999 ^ n1776 ;
  assign n4001 = n4000 ^ n1778 ;
  assign n4002 = n4001 ^ n3998 ;
  assign n4003 = ~n3985 & n4002 ;
  assign n4004 = n4003 ^ n3999 ;
  assign n4013 = n4012 ^ n4004 ;
  assign n3979 = n1774 & n1779 ;
  assign n9764 = n4013 ^ n3979 ;
  assign n3981 = n1763 & n1768 ;
  assign n9766 = n9764 ^ n3981 ;
  assign n3978 = n1769 & n1780 ;
  assign n9767 = n9766 ^ n3978 ;
  assign n3931 = x513 & x514 ;
  assign n3930 = x515 & x516 ;
  assign n3932 = n3931 ^ n3930 ;
  assign n3936 = n3930 ^ n1767 ;
  assign n3937 = n3931 ^ n1764 ;
  assign n3938 = n3936 & n3937 ;
  assign n3940 = n3938 ^ n3930 ;
  assign n3941 = n3940 ^ n1765 ;
  assign n3942 = ~n3932 & ~n3941 ;
  assign n3933 = n3932 ^ n1767 ;
  assign n3934 = n3933 ^ n1764 ;
  assign n3935 = n3934 ^ x512 ;
  assign n3939 = n3938 ^ n3935 ;
  assign n3943 = n3942 ^ n3939 ;
  assign n3944 = n3943 ^ n3935 ;
  assign n3946 = n3938 ^ x512 ;
  assign n3947 = n3946 ^ n3935 ;
  assign n3948 = n3944 & ~n3947 ;
  assign n3949 = n3948 ^ n3935 ;
  assign n3976 = n1765 & n3949 ;
  assign n3973 = n3942 ^ x511 ;
  assign n3952 = x521 & x522 ;
  assign n3954 = n3952 ^ n1762 ;
  assign n3951 = x519 & x520 ;
  assign n3955 = n3951 ^ n1760 ;
  assign n3956 = n3954 & n3955 ;
  assign n3965 = n3956 ^ x518 ;
  assign n3953 = n3952 ^ n3951 ;
  assign n3957 = n3956 ^ n3952 ;
  assign n3958 = n3957 ^ n1759 ;
  assign n3959 = ~n3953 & ~n3958 ;
  assign n3960 = n3959 ^ n3956 ;
  assign n3961 = n3953 ^ n1760 ;
  assign n3962 = n3961 ^ n1762 ;
  assign n3963 = n3962 ^ n3959 ;
  assign n3964 = ~n3960 & ~n3963 ;
  assign n3966 = n3965 ^ n3964 ;
  assign n3970 = n1759 & ~n3966 ;
  assign n3968 = n3959 ^ x517 ;
  assign n3971 = n3970 ^ n3968 ;
  assign n3974 = n3973 ^ n3971 ;
  assign n3977 = n3976 ^ n3974 ;
  assign n9768 = n9767 ^ n3977 ;
  assign n4110 = n1802 ^ n1786 ;
  assign n4111 = ~n1803 & ~n4110 ;
  assign n4112 = n4110 ^ n1791 ;
  assign n4113 = n4111 & n4112 ;
  assign n4114 = n4113 ^ n1791 ;
  assign n4117 = n1786 & n1791 ;
  assign n4118 = n4117 ^ n4111 ;
  assign n4115 = n1803 ^ n1786 ;
  assign n4116 = ~n4114 & n4115 ;
  assign n4119 = n4118 ^ n4116 ;
  assign n4120 = ~n4114 & n4119 ;
  assign n4084 = ~x555 & ~x556 ;
  assign n4085 = n4084 ^ n1783 ;
  assign n4081 = x557 & x558 ;
  assign n4086 = n4081 ^ n1785 ;
  assign n4087 = n4085 & ~n4086 ;
  assign n4082 = n4081 ^ x556 ;
  assign n4083 = ~n1783 & ~n4082 ;
  assign n4088 = n4087 ^ n4083 ;
  assign n4104 = n4083 ^ n1782 ;
  assign n4105 = ~n4088 & ~n4104 ;
  assign n4107 = x554 & ~n1782 ;
  assign n4108 = ~n4105 & n4107 ;
  assign n4097 = x554 & ~n4088 ;
  assign n4098 = ~n4083 & n4097 ;
  assign n4099 = n4098 ^ n4083 ;
  assign n4089 = n1785 ^ n1783 ;
  assign n4090 = n4089 ^ n4088 ;
  assign n4091 = n4090 ^ n4083 ;
  assign n4100 = n4099 ^ n4091 ;
  assign n4101 = ~n1782 & n4100 ;
  assign n4102 = n4101 ^ n4090 ;
  assign n4076 = x547 & x548 ;
  assign n4074 = n1789 & n1790 ;
  assign n4063 = ~x551 & ~x552 ;
  assign n4064 = x549 & ~x550 ;
  assign n4065 = n4063 & n4064 ;
  assign n4066 = n4065 ^ x549 ;
  assign n4075 = n4074 ^ n4066 ;
  assign n4077 = n4076 ^ n4075 ;
  assign n4071 = x549 & x550 ;
  assign n4072 = n4063 ^ n1788 ;
  assign n4073 = n4071 & ~n4072 ;
  assign n4078 = n4077 ^ n4073 ;
  assign n4067 = x551 ^ x550 ;
  assign n4068 = ~n1788 & n4067 ;
  assign n4069 = n4068 ^ x550 ;
  assign n4070 = ~n4066 & n4069 ;
  assign n4079 = n4078 ^ n4070 ;
  assign n4080 = n4079 ^ n1782 ;
  assign n4103 = n4102 ^ n4080 ;
  assign n4106 = n4105 ^ n4103 ;
  assign n4109 = n4108 ^ n4106 ;
  assign n4121 = n4120 ^ n4109 ;
  assign n4017 = x537 & x538 ;
  assign n4015 = x539 & x540 ;
  assign n4020 = n4017 ^ n4015 ;
  assign n4016 = n4015 ^ n1796 ;
  assign n4018 = n4017 ^ n1793 ;
  assign n4019 = n4016 & n4018 ;
  assign n4025 = n4019 ^ n4015 ;
  assign n4026 = n4025 ^ n1794 ;
  assign n4027 = ~n4020 & ~n4026 ;
  assign n4021 = n1796 ^ n1793 ;
  assign n4022 = n4021 ^ n4020 ;
  assign n4023 = n4022 ^ x536 ;
  assign n4024 = n4023 ^ n4019 ;
  assign n4028 = n4027 ^ n4024 ;
  assign n4029 = n4028 ^ n4023 ;
  assign n4031 = n4019 ^ x536 ;
  assign n4032 = n4031 ^ n4023 ;
  assign n4033 = n4029 & ~n4032 ;
  assign n4034 = n4033 ^ n4023 ;
  assign n4061 = n1794 & n4034 ;
  assign n4058 = n4027 ^ x535 ;
  assign n4036 = ~x545 & ~x546 ;
  assign n4037 = x543 & x544 ;
  assign n4054 = n4036 & ~n4037 ;
  assign n4055 = ~x542 & n4054 ;
  assign n4048 = n1802 ^ x541 ;
  assign n4038 = n4036 ^ n1800 ;
  assign n4040 = n4038 ^ x544 ;
  assign n4039 = n4037 & ~n4038 ;
  assign n4049 = n4040 ^ n4039 ;
  assign n4041 = n1799 & n4040 ;
  assign n4050 = n4049 ^ n4041 ;
  assign n4051 = n4050 ^ n1802 ;
  assign n4052 = n4048 & ~n4051 ;
  assign n4042 = n4041 ^ x543 ;
  assign n4043 = ~n4039 & n4042 ;
  assign n4044 = x542 & n4043 ;
  assign n4045 = ~n4036 & n4044 ;
  assign n4046 = n4045 ^ n4043 ;
  assign n4047 = n4046 ^ n4042 ;
  assign n4053 = n4052 ^ n4047 ;
  assign n4056 = n4055 ^ n4053 ;
  assign n4059 = n4058 ^ n4056 ;
  assign n4062 = n4061 ^ n4059 ;
  assign n4122 = n4121 ^ n4062 ;
  assign n4123 = n9768 ^ n4122 ;
  assign n9750 = n9749 ^ n4123 ;
  assign n3611 = ~x651 & ~x652 ;
  assign n1693 = x652 ^ x651 ;
  assign n3620 = n3611 ^ n1693 ;
  assign n3618 = ~x653 & ~x654 ;
  assign n1695 = x654 ^ x653 ;
  assign n3619 = n3618 ^ n1695 ;
  assign n3621 = n3620 ^ n3619 ;
  assign n3622 = ~n3611 & ~n3618 ;
  assign n3627 = x650 & n3622 ;
  assign n3628 = n3627 ^ n3619 ;
  assign n3629 = n3621 & n3628 ;
  assign n3630 = n3629 ^ n3620 ;
  assign n3612 = x653 ^ x650 ;
  assign n3615 = n1695 & n3612 ;
  assign n3616 = n3615 ^ x653 ;
  assign n3617 = n3611 & ~n3616 ;
  assign n3631 = n3630 ^ n3617 ;
  assign n3632 = ~x649 & ~n3631 ;
  assign n1692 = x650 ^ x649 ;
  assign n1694 = n1693 ^ n1692 ;
  assign n3641 = n1694 & n3618 ;
  assign n3642 = ~x650 & n3641 ;
  assign n3643 = n3642 ^ x650 ;
  assign n3633 = x649 & x650 ;
  assign n3634 = ~x653 & n3633 ;
  assign n3635 = n3634 ^ x650 ;
  assign n3644 = n3643 ^ n3635 ;
  assign n3645 = n3620 & n3644 ;
  assign n3646 = n3645 ^ n3634 ;
  assign n3647 = x654 & ~n3620 ;
  assign n3648 = n3633 & n3647 ;
  assign n3649 = n3648 ^ n3633 ;
  assign n3650 = n3649 ^ n3622 ;
  assign n3655 = n3619 & n3620 ;
  assign n3656 = n3655 ^ n3649 ;
  assign n3657 = n3650 & ~n3656 ;
  assign n3658 = n3657 ^ n3649 ;
  assign n3659 = ~n1692 & n3658 ;
  assign n3660 = n3657 & n3659 ;
  assign n3661 = n3660 ^ n3658 ;
  assign n3662 = ~n3646 & ~n3661 ;
  assign n3663 = ~n3632 & n3662 ;
  assign n3587 = ~x645 & ~x646 ;
  assign n3585 = ~x647 & ~x648 ;
  assign n3596 = n3587 ^ n3585 ;
  assign n3595 = n3585 & n3587 ;
  assign n3597 = n3596 ^ n3595 ;
  assign n1688 = x648 ^ x647 ;
  assign n3586 = n3585 ^ n1688 ;
  assign n1690 = x646 ^ x645 ;
  assign n3588 = n3587 ^ n1690 ;
  assign n3590 = n3586 & n3588 ;
  assign n3598 = n3597 ^ n3590 ;
  assign n1687 = x644 ^ x643 ;
  assign n3606 = n3585 ^ n1687 ;
  assign n3607 = n3606 ^ n3587 ;
  assign n3608 = ~n3595 & ~n3607 ;
  assign n3609 = ~n3598 & ~n3608 ;
  assign n3589 = n3588 ^ n3586 ;
  assign n3591 = n3590 ^ n3589 ;
  assign n3592 = x643 & x644 ;
  assign n3593 = n3591 & n3592 ;
  assign n3594 = n3593 ^ n1687 ;
  assign n3599 = n3590 ^ n1687 ;
  assign n3600 = ~n3598 & n3599 ;
  assign n3601 = n3594 & n3600 ;
  assign n3602 = n3601 ^ n3593 ;
  assign n3603 = n3591 & ~n3602 ;
  assign n3604 = n3603 ^ n3602 ;
  assign n3605 = n3604 ^ n3592 ;
  assign n3610 = n3609 ^ n3605 ;
  assign n3664 = n3663 ^ n3610 ;
  assign n1696 = n1695 ^ n1694 ;
  assign n1706 = x642 ^ x641 ;
  assign n1704 = x640 ^ x639 ;
  assign n1703 = x638 ^ x637 ;
  assign n1705 = n1704 ^ n1703 ;
  assign n1707 = n1706 ^ n1705 ;
  assign n1689 = n1688 ^ n1687 ;
  assign n1691 = n1690 ^ n1689 ;
  assign n3579 = n1707 ^ n1691 ;
  assign n1701 = x636 ^ x635 ;
  assign n1699 = x634 ^ x633 ;
  assign n1698 = x632 ^ x631 ;
  assign n1700 = n1699 ^ n1698 ;
  assign n1702 = n1701 ^ n1700 ;
  assign n3582 = n3579 ^ n1702 ;
  assign n3583 = ~n1696 & n3582 ;
  assign n3580 = n1702 ^ n1691 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3584 = n3583 ^ n3581 ;
  assign n3665 = n3664 ^ n3584 ;
  assign n3531 = x639 & x640 ;
  assign n3532 = n3531 ^ x638 ;
  assign n3535 = n1704 ^ x637 ;
  assign n3536 = ~x642 & n3535 ;
  assign n3537 = n3536 ^ x637 ;
  assign n3538 = ~n3531 & n3537 ;
  assign n3539 = n3538 ^ x637 ;
  assign n3540 = ~n3532 & n3539 ;
  assign n3541 = ~x641 & n3540 ;
  assign n3542 = x641 & x642 ;
  assign n3543 = n3542 ^ n1706 ;
  assign n3548 = n3531 & n3542 ;
  assign n3544 = n3542 ^ x640 ;
  assign n3549 = n3548 ^ n3544 ;
  assign n3545 = n1704 & ~n3544 ;
  assign n3550 = n3549 ^ n3545 ;
  assign n3546 = n3545 ^ x639 ;
  assign n3547 = n3546 ^ n3531 ;
  assign n3551 = n3550 ^ n3547 ;
  assign n3552 = n3551 ^ n3546 ;
  assign n3555 = x638 & n3552 ;
  assign n3556 = n3555 ^ n3546 ;
  assign n3557 = ~n1703 & n3556 ;
  assign n3558 = n3557 ^ n3546 ;
  assign n3559 = n3543 & n3558 ;
  assign n3560 = x637 & x638 ;
  assign n3561 = ~x642 & n3531 ;
  assign n3562 = n3560 & n3561 ;
  assign n3563 = ~n3559 & ~n3562 ;
  assign n3564 = ~x637 & n3563 ;
  assign n3565 = x638 & n3543 ;
  assign n3573 = ~n3550 & ~n3565 ;
  assign n3566 = n3546 & ~n3548 ;
  assign n3567 = ~n3565 & n3566 ;
  assign n3568 = n3567 ^ n3546 ;
  assign n3574 = n3573 ^ n3568 ;
  assign n3575 = n3564 & n3574 ;
  assign n3576 = n3575 ^ n3563 ;
  assign n3577 = ~n3541 & n3576 ;
  assign n3493 = x635 ^ x634 ;
  assign n3497 = ~n1701 & ~n3493 ;
  assign n3492 = x633 ^ x632 ;
  assign n3494 = n3493 ^ x633 ;
  assign n3495 = n3494 ^ x636 ;
  assign n3496 = ~n3492 & n3495 ;
  assign n3498 = n3497 ^ n3496 ;
  assign n3499 = ~x631 & n3498 ;
  assign n3500 = ~n1699 & ~n3492 ;
  assign n3501 = x636 ^ x631 ;
  assign n3504 = ~x634 & ~n3501 ;
  assign n3505 = n3504 ^ x631 ;
  assign n3506 = n3500 & n3505 ;
  assign n3507 = ~x635 & n3506 ;
  assign n3508 = ~x633 & ~x634 ;
  assign n3511 = n3508 ^ n1699 ;
  assign n3512 = x631 & x632 ;
  assign n3513 = x636 & n3512 ;
  assign n3514 = ~n3511 & n3513 ;
  assign n3515 = n3514 ^ n3512 ;
  assign n3509 = ~x635 & ~x636 ;
  assign n3510 = ~n3508 & ~n3509 ;
  assign n3516 = n3515 ^ n3510 ;
  assign n3517 = n3509 ^ n1701 ;
  assign n3522 = n3511 & n3517 ;
  assign n3523 = n3522 ^ n3510 ;
  assign n3524 = n3516 & n3523 ;
  assign n3525 = n3524 ^ n3515 ;
  assign n3526 = ~n1698 & n3525 ;
  assign n3527 = n3524 & n3526 ;
  assign n3528 = n3527 ^ n3525 ;
  assign n3529 = ~n3507 & ~n3528 ;
  assign n3530 = ~n3499 & n3529 ;
  assign n3578 = n3577 ^ n3530 ;
  assign n3666 = n3665 ^ n3578 ;
  assign n1683 = x618 ^ x617 ;
  assign n3452 = x617 ^ x616 ;
  assign n3456 = ~n1683 & ~n3452 ;
  assign n3451 = x615 ^ x614 ;
  assign n3453 = n3452 ^ x615 ;
  assign n3454 = n3453 ^ x618 ;
  assign n3455 = ~n3451 & n3454 ;
  assign n3457 = n3456 ^ n3455 ;
  assign n3458 = ~x613 & n3457 ;
  assign n1681 = x616 ^ x615 ;
  assign n3459 = ~n1681 & ~n3451 ;
  assign n3460 = x618 ^ x613 ;
  assign n3463 = ~x616 & ~n3460 ;
  assign n3464 = n3463 ^ x613 ;
  assign n3465 = n3459 & n3464 ;
  assign n3466 = ~x617 & n3465 ;
  assign n3467 = ~x615 & ~x616 ;
  assign n3470 = n3467 ^ n1681 ;
  assign n3471 = x613 & x614 ;
  assign n3472 = x618 & n3471 ;
  assign n3473 = ~n3470 & n3472 ;
  assign n3474 = n3473 ^ n3471 ;
  assign n3468 = ~x617 & ~x618 ;
  assign n3469 = ~n3467 & ~n3468 ;
  assign n3475 = n3474 ^ n3469 ;
  assign n3476 = n3468 ^ n1683 ;
  assign n3481 = n3470 & n3476 ;
  assign n3482 = n3481 ^ n3469 ;
  assign n3483 = n3475 & n3482 ;
  assign n1680 = x614 ^ x613 ;
  assign n3484 = n3483 ^ n3474 ;
  assign n3485 = ~n1680 & n3484 ;
  assign n3486 = n3483 & n3485 ;
  assign n3487 = n3486 ^ n3484 ;
  assign n3488 = ~n3466 & ~n3487 ;
  assign n3489 = ~n3458 & n3488 ;
  assign n3397 = ~x609 & ~x610 ;
  assign n1676 = x610 ^ x609 ;
  assign n3406 = n3397 ^ n1676 ;
  assign n3404 = ~x611 & ~x612 ;
  assign n1678 = x612 ^ x611 ;
  assign n3405 = n3404 ^ n1678 ;
  assign n3407 = n3406 ^ n3405 ;
  assign n3408 = ~n3397 & ~n3404 ;
  assign n3413 = x608 & n3408 ;
  assign n3414 = n3413 ^ n3405 ;
  assign n3415 = n3407 & n3414 ;
  assign n3416 = n3415 ^ n3406 ;
  assign n3398 = x611 ^ x608 ;
  assign n3401 = n1678 & n3398 ;
  assign n3402 = n3401 ^ x611 ;
  assign n3403 = n3397 & ~n3402 ;
  assign n3417 = n3416 ^ n3403 ;
  assign n3418 = ~x607 & ~n3417 ;
  assign n1675 = x608 ^ x607 ;
  assign n1677 = n1676 ^ n1675 ;
  assign n3419 = x607 & x608 ;
  assign n3420 = ~x611 & n3419 ;
  assign n3425 = n3420 ^ n3404 ;
  assign n3428 = n1677 & n3425 ;
  assign n3429 = ~x608 & n3428 ;
  assign n3430 = n3429 ^ x608 ;
  assign n3421 = n3420 ^ x608 ;
  assign n3431 = n3430 ^ n3421 ;
  assign n3432 = n3406 & n3431 ;
  assign n3433 = n3432 ^ n3420 ;
  assign n3434 = x612 & ~n3406 ;
  assign n3435 = n3419 & n3434 ;
  assign n3436 = n3435 ^ n3419 ;
  assign n3437 = n3436 ^ n3408 ;
  assign n3442 = n3405 & n3406 ;
  assign n3443 = n3442 ^ n3436 ;
  assign n3444 = n3437 & ~n3443 ;
  assign n3445 = n3444 ^ n3436 ;
  assign n3446 = ~n1675 & n3445 ;
  assign n3447 = n3444 & n3446 ;
  assign n3448 = n3447 ^ n3445 ;
  assign n3449 = ~n3433 & ~n3448 ;
  assign n3450 = ~n3418 & n3449 ;
  assign n3490 = n3489 ^ n3450 ;
  assign n1665 = x626 ^ x625 ;
  assign n3373 = ~x627 & ~x628 ;
  assign n1667 = x628 ^ x627 ;
  assign n3374 = n3373 ^ n1667 ;
  assign n3375 = x629 & x630 ;
  assign n1664 = x630 ^ x629 ;
  assign n3376 = n3375 ^ n1664 ;
  assign n3378 = ~n3374 & n3376 ;
  assign n3390 = ~n3373 & n3375 ;
  assign n3391 = ~n3378 & ~n3390 ;
  assign n3392 = n1665 & ~n3391 ;
  assign n3377 = n3376 ^ n3374 ;
  assign n3379 = n3378 ^ n3377 ;
  assign n3383 = n3379 ^ x626 ;
  assign n3380 = n3375 ^ x628 ;
  assign n3381 = ~n1667 & ~n3380 ;
  assign n3384 = n3383 ^ n3381 ;
  assign n3385 = n1665 & ~n3384 ;
  assign n3386 = n3385 ^ x625 ;
  assign n3382 = ~n3379 & ~n3381 ;
  assign n3388 = n3386 ^ n3382 ;
  assign n3387 = ~n3382 & ~n3386 ;
  assign n3389 = n3388 ^ n3387 ;
  assign n3393 = n3392 ^ n3389 ;
  assign n3394 = n3393 ^ n3387 ;
  assign n1670 = x620 ^ x619 ;
  assign n3351 = ~x621 & ~x622 ;
  assign n1672 = x622 ^ x621 ;
  assign n3352 = n3351 ^ n1672 ;
  assign n3353 = x623 & x624 ;
  assign n1669 = x624 ^ x623 ;
  assign n3354 = n3353 ^ n1669 ;
  assign n3356 = ~n3352 & n3354 ;
  assign n3368 = ~n3351 & n3353 ;
  assign n3369 = ~n3356 & ~n3368 ;
  assign n3370 = n1670 & ~n3369 ;
  assign n3355 = n3354 ^ n3352 ;
  assign n3357 = n3356 ^ n3355 ;
  assign n3361 = n3357 ^ x620 ;
  assign n3358 = n3353 ^ x622 ;
  assign n3359 = ~n1672 & ~n3358 ;
  assign n3362 = n3361 ^ n3359 ;
  assign n3363 = n1670 & ~n3362 ;
  assign n3364 = n3363 ^ x619 ;
  assign n3360 = ~n3357 & ~n3359 ;
  assign n3366 = n3364 ^ n3360 ;
  assign n3365 = ~n3360 & ~n3364 ;
  assign n3367 = n3366 ^ n3365 ;
  assign n3371 = n3370 ^ n3367 ;
  assign n3372 = n3371 ^ n3365 ;
  assign n3395 = n3394 ^ n3372 ;
  assign n1679 = n1678 ^ n1677 ;
  assign n1682 = n1681 ^ n1680 ;
  assign n1684 = n1683 ^ n1682 ;
  assign n3349 = n1679 & n1684 ;
  assign n1666 = n1665 ^ n1664 ;
  assign n1668 = n1667 ^ n1666 ;
  assign n1671 = n1670 ^ n1669 ;
  assign n1673 = n1672 ^ n1671 ;
  assign n3347 = n1668 & n1673 ;
  assign n1674 = n1673 ^ n1668 ;
  assign n1685 = n1684 ^ n1679 ;
  assign n3346 = n1674 & n1685 ;
  assign n3348 = n3347 ^ n3346 ;
  assign n3350 = n3349 ^ n3348 ;
  assign n3396 = n3395 ^ n3350 ;
  assign n3491 = n3490 ^ n3396 ;
  assign n3667 = n3666 ^ n3491 ;
  assign n3284 = x587 & x588 ;
  assign n1647 = x588 ^ x587 ;
  assign n3286 = n3284 ^ n1647 ;
  assign n3287 = n3286 ^ x584 ;
  assign n3282 = ~x585 & ~x586 ;
  assign n3288 = n3287 ^ n3282 ;
  assign n3290 = n3286 ^ n3282 ;
  assign n3289 = n3282 & ~n3286 ;
  assign n3291 = n3290 ^ n3289 ;
  assign n3292 = ~n3288 & ~n3291 ;
  assign n3341 = n3289 ^ x583 ;
  assign n3342 = ~n3292 & ~n3341 ;
  assign n1646 = x586 ^ x585 ;
  assign n3283 = n3282 ^ n1646 ;
  assign n3299 = x587 ^ x584 ;
  assign n3300 = n3299 ^ x586 ;
  assign n3301 = n3300 ^ x588 ;
  assign n3297 = x587 ^ x585 ;
  assign n3302 = n3301 ^ n3297 ;
  assign n3303 = n3302 ^ x588 ;
  assign n3304 = n3303 ^ x587 ;
  assign n3305 = n3304 ^ n3297 ;
  assign n1648 = n1647 ^ n1646 ;
  assign n3311 = n3297 ^ n1648 ;
  assign n3312 = ~n3305 & ~n3311 ;
  assign n3313 = ~x587 & n3312 ;
  assign n3316 = n3313 ^ n3312 ;
  assign n3314 = n3313 ^ n3297 ;
  assign n3315 = n3302 & n3314 ;
  assign n3317 = n3316 ^ n3315 ;
  assign n3318 = n3317 ^ x587 ;
  assign n3336 = n3318 ^ x583 ;
  assign n3335 = x583 & n3318 ;
  assign n3337 = n3336 ^ n3335 ;
  assign n3338 = ~n3284 & ~n3337 ;
  assign n3339 = n3283 & n3338 ;
  assign n1641 = x590 ^ x589 ;
  assign n3329 = x589 & ~n1641 ;
  assign n1643 = x594 ^ x593 ;
  assign n3328 = x593 & ~n1643 ;
  assign n3330 = n3329 ^ n3328 ;
  assign n1640 = x592 ^ x591 ;
  assign n1642 = n1641 ^ n1640 ;
  assign n3326 = n1643 ^ n1641 ;
  assign n3327 = n1642 & ~n3326 ;
  assign n3331 = n3330 ^ n3327 ;
  assign n3325 = ~x591 & ~x592 ;
  assign n3332 = n3331 ^ n3325 ;
  assign n3333 = n3332 ^ n3318 ;
  assign n3285 = n3284 ^ n3283 ;
  assign n3293 = n3292 ^ n3288 ;
  assign n3294 = n3293 ^ n3283 ;
  assign n3295 = ~n3285 & ~n3294 ;
  assign n3296 = n3295 ^ n3284 ;
  assign n3322 = ~x583 & ~n3317 ;
  assign n3323 = n3322 ^ x587 ;
  assign n3324 = n3296 & ~n3323 ;
  assign n3334 = n3333 ^ n3324 ;
  assign n3340 = n3339 ^ n3334 ;
  assign n3343 = n3342 ^ n3340 ;
  assign n1659 = x600 ^ x599 ;
  assign n3242 = x599 ^ x598 ;
  assign n3246 = ~n1659 & ~n3242 ;
  assign n3241 = x597 ^ x596 ;
  assign n3243 = n3242 ^ x597 ;
  assign n3244 = n3243 ^ x600 ;
  assign n3245 = ~n3241 & n3244 ;
  assign n3247 = n3246 ^ n3245 ;
  assign n3248 = ~x595 & n3247 ;
  assign n1657 = x598 ^ x597 ;
  assign n3249 = ~n1657 & ~n3241 ;
  assign n3250 = x600 ^ x595 ;
  assign n3253 = ~x598 & ~n3250 ;
  assign n3254 = n3253 ^ x595 ;
  assign n3255 = n3249 & n3254 ;
  assign n3256 = ~x599 & n3255 ;
  assign n3257 = ~x597 & ~x598 ;
  assign n3260 = n3257 ^ n1657 ;
  assign n3261 = x595 & x596 ;
  assign n3262 = x600 & n3261 ;
  assign n3263 = ~n3260 & n3262 ;
  assign n3264 = n3263 ^ n3261 ;
  assign n3258 = ~x599 & ~x600 ;
  assign n3259 = ~n3257 & ~n3258 ;
  assign n3265 = n3264 ^ n3259 ;
  assign n3266 = n3258 ^ n1659 ;
  assign n3271 = n3260 & n3266 ;
  assign n3272 = n3271 ^ n3259 ;
  assign n3273 = n3265 & n3272 ;
  assign n1656 = x596 ^ x595 ;
  assign n3274 = n3273 ^ n3264 ;
  assign n3275 = ~n1656 & n3274 ;
  assign n3276 = n3273 & n3275 ;
  assign n3277 = n3276 ^ n3274 ;
  assign n3278 = ~n3256 & ~n3277 ;
  assign n3279 = ~n3248 & n3278 ;
  assign n1654 = x606 ^ x605 ;
  assign n3203 = x605 ^ x604 ;
  assign n3207 = ~n1654 & ~n3203 ;
  assign n3202 = x603 ^ x602 ;
  assign n3204 = n3203 ^ x603 ;
  assign n3205 = n3204 ^ x606 ;
  assign n3206 = ~n3202 & n3205 ;
  assign n3208 = n3207 ^ n3206 ;
  assign n3209 = ~x601 & n3208 ;
  assign n1652 = x604 ^ x603 ;
  assign n3210 = ~n1652 & ~n3202 ;
  assign n3211 = x606 ^ x601 ;
  assign n3214 = ~x604 & ~n3211 ;
  assign n3215 = n3214 ^ x601 ;
  assign n3216 = n3210 & n3215 ;
  assign n3217 = ~x605 & n3216 ;
  assign n3218 = ~x603 & ~x604 ;
  assign n3221 = n3218 ^ n1652 ;
  assign n3222 = x601 & x602 ;
  assign n3223 = x606 & n3222 ;
  assign n3224 = ~n3221 & n3223 ;
  assign n3225 = n3224 ^ n3222 ;
  assign n3219 = ~x605 & ~x606 ;
  assign n3220 = ~n3218 & ~n3219 ;
  assign n3226 = n3225 ^ n3220 ;
  assign n3227 = n3219 ^ n1654 ;
  assign n3232 = n3221 & n3227 ;
  assign n3233 = n3232 ^ n3220 ;
  assign n3234 = n3226 & n3233 ;
  assign n1651 = x602 ^ x601 ;
  assign n3235 = n3234 ^ n3225 ;
  assign n3236 = ~n1651 & n3235 ;
  assign n3237 = n3234 & n3236 ;
  assign n3238 = n3237 ^ n3235 ;
  assign n3239 = ~n3217 & ~n3238 ;
  assign n3240 = ~n3209 & n3239 ;
  assign n3280 = n3279 ^ n3240 ;
  assign n1644 = n1643 ^ n1642 ;
  assign n1645 = x584 ^ x583 ;
  assign n1649 = n1648 ^ n1645 ;
  assign n3199 = n1644 & n1649 ;
  assign n1635 = x560 ^ x559 ;
  assign n1634 = x564 ^ x563 ;
  assign n1636 = n1635 ^ n1634 ;
  assign n1633 = x562 ^ x561 ;
  assign n1637 = n1636 ^ n1633 ;
  assign n1630 = x566 ^ x565 ;
  assign n1629 = x568 ^ x567 ;
  assign n1631 = n1630 ^ n1629 ;
  assign n1628 = x570 ^ x569 ;
  assign n1632 = n1631 ^ n1628 ;
  assign n1638 = n1637 ^ n1632 ;
  assign n1625 = x576 ^ x575 ;
  assign n1623 = x574 ^ x573 ;
  assign n1622 = x572 ^ x571 ;
  assign n1624 = n1623 ^ n1622 ;
  assign n1626 = n1625 ^ n1624 ;
  assign n1620 = x582 ^ x581 ;
  assign n1618 = x580 ^ x579 ;
  assign n1617 = x578 ^ x577 ;
  assign n1619 = n1618 ^ n1617 ;
  assign n1621 = n1620 ^ n1619 ;
  assign n1627 = n1626 ^ n1621 ;
  assign n1639 = n1638 ^ n1627 ;
  assign n1658 = n1657 ^ n1656 ;
  assign n1660 = n1659 ^ n1658 ;
  assign n1653 = n1652 ^ n1651 ;
  assign n1655 = n1654 ^ n1653 ;
  assign n1661 = n1660 ^ n1655 ;
  assign n1650 = n1649 ^ n1644 ;
  assign n1662 = n1661 ^ n1650 ;
  assign n3198 = n1639 & n1662 ;
  assign n3200 = n3199 ^ n3198 ;
  assign n3195 = n1655 ^ n1650 ;
  assign n3196 = n1661 & ~n3195 ;
  assign n3197 = n3196 ^ n1660 ;
  assign n3201 = n3200 ^ n3197 ;
  assign n3281 = n3280 ^ n3201 ;
  assign n3344 = n3343 ^ n3281 ;
  assign n3185 = x581 & x582 ;
  assign n3184 = x579 & x580 ;
  assign n3186 = n3185 ^ n3184 ;
  assign n3187 = n3184 ^ n1618 ;
  assign n3188 = n3185 ^ n1620 ;
  assign n3189 = n3187 & n3188 ;
  assign n3190 = n3189 ^ n3184 ;
  assign n3191 = ~n3186 & ~n3190 ;
  assign n3163 = n1620 ^ x578 ;
  assign n3164 = n3163 ^ n1618 ;
  assign n3170 = x575 & x576 ;
  assign n3169 = x573 & x574 ;
  assign n3171 = n3170 ^ n3169 ;
  assign n3172 = n3169 ^ n1623 ;
  assign n3173 = n3170 ^ n1625 ;
  assign n3174 = n3172 & n3173 ;
  assign n3175 = n3174 ^ n3169 ;
  assign n3176 = ~n3171 & ~n3175 ;
  assign n3165 = n1625 ^ x572 ;
  assign n3166 = n3165 ^ n1623 ;
  assign n3167 = n1622 & ~n3166 ;
  assign n3168 = n3167 ^ x571 ;
  assign n3177 = n3176 ^ n3168 ;
  assign n3178 = n3177 ^ x577 ;
  assign n3179 = n3178 ^ n1620 ;
  assign n3180 = n3179 ^ n1618 ;
  assign n3181 = n3180 ^ n3177 ;
  assign n3182 = ~n3164 & n3181 ;
  assign n3183 = n3182 ^ n3178 ;
  assign n3192 = n3191 ^ n3183 ;
  assign n3158 = n1632 ^ n1626 ;
  assign n3161 = ~n1627 & ~n3158 ;
  assign n3159 = n3158 ^ n1621 ;
  assign n3160 = ~n1637 & n3159 ;
  assign n3162 = n3161 ^ n3160 ;
  assign n3193 = n3192 ^ n3162 ;
  assign n3122 = ~x563 & ~x564 ;
  assign n3121 = ~x561 & ~x562 ;
  assign n3123 = n3122 ^ n3121 ;
  assign n3125 = n3122 ^ n1634 ;
  assign n3124 = n3121 ^ n1633 ;
  assign n3128 = n3125 ^ n3124 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = n3126 ^ n3121 ;
  assign n3129 = n3128 ^ n3127 ;
  assign n3130 = n3129 ^ n3121 ;
  assign n3133 = ~n1635 & ~n3130 ;
  assign n3134 = n3133 ^ n3121 ;
  assign n3135 = n3123 & ~n3134 ;
  assign n3136 = n3135 ^ n3122 ;
  assign n3137 = ~n3121 & ~n3122 ;
  assign n3142 = n1635 & n3137 ;
  assign n3143 = n3142 ^ n3125 ;
  assign n3152 = n3128 & n3143 ;
  assign n3144 = x559 & x560 ;
  assign n3145 = ~n3126 & n3144 ;
  assign n3146 = ~n3128 & ~n3137 ;
  assign n3147 = n3145 & n3146 ;
  assign n3148 = n3147 ^ n3145 ;
  assign n3149 = n3148 ^ n3124 ;
  assign n3153 = n3152 ^ n3149 ;
  assign n3154 = ~n3136 & n3153 ;
  assign n3155 = n3148 ^ n3144 ;
  assign n3156 = ~n3154 & ~n3155 ;
  assign n3066 = ~x567 & ~x568 ;
  assign n3065 = x569 & x570 ;
  assign n3075 = n3066 ^ n3065 ;
  assign n3067 = n3065 & ~n3066 ;
  assign n3076 = n3075 ^ n3067 ;
  assign n3068 = n3066 ^ n1629 ;
  assign n3069 = n3065 ^ n1628 ;
  assign n3070 = ~n3068 & n3069 ;
  assign n3072 = n3070 ^ n3067 ;
  assign n3071 = ~n3067 & ~n3070 ;
  assign n3073 = n3072 ^ n3071 ;
  assign n3077 = n3076 ^ n3073 ;
  assign n3074 = n3073 ^ x566 ;
  assign n3078 = n3077 ^ n3074 ;
  assign n3079 = n3069 ^ n3068 ;
  assign n3080 = n3079 ^ n3070 ;
  assign n3081 = n3080 ^ x566 ;
  assign n3082 = ~n3078 & ~n3081 ;
  assign n3083 = n3082 ^ n3074 ;
  assign n3084 = ~x565 & n3083 ;
  assign n3116 = ~x566 & n3066 ;
  assign n3117 = n3080 & n3116 ;
  assign n3118 = n3117 ^ n3080 ;
  assign n3085 = x567 ^ x566 ;
  assign n3086 = n3085 ^ x568 ;
  assign n3087 = n3086 ^ x569 ;
  assign n3088 = n3087 ^ x570 ;
  assign n3089 = n3088 ^ x566 ;
  assign n3090 = n3088 ^ x569 ;
  assign n3091 = n3090 ^ x566 ;
  assign n3092 = ~n3089 & ~n3091 ;
  assign n3093 = n3092 ^ x566 ;
  assign n3102 = x569 ^ x566 ;
  assign n3095 = n3088 ^ x567 ;
  assign n3096 = n3095 ^ n3087 ;
  assign n3100 = ~n1629 & ~n3096 ;
  assign n3103 = n3102 ^ n3100 ;
  assign n3104 = ~n3093 & ~n3103 ;
  assign n3105 = n3104 ^ x566 ;
  assign n3106 = n3105 ^ n3088 ;
  assign n3107 = n3106 ^ x566 ;
  assign n3108 = ~n1630 & n3107 ;
  assign n3109 = n3108 ^ n3071 ;
  assign n3110 = n3109 ^ n3080 ;
  assign n3119 = n3118 ^ n3110 ;
  assign n3120 = ~n3084 & n3119 ;
  assign n3157 = n3156 ^ n3120 ;
  assign n3194 = n3193 ^ n3157 ;
  assign n3345 = n3344 ^ n3194 ;
  assign n3668 = n3667 ^ n3345 ;
  assign n1686 = n1685 ^ n1674 ;
  assign n1663 = n1662 ^ n1639 ;
  assign n3049 = n1686 ^ n1663 ;
  assign n1806 = n1805 ^ n1758 ;
  assign n3050 = n3049 ^ n1806 ;
  assign n1708 = n1707 ^ n1702 ;
  assign n1697 = n1696 ^ n1691 ;
  assign n1709 = n1708 ^ n1697 ;
  assign n3051 = n1806 ^ n1709 ;
  assign n3052 = n3050 & ~n3051 ;
  assign n3053 = n3052 ^ n1663 ;
  assign n3054 = n1686 & n3053 ;
  assign n3055 = ~n3052 & n3054 ;
  assign n3056 = n3055 ^ n3053 ;
  assign n9730 = n3056 ^ n1686 ;
  assign n1710 = n1709 ^ n1686 ;
  assign n3058 = n1709 ^ n1663 ;
  assign n3059 = n1710 & ~n3058 ;
  assign n1711 = n1710 ^ n1663 ;
  assign n3057 = n1711 & n1806 ;
  assign n3060 = n3059 ^ n3057 ;
  assign n3061 = n3060 ^ n3056 ;
  assign n3064 = n9730 ^ n3061 ;
  assign n3669 = n3668 ^ n3064 ;
  assign n4125 = n9750 ^ n3669 ;
  assign n10994 = n10993 ^ n4125 ;
  assign n3047 = n3046 ^ n2487 ;
  assign n1807 = n1806 ^ n1711 ;
  assign n2008 = n1807 & ~n2001 ;
  assign n2009 = n2008 ^ n2003 ;
  assign n2010 = n2002 & ~n2009 ;
  assign n3048 = n3047 ^ n2010 ;
  assign n10351 = n4125 ^ n2002 ;
  assign n10352 = n10351 ^ n2003 ;
  assign n10353 = n10352 ^ n2010 ;
  assign n10354 = n3048 & n10353 ;
  assign n10995 = n10994 ^ n10354 ;
  assign n10150 = n1686 & n1709 ;
  assign n10317 = n10150 ^ n3666 ;
  assign n10318 = ~n3667 & ~n10317 ;
  assign n10306 = n3476 ^ n3470 ;
  assign n10307 = x614 & n3469 ;
  assign n10308 = n10307 ^ n3470 ;
  assign n10309 = n10306 & ~n10308 ;
  assign n10310 = n10309 ^ n3470 ;
  assign n10311 = ~n3487 & ~n10310 ;
  assign n10312 = n10311 ^ n3487 ;
  assign n10299 = n3395 ^ n3347 ;
  assign n10301 = n3349 ^ n3346 ;
  assign n10304 = n10299 & n10301 ;
  assign n10300 = n10299 ^ n3349 ;
  assign n10302 = n10301 ^ n10300 ;
  assign n10303 = n3490 & n10302 ;
  assign n10305 = n10304 ^ n10303 ;
  assign n10313 = n10312 ^ n10305 ;
  assign n10296 = n3416 & ~n3448 ;
  assign n10293 = n3450 ^ n3349 ;
  assign n10294 = n3490 & n10293 ;
  assign n10295 = n10294 ^ n3450 ;
  assign n10297 = n10296 ^ n10295 ;
  assign n10288 = n3390 ^ n3378 ;
  assign n10289 = n10288 ^ n3391 ;
  assign n10290 = n3393 & n10289 ;
  assign n10285 = n3368 ^ n3356 ;
  assign n10286 = n10285 ^ n3369 ;
  assign n10287 = n3371 & n10286 ;
  assign n10291 = n10290 ^ n10287 ;
  assign n10282 = n3372 ^ n3347 ;
  assign n10283 = n3395 & n10282 ;
  assign n10284 = n10283 ^ n3372 ;
  assign n10292 = n10291 ^ n10284 ;
  assign n10298 = n10297 ^ n10292 ;
  assign n10314 = n10313 ^ n10298 ;
  assign n10315 = n10314 ^ n3666 ;
  assign n10319 = n10318 ^ n10315 ;
  assign n10342 = n3630 & ~n3661 ;
  assign n10343 = n10342 ^ n3603 ;
  assign n10321 = n1691 & n1696 ;
  assign n10339 = n10321 ^ n3610 ;
  assign n10340 = n3664 & ~n10339 ;
  assign n10341 = n10340 ^ n3663 ;
  assign n10344 = n10343 ^ n10341 ;
  assign n10324 = n1702 & n1707 ;
  assign n10336 = n10324 ^ n3530 ;
  assign n10337 = n3578 & ~n10336 ;
  assign n10338 = n10337 ^ n3577 ;
  assign n10345 = n10344 ^ n10338 ;
  assign n10328 = n3517 ^ n3511 ;
  assign n10329 = x632 & n3510 ;
  assign n10330 = n10329 ^ n3511 ;
  assign n10331 = n10328 & ~n10330 ;
  assign n10332 = n10331 ^ n3511 ;
  assign n10333 = ~n3528 & ~n10332 ;
  assign n10334 = n10333 ^ n3528 ;
  assign n10327 = n3563 & ~n3568 ;
  assign n10335 = n10334 ^ n10327 ;
  assign n10346 = n10345 ^ n10335 ;
  assign n10325 = n3578 & ~n10324 ;
  assign n10320 = n3664 ^ n3578 ;
  assign n10322 = n10321 ^ n10320 ;
  assign n10323 = n3665 & n10322 ;
  assign n10326 = n10325 ^ n10323 ;
  assign n10347 = n10346 ^ n10326 ;
  assign n11220 = n10347 ^ n10314 ;
  assign n11221 = n10319 & n11220 ;
  assign n11222 = n11221 ^ n10314 ;
  assign n11216 = n10290 ^ n10284 ;
  assign n11217 = n10291 & ~n11216 ;
  assign n11218 = n11217 ^ n10290 ;
  assign n11207 = ~n10295 & n10296 ;
  assign n11206 = ~n10305 & ~n10312 ;
  assign n11208 = n11207 ^ n11206 ;
  assign n11209 = n11206 ^ n10292 ;
  assign n11210 = ~n11208 & ~n11209 ;
  assign n11211 = n10314 & ~n11210 ;
  assign n11212 = n11210 ^ n10292 ;
  assign n11213 = n11212 ^ n11208 ;
  assign n11214 = n11211 & n11213 ;
  assign n11215 = n11214 ^ n11212 ;
  assign n11219 = n11218 ^ n11215 ;
  assign n11223 = n11222 ^ n11219 ;
  assign n11201 = n10341 ^ n3603 ;
  assign n11202 = n10343 & ~n11201 ;
  assign n11203 = n11202 ^ n3603 ;
  assign n11197 = n10344 ^ n10327 ;
  assign n11198 = n10335 ^ n10326 ;
  assign n11199 = n11198 ^ n10338 ;
  assign n11200 = n11197 & ~n11199 ;
  assign n11204 = n11203 ^ n11200 ;
  assign n11194 = n10338 ^ n10326 ;
  assign n11195 = n10334 ^ n10326 ;
  assign n11196 = ~n11194 & ~n11195 ;
  assign n11205 = n11204 ^ n11196 ;
  assign n11224 = n11223 ^ n11205 ;
  assign n10151 = n10150 ^ n3668 ;
  assign n10152 = n10150 ^ n3667 ;
  assign n10278 = n10152 ^ n3668 ;
  assign n9741 = n3059 ^ n1686 ;
  assign n10279 = n10278 ^ n9741 ;
  assign n10280 = ~n10151 & ~n10279 ;
  assign n10263 = n3227 ^ n3221 ;
  assign n10264 = x602 & n3220 ;
  assign n10265 = n10264 ^ n3221 ;
  assign n10266 = n10263 & ~n10265 ;
  assign n10267 = n10266 ^ n3221 ;
  assign n10268 = ~n3238 & ~n10267 ;
  assign n10269 = n10268 ^ n3238 ;
  assign n10257 = n3266 ^ n3260 ;
  assign n10258 = x596 & n3259 ;
  assign n10259 = n10258 ^ n3260 ;
  assign n10260 = n10257 & ~n10259 ;
  assign n10261 = n10260 ^ n3260 ;
  assign n10262 = ~n3277 & n10261 ;
  assign n10270 = n10269 ^ n10262 ;
  assign n10214 = n1655 & n1660 ;
  assign n10254 = n10214 ^ n3240 ;
  assign n10255 = n3280 & ~n10254 ;
  assign n10256 = n10255 ^ n3279 ;
  assign n10271 = n10270 ^ n10256 ;
  assign n10230 = n3325 ^ n1640 ;
  assign n10231 = x594 & n3329 ;
  assign n10232 = ~n10230 & n10231 ;
  assign n10233 = n10232 ^ n3329 ;
  assign n10227 = n3328 ^ n1643 ;
  assign n10228 = ~n3325 & n10227 ;
  assign n10234 = n10233 ^ n10228 ;
  assign n10239 = ~n3328 & n10230 ;
  assign n10240 = n10239 ^ n10228 ;
  assign n10241 = n10234 & n10240 ;
  assign n10243 = n10241 ^ n10233 ;
  assign n10229 = ~n1641 & n10228 ;
  assign n10242 = n10229 & n10241 ;
  assign n10244 = n10243 ^ n10242 ;
  assign n10245 = n10230 ^ n3328 ;
  assign n10246 = x590 & n10228 ;
  assign n10247 = n10246 ^ n3328 ;
  assign n10248 = ~n10245 & n10247 ;
  assign n10249 = n10248 ^ n3328 ;
  assign n10250 = ~n10244 & n10249 ;
  assign n10251 = n10250 ^ n10244 ;
  assign n10226 = ~n3296 & ~n3335 ;
  assign n10252 = n10251 ^ n10226 ;
  assign n10223 = n3332 ^ n3199 ;
  assign n10224 = n3343 & ~n10223 ;
  assign n10225 = n10224 ^ n3332 ;
  assign n10253 = n10252 ^ n10225 ;
  assign n10272 = n10271 ^ n10253 ;
  assign n10215 = n3280 ^ n3199 ;
  assign n10217 = n10214 ^ n3199 ;
  assign n10221 = n10215 & ~n10217 ;
  assign n10213 = n3343 ^ n3280 ;
  assign n10219 = n3280 ^ n3197 ;
  assign n10220 = n10213 & n10219 ;
  assign n10222 = n10221 ^ n10220 ;
  assign n10273 = n10272 ^ n10222 ;
  assign n10192 = ~n3120 & n3156 ;
  assign n10206 = ~n3193 & n10192 ;
  assign n10193 = n10192 ^ n3157 ;
  assign n10207 = n10206 ^ n10193 ;
  assign n10195 = n1632 & n1637 ;
  assign n10196 = n10195 ^ n1621 ;
  assign n10197 = n10196 ^ n1638 ;
  assign n10198 = n10197 ^ n1621 ;
  assign n10201 = ~n3192 & n10198 ;
  assign n10202 = n10201 ^ n1621 ;
  assign n10203 = n1627 & n10202 ;
  assign n10199 = n3192 ^ n1621 ;
  assign n10204 = n10203 ^ n10199 ;
  assign n10208 = ~n10195 & ~n10204 ;
  assign n10209 = ~n10207 & n10208 ;
  assign n10210 = n10209 ^ n10206 ;
  assign n10194 = n3193 & n10193 ;
  assign n10205 = n10194 & n10204 ;
  assign n10211 = n10210 ^ n10205 ;
  assign n10186 = n1621 & n1626 ;
  assign n10187 = n10186 ^ n3177 ;
  assign n10188 = n3192 & ~n10187 ;
  assign n10189 = n10188 ^ n3177 ;
  assign n10158 = n3189 ^ x578 ;
  assign n10159 = n3186 ^ x577 ;
  assign n10160 = n10159 ^ n3189 ;
  assign n10161 = n10158 & ~n10160 ;
  assign n10162 = n10161 ^ n3190 ;
  assign n10163 = ~n3186 & n10162 ;
  assign n10164 = x577 & n10163 ;
  assign n10165 = n10161 ^ n3189 ;
  assign n10166 = n10165 ^ n10163 ;
  assign n10180 = n10164 & ~n10166 ;
  assign n10167 = n3174 ^ x572 ;
  assign n10168 = n3171 ^ x571 ;
  assign n10169 = n10168 ^ n3174 ;
  assign n10170 = n10167 & ~n10169 ;
  assign n10173 = n10170 ^ n3174 ;
  assign n10171 = n10170 ^ n3175 ;
  assign n10172 = ~n3171 & n10171 ;
  assign n10174 = n10173 ^ n10172 ;
  assign n10175 = x571 & n10172 ;
  assign n10176 = ~n10174 & n10175 ;
  assign n10177 = n10176 ^ n10174 ;
  assign n10178 = n10177 ^ n10166 ;
  assign n10181 = n10180 ^ n10178 ;
  assign n10190 = n10189 ^ n10181 ;
  assign n10156 = n3073 & n3109 ;
  assign n10157 = n10156 ^ n3153 ;
  assign n10191 = n10190 ^ n10157 ;
  assign n10212 = n10211 ^ n10191 ;
  assign n10274 = n10273 ^ n10212 ;
  assign n10153 = n3198 ^ n3194 ;
  assign n10154 = n3344 & n10153 ;
  assign n10155 = n10154 ^ n3198 ;
  assign n10275 = n10274 ^ n10155 ;
  assign n10276 = n10275 ^ n10152 ;
  assign n10281 = n10280 ^ n10276 ;
  assign n10348 = n10347 ^ n10319 ;
  assign n11191 = n10348 ^ n10275 ;
  assign n11192 = ~n10281 & n11191 ;
  assign n11193 = n11192 ^ n10348 ;
  assign n11225 = n11224 ^ n11193 ;
  assign n11159 = n10189 ^ n10177 ;
  assign n11160 = n10181 & ~n11159 ;
  assign n11161 = n11160 ^ n10177 ;
  assign n11167 = ~n10156 & ~n11161 ;
  assign n11168 = n10211 & n11167 ;
  assign n11162 = n10190 & n11161 ;
  assign n11163 = ~n3153 & ~n10156 ;
  assign n11164 = n11163 ^ n3153 ;
  assign n11165 = n11162 & n11164 ;
  assign n11166 = n11165 ^ n11163 ;
  assign n11169 = n11168 ^ n11166 ;
  assign n11179 = n11161 ^ n10210 ;
  assign n11180 = n11179 ^ n10190 ;
  assign n11181 = n11180 ^ n11161 ;
  assign n11171 = n11169 & ~n11181 ;
  assign n11172 = n11171 ^ n11167 ;
  assign n11177 = n3153 & ~n10205 ;
  assign n11178 = n11177 ^ n10190 ;
  assign n11182 = ~n11178 & n11181 ;
  assign n11183 = n11182 ^ n11179 ;
  assign n11184 = n3126 & n10181 ;
  assign n11185 = n10205 & n11184 ;
  assign n11186 = n11185 ^ n10156 ;
  assign n11188 = ~n11183 & n11186 ;
  assign n11189 = ~n11172 & ~n11188 ;
  assign n11156 = n10212 ^ n10155 ;
  assign n11157 = ~n10274 & n11156 ;
  assign n11150 = n10269 ^ n10256 ;
  assign n11151 = ~n10270 & n11150 ;
  assign n11152 = n11151 ^ n10269 ;
  assign n12246 = n10226 ^ n10222 ;
  assign n12247 = n12246 ^ n10251 ;
  assign n11132 = n12247 ^ n10225 ;
  assign n11139 = n10251 ^ n10222 ;
  assign n12245 = n10225 ^ n10222 ;
  assign n11140 = ~n11139 & n12245 ;
  assign n11146 = n10225 & n11140 ;
  assign n11133 = n10271 ^ n10226 ;
  assign n11141 = n11140 ^ n11133 ;
  assign n11147 = n11146 ^ n11141 ;
  assign n11148 = ~n11132 & ~n11147 ;
  assign n11149 = n11148 ^ n11141 ;
  assign n11153 = n11152 ^ n11149 ;
  assign n11154 = n11153 ^ n10212 ;
  assign n11158 = n11157 ^ n11154 ;
  assign n11190 = n11189 ^ n11158 ;
  assign n11226 = n11225 ^ n11190 ;
  assign n10076 = n1727 & n1732 ;
  assign n10125 = n10124 ^ n10076 ;
  assign n10131 = n10125 ^ n10121 ;
  assign n10134 = n3726 & n10131 ;
  assign n10135 = n10134 ^ n10076 ;
  assign n10137 = n10134 ^ n10131 ;
  assign n10138 = n3796 & n10137 ;
  assign n10139 = n10138 ^ n3730 ;
  assign n10140 = n10139 ^ n3796 ;
  assign n10141 = n10135 & ~n10140 ;
  assign n10142 = n10141 ^ n10138 ;
  assign n10143 = n10142 ^ n10121 ;
  assign n10144 = n10143 ^ n3709 ;
  assign n10116 = n3795 ^ n3730 ;
  assign n10117 = n3796 & ~n10116 ;
  assign n10118 = n10117 ^ n3730 ;
  assign n10110 = n3776 ^ x500 ;
  assign n10089 = n3781 ^ n3777 ;
  assign n10095 = n10110 ^ n10089 ;
  assign n10099 = n1717 & n10095 ;
  assign n10093 = n3776 & ~n3780 ;
  assign n10100 = n10099 ^ n10093 ;
  assign n10086 = n3776 ^ x499 ;
  assign n10087 = n10086 ^ n3781 ;
  assign n10091 = n10087 ^ n3777 ;
  assign n10101 = n10100 ^ n10091 ;
  assign n10102 = n10099 ^ n10089 ;
  assign n10103 = n10102 ^ n10091 ;
  assign n10104 = n10101 & n10103 ;
  assign n10105 = ~n3777 & n10104 ;
  assign n10106 = n10105 ^ n10099 ;
  assign n10107 = n10106 ^ n1717 ;
  assign n10113 = n10107 ^ n3776 ;
  assign n10114 = n10113 ^ n10110 ;
  assign n10082 = n3737 & ~n3767 ;
  assign n10115 = n10114 ^ n10082 ;
  assign n10119 = n10118 ^ n10115 ;
  assign n10080 = n3719 ^ n3684 ;
  assign n10077 = n10076 ^ n3713 ;
  assign n10078 = n3726 & n10077 ;
  assign n10079 = n10078 ^ n10076 ;
  assign n10081 = n10080 ^ n10079 ;
  assign n10120 = n10119 ^ n10081 ;
  assign n10145 = n10144 ^ n10120 ;
  assign n10031 = n3798 ^ x476 ;
  assign n10029 = n3798 ^ x475 ;
  assign n10030 = n10029 ^ n3800 ;
  assign n10032 = n10031 ^ n10030 ;
  assign n10052 = n3814 & n10032 ;
  assign n10037 = n10029 ^ n3808 ;
  assign n10042 = n10037 ^ n3798 ;
  assign n10045 = n10037 ^ n3800 ;
  assign n10046 = n10045 ^ x475 ;
  assign n10047 = n10042 & ~n10046 ;
  assign n10053 = n10052 ^ n10047 ;
  assign n10054 = n10053 ^ n10045 ;
  assign n10055 = n10052 ^ n10029 ;
  assign n10056 = n10055 ^ n10045 ;
  assign n10057 = n10054 & n10056 ;
  assign n10058 = ~n3800 & n10057 ;
  assign n10059 = n10058 ^ n10052 ;
  assign n10060 = n10059 ^ n3814 ;
  assign n10063 = n10060 ^ x476 ;
  assign n10023 = n3844 ^ n3838 ;
  assign n10024 = x482 & n3837 ;
  assign n10025 = n10024 ^ n3838 ;
  assign n10026 = n10023 & ~n10025 ;
  assign n10027 = n10026 ^ n3838 ;
  assign n10028 = ~n3855 & n10027 ;
  assign n10072 = n10063 ^ n10028 ;
  assign n10020 = n3867 ^ n3857 ;
  assign n10021 = n3863 & n10020 ;
  assign n10022 = n10021 ^ n3867 ;
  assign n10073 = n10072 ^ n10022 ;
  assign n10009 = n3872 ^ n1746 ;
  assign n10010 = n3884 & n10009 ;
  assign n10013 = n10010 ^ n3875 ;
  assign n10011 = n10010 ^ n3876 ;
  assign n10012 = ~n3872 & n10011 ;
  assign n10014 = n10013 ^ n10012 ;
  assign n10015 = x463 & n10012 ;
  assign n10016 = ~n10014 & n10015 ;
  assign n10017 = n10016 ^ n10014 ;
  assign n10008 = ~n3909 & ~n3915 ;
  assign n10018 = n10017 ^ n10008 ;
  assign n10005 = n3890 ^ n3865 ;
  assign n10006 = n3926 & ~n10005 ;
  assign n10007 = n10006 ^ n3865 ;
  assign n10019 = n10018 ^ n10007 ;
  assign n10074 = n10073 ^ n10019 ;
  assign n9995 = n3863 & n3864 ;
  assign n9986 = n9985 ^ n3864 ;
  assign n9990 = n9989 ^ n9986 ;
  assign n9996 = n9995 ^ n9990 ;
  assign n9998 = n9995 ^ n3864 ;
  assign n9999 = n3926 & n9998 ;
  assign n10000 = n9999 ^ n3865 ;
  assign n10001 = n10000 ^ n3926 ;
  assign n10002 = n9996 & ~n10001 ;
  assign n10003 = n10002 ^ n9999 ;
  assign n10004 = n10003 ^ n9985 ;
  assign n10075 = n10074 ^ n10004 ;
  assign n10146 = n10145 ^ n10075 ;
  assign n9982 = n10124 ^ n3671 ;
  assign n9983 = n3928 & n9982 ;
  assign n9984 = n10124 ^ n9983 ;
  assign n10147 = n10146 ^ n9984 ;
  assign n9962 = ~n4073 & ~n4076 ;
  assign n9961 = n4073 ^ n4069 ;
  assign n9963 = n9962 ^ n9961 ;
  assign n9968 = n4069 & ~n4075 ;
  assign n9969 = n9968 ^ n4066 ;
  assign n9970 = ~n9963 & ~n9969 ;
  assign n9971 = n9970 ^ n9962 ;
  assign n9958 = ~n4081 & n4084 ;
  assign n9959 = n9958 ^ n4083 ;
  assign n9960 = ~n4102 & ~n9959 ;
  assign n9972 = n9971 ^ n9960 ;
  assign n9951 = n4117 ^ n4079 ;
  assign n9952 = n4109 & n9951 ;
  assign n9953 = n9952 ^ n4079 ;
  assign n9973 = n9972 ^ n9953 ;
  assign n9941 = n1797 & n1802 ;
  assign n9948 = n9941 ^ n4056 ;
  assign n9949 = ~n4062 & ~n9948 ;
  assign n9950 = n9949 ^ n9941 ;
  assign n9974 = n9973 ^ n9950 ;
  assign n9939 = ~n4109 & n4119 ;
  assign n9940 = n9939 ^ n4117 ;
  assign n9942 = n9941 ^ n4121 ;
  assign n9945 = ~n4062 & ~n9942 ;
  assign n9946 = n9945 ^ n9941 ;
  assign n9947 = ~n9940 & ~n9946 ;
  assign n9975 = n9974 ^ n9947 ;
  assign n9932 = x541 & ~n4036 ;
  assign n9933 = n4042 & n9932 ;
  assign n9929 = ~n4050 & ~n4054 ;
  assign n9930 = n9929 ^ n4039 ;
  assign n9931 = x541 & n9930 ;
  assign n9934 = n9933 ^ n9931 ;
  assign n9935 = x542 & n9934 ;
  assign n9936 = n9935 ^ n9933 ;
  assign n9937 = ~n4047 & ~n9936 ;
  assign n9912 = n4019 ^ n4017 ;
  assign n9894 = n4015 ^ x535 ;
  assign n9895 = n9894 ^ n4020 ;
  assign n9893 = n4015 ^ x536 ;
  assign n9896 = n9895 ^ n9893 ;
  assign n9910 = n4031 & n9896 ;
  assign n9913 = n9912 ^ n9910 ;
  assign n9914 = ~n4020 & n9913 ;
  assign n9916 = n4019 & n9894 ;
  assign n9917 = n9914 & n9916 ;
  assign n9911 = n9910 ^ n4031 ;
  assign n9915 = n9914 ^ n9911 ;
  assign n9918 = n9917 ^ n9915 ;
  assign n9923 = n9918 ^ n4015 ;
  assign n9924 = n9923 ^ n9893 ;
  assign n9938 = n9937 ^ n9924 ;
  assign n9976 = n9975 ^ n9938 ;
  assign n9864 = n4010 ^ x530 ;
  assign n9865 = n4007 ^ x529 ;
  assign n9866 = n9865 ^ n4010 ;
  assign n9867 = n9864 & ~n9866 ;
  assign n9868 = n9867 ^ n4011 ;
  assign n9869 = ~n4007 & n9868 ;
  assign n9870 = x529 & n9869 ;
  assign n9871 = n9867 ^ n4010 ;
  assign n9872 = n9871 ^ n9869 ;
  assign n9886 = n9870 & ~n9872 ;
  assign n9873 = n3995 ^ x524 ;
  assign n9874 = n3992 ^ x523 ;
  assign n9875 = n9874 ^ n3995 ;
  assign n9876 = n9873 & ~n9875 ;
  assign n9879 = n9876 ^ n3995 ;
  assign n9877 = n9876 ^ n3996 ;
  assign n9878 = ~n3992 & n9877 ;
  assign n9880 = n9879 ^ n9878 ;
  assign n9881 = x523 & n9878 ;
  assign n9882 = ~n9880 & n9881 ;
  assign n9883 = n9882 ^ n9880 ;
  assign n9884 = n9883 ^ n9872 ;
  assign n9887 = n9886 ^ n9884 ;
  assign n9861 = n3998 ^ n3979 ;
  assign n9862 = n4013 & ~n9861 ;
  assign n9863 = n9862 ^ n3998 ;
  assign n9888 = n9887 ^ n9863 ;
  assign n9857 = n3981 ^ n3971 ;
  assign n9858 = ~n3977 & ~n9857 ;
  assign n9859 = n9858 ^ n3981 ;
  assign n9820 = n3930 ^ x512 ;
  assign n9818 = n3930 ^ x511 ;
  assign n9819 = n9818 ^ n3932 ;
  assign n9821 = n9820 ^ n9819 ;
  assign n9841 = n3946 & n9821 ;
  assign n9826 = n9818 ^ n3940 ;
  assign n9831 = n9826 ^ n3930 ;
  assign n9834 = n9826 ^ n3932 ;
  assign n9835 = n9834 ^ x511 ;
  assign n9836 = n9831 & ~n9835 ;
  assign n9842 = n9841 ^ n9836 ;
  assign n9843 = n9842 ^ n9834 ;
  assign n9844 = n9841 ^ n9818 ;
  assign n9845 = n9844 ^ n9834 ;
  assign n9846 = n9843 & n9845 ;
  assign n9847 = ~n3932 & n9846 ;
  assign n9848 = n9847 ^ n9841 ;
  assign n9849 = n9848 ^ n3946 ;
  assign n9854 = n9849 ^ n3930 ;
  assign n9855 = n9854 ^ n9820 ;
  assign n9811 = n3952 ^ x518 ;
  assign n9790 = n3957 ^ n3953 ;
  assign n9796 = n9811 ^ n9790 ;
  assign n9800 = n1759 & n9796 ;
  assign n9794 = n3952 & ~n3956 ;
  assign n9801 = n9800 ^ n9794 ;
  assign n9787 = n3952 ^ x517 ;
  assign n9788 = n9787 ^ n3957 ;
  assign n9792 = n9788 ^ n3953 ;
  assign n9802 = n9801 ^ n9792 ;
  assign n9803 = n9800 ^ n9790 ;
  assign n9804 = n9803 ^ n9792 ;
  assign n9805 = n9802 & n9804 ;
  assign n9806 = ~n3953 & n9805 ;
  assign n9807 = n9806 ^ n9800 ;
  assign n9808 = n9807 ^ n1759 ;
  assign n9814 = n9808 ^ n3952 ;
  assign n9815 = n9814 ^ n9811 ;
  assign n9856 = n9855 ^ n9815 ;
  assign n9860 = n9859 ^ n9856 ;
  assign n9889 = n9888 ^ n9860 ;
  assign n9774 = ~n3977 & n3978 ;
  assign n9765 = n9764 ^ n3978 ;
  assign n9769 = n9768 ^ n9765 ;
  assign n9775 = n9774 ^ n9769 ;
  assign n9777 = n9774 ^ n3978 ;
  assign n9778 = ~n4013 & n9777 ;
  assign n9779 = n9778 ^ n3979 ;
  assign n9780 = n9779 ^ n4013 ;
  assign n9781 = ~n9775 & n9780 ;
  assign n9782 = n9781 ^ n9778 ;
  assign n9783 = n9782 ^ n9764 ;
  assign n9890 = n9889 ^ n9783 ;
  assign n9977 = n9976 ^ n9890 ;
  assign n9761 = n4122 ^ n3670 ;
  assign n9762 = ~n4123 & ~n9761 ;
  assign n9763 = n9762 ^ n4122 ;
  assign n9978 = n9977 ^ n9763 ;
  assign n9979 = n9978 ^ n9750 ;
  assign n9755 = ~n3928 & n4123 ;
  assign n9756 = n9755 ^ n9750 ;
  assign n9757 = n3673 & ~n9756 ;
  assign n9980 = n9979 ^ n9757 ;
  assign n9758 = ~n9748 & ~n9757 ;
  assign n9759 = n9750 ^ n3673 ;
  assign n9760 = n9758 & n9759 ;
  assign n9981 = n9980 ^ n9760 ;
  assign n10148 = n10147 ^ n9981 ;
  assign n9734 = n1663 & n1686 ;
  assign n9735 = n9734 ^ n9730 ;
  assign n9736 = n9735 & n9750 ;
  assign n9737 = n9736 ^ n9730 ;
  assign n9738 = n3668 & n9737 ;
  assign n9739 = n9738 ^ n3668 ;
  assign n9740 = n9750 ^ n3057 ;
  assign n9742 = ~n3668 & n9741 ;
  assign n9743 = n9750 ^ n9742 ;
  assign n9744 = ~n9740 & n9743 ;
  assign n9745 = n9750 ^ n9744 ;
  assign n9746 = ~n9739 & ~n9745 ;
  assign n10149 = n10148 ^ n9746 ;
  assign n10349 = n10348 ^ n10281 ;
  assign n11128 = n10349 ^ n10148 ;
  assign n11129 = n10149 & n11128 ;
  assign n11130 = n11129 ^ n10349 ;
  assign n11227 = n11226 ^ n11130 ;
  assign n11106 = n10080 ^ n3709 ;
  assign n11107 = n11106 ^ n10079 ;
  assign n11108 = n11107 ^ n10143 ;
  assign n11112 = n10143 ^ n10079 ;
  assign n11113 = ~n10144 & n11112 ;
  assign n11121 = ~n10143 & n11113 ;
  assign n11114 = n10119 ^ n10080 ;
  assign n11122 = n11121 ^ n11114 ;
  assign n11123 = ~n11108 & n11122 ;
  assign n11109 = n10118 ^ n10114 ;
  assign n11110 = n10115 & n11109 ;
  assign n11111 = n11110 ^ n10118 ;
  assign n11115 = n11114 ^ n11111 ;
  assign n11116 = n11115 ^ n11113 ;
  assign n11124 = n11123 ^ n11116 ;
  assign n11103 = n10145 ^ n9984 ;
  assign n11104 = n10146 & ~n11103 ;
  assign n11065 = ~n10008 & n10017 ;
  assign n11066 = n11065 ^ n10018 ;
  assign n11067 = n10073 ^ n10004 ;
  assign n11070 = n11067 ^ n10017 ;
  assign n11071 = n11070 ^ n10004 ;
  assign n11068 = n11067 ^ n10007 ;
  assign n11069 = n11068 ^ n10004 ;
  assign n11072 = n11071 ^ n11069 ;
  assign n11073 = n11072 ^ n11067 ;
  assign n11079 = ~n10018 & n11073 ;
  assign n11080 = n11079 ^ n11071 ;
  assign n11081 = n11073 ^ n11069 ;
  assign n11082 = n11081 ^ n11079 ;
  assign n11083 = n11082 ^ n11069 ;
  assign n11086 = ~n10004 & n11083 ;
  assign n11087 = n11086 ^ n11069 ;
  assign n11088 = n11080 & n11087 ;
  assign n11094 = ~n10004 & n10074 ;
  assign n11095 = n10007 & ~n10073 ;
  assign n11096 = ~n11094 & n11095 ;
  assign n11097 = n11096 ^ n11094 ;
  assign n11098 = ~n11088 & ~n11097 ;
  assign n11099 = n11066 & n11098 ;
  assign n11089 = n10063 ^ n10022 ;
  assign n11090 = ~n10072 & n11089 ;
  assign n11091 = n11090 ^ n10063 ;
  assign n11092 = n11091 ^ n11088 ;
  assign n11100 = n11099 ^ n11092 ;
  assign n11101 = n11100 ^ n10145 ;
  assign n11105 = n11104 ^ n11101 ;
  assign n11125 = n11124 ^ n11105 ;
  assign n11062 = n10147 ^ n9978 ;
  assign n11063 = n9981 & ~n11062 ;
  assign n11064 = n11063 ^ n10147 ;
  assign n11126 = n11125 ^ n11064 ;
  assign n11034 = ~n9924 & n9937 ;
  assign n11038 = n9975 & n11034 ;
  assign n11033 = ~n9950 & ~n9973 ;
  assign n11035 = n11034 ^ n9938 ;
  assign n11036 = n11033 & ~n11035 ;
  assign n11037 = ~n9947 & n11036 ;
  assign n11039 = n11038 ^ n11037 ;
  assign n11040 = n9971 ^ n9953 ;
  assign n11041 = n9972 & ~n11040 ;
  assign n11042 = n11041 ^ n9971 ;
  assign n11043 = n11033 ^ n9974 ;
  assign n11044 = n11043 ^ n11035 ;
  assign n11045 = n9947 & ~n11033 ;
  assign n11046 = n11045 ^ n11035 ;
  assign n11047 = ~n11044 & n11046 ;
  assign n11048 = n11047 ^ n11035 ;
  assign n11049 = n11042 & ~n11048 ;
  assign n11050 = ~n11039 & ~n11049 ;
  assign n11051 = n9973 & n11050 ;
  assign n11053 = n11038 & ~n11045 ;
  assign n11052 = n11035 & ~n11043 ;
  assign n11054 = n11053 ^ n11052 ;
  assign n11055 = n11054 ^ n11037 ;
  assign n11058 = n9947 & ~n11055 ;
  assign n11059 = n11051 & n11058 ;
  assign n11056 = n11055 ^ n11042 ;
  assign n11060 = n11059 ^ n11056 ;
  assign n11026 = n9883 ^ n9863 ;
  assign n11027 = n9887 & ~n11026 ;
  assign n11028 = n11027 ^ n9883 ;
  assign n11017 = n9888 ^ n9855 ;
  assign n11018 = ~n9856 & n11017 ;
  assign n11029 = n11028 ^ n11018 ;
  assign n11011 = n9859 ^ n9783 ;
  assign n11010 = n9783 & n9859 ;
  assign n11012 = n11011 ^ n11010 ;
  assign n11013 = n11012 ^ n9855 ;
  assign n11014 = n11013 ^ n9815 ;
  assign n11015 = n11014 ^ n9888 ;
  assign n11016 = n11012 ^ n9888 ;
  assign n11019 = n11018 ^ n11016 ;
  assign n11020 = n11019 ^ n11012 ;
  assign n11023 = n11010 & ~n11020 ;
  assign n11024 = n11023 ^ n11012 ;
  assign n11025 = ~n11015 & ~n11024 ;
  assign n11030 = n11029 ^ n11025 ;
  assign n11031 = n11030 ^ n9890 ;
  assign n11008 = n9890 ^ n9763 ;
  assign n11009 = n9977 & n11008 ;
  assign n11032 = n11031 ^ n11009 ;
  assign n11061 = n11060 ^ n11032 ;
  assign n11127 = n11126 ^ n11061 ;
  assign n11228 = n11227 ^ n11127 ;
  assign n11229 = n11228 ^ n10993 ;
  assign n11230 = n11229 ^ n11228 ;
  assign n10350 = n10349 ^ n10149 ;
  assign n11231 = n11230 ^ n10350 ;
  assign n11232 = n10995 & n11231 ;
  assign n11233 = n11232 ^ n11229 ;
  assign n12256 = n11149 & ~n11152 ;
  assign n12242 = n10271 ^ n10251 ;
  assign n12243 = n11133 & ~n12242 ;
  assign n12244 = n12243 ^ n10271 ;
  assign n12251 = n10271 ^ n10252 ;
  assign n12248 = n12247 ^ n10271 ;
  assign n12249 = n12245 & n12248 ;
  assign n12252 = n12251 ^ n12249 ;
  assign n12253 = n12244 & ~n12252 ;
  assign n12257 = n12256 ^ n12253 ;
  assign n12235 = n11189 ^ n11153 ;
  assign n12236 = n11158 & ~n12235 ;
  assign n12237 = n12236 ^ n11153 ;
  assign n12221 = n11189 ^ n11163 ;
  assign n12226 = ~n10190 & ~n10210 ;
  assign n12227 = n12226 ^ n12221 ;
  assign n12228 = ~n11161 & ~n12227 ;
  assign n12229 = ~n12221 & ~n12228 ;
  assign n12230 = n12221 ^ n11161 ;
  assign n12231 = n12230 ^ n12228 ;
  assign n12232 = n12231 ^ n11189 ;
  assign n12233 = n12229 & ~n12232 ;
  assign n12234 = n12233 ^ n12231 ;
  assign n12238 = n12237 ^ n12234 ;
  assign n12258 = n12257 ^ n12238 ;
  assign n12218 = n11222 ^ n11205 ;
  assign n12219 = n11223 & ~n12218 ;
  assign n12220 = n12219 ^ n11222 ;
  assign n12259 = n12258 ^ n12220 ;
  assign n12214 = n11193 ^ n11190 ;
  assign n12215 = n11225 & n12214 ;
  assign n12216 = n12215 ^ n11190 ;
  assign n12211 = n11215 & n11218 ;
  assign n12207 = ~n10292 & ~n10314 ;
  assign n12208 = n12207 ^ n11206 ;
  assign n12209 = n11208 & ~n12208 ;
  assign n12210 = n12209 ^ n11207 ;
  assign n12212 = n12211 ^ n12210 ;
  assign n12193 = n10344 ^ n10326 ;
  assign n12196 = ~n11194 & n12193 ;
  assign n12197 = n12196 ^ n10344 ;
  assign n12198 = n11203 & ~n12197 ;
  assign n12199 = n11205 & ~n12198 ;
  assign n12200 = n10334 & n12199 ;
  assign n12201 = ~n10327 & n12200 ;
  assign n12202 = n12201 ^ n12199 ;
  assign n12203 = n12202 ^ n12198 ;
  assign n12213 = n12212 ^ n12203 ;
  assign n12217 = n12216 ^ n12213 ;
  assign n12260 = n12259 ^ n12217 ;
  assign n12182 = ~n11065 & ~n11100 ;
  assign n12183 = ~n11091 & ~n11097 ;
  assign n12184 = ~n12182 & n12183 ;
  assign n12185 = n12184 ^ n12182 ;
  assign n12157 = n11124 ^ n10080 ;
  assign n12170 = n10079 & ~n12157 ;
  assign n12171 = ~n10119 & n11124 ;
  assign n12172 = n10145 & n12171 ;
  assign n12173 = n12172 ^ n10080 ;
  assign n12174 = n12170 & n12173 ;
  assign n12175 = n12174 ^ n12172 ;
  assign n12186 = n12185 ^ n12175 ;
  assign n12156 = n11124 ^ n11111 ;
  assign n12162 = ~n10079 & n10119 ;
  assign n12163 = n12162 ^ n12157 ;
  assign n12164 = n11111 & ~n12163 ;
  assign n12165 = n12164 ^ n12157 ;
  assign n12166 = ~n12164 & ~n12165 ;
  assign n12167 = ~n12156 & n12166 ;
  assign n12168 = n12167 ^ n12165 ;
  assign n12176 = n12168 ^ n11111 ;
  assign n12177 = n12176 ^ n3709 ;
  assign n12178 = n10144 & n12177 ;
  assign n12179 = n12178 ^ n3709 ;
  assign n12180 = ~n12175 & ~n12179 ;
  assign n12187 = n12186 ^ n12180 ;
  assign n12169 = ~n11111 & n12168 ;
  assign n12181 = n12169 & n12180 ;
  assign n12188 = n12187 ^ n12181 ;
  assign n12153 = n11124 ^ n11100 ;
  assign n12154 = ~n11105 & n12153 ;
  assign n12155 = n12154 ^ n11124 ;
  assign n12189 = n12188 ^ n12155 ;
  assign n12141 = n9815 & n9855 ;
  assign n12142 = ~n11030 & n12141 ;
  assign n12143 = n12142 ^ n11030 ;
  assign n12144 = ~n11028 & n12143 ;
  assign n12145 = n11012 & n12144 ;
  assign n12146 = ~n9888 & n12145 ;
  assign n12147 = n12146 ^ n12144 ;
  assign n12148 = n12147 ^ n12143 ;
  assign n12149 = n12148 ^ n11050 ;
  assign n12138 = n11060 ^ n11030 ;
  assign n12139 = ~n11032 & ~n12138 ;
  assign n12140 = n12139 ^ n11060 ;
  assign n12150 = n12149 ^ n12140 ;
  assign n12151 = n12150 ^ n11061 ;
  assign n12136 = n11064 ^ n11061 ;
  assign n12137 = n11126 & n12136 ;
  assign n12152 = n12151 ^ n12137 ;
  assign n12190 = n12189 ^ n12152 ;
  assign n12191 = n12190 ^ n11127 ;
  assign n12134 = n11130 ^ n11127 ;
  assign n12135 = n11227 & n12134 ;
  assign n12192 = n12191 ^ n12135 ;
  assign n12261 = n12260 ^ n12192 ;
  assign n12263 = n12261 ^ n11228 ;
  assign n11441 = ~n10523 & ~n10530 ;
  assign n11443 = n11441 ^ n10531 ;
  assign n11450 = n11443 ^ n10553 ;
  assign n11444 = ~n10553 & n11443 ;
  assign n11451 = n11450 ^ n11444 ;
  assign n11452 = ~n10573 & ~n11451 ;
  assign n11453 = ~n10549 & ~n11452 ;
  assign n11437 = n10548 ^ n10544 ;
  assign n11438 = ~n10545 & n11437 ;
  assign n11439 = n11438 ^ n10544 ;
  assign n11442 = ~n10574 & n11441 ;
  assign n11457 = ~n11439 & ~n11442 ;
  assign n11458 = ~n11444 & n11457 ;
  assign n11459 = n11453 & n11458 ;
  assign n11460 = n11459 ^ n11457 ;
  assign n11461 = n11460 ^ n11442 ;
  assign n11462 = n11453 & n11461 ;
  assign n11445 = ~n10573 & ~n11442 ;
  assign n11446 = n11444 & n11445 ;
  assign n11447 = n10549 & n11446 ;
  assign n11448 = n11447 ^ n11445 ;
  assign n11449 = n11448 ^ n10573 ;
  assign n11454 = n11453 ^ n11449 ;
  assign n11455 = ~n11442 & n11454 ;
  assign n11418 = n10597 ^ n10584 ;
  assign n11434 = n10646 & n11418 ;
  assign n11427 = n10595 & ~n10596 ;
  assign n11420 = n10597 ^ n2561 ;
  assign n11419 = n10597 ^ n2553 ;
  assign n11421 = n11420 ^ n11419 ;
  assign n11424 = n2559 & n11421 ;
  assign n11425 = n11424 ^ n11420 ;
  assign n11426 = n10584 & n11425 ;
  assign n11428 = n11427 ^ n11426 ;
  assign n11435 = n11434 ^ n11428 ;
  assign n11415 = n10645 ^ n10638 ;
  assign n11416 = ~n10642 & ~n11415 ;
  assign n11417 = n11416 ^ n10645 ;
  assign n11436 = n11435 ^ n11417 ;
  assign n11440 = n11439 ^ n11436 ;
  assign n11456 = n11455 ^ n11440 ;
  assign n11463 = n11462 ^ n11456 ;
  assign n11412 = n10648 ^ n10574 ;
  assign n11413 = ~n10576 & n11412 ;
  assign n11414 = n11413 ^ n10574 ;
  assign n11464 = n11463 ^ n11414 ;
  assign n11388 = ~n10366 & n10433 ;
  assign n11390 = n11388 ^ n10434 ;
  assign n11391 = n10437 & ~n11390 ;
  assign n11389 = ~n10438 & ~n10439 ;
  assign n11397 = n11389 ^ n11388 ;
  assign n11398 = n11389 ^ n10440 ;
  assign n11399 = n10442 & n11398 ;
  assign n11402 = n11397 & n11399 ;
  assign n11403 = n11402 ^ n11389 ;
  assign n11404 = ~n11391 & ~n11403 ;
  assign n11405 = n11404 ^ n11399 ;
  assign n11394 = n10431 ^ n10369 ;
  assign n11395 = ~n10432 & ~n11394 ;
  assign n11396 = n11395 ^ n10369 ;
  assign n11406 = n11405 ^ n11396 ;
  assign n11392 = ~n11389 & ~n11391 ;
  assign n11393 = n11388 & n11392 ;
  assign n11408 = n11406 ^ n11393 ;
  assign n12324 = n10504 ^ n10492 ;
  assign n10485 = n10484 ^ n10477 ;
  assign n11359 = n11346 ^ n10484 ;
  assign n11351 = n11346 ^ n10504 ;
  assign n11358 = ~n11344 & ~n11351 ;
  assign n11360 = n11359 ^ n11358 ;
  assign n11361 = ~n10485 & n11360 ;
  assign n11362 = n11361 ^ n10492 ;
  assign n11363 = n11346 & ~n11362 ;
  assign n11364 = n11358 ^ n10505 ;
  assign n11365 = n11364 ^ n11361 ;
  assign n11366 = n11363 & ~n11365 ;
  assign n11367 = n11366 ^ n11361 ;
  assign n11357 = n12324 ^ n11344 ;
  assign n11368 = n11367 ^ n11357 ;
  assign n11369 = n11368 ^ n10504 ;
  assign n11381 = n12324 ^ n11369 ;
  assign n11331 = n10490 ^ n10488 ;
  assign n11332 = n10491 & ~n11331 ;
  assign n11333 = n11332 ^ n10490 ;
  assign n11382 = n11381 ^ n11333 ;
  assign n11384 = n11382 ^ n10442 ;
  assign n11383 = n11382 ^ n11346 ;
  assign n11385 = n11384 ^ n11383 ;
  assign n11386 = n10447 & n11385 ;
  assign n11387 = n11386 ^ n11384 ;
  assign n11409 = n11408 ^ n11387 ;
  assign n11410 = n11409 ^ n10507 ;
  assign n11329 = n10510 ^ n10507 ;
  assign n11330 = ~n10650 & ~n11329 ;
  assign n11411 = n11410 ^ n11330 ;
  assign n11465 = n11464 ^ n11411 ;
  assign n11319 = n10980 ^ n10955 ;
  assign n11320 = n10981 & ~n11319 ;
  assign n11321 = n11320 ^ n10980 ;
  assign n11304 = n10986 ^ n10950 ;
  assign n11308 = n10950 ^ n10931 ;
  assign n11309 = n11304 & ~n11308 ;
  assign n11315 = ~n10950 & n11309 ;
  assign n11307 = n10982 ^ n10939 ;
  assign n11310 = n11309 ^ n11307 ;
  assign n11316 = n11315 ^ n11310 ;
  assign n12295 = n11304 ^ n10939 ;
  assign n12296 = n12295 ^ n10931 ;
  assign n11317 = n11316 & ~n12296 ;
  assign n11318 = n11317 ^ n11310 ;
  assign n11322 = n11321 ^ n11318 ;
  assign n11323 = n11322 ^ n10927 ;
  assign n11302 = n10930 ^ n10927 ;
  assign n11303 = ~n10988 & n11302 ;
  assign n11324 = n11323 ^ n11303 ;
  assign n11293 = n10925 ^ n10879 ;
  assign n11294 = n10926 & n11293 ;
  assign n11295 = n11294 ^ n10925 ;
  assign n11289 = n10915 ^ n10887 ;
  assign n11290 = ~n10924 & ~n11289 ;
  assign n11291 = n11290 ^ n10915 ;
  assign n12285 = n11295 ^ n11291 ;
  assign n12286 = n12285 ^ n10867 ;
  assign n11287 = n10926 ^ n10879 ;
  assign n11288 = n11287 ^ n10866 ;
  assign n11300 = n10868 & n11288 ;
  assign n11301 = n12286 ^ n11300 ;
  assign n11325 = n11324 ^ n11301 ;
  assign n11280 = n10814 ^ n2364 ;
  assign n11281 = ~n10818 & ~n11280 ;
  assign n11282 = n11281 ^ n2364 ;
  assign n11272 = n10861 ^ n10811 ;
  assign n11273 = n10819 & n11272 ;
  assign n11274 = n10859 ^ n10827 ;
  assign n11275 = n10859 ^ n10811 ;
  assign n11276 = n11274 & n11275 ;
  assign n11277 = n11276 ^ n10859 ;
  assign n11278 = n11273 & n11277 ;
  assign n11258 = n10859 ^ n10819 ;
  assign n11259 = n10860 & n11258 ;
  assign n11260 = n11259 ^ n10859 ;
  assign n11266 = n11258 ^ n10860 ;
  assign n11267 = n11266 ^ n10859 ;
  assign n11261 = n10827 ^ n10811 ;
  assign n11262 = n10827 ^ n10819 ;
  assign n11263 = n11262 ^ n10856 ;
  assign n11264 = n11263 ^ n10859 ;
  assign n11265 = ~n11261 & n11264 ;
  assign n11268 = n11267 ^ n11265 ;
  assign n11269 = ~n11260 & ~n11268 ;
  assign n11279 = n11278 ^ n11269 ;
  assign n11283 = n11282 ^ n11279 ;
  assign n11241 = n10795 ^ n10664 ;
  assign n11243 = n10793 ^ n10733 ;
  assign n11244 = ~n10794 & ~n11243 ;
  assign n11245 = n11244 ^ n10793 ;
  assign n11248 = n10664 & ~n11245 ;
  assign n11249 = n11248 ^ n10729 ;
  assign n11250 = ~n11241 & ~n11249 ;
  assign n11246 = n11245 ^ n10729 ;
  assign n11251 = n11250 ^ n11246 ;
  assign n11238 = n10727 ^ n10667 ;
  assign n11239 = ~n10728 & n11238 ;
  assign n11240 = n11239 ^ n10727 ;
  assign n11252 = n11251 ^ n11240 ;
  assign n11254 = n11252 ^ n10796 ;
  assign n11253 = n11252 ^ n10862 ;
  assign n11255 = n11254 ^ n11253 ;
  assign n11256 = ~n10801 & ~n11255 ;
  assign n11257 = n11256 ^ n11254 ;
  assign n11284 = n11283 ^ n11257 ;
  assign n11285 = n11284 ^ n10863 ;
  assign n11236 = n10863 ^ n10656 ;
  assign n11237 = ~n10990 & n11236 ;
  assign n11286 = n11285 ^ n11237 ;
  assign n11326 = n11325 ^ n11286 ;
  assign n11327 = n11326 ^ n10651 ;
  assign n11234 = n10651 ^ n10363 ;
  assign n11235 = ~n10992 & n11234 ;
  assign n11328 = n11327 ^ n11235 ;
  assign n11466 = n11465 ^ n11328 ;
  assign n12262 = n12261 ^ n11466 ;
  assign n12264 = n12263 ^ n12262 ;
  assign n12265 = n11233 & n12264 ;
  assign n12266 = n12265 ^ n12263 ;
  assign n12337 = n11392 & ~n11399 ;
  assign n12336 = ~n11396 & ~n11405 ;
  assign n12338 = n12337 ^ n12336 ;
  assign n12320 = n11408 ^ n11382 ;
  assign n12321 = ~n11387 & ~n12320 ;
  assign n12322 = n12321 ^ n11382 ;
  assign n12775 = n12338 ^ n12322 ;
  assign n12323 = ~n10505 & ~n11343 ;
  assign n12325 = n12324 ^ n12323 ;
  assign n12326 = n11333 & ~n12325 ;
  assign n12327 = ~n10504 & n12326 ;
  assign n12328 = ~n12323 & n12327 ;
  assign n12329 = n12328 ^ n12326 ;
  assign n12330 = n12329 ^ n11333 ;
  assign n12331 = n11382 & ~n12330 ;
  assign n12332 = n10484 & n12331 ;
  assign n12333 = n10477 & n12332 ;
  assign n12334 = n12333 ^ n12331 ;
  assign n12335 = n12334 ^ n12330 ;
  assign n12776 = n12335 ^ n12322 ;
  assign n12777 = ~n12775 & n12776 ;
  assign n12778 = n12777 ^ n12338 ;
  assign n12339 = n12338 ^ n12335 ;
  assign n12340 = n12339 ^ n12322 ;
  assign n12779 = n12778 ^ n12340 ;
  assign n12350 = n11449 & ~n11461 ;
  assign n12346 = n11427 ^ n10597 ;
  assign n12347 = ~n10646 & n11428 ;
  assign n12348 = ~n12346 & n12347 ;
  assign n12345 = ~n11417 & ~n11435 ;
  assign n12349 = n12348 ^ n12345 ;
  assign n12351 = n12350 ^ n12349 ;
  assign n12342 = n11464 ^ n11409 ;
  assign n12343 = n11411 & ~n12342 ;
  assign n12344 = n12343 ^ n11464 ;
  assign n12317 = n11436 ^ n11414 ;
  assign n12318 = n11463 & ~n12317 ;
  assign n12319 = n12318 ^ n11436 ;
  assign n12765 = n12349 ^ n12319 ;
  assign n12766 = n12765 ^ n12349 ;
  assign n12769 = ~n12344 & n12766 ;
  assign n12770 = n12340 & n12769 ;
  assign n12771 = n12770 ^ n12340 ;
  assign n12763 = n12349 ^ n12340 ;
  assign n12772 = n12771 ^ n12763 ;
  assign n12773 = n12351 & ~n12772 ;
  assign n12774 = n12773 ^ n12350 ;
  assign n12780 = n12779 ^ n12774 ;
  assign n12758 = ~n12349 & ~n12350 ;
  assign n12759 = ~n12340 & n12758 ;
  assign n12760 = n12344 & n12759 ;
  assign n12761 = n12760 ^ n12759 ;
  assign n12762 = n12319 & n12761 ;
  assign n12781 = n12780 ^ n12762 ;
  assign n12754 = n12351 ^ n12340 ;
  assign n12755 = ~n12319 & n12344 ;
  assign n12756 = n12755 ^ n12340 ;
  assign n12757 = n12754 & ~n12756 ;
  assign n12782 = n12781 ^ n12757 ;
  assign n12352 = n12351 ^ n12344 ;
  assign n12341 = n12340 ^ n12319 ;
  assign n12353 = n12352 ^ n12341 ;
  assign n12311 = n11322 ^ n11301 ;
  assign n12312 = n11324 & ~n12311 ;
  assign n12313 = n12312 ^ n11322 ;
  assign n12290 = ~n10866 & ~n10867 ;
  assign n12291 = n12290 ^ n12285 ;
  assign n12292 = ~n11301 & ~n12291 ;
  assign n12293 = n11301 ^ n11295 ;
  assign n12294 = ~n12292 & ~n12293 ;
  assign n12301 = ~n11318 & ~n11321 ;
  assign n12297 = n10982 & n12296 ;
  assign n12298 = ~n10951 & n11308 ;
  assign n12299 = n12298 ^ n10950 ;
  assign n12300 = n12297 & n12299 ;
  assign n12302 = n12301 ^ n12300 ;
  assign n12304 = n12302 ^ n11291 ;
  assign n12305 = n12304 ^ n11295 ;
  assign n12306 = n12305 ^ n11301 ;
  assign n12307 = n12306 ^ n12292 ;
  assign n12303 = n12302 ^ n11301 ;
  assign n12308 = n12307 ^ n12303 ;
  assign n12309 = n12294 & ~n12308 ;
  assign n12310 = n12309 ^ n12307 ;
  assign n12314 = n12313 ^ n12310 ;
  assign n12281 = n11283 ^ n11252 ;
  assign n12282 = n11257 & n12281 ;
  assign n12283 = n12282 ^ n11252 ;
  assign n12278 = n11245 ^ n11240 ;
  assign n12279 = ~n11251 & n12278 ;
  assign n12273 = ~n11278 & ~n11282 ;
  assign n12274 = ~n11269 & n12273 ;
  assign n12275 = n12274 ^ n11269 ;
  assign n12276 = n12275 ^ n11245 ;
  assign n12280 = n12279 ^ n12276 ;
  assign n12284 = n12283 ^ n12280 ;
  assign n12315 = n12314 ^ n12284 ;
  assign n12270 = n11325 ^ n11284 ;
  assign n12271 = ~n11286 & n12270 ;
  assign n12272 = n12271 ^ n11325 ;
  assign n12316 = n12315 ^ n12272 ;
  assign n12354 = n12353 ^ n12316 ;
  assign n12267 = n11465 ^ n11326 ;
  assign n12268 = ~n11328 & ~n12267 ;
  assign n12269 = n12268 ^ n11465 ;
  assign n12751 = n12316 ^ n12269 ;
  assign n12752 = ~n12354 & ~n12751 ;
  assign n12753 = n12752 ^ n12353 ;
  assign n12783 = n12782 ^ n12753 ;
  assign n12747 = n12284 ^ n12272 ;
  assign n12748 = ~n12315 & ~n12747 ;
  assign n12749 = n12748 ^ n12284 ;
  assign n12743 = n12283 ^ n12275 ;
  assign n12744 = ~n12280 & n12743 ;
  assign n12745 = n12744 ^ n12275 ;
  assign n12740 = n12313 ^ n12302 ;
  assign n12741 = ~n12310 & n12740 ;
  assign n12742 = n12741 ^ n12302 ;
  assign n12746 = n12745 ^ n12742 ;
  assign n12750 = n12749 ^ n12746 ;
  assign n12784 = n12783 ^ n12750 ;
  assign n12786 = n12784 ^ n12261 ;
  assign n12355 = n12354 ^ n12269 ;
  assign n12785 = n12784 ^ n12355 ;
  assign n12787 = n12786 ^ n12785 ;
  assign n12788 = ~n12266 & n12787 ;
  assign n12789 = n12788 ^ n12786 ;
  assign n13072 = n12782 ^ n12742 ;
  assign n13073 = n12746 & ~n13072 ;
  assign n13067 = n12753 ^ n12749 ;
  assign n13068 = n12782 ^ n12746 ;
  assign n13069 = n13068 ^ n12753 ;
  assign n13070 = n13067 & ~n13069 ;
  assign n13052 = ~n12322 & n12338 ;
  assign n13053 = n12335 & ~n12760 ;
  assign n13054 = n13052 & n13053 ;
  assign n13055 = n13054 ^ n12760 ;
  assign n13056 = ~n12353 & ~n13055 ;
  assign n13057 = ~n12319 & ~n12774 ;
  assign n13058 = n13056 & n13057 ;
  assign n13059 = n13058 ^ n13055 ;
  assign n13060 = n12778 & ~n13059 ;
  assign n13061 = n12774 & n13060 ;
  assign n13062 = ~n12755 & n13061 ;
  assign n13063 = n13062 ^ n13060 ;
  assign n13064 = n13063 ^ n13059 ;
  assign n13065 = n13064 ^ n12742 ;
  assign n13066 = n13065 ^ n12745 ;
  assign n13071 = n13070 ^ n13066 ;
  assign n13074 = n13073 ^ n13071 ;
  assign n13075 = n13074 ^ n13065 ;
  assign n13076 = n13070 & n13073 ;
  assign n13077 = ~n13075 & n13076 ;
  assign n13078 = n13077 ^ n13074 ;
  assign n13080 = n13078 ^ n12784 ;
  assign n12806 = n12220 ^ n12212 ;
  assign n12807 = n12806 ^ n12216 ;
  assign n12808 = n12807 ^ n12203 ;
  assign n12814 = n12216 ^ n12212 ;
  assign n12815 = ~n12213 & ~n12814 ;
  assign n12821 = ~n12203 & n12815 ;
  assign n12822 = n12821 ^ n12259 ;
  assign n12823 = ~n12808 & n12822 ;
  assign n12810 = n12234 & ~n12237 ;
  assign n12809 = ~n12238 & n12257 ;
  assign n12811 = n12810 ^ n12809 ;
  assign n12812 = n12811 ^ n12259 ;
  assign n12816 = n12815 ^ n12812 ;
  assign n12824 = n12823 ^ n12816 ;
  assign n12800 = n12185 ^ n12155 ;
  assign n12801 = ~n12188 & n12800 ;
  assign n12802 = n12801 ^ n12185 ;
  assign n12796 = n12140 ^ n11050 ;
  assign n12797 = n12148 ^ n12140 ;
  assign n12798 = n12796 & ~n12797 ;
  assign n12799 = n12798 ^ n11050 ;
  assign n12803 = n12802 ^ n12799 ;
  assign n12793 = n12189 ^ n12150 ;
  assign n12794 = ~n12152 & n12793 ;
  assign n12795 = n12794 ^ n12189 ;
  assign n12804 = n12803 ^ n12795 ;
  assign n12790 = n12260 ^ n12190 ;
  assign n12791 = n12192 & n12790 ;
  assign n12792 = n12791 ^ n12260 ;
  assign n12805 = n12804 ^ n12792 ;
  assign n12825 = n12824 ^ n12805 ;
  assign n13079 = n13078 ^ n12825 ;
  assign n13081 = n13080 ^ n13079 ;
  assign n13082 = n12789 & n13081 ;
  assign n13083 = n13082 ^ n13080 ;
  assign n13084 = ~n12799 & n12802 ;
  assign n13085 = ~n12795 & n13084 ;
  assign n13086 = ~n12260 & n12811 ;
  assign n13087 = n12216 & n13086 ;
  assign n13088 = n12220 & n13087 ;
  assign n13089 = n13088 ^ n13086 ;
  assign n13090 = n13089 ^ n12811 ;
  assign n13091 = n12824 & ~n13090 ;
  assign n13092 = ~n12212 & n13091 ;
  assign n13093 = ~n12203 & n13092 ;
  assign n13094 = n13093 ^ n13091 ;
  assign n13095 = n13094 ^ n13090 ;
  assign n13096 = ~n13085 & ~n13095 ;
  assign n13097 = n13096 ^ n13095 ;
  assign n13112 = n12802 ^ n12795 ;
  assign n13113 = n12803 & ~n13112 ;
  assign n13114 = n13113 ^ n12795 ;
  assign n13115 = ~n12792 & ~n13114 ;
  assign n13116 = ~n13085 & ~n13115 ;
  assign n13098 = n12258 ^ n12216 ;
  assign n13099 = n12814 & ~n13098 ;
  assign n13100 = n13099 ^ n12216 ;
  assign n13106 = n13098 ^ n12814 ;
  assign n13107 = n13106 ^ n12216 ;
  assign n13101 = n12220 ^ n12203 ;
  assign n13102 = n12258 ^ n12203 ;
  assign n13103 = n13102 ^ n12212 ;
  assign n13104 = n13103 ^ n12216 ;
  assign n13105 = ~n13101 & ~n13104 ;
  assign n13108 = n13107 ^ n13105 ;
  assign n13109 = n13100 & ~n13108 ;
  assign n13117 = n13116 ^ n13109 ;
  assign n13118 = ~n12824 & ~n13117 ;
  assign n13119 = n13085 ^ n12803 ;
  assign n13120 = n13119 ^ n13113 ;
  assign n13121 = n13114 ^ n12792 ;
  assign n13122 = n13121 ^ n13115 ;
  assign n13123 = n13095 & n13122 ;
  assign n13124 = n13120 & n13123 ;
  assign n13125 = n13124 ^ n13122 ;
  assign n13126 = n12824 & ~n13120 ;
  assign n13127 = n13096 ^ n13085 ;
  assign n13128 = ~n12792 & n13127 ;
  assign n13129 = n13126 & n13128 ;
  assign n13130 = n13129 ^ n12824 ;
  assign n13131 = n13125 & n13130 ;
  assign n13132 = ~n13118 & ~n13131 ;
  assign n13133 = n13097 & n13132 ;
  assign n13245 = n13133 ^ n13078 ;
  assign n13246 = n13083 & ~n13245 ;
  assign n13247 = n13246 ^ n13133 ;
  assign n13217 = n12749 ^ n12745 ;
  assign n13216 = ~n12745 & n12749 ;
  assign n13218 = n13217 ^ n13216 ;
  assign n13219 = n13218 ^ n13064 ;
  assign n13220 = n12782 & n13219 ;
  assign n13221 = n13064 & n13220 ;
  assign n13222 = n13221 ^ n13219 ;
  assign n13223 = n13065 ^ n12783 ;
  assign n13224 = n13223 ^ n13219 ;
  assign n13225 = n13222 & n13224 ;
  assign n13226 = n13065 & n13225 ;
  assign n13227 = n13226 ^ n13221 ;
  assign n13228 = n13227 ^ n13218 ;
  assign n13229 = n12753 & ~n13216 ;
  assign n13230 = n13064 & n13229 ;
  assign n13231 = n13230 ^ n13216 ;
  assign n13232 = n13230 ^ n12783 ;
  assign n13233 = n13230 ^ n12742 ;
  assign n13234 = n13233 ^ n13230 ;
  assign n13235 = ~n13232 & ~n13234 ;
  assign n13236 = ~n13231 & n13235 ;
  assign n13237 = n13236 ^ n13231 ;
  assign n13238 = n13237 ^ n13216 ;
  assign n13239 = ~n13228 & ~n13238 ;
  assign n13240 = n13239 ^ n13118 ;
  assign n13241 = n13240 ^ n13239 ;
  assign n13242 = ~n13096 & n13125 ;
  assign n13243 = ~n13241 & n13242 ;
  assign n13244 = n13243 ^ n13240 ;
  assign n13248 = n13247 ^ n13244 ;
  assign n13343 = n13342 ^ n13248 ;
  assign n13212 = n13211 ^ n13181 ;
  assign n13351 = n13342 ^ n13212 ;
  assign n13134 = n13133 ^ n13083 ;
  assign n13213 = n13212 ^ n13134 ;
  assign n13352 = n13351 ^ n13213 ;
  assign n13353 = n13352 ^ n13351 ;
  assign n13045 = n13044 ^ n12983 ;
  assign n12826 = n12825 ^ n12789 ;
  assign n13046 = n13045 ^ n12826 ;
  assign n12356 = n12355 ^ n12266 ;
  assign n12123 = n12122 ^ n11757 ;
  assign n12357 = n12356 ^ n12123 ;
  assign n11467 = n11466 ^ n11233 ;
  assign n12124 = n12123 ^ n11467 ;
  assign n10996 = n10995 ^ n10350 ;
  assign n12131 = n12123 ^ n10996 ;
  assign n9729 = n9728 ^ n8976 ;
  assign n10997 = n10996 ^ n9729 ;
  assign n4129 = n4128 ^ n4127 ;
  assign n4131 = n4130 ^ n4129 ;
  assign n5416 = n5415 ^ n4131 ;
  assign n7942 = n7941 ^ n5416 ;
  assign n4126 = n4125 ^ n3048 ;
  assign n7943 = n7942 ^ n4126 ;
  assign n1384 = n1383 ^ n1192 ;
  assign n1616 = n1615 ^ n1384 ;
  assign n10998 = n4126 ^ n1616 ;
  assign n10999 = n10998 ^ n4126 ;
  assign n1999 = n1998 ^ n1807 ;
  assign n11000 = n4126 ^ n1999 ;
  assign n11001 = n11000 ^ n4126 ;
  assign n11002 = n10999 & n11001 ;
  assign n11003 = n11002 ^ n4126 ;
  assign n11004 = ~n7943 & n11003 ;
  assign n11005 = n11004 ^ n7942 ;
  assign n11006 = n11005 ^ n9729 ;
  assign n11007 = ~n10997 & n11006 ;
  assign n12132 = n12131 ^ n11007 ;
  assign n12133 = ~n12124 & ~n12132 ;
  assign n12358 = n12357 ^ n12133 ;
  assign n12734 = n12733 ^ n12535 ;
  assign n12737 = n12734 ^ n12356 ;
  assign n12738 = n12358 & n12737 ;
  assign n12739 = n12738 ^ n12734 ;
  assign n13049 = n12826 ^ n12739 ;
  assign n13050 = n13046 & n13049 ;
  assign n13051 = n13050 ^ n13045 ;
  assign n13354 = n13248 ^ n13051 ;
  assign n13355 = n13354 ^ n13351 ;
  assign n13356 = n13353 & n13355 ;
  assign n13357 = n13356 ^ n13351 ;
  assign n13358 = n13343 & n13357 ;
  assign n13359 = n13358 ^ n13342 ;
  assign n2000 = n1999 ^ n1616 ;
  assign n7944 = n7943 ^ n1616 ;
  assign n7945 = ~x1000 & n7944 ;
  assign n7946 = ~n2000 & n7945 ;
  assign n12125 = n12124 ^ n10996 ;
  assign n12126 = n12125 ^ n11007 ;
  assign n12127 = ~n7946 & n12126 ;
  assign n12128 = n11005 ^ n10997 ;
  assign n12129 = n12127 & ~n12128 ;
  assign n12130 = n12129 ^ n12126 ;
  assign n12735 = n12734 ^ n12358 ;
  assign n12736 = ~n12130 & ~n12735 ;
  assign n13047 = n13046 ^ n12739 ;
  assign n13048 = n12736 & n13047 ;
  assign n13214 = n13213 ^ n13051 ;
  assign n13215 = n13048 & ~n13214 ;
  assign n13344 = n13343 ^ n13212 ;
  assign n13345 = n13344 ^ n13343 ;
  assign n13346 = n13343 ^ n13051 ;
  assign n13347 = n13346 ^ n13343 ;
  assign n13348 = n13345 & ~n13347 ;
  assign n13349 = n13348 ^ n13343 ;
  assign n13350 = n13215 & n13349 ;
  assign n13360 = n13359 ^ n13350 ;
  assign n13370 = n13148 ^ n13144 ;
  assign n13371 = n13180 & n13370 ;
  assign n13369 = n13268 ^ n13144 ;
  assign n13372 = n13371 ^ n13369 ;
  assign n13374 = ~n13137 & ~n13140 ;
  assign n13373 = n13268 ^ n13141 ;
  assign n13375 = n13374 ^ n13373 ;
  assign n13376 = ~n13372 & ~n13375 ;
  assign n13377 = n13376 ^ n13268 ;
  assign n13380 = n13268 ^ n13180 ;
  assign n13381 = n13380 ^ n13268 ;
  assign n13382 = n13369 ^ n13268 ;
  assign n13383 = n13382 ^ n13268 ;
  assign n13384 = n13381 & ~n13383 ;
  assign n13385 = ~n13370 & n13384 ;
  assign n13386 = n13385 ^ n13370 ;
  assign n13378 = n13370 ^ n13268 ;
  assign n13387 = n13386 ^ n13378 ;
  assign n13388 = ~n13374 & n13387 ;
  assign n13389 = ~n13377 & ~n13388 ;
  assign n13361 = n13341 ^ n13252 ;
  assign n13362 = ~n13260 & n13361 ;
  assign n13363 = n13362 ^ n13341 ;
  assign n13365 = n13363 ^ n13247 ;
  assign n13364 = n13363 ^ n13239 ;
  assign n13366 = n13365 ^ n13364 ;
  assign n13367 = n13244 & ~n13366 ;
  assign n13368 = n13367 ^ n13365 ;
  assign n13390 = n13389 ^ n13368 ;
  assign n13391 = n13390 ^ n13359 ;
  assign n13392 = ~n13360 & ~n13391 ;
  assign n13393 = n13392 ^ n13390 ;
  assign n13394 = n13392 ^ n13363 ;
  assign n13397 = ~n13368 & ~n13394 ;
  assign n13398 = n13397 ^ n13363 ;
  assign n13399 = n13393 & ~n13398 ;
  assign y0 = ~n13399 ;
endmodule
