module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n61 = x6 & x7 ;
  assign n62 = x0 & x1 ;
  assign n63 = x2 & x3 ;
  assign n64 = x4 & x5 ;
  assign n65 = n63 & n64 ;
  assign n66 = n62 & n65 ;
  assign n67 = x8 & n66 ;
  assign n68 = n61 & n67 ;
  assign n69 = ~x9 & ~n68 ;
  assign n70 = ~x26 & ~n69 ;
  assign n71 = ~x5 & ~x6 ;
  assign n72 = ~x7 & ~x8 ;
  assign n73 = n71 & n72 ;
  assign n74 = ~x1 & ~x2 ;
  assign n75 = ~x3 & ~x4 ;
  assign n76 = n74 & n75 ;
  assign n77 = n73 & n76 ;
  assign n78 = x9 & ~n77 ;
  assign n79 = x14 & x15 ;
  assign n80 = ~x12 & ~x13 ;
  assign n81 = n79 & ~n80 ;
  assign n82 = ~x21 & ~x22 ;
  assign n83 = ~x16 & ~x18 ;
  assign n84 = n82 & n83 ;
  assign n85 = ~n81 & n84 ;
  assign n86 = ~x10 & n85 ;
  assign n87 = ~n78 & n86 ;
  assign n88 = x11 & n79 ;
  assign n89 = n85 & ~n88 ;
  assign n90 = ~x17 & ~x18 ;
  assign n91 = x19 & x20 ;
  assign n92 = ~n90 & n91 ;
  assign n93 = n82 & ~n92 ;
  assign n94 = x27 & x28 ;
  assign n95 = x29 & n94 ;
  assign n96 = x23 & x24 ;
  assign n97 = x25 & n96 ;
  assign n98 = n95 & n97 ;
  assign n99 = ~n93 & n98 ;
  assign n100 = ~n89 & n99 ;
  assign n101 = n87 & n100 ;
  assign n102 = n70 & n101 ;
  assign n103 = x26 & n95 ;
  assign n104 = x57 & x58 ;
  assign n105 = x59 & n104 ;
  assign n106 = x53 & x54 ;
  assign n107 = x55 & n106 ;
  assign n108 = x49 & x50 ;
  assign n109 = x46 & x47 ;
  assign n110 = ~x48 & ~n109 ;
  assign n111 = n108 & ~n110 ;
  assign n112 = ~x51 & ~x52 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = n107 & ~n113 ;
  assign n115 = ~x56 & ~n114 ;
  assign n116 = ~x37 & ~x38 ;
  assign n117 = ~x31 & ~x36 ;
  assign n118 = n116 & n117 ;
  assign n120 = ~x0 & ~x30 ;
  assign n119 = x30 ^ x0 ;
  assign n121 = n120 ^ n119 ;
  assign n122 = n118 & n121 ;
  assign n124 = x32 & x33 ;
  assign n123 = x33 ^ x32 ;
  assign n125 = n124 ^ n123 ;
  assign n127 = x34 & x35 ;
  assign n126 = x35 ^ x34 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = ~n125 & ~n128 ;
  assign n130 = n122 & n129 ;
  assign n131 = x39 & ~n130 ;
  assign n132 = ~x42 & ~x43 ;
  assign n133 = ~x40 & n132 ;
  assign n134 = ~n131 & n133 ;
  assign n135 = ~x41 & n132 ;
  assign n136 = x44 & x47 ;
  assign n137 = ~n135 & n136 ;
  assign n138 = x45 & n108 ;
  assign n139 = n107 & n138 ;
  assign n140 = n137 & n139 ;
  assign n141 = ~n134 & n140 ;
  assign n142 = n115 & ~n141 ;
  assign n143 = x36 & x37 ;
  assign n144 = ~x0 & x31 ;
  assign n145 = n124 & n127 ;
  assign n146 = n144 & n145 ;
  assign n147 = x38 & n146 ;
  assign n148 = n143 & n147 ;
  assign n149 = ~x39 & ~n148 ;
  assign n150 = ~n120 & n140 ;
  assign n151 = ~n149 & n150 ;
  assign n152 = n142 & ~n151 ;
  assign n153 = ~n69 & ~n152 ;
  assign n154 = n105 & n153 ;
  assign n155 = n87 & ~n154 ;
  assign n156 = n100 & ~n155 ;
  assign n157 = n103 & ~n156 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n102 & n105 ;
  assign n160 = ~n142 & n159 ;
  assign y0 = ~n102 ;
  assign y1 = ~n158 ;
  assign y2 = n160 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
