module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n193 , n194 , n195 , n196 , n197 , n198 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n557 , n558 , n559 , n561 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n686 , n687 , n688 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n861 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n890 , n891 , n892 , n893 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n928 , n929 , n930 , n931 , n934 , n935 , n936 , n938 , n939 , n940 , n941 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1014 , n1015 , n1016 , n1018 , n1021 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1033 , n1034 , n1035 , n1036 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1058 , n1059 , n1060 , n1061 , n1064 , n1065 , n1066 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1099 , n1100 , n1101 , n1102 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1130 , n1131 , n1132 , n1133 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1265 , n1266 , n1267 , n1268 , n1269 , n1274 , n1275 , n1276 , n1277 , n1282 , n1283 , n1284 , n1285 , n1286 , n1289 , n1290 , n1291 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1316 , n1317 , n1318 , n1319 , n1320 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1363 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1476 , n1479 , n1480 , n1481 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1623 , n1624 , n1625 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1847 , n1848 , n1849 , n1850 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1990 , n1991 , n1992 , n1993 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2451 , n2452 , n2453 , n2454 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2470 , n2471 , n2472 , n2473 , n2476 , n2477 , n2478 , n2479 , n2484 , n2485 , n2486 , n2487 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2715 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2847 , n2848 , n2849 , n2850 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2934 , n2935 , n2936 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2964 , n2965 , n2966 , n2967 , n2968 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2982 , n2983 , n2984 , n2985 , n2986 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4850 , n4851 , n4852 , n4853 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4911 , n4912 , n4913 , n4914 , n4915 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5451 , n5452 , n5455 , n5456 , n5457 , n5458 , n5459 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5847 , n5848 , n5849 , n5850 , n5851 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7798 , n7799 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7938 , n7939 , n7940 , n7941 , n7942 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9251 , n9252 , n9253 , n9254 , n9255 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9930 , n9931 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9974 , n9975 , n9976 , n9977 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10024 , n10025 , n10026 , n10027 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10655 , n10656 , n10657 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11358 , n11359 , n11360 , n11361 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11628 , n11629 , n11630 , n11631 , n11632 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12060 , n12061 , n12062 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13379 , n13380 , n13381 , n13382 , n13383 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13943 , n13944 , n13945 , n13946 , n13947 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15355 , n15356 , n15357 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15427 , n15428 , n15429 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16660 , n16661 , n16662 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17238 , n17239 , n17240 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17308 , n17309 , n17310 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17467 , n17468 , n17469 , n17470 , n17471 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17523 , n17524 , n17525 , n17528 , n17529 , n17530 , n17531 , n17532 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17591 , n17592 , n17593 , n17594 , n17595 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17748 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18021 , n18022 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18230 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19191 , n19192 , n19193 , n19194 , n19195 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19711 , n19712 , n19713 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19735 , n19736 , n19737 , n19738 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22427 , n22428 , n22429 , n22430 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23991 , n23992 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24828 , n24829 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24849 , n24850 , n24851 , n24852 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 ;
  assign n325 = x125 ^ x14 ;
  assign n326 = x77 ^ x30 ;
  assign n344 = n325 & n326 ;
  assign n330 = x118 ^ x6 ;
  assign n327 = x76 ^ x22 ;
  assign n345 = n330 ^ n327 ;
  assign n346 = n344 & n345 ;
  assign n332 = ~n327 & n330 ;
  assign n333 = n326 & n332 ;
  assign n358 = n346 ^ n333 ;
  assign n352 = n327 & n344 ;
  assign n328 = ~n326 & n327 ;
  assign n351 = n328 ^ n327 ;
  assign n353 = n352 ^ n351 ;
  assign n354 = ~n330 & n353 ;
  assign n355 = n354 ^ n352 ;
  assign n329 = n325 & n328 ;
  assign n337 = n329 ^ n328 ;
  assign n349 = ~n330 & n337 ;
  assign n334 = n333 ^ n332 ;
  assign n335 = ~n325 & n334 ;
  assign n348 = n335 ^ n334 ;
  assign n350 = n349 ^ n348 ;
  assign n356 = n355 ^ n350 ;
  assign n340 = n329 ^ n325 ;
  assign n339 = n329 ^ n327 ;
  assign n341 = n340 ^ n339 ;
  assign n342 = ~n330 & n341 ;
  assign n343 = n342 ^ n340 ;
  assign n347 = n346 ^ n343 ;
  assign n357 = n356 ^ n347 ;
  assign n359 = n358 ^ n357 ;
  assign n2082 = n359 ^ n354 ;
  assign n322 = x108 ^ x38 ;
  assign n372 = n328 ^ n326 ;
  assign n373 = n372 ^ n334 ;
  assign n374 = n325 & ~n373 ;
  assign n390 = n374 ^ n373 ;
  assign n2078 = n390 ^ n354 ;
  assign n2079 = n2078 ^ n348 ;
  assign n2080 = n2079 ^ n357 ;
  assign n2081 = n322 & ~n2080 ;
  assign n2083 = n2082 ^ n2081 ;
  assign n331 = n329 & ~n330 ;
  assign n779 = n331 ^ n329 ;
  assign n780 = n779 ^ n374 ;
  assign n778 = n346 ^ n344 ;
  assign n781 = n780 ^ n778 ;
  assign n782 = ~n322 & n781 ;
  assign n783 = n782 ^ n780 ;
  assign n2089 = n2083 ^ n783 ;
  assign n323 = x94 ^ x56 ;
  assign n324 = n323 ^ n322 ;
  assign n376 = n355 ^ n351 ;
  assign n360 = n344 ^ n326 ;
  assign n361 = n360 ^ n353 ;
  assign n362 = n361 ^ n359 ;
  assign n1571 = n376 ^ n362 ;
  assign n391 = n349 ^ n337 ;
  assign n392 = n391 ^ n390 ;
  assign n1572 = n1571 ^ n392 ;
  assign n1575 = n322 & ~n1572 ;
  assign n1576 = n1575 ^ n392 ;
  assign n1577 = n324 & ~n1576 ;
  assign n2090 = n2089 ^ n1577 ;
  assign n2091 = n2090 ^ x25 ;
  assign n2084 = n2083 ^ n353 ;
  assign n809 = n779 ^ n350 ;
  assign n1568 = n809 ^ n335 ;
  assign n2077 = n1568 ^ n783 ;
  assign n2085 = n2084 ^ n2077 ;
  assign n2075 = n779 ^ n390 ;
  assign n2076 = n322 & ~n2075 ;
  assign n2086 = n2085 ^ n2076 ;
  assign n2087 = ~n324 & n2086 ;
  assign n2092 = n2091 ^ n2087 ;
  assign n370 = n322 & n323 ;
  assign n399 = n370 ^ n324 ;
  assign n2074 = ~n399 & n778 ;
  assign n2093 = n2092 ^ n2074 ;
  assign n2068 = n346 ^ n329 ;
  assign n2071 = n322 & n2068 ;
  assign n2072 = n2071 ^ n329 ;
  assign n2073 = n323 & n2072 ;
  assign n2094 = n2093 ^ n2073 ;
  assign n2337 = n2094 ^ x112 ;
  assign n409 = x83 ^ x30 ;
  assign n410 = x124 ^ x4 ;
  assign n475 = n409 & n410 ;
  assign n487 = n475 ^ n410 ;
  assign n416 = x101 ^ x54 ;
  assign n417 = x126 ^ x46 ;
  assign n418 = ~n416 & n417 ;
  assign n419 = n418 ^ n416 ;
  assign n421 = n419 ^ n417 ;
  assign n412 = x78 ^ x38 ;
  assign n413 = x84 ^ x62 ;
  assign n414 = n412 & ~n413 ;
  assign n415 = n414 ^ n413 ;
  assign n441 = n415 ^ n412 ;
  assign n443 = n441 ^ n413 ;
  assign n444 = n421 & n443 ;
  assign n435 = ~n415 & n421 ;
  assign n431 = n418 ^ n417 ;
  assign n432 = n414 & n431 ;
  assign n425 = ~n415 & n418 ;
  assign n422 = n414 & n421 ;
  assign n430 = n425 ^ n422 ;
  assign n433 = n432 ^ n430 ;
  assign n424 = n414 & n418 ;
  assign n426 = n425 ^ n424 ;
  assign n429 = n426 ^ n414 ;
  assign n434 = n433 ^ n429 ;
  assign n436 = n435 ^ n434 ;
  assign n437 = n436 ^ n432 ;
  assign n420 = ~n415 & ~n419 ;
  assign n423 = n422 ^ n420 ;
  assign n427 = n426 ^ n423 ;
  assign n428 = n427 ^ n413 ;
  assign n438 = n437 ^ n428 ;
  assign n2360 = n444 ^ n438 ;
  assign n2361 = n487 & ~n2360 ;
  assign n449 = n431 & n443 ;
  assign n450 = n449 ^ n432 ;
  assign n451 = n450 ^ n431 ;
  assign n452 = n451 ^ n438 ;
  assign n460 = n452 ^ n441 ;
  assign n457 = n418 & n443 ;
  assign n456 = n426 ^ n418 ;
  assign n458 = n457 ^ n456 ;
  assign n446 = n421 & n441 ;
  assign n459 = n458 ^ n446 ;
  assign n461 = n460 ^ n459 ;
  assign n478 = n461 ^ n419 ;
  assign n477 = n434 ^ n420 ;
  assign n479 = n478 ^ n477 ;
  assign n1310 = n479 ^ n452 ;
  assign n2357 = n1310 ^ x9 ;
  assign n469 = n438 ^ n435 ;
  assign n472 = ~n410 & ~n469 ;
  assign n473 = n472 ^ n435 ;
  assign n474 = n409 & n473 ;
  assign n411 = n410 ^ n409 ;
  assign n2350 = n437 ^ n427 ;
  assign n2351 = n2350 ^ n461 ;
  assign n2349 = n425 & n475 ;
  assign n2352 = n2351 ^ n2349 ;
  assign n2353 = ~n411 & ~n2352 ;
  assign n2354 = n2353 ^ n427 ;
  assign n476 = n475 ^ n409 ;
  assign n2346 = n458 ^ n444 ;
  assign n2347 = n2346 ^ n479 ;
  assign n2348 = n476 & n2347 ;
  assign n2355 = n2354 ^ n2348 ;
  assign n2356 = ~n474 & ~n2355 ;
  assign n2358 = n2357 ^ n2356 ;
  assign n2345 = ~n411 & n457 ;
  assign n2359 = n2358 ^ n2345 ;
  assign n2362 = n2361 ^ n2359 ;
  assign n1334 = n459 ^ n449 ;
  assign n2342 = ~n409 & n1334 ;
  assign n2343 = n2342 ^ n1310 ;
  assign n2344 = ~n410 & ~n2343 ;
  assign n2363 = n2362 ^ n2344 ;
  assign n2364 = n2363 ^ x64 ;
  assign n2365 = ~n2337 & n2364 ;
  assign n603 = x85 ^ x2 ;
  assign n614 = x102 ^ x52 ;
  assign n606 = x117 ^ x44 ;
  assign n607 = x100 ^ x36 ;
  assign n608 = x91 ^ x60 ;
  assign n634 = n607 & n608 ;
  assign n635 = ~n606 & n634 ;
  assign n636 = n614 & n635 ;
  assign n637 = n636 ^ n635 ;
  assign n621 = n606 & ~n614 ;
  assign n626 = n607 & n621 ;
  assign n627 = n626 ^ n621 ;
  assign n612 = n606 & ~n607 ;
  assign n628 = n627 ^ n612 ;
  assign n623 = n607 ^ n606 ;
  assign n624 = n614 ^ n606 ;
  assign n625 = n623 & ~n624 ;
  assign n629 = n628 ^ n625 ;
  assign n638 = n637 ^ n629 ;
  assign n615 = ~n608 & n614 ;
  assign n618 = n607 & n615 ;
  assign n632 = n606 & n618 ;
  assign n633 = n632 ^ n618 ;
  assign n639 = n638 ^ n633 ;
  assign n622 = n621 ^ n614 ;
  assign n630 = n629 ^ n622 ;
  assign n616 = n612 & n615 ;
  assign n617 = n616 ^ n615 ;
  assign n619 = n618 ^ n617 ;
  assign n613 = n612 ^ n607 ;
  assign n620 = n619 ^ n613 ;
  assign n631 = n630 ^ n620 ;
  assign n640 = n639 ^ n631 ;
  assign n609 = n608 ^ n607 ;
  assign n610 = n609 ^ n606 ;
  assign n611 = ~n606 & n610 ;
  assign n641 = n640 ^ n611 ;
  assign n678 = n641 ^ n633 ;
  assign n643 = n628 ^ n616 ;
  assign n1746 = n678 ^ n643 ;
  assign n647 = ~n608 & n627 ;
  assign n679 = n647 ^ n627 ;
  assign n680 = n679 ^ n678 ;
  assign n681 = n680 ^ n632 ;
  assign n1747 = n1746 ^ n681 ;
  assign n645 = ~n608 & n626 ;
  assign n699 = n645 ^ n619 ;
  assign n661 = n645 ^ n626 ;
  assign n660 = n635 ^ n634 ;
  assign n662 = n661 ^ n660 ;
  assign n700 = n699 ^ n662 ;
  assign n1748 = n1747 ^ n700 ;
  assign n1749 = n603 & n1748 ;
  assign n1750 = n1749 ^ n1746 ;
  assign n604 = x67 ^ x28 ;
  assign n655 = n603 & ~n604 ;
  assign n656 = n655 ^ n604 ;
  assign n698 = n656 ^ n603 ;
  assign n1520 = n698 ^ n604 ;
  assign n1521 = n647 ^ n638 ;
  assign n1522 = n1520 & n1521 ;
  assign n707 = n616 & n698 ;
  assign n1523 = n1522 ^ n707 ;
  assign n1765 = n1750 ^ n1523 ;
  assign n605 = n604 ^ n603 ;
  assign n693 = n604 & n639 ;
  assign n694 = n693 ^ n638 ;
  assign n695 = ~n605 & n694 ;
  assign n1766 = n1765 ^ n695 ;
  assign n1532 = n603 & n637 ;
  assign n663 = n662 ^ n631 ;
  assign n664 = n663 ^ n661 ;
  assign n1526 = ~n604 & n664 ;
  assign n1527 = n1526 ^ n661 ;
  assign n1533 = n1532 ^ n1527 ;
  assign n1534 = n605 & n1533 ;
  assign n1535 = n1534 ^ n1527 ;
  assign n1767 = n1766 ^ n1535 ;
  assign n1760 = n661 ^ n616 ;
  assign n1761 = n1760 ^ n638 ;
  assign n1762 = ~n604 & n1761 ;
  assign n1763 = n1762 ^ n638 ;
  assign n1764 = ~n603 & n1763 ;
  assign n1768 = n1767 ^ n1764 ;
  assign n1769 = n1768 ^ x1 ;
  assign n1752 = n645 ^ n636 ;
  assign n670 = n661 ^ n643 ;
  assign n1553 = n679 ^ n670 ;
  assign n701 = n641 ^ n630 ;
  assign n1554 = n1553 ^ n701 ;
  assign n1751 = n1750 ^ n1554 ;
  assign n1753 = n1752 ^ n1751 ;
  assign n1754 = n1753 ^ n1750 ;
  assign n1757 = ~n603 & ~n1754 ;
  assign n1758 = n1757 ^ n1750 ;
  assign n1759 = n604 & n1758 ;
  assign n1770 = n1769 ^ n1759 ;
  assign n1743 = n632 ^ n631 ;
  assign n1742 = n701 ^ n637 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1745 = n1520 & ~n1744 ;
  assign n1771 = n1770 ^ n1745 ;
  assign n2366 = n1771 ^ x74 ;
  assign n237 = x98 ^ x58 ;
  assign n238 = x89 ^ x50 ;
  assign n239 = n237 & n238 ;
  assign n234 = x107 ^ x34 ;
  assign n235 = x88 ^ x42 ;
  assign n236 = n234 & ~n235 ;
  assign n245 = n236 ^ n234 ;
  assign n259 = n245 ^ n235 ;
  assign n265 = n239 & n259 ;
  assign n248 = n239 ^ n237 ;
  assign n249 = n245 & n248 ;
  assign n266 = n265 ^ n249 ;
  assign n263 = n236 ^ n235 ;
  assign n264 = n239 & ~n263 ;
  assign n267 = n266 ^ n264 ;
  assign n261 = n238 ^ n234 ;
  assign n262 = n237 & n261 ;
  assign n268 = n267 ^ n262 ;
  assign n1240 = n268 ^ n264 ;
  assign n1250 = n1240 ^ n249 ;
  assign n240 = n239 ^ n238 ;
  assign n241 = n236 & n240 ;
  assign n2374 = n1250 ^ n241 ;
  assign n270 = n268 ^ n236 ;
  assign n242 = n240 ^ n237 ;
  assign n243 = n236 & ~n242 ;
  assign n244 = n243 ^ n241 ;
  assign n271 = n270 ^ n244 ;
  assign n2383 = n2374 ^ n271 ;
  assign n233 = x66 ^ x0 ;
  assign n252 = x121 ^ x26 ;
  assign n286 = n240 & ~n263 ;
  assign n1644 = n252 & n286 ;
  assign n277 = n240 & n259 ;
  assign n1241 = n1240 ^ n277 ;
  assign n274 = n240 & n245 ;
  assign n1637 = n1241 ^ n274 ;
  assign n1638 = n252 & n1637 ;
  assign n1639 = n1638 ^ n1241 ;
  assign n1645 = n1644 ^ n1639 ;
  assign n1646 = ~n233 & n1645 ;
  assign n1647 = n1646 ^ n1639 ;
  assign n2384 = n2383 ^ n1647 ;
  assign n258 = n252 ^ n233 ;
  assign n287 = n286 ^ n266 ;
  assign n260 = n248 & n259 ;
  assign n285 = n260 ^ n243 ;
  assign n288 = n287 ^ n285 ;
  assign n283 = n237 ^ n235 ;
  assign n246 = n239 & n245 ;
  assign n282 = n246 ^ n241 ;
  assign n284 = n283 ^ n282 ;
  assign n289 = n288 ^ n284 ;
  assign n275 = n274 ^ n245 ;
  assign n250 = n249 ^ n246 ;
  assign n276 = n275 ^ n250 ;
  assign n290 = n289 ^ n276 ;
  assign n1274 = n233 & ~n290 ;
  assign n281 = n243 ^ n242 ;
  assign n291 = n290 ^ n281 ;
  assign n1275 = n1274 ^ n291 ;
  assign n1276 = n258 & n1275 ;
  assign n1277 = n1276 ^ n291 ;
  assign n2385 = n2384 ^ n1277 ;
  assign n1265 = n252 & ~n289 ;
  assign n1257 = n260 ^ n246 ;
  assign n1258 = n1257 ^ n274 ;
  assign n1259 = n252 & n1258 ;
  assign n1260 = n1259 ^ n274 ;
  assign n1266 = n1265 ^ n1260 ;
  assign n1267 = n233 & n1266 ;
  assign n1268 = n1267 ^ n1260 ;
  assign n307 = n233 & ~n252 ;
  assign n308 = n307 ^ n252 ;
  assign n309 = n308 ^ n233 ;
  assign n1256 = ~n290 & n309 ;
  assign n1269 = n1268 ^ n1256 ;
  assign n2386 = n2385 ^ n1269 ;
  assign n2387 = n2386 ^ x17 ;
  assign n2375 = n2374 ^ n265 ;
  assign n2376 = n2375 ^ n243 ;
  assign n2377 = n2376 ^ n2374 ;
  assign n2380 = ~n233 & n2377 ;
  assign n2381 = n2380 ^ n2374 ;
  assign n2382 = n258 & n2381 ;
  assign n2388 = n2387 ^ n2382 ;
  assign n279 = n249 ^ n248 ;
  assign n269 = n268 ^ n260 ;
  assign n280 = n279 ^ n269 ;
  assign n1623 = n280 ^ n277 ;
  assign n2373 = ~n308 & n1623 ;
  assign n2389 = n2388 ^ n2373 ;
  assign n2367 = n282 ^ n271 ;
  assign n2368 = n2367 ^ n280 ;
  assign n2369 = n2368 ^ n271 ;
  assign n2370 = n233 & n2369 ;
  assign n2371 = n2370 ^ n271 ;
  assign n2372 = ~n252 & n2371 ;
  assign n2390 = n2389 ^ n2372 ;
  assign n2391 = n2390 ^ x122 ;
  assign n2392 = n2366 & ~n2391 ;
  assign n2414 = n2365 & n2392 ;
  assign n2393 = n2392 ^ n2366 ;
  assign n2394 = n2393 ^ n2391 ;
  assign n2395 = n2365 & n2394 ;
  assign n2415 = n2414 ^ n2395 ;
  assign n2412 = n2365 & n2393 ;
  assign n2413 = n2412 ^ n2365 ;
  assign n2416 = n2415 ^ n2413 ;
  assign n2400 = n2392 ^ n2391 ;
  assign n2417 = n2416 ^ n2400 ;
  assign n2405 = n2365 ^ n2337 ;
  assign n2410 = ~n2400 & ~n2405 ;
  assign n2397 = n2365 ^ n2364 ;
  assign n2401 = n2397 & ~n2400 ;
  assign n2411 = n2410 ^ n2401 ;
  assign n2418 = n2417 ^ n2411 ;
  assign n2406 = n2405 ^ n2364 ;
  assign n2409 = n2393 & n2406 ;
  assign n2419 = n2418 ^ n2409 ;
  assign n2407 = n2392 & n2406 ;
  assign n2408 = n2407 ^ n2406 ;
  assign n2420 = n2419 ^ n2408 ;
  assign n2398 = n2392 & n2397 ;
  assign n2444 = n2420 ^ n2398 ;
  assign n133 = x114 ^ x56 ;
  assign n134 = x123 ^ x40 ;
  assign n135 = n133 & n134 ;
  assign n137 = x112 ^ x32 ;
  assign n138 = x97 ^ x48 ;
  assign n139 = ~n137 & n138 ;
  assign n185 = n135 & n139 ;
  assign n129 = x80 ^ x24 ;
  assign n130 = x73 ^ x6 ;
  assign n131 = ~n129 & n130 ;
  assign n145 = n138 ^ n133 ;
  assign n147 = n138 ^ n137 ;
  assign n148 = n134 & n147 ;
  assign n146 = n137 ^ n134 ;
  assign n149 = n148 ^ n146 ;
  assign n150 = ~n145 & n149 ;
  assign n187 = n150 ^ n145 ;
  assign n158 = n138 ^ n134 ;
  assign n159 = ~n137 & n158 ;
  assign n160 = n159 ^ n134 ;
  assign n161 = ~n133 & n160 ;
  assign n174 = n161 ^ n160 ;
  assign n188 = n187 ^ n174 ;
  assign n151 = n135 & n147 ;
  assign n186 = n185 ^ n151 ;
  assign n189 = n188 ^ n186 ;
  assign n140 = n139 ^ n137 ;
  assign n141 = n140 ^ n138 ;
  assign n136 = n135 ^ n133 ;
  assign n153 = n136 ^ n134 ;
  assign n157 = n141 & ~n153 ;
  assign n1831 = n189 ^ n157 ;
  assign n1832 = n131 & ~n1831 ;
  assign n154 = n153 ^ n133 ;
  assign n152 = n151 ^ n148 ;
  assign n177 = n154 ^ n152 ;
  assign n162 = n139 & ~n153 ;
  assign n163 = n162 ^ n154 ;
  assign n164 = n163 ^ n161 ;
  assign n178 = n177 ^ n164 ;
  assign n165 = n164 ^ n157 ;
  assign n155 = n139 & n154 ;
  assign n156 = n155 ^ n152 ;
  assign n166 = n165 ^ n156 ;
  assign n167 = n166 ^ n150 ;
  assign n144 = n136 & ~n140 ;
  assign n168 = n167 ^ n144 ;
  assign n142 = n136 & n141 ;
  assign n143 = n142 ^ n136 ;
  assign n169 = n168 ^ n143 ;
  assign n172 = n169 ^ n151 ;
  assign n176 = n172 ^ n167 ;
  assign n179 = n178 ^ n176 ;
  assign n175 = n174 ^ n172 ;
  assign n180 = n179 ^ n175 ;
  assign n171 = n139 ^ n138 ;
  assign n173 = n172 ^ n171 ;
  assign n181 = n180 ^ n173 ;
  assign n1816 = n181 ^ n155 ;
  assign n182 = n181 ^ n164 ;
  assign n1813 = n182 ^ n156 ;
  assign n1814 = n1813 ^ n142 ;
  assign n1815 = n1814 ^ n174 ;
  assign n1817 = n1816 ^ n1815 ;
  assign n1818 = n130 & n1817 ;
  assign n1819 = n1818 ^ n1814 ;
  assign n1833 = n1832 ^ n1819 ;
  assign n205 = n131 ^ n129 ;
  assign n1828 = n157 ^ n144 ;
  assign n196 = n169 ^ n135 ;
  assign n197 = n196 ^ n174 ;
  assign n210 = n197 ^ n169 ;
  assign n211 = n210 ^ n175 ;
  assign n1829 = n1828 ^ n211 ;
  assign n1830 = ~n205 & n1829 ;
  assign n1834 = n1833 ^ n1830 ;
  assign n1812 = n130 ^ n129 ;
  assign n1821 = n1819 ^ n162 ;
  assign n1820 = n1819 ^ n161 ;
  assign n1822 = n1821 ^ n1820 ;
  assign n1825 = n130 & n1822 ;
  assign n1826 = n1825 ^ n1821 ;
  assign n1827 = ~n1812 & n1826 ;
  assign n1835 = n1834 ^ n1827 ;
  assign n132 = n131 ^ n130 ;
  assign n1369 = n132 & n144 ;
  assign n1836 = n1835 ^ n1369 ;
  assign n198 = n197 ^ n178 ;
  assign n201 = n130 & n198 ;
  assign n202 = n201 ^ n178 ;
  assign n203 = n129 & n202 ;
  assign n1837 = n1836 ^ n203 ;
  assign n1363 = n167 ^ n156 ;
  assign n1366 = n129 & n1363 ;
  assign n1367 = n1366 ^ n156 ;
  assign n1368 = ~n130 & n1367 ;
  assign n1838 = n1837 ^ n1368 ;
  assign n190 = n189 ^ n167 ;
  assign n193 = ~n130 & ~n190 ;
  assign n194 = n193 ^ n167 ;
  assign n195 = n129 & n194 ;
  assign n1839 = n1838 ^ n195 ;
  assign n1840 = ~n185 & ~n1839 ;
  assign n1841 = n1840 ^ x59 ;
  assign n2334 = n1841 ^ x97 ;
  assign n861 = x110 ^ x36 ;
  assign n822 = x92 ^ x62 ;
  assign n893 = n861 ^ n822 ;
  assign n823 = x68 ^ x20 ;
  assign n824 = x93 ^ x28 ;
  assign n825 = x116 ^ x12 ;
  assign n826 = n824 & n825 ;
  assign n827 = n826 ^ n824 ;
  assign n828 = n823 & ~n827 ;
  assign n830 = x86 ^ x4 ;
  assign n831 = n823 & ~n830 ;
  assign n833 = n831 ^ n830 ;
  assign n836 = n833 ^ n823 ;
  assign n850 = n836 ^ n830 ;
  assign n852 = n824 & n850 ;
  assign n851 = n827 & n850 ;
  assign n853 = n852 ^ n851 ;
  assign n840 = n830 ^ n823 ;
  assign n841 = n840 ^ n824 ;
  assign n842 = ~n823 & n841 ;
  assign n837 = n826 & n836 ;
  assign n838 = n837 ^ n826 ;
  assign n834 = ~n824 & ~n833 ;
  assign n835 = n834 ^ n833 ;
  assign n839 = n838 ^ n835 ;
  assign n843 = n842 ^ n839 ;
  assign n844 = n843 ^ n824 ;
  assign n845 = n844 ^ n840 ;
  assign n829 = n828 ^ n823 ;
  assign n832 = n831 ^ n829 ;
  assign n846 = n845 ^ n832 ;
  assign n847 = n846 ^ n837 ;
  assign n848 = n847 ^ n826 ;
  assign n849 = n848 ^ n839 ;
  assign n854 = n853 ^ n849 ;
  assign n855 = n854 ^ n838 ;
  assign n856 = n855 ^ n851 ;
  assign n918 = n856 ^ n849 ;
  assign n1993 = n918 ^ n837 ;
  assign n1382 = n851 ^ n829 ;
  assign n1996 = n1993 ^ n1382 ;
  assign n1997 = ~n828 & n1996 ;
  assign n1998 = n1997 ^ n1993 ;
  assign n1999 = n861 & n1998 ;
  assign n2000 = n1999 ^ n1993 ;
  assign n2001 = ~n893 & n2000 ;
  assign n2002 = n2001 ^ x33 ;
  assign n857 = n826 ^ n825 ;
  assign n872 = n850 & n857 ;
  assign n873 = n872 ^ n850 ;
  assign n874 = n873 ^ n852 ;
  assign n875 = n874 ^ n834 ;
  assign n868 = n830 ^ n825 ;
  assign n876 = n875 ^ n868 ;
  assign n869 = ~n825 & ~n868 ;
  assign n870 = n869 ^ n824 ;
  assign n871 = ~n823 & n870 ;
  assign n877 = n876 ^ n871 ;
  assign n1990 = ~n822 & ~n877 ;
  assign n1991 = n1990 ^ n875 ;
  assign n1992 = n861 & n1991 ;
  assign n2003 = n2002 ^ n1992 ;
  assign n917 = n822 & ~n861 ;
  assign n1983 = n845 ^ n825 ;
  assign n1984 = n1983 ^ n824 ;
  assign n1985 = n917 & ~n1984 ;
  assign n2004 = n2003 ^ n1985 ;
  assign n1982 = ~n846 & ~n861 ;
  assign n2005 = n2004 ^ n1982 ;
  assign n879 = n877 ^ n837 ;
  assign n858 = n831 & n857 ;
  assign n859 = n858 ^ n856 ;
  assign n880 = n879 ^ n859 ;
  assign n1974 = n880 ^ n874 ;
  assign n1975 = n1974 ^ n858 ;
  assign n1976 = n1975 ^ n880 ;
  assign n1979 = ~n861 & n1976 ;
  assign n1980 = n1979 ^ n880 ;
  assign n1981 = ~n893 & n1980 ;
  assign n2006 = n2005 ^ n1981 ;
  assign n2335 = n2006 ^ x88 ;
  assign n2493 = ~n2334 & ~n2335 ;
  assign n2494 = n2493 ^ n2335 ;
  assign n3232 = ~n2444 & ~n2494 ;
  assign n2495 = n2494 ^ n2334 ;
  assign n2496 = n2416 & ~n2495 ;
  assign n3233 = n3232 ^ n2496 ;
  assign n2446 = n2391 ^ n2366 ;
  assign n2447 = n2446 ^ n2337 ;
  assign n2461 = n2447 ^ n2364 ;
  assign n2431 = n2415 ^ n2407 ;
  assign n2402 = n2393 & n2397 ;
  assign n2403 = n2402 ^ n2401 ;
  assign n2430 = n2410 ^ n2403 ;
  assign n2432 = n2431 ^ n2430 ;
  assign n2462 = n2461 ^ n2432 ;
  assign n2463 = n2462 ^ n2420 ;
  assign n3227 = n2463 ^ n2395 ;
  assign n3228 = n2493 & n3227 ;
  assign n2399 = n2398 ^ n2397 ;
  assign n2404 = n2403 ^ n2399 ;
  assign n2421 = n2420 ^ n2404 ;
  assign n2396 = n2395 ^ n2394 ;
  assign n2422 = n2421 ^ n2396 ;
  assign n2931 = n2422 ^ n2409 ;
  assign n2934 = ~n2335 & ~n2931 ;
  assign n2935 = n2934 ^ n2409 ;
  assign n2936 = n2334 & n2935 ;
  assign n3229 = n3228 ^ n2936 ;
  assign n3209 = n2463 ^ n2415 ;
  assign n3210 = n3209 ^ n2418 ;
  assign n3211 = n3210 ^ n2409 ;
  assign n2443 = n2416 ^ n2401 ;
  assign n2445 = n2444 ^ n2443 ;
  assign n2448 = n2447 ^ n2445 ;
  assign n3212 = n3211 ^ n2448 ;
  assign n3213 = ~n2334 & ~n3212 ;
  assign n3214 = n3213 ^ n3210 ;
  assign n2479 = n2407 ^ n2402 ;
  assign n2484 = ~n2334 & n2479 ;
  assign n2485 = n2484 ^ n2407 ;
  assign n2486 = ~n2335 & n2485 ;
  assign n3224 = n3214 ^ n2486 ;
  assign n2336 = n2335 ^ n2334 ;
  assign n2941 = n2334 & ~n2421 ;
  assign n2942 = n2941 ^ n2420 ;
  assign n2943 = ~n2336 & ~n2942 ;
  assign n3225 = n3224 ^ n2943 ;
  assign n2464 = n2463 ^ n2422 ;
  assign n2460 = n2410 ^ n2405 ;
  assign n2465 = n2464 ^ n2460 ;
  assign n2473 = n2465 ^ n2412 ;
  assign n2476 = n2335 & n2473 ;
  assign n2477 = n2476 ^ n2412 ;
  assign n2478 = n2334 & n2477 ;
  assign n3226 = n3225 ^ n2478 ;
  assign n3230 = n3229 ^ n3226 ;
  assign n2927 = n2495 ^ n2335 ;
  assign n2945 = n2416 & ~n2927 ;
  assign n2944 = n2402 & ~n2494 ;
  assign n2946 = n2945 ^ n2944 ;
  assign n3231 = n3230 ^ n2946 ;
  assign n3234 = n3233 ^ n3231 ;
  assign n3235 = n3234 ^ x38 ;
  assign n3217 = n3214 ^ n2411 ;
  assign n2952 = n2465 ^ n2422 ;
  assign n2435 = n2418 ^ n2398 ;
  assign n3215 = n2952 ^ n2435 ;
  assign n3216 = n3215 ^ n3214 ;
  assign n3218 = n3217 ^ n3216 ;
  assign n3221 = ~n2334 & n3218 ;
  assign n3222 = n3221 ^ n3217 ;
  assign n3223 = ~n2335 & ~n3222 ;
  assign n3236 = n3235 ^ n3223 ;
  assign n3443 = n3236 ^ x84 ;
  assign n226 = n142 & ~n1812 ;
  assign n221 = n185 ^ n168 ;
  assign n217 = n185 ^ n167 ;
  assign n218 = n217 ^ n174 ;
  assign n219 = n218 ^ n181 ;
  assign n220 = n129 & n219 ;
  assign n222 = n221 ^ n220 ;
  assign n223 = ~n130 & n222 ;
  assign n206 = n162 & n205 ;
  assign n204 = n161 ^ n157 ;
  assign n207 = n206 ^ n204 ;
  assign n208 = n207 ^ n131 ;
  assign n212 = n211 ^ n167 ;
  assign n213 = n212 ^ n207 ;
  assign n209 = n161 & ~n205 ;
  assign n214 = n213 ^ n209 ;
  assign n215 = n208 & ~n214 ;
  assign n216 = n215 ^ n131 ;
  assign n224 = n223 ^ n216 ;
  assign n227 = n226 ^ n224 ;
  assign n228 = n227 ^ n203 ;
  assign n229 = n228 ^ n195 ;
  assign n230 = n229 ^ x61 ;
  assign n170 = n169 ^ n152 ;
  assign n183 = n182 ^ n170 ;
  assign n184 = n132 & n183 ;
  assign n231 = n230 ^ n184 ;
  assign n232 = n231 ^ x96 ;
  assign n319 = n267 & n307 ;
  assign n310 = n286 ^ n249 ;
  assign n311 = n310 ^ n234 ;
  assign n292 = n291 ^ n280 ;
  assign n312 = n311 ^ n292 ;
  assign n313 = n309 & ~n312 ;
  assign n301 = n242 ^ n241 ;
  assign n302 = n301 ^ n276 ;
  assign n303 = ~n252 & ~n302 ;
  assign n298 = n292 ^ n274 ;
  assign n278 = n277 ^ n276 ;
  assign n293 = n292 ^ n278 ;
  assign n294 = n278 ^ n233 ;
  assign n295 = n258 & n294 ;
  assign n296 = n295 ^ n233 ;
  assign n297 = n293 & ~n296 ;
  assign n299 = n298 ^ n297 ;
  assign n300 = n299 ^ n286 ;
  assign n304 = n303 ^ n300 ;
  assign n305 = ~n258 & n304 ;
  assign n306 = n305 ^ n303 ;
  assign n314 = n313 ^ n306 ;
  assign n272 = n271 ^ n269 ;
  assign n273 = ~n258 & n272 ;
  assign n315 = n314 ^ n273 ;
  assign n316 = n315 ^ n246 ;
  assign n317 = n316 ^ x3 ;
  assign n247 = n246 ^ n244 ;
  assign n251 = n250 ^ n247 ;
  assign n253 = n252 ^ n250 ;
  assign n254 = n253 ^ n250 ;
  assign n255 = n251 & n254 ;
  assign n256 = n255 ^ n250 ;
  assign n257 = ~n233 & n256 ;
  assign n318 = n317 ^ n257 ;
  assign n320 = n319 ^ n318 ;
  assign n321 = n320 ^ x73 ;
  assign n378 = n357 ^ n344 ;
  assign n400 = n378 & ~n399 ;
  assign n393 = n370 & ~n392 ;
  assign n394 = n393 ^ n362 ;
  assign n381 = n327 ^ n326 ;
  assign n382 = n381 ^ n325 ;
  assign n383 = n382 ^ n333 ;
  assign n336 = n335 ^ n331 ;
  assign n338 = n337 ^ n336 ;
  assign n384 = n383 ^ n338 ;
  assign n385 = n322 & ~n384 ;
  assign n386 = n385 ^ n338 ;
  assign n395 = n394 ^ n386 ;
  assign n396 = n395 ^ x11 ;
  assign n375 = n374 ^ n348 ;
  assign n387 = n386 ^ n375 ;
  assign n377 = n376 ^ n375 ;
  assign n379 = n378 ^ n377 ;
  assign n380 = ~n322 & n379 ;
  assign n388 = n387 ^ n380 ;
  assign n389 = n323 & n388 ;
  assign n397 = n396 ^ n389 ;
  assign n371 = n355 & n370 ;
  assign n398 = n397 ^ n371 ;
  assign n401 = n400 ^ n398 ;
  assign n363 = n362 ^ n338 ;
  assign n364 = n363 ^ n362 ;
  assign n365 = n362 ^ n322 ;
  assign n366 = n365 ^ n362 ;
  assign n367 = n364 & ~n366 ;
  assign n368 = n367 ^ n362 ;
  assign n369 = n324 & n368 ;
  assign n402 = n401 ^ n369 ;
  assign n403 = n402 ^ x82 ;
  assign n404 = n321 & ~n403 ;
  assign n405 = n404 ^ n403 ;
  assign n406 = n405 ^ n321 ;
  assign n407 = n232 & n406 ;
  assign n490 = n436 ^ n424 ;
  assign n491 = n490 ^ n413 ;
  assign n453 = n452 ^ n429 ;
  assign n492 = n491 ^ n453 ;
  assign n488 = n417 ^ n413 ;
  assign n489 = n488 ^ n412 ;
  assign n493 = n492 ^ n489 ;
  assign n494 = n487 & n493 ;
  assign n480 = n479 ^ n446 ;
  assign n481 = n476 & n480 ;
  assign n462 = n461 ^ n449 ;
  assign n463 = n462 ^ n458 ;
  assign n454 = n453 ^ n430 ;
  assign n455 = n454 ^ n444 ;
  assign n464 = n463 ^ n455 ;
  assign n465 = ~n409 & n464 ;
  assign n466 = n465 ^ n453 ;
  assign n482 = n481 ^ n466 ;
  assign n483 = n482 ^ n474 ;
  assign n484 = n483 ^ x35 ;
  assign n442 = n441 ^ n424 ;
  assign n445 = n444 ^ n442 ;
  assign n447 = n446 ^ n445 ;
  assign n448 = n409 & n447 ;
  assign n467 = n466 ^ n448 ;
  assign n468 = n410 & ~n467 ;
  assign n485 = n484 ^ n468 ;
  assign n439 = n438 ^ n434 ;
  assign n440 = ~n411 & ~n439 ;
  assign n486 = n485 ^ n440 ;
  assign n495 = n494 ^ n486 ;
  assign n496 = n495 ^ x114 ;
  assign n702 = n701 ^ n700 ;
  assign n703 = n698 & ~n702 ;
  assign n686 = ~n603 & n681 ;
  assign n687 = n686 ^ n632 ;
  assign n688 = n604 & n687 ;
  assign n696 = n695 ^ n688 ;
  assign n659 = n615 ^ n610 ;
  assign n665 = n664 ^ n659 ;
  assign n642 = n641 ^ n635 ;
  assign n644 = n643 ^ n642 ;
  assign n646 = n645 ^ n644 ;
  assign n666 = n665 ^ n646 ;
  assign n667 = n655 & ~n666 ;
  assign n668 = n667 ^ n656 ;
  assign n669 = n637 ^ n631 ;
  assign n671 = n670 ^ n669 ;
  assign n672 = n671 ^ n637 ;
  assign n675 = ~n655 & ~n672 ;
  assign n676 = n675 ^ n637 ;
  assign n677 = ~n668 & ~n676 ;
  assign n697 = n696 ^ n677 ;
  assign n704 = n703 ^ n697 ;
  assign n657 = n632 ^ n619 ;
  assign n658 = ~n656 & n657 ;
  assign n705 = n704 ^ n658 ;
  assign n652 = n603 & n646 ;
  assign n653 = n652 ^ n647 ;
  assign n654 = ~n605 & n653 ;
  assign n706 = n705 ^ n654 ;
  assign n708 = n707 ^ n706 ;
  assign n709 = n708 ^ x19 ;
  assign n710 = n709 ^ x120 ;
  assign n2570 = ~n496 & ~n710 ;
  assign n2571 = n407 & n2570 ;
  assign n500 = x72 ^ x8 ;
  assign n501 = x82 ^ x0 ;
  assign n502 = n500 & n501 ;
  assign n497 = x65 ^ x16 ;
  assign n498 = x120 ^ x24 ;
  assign n499 = ~n497 & ~n498 ;
  assign n511 = n499 ^ n497 ;
  assign n512 = n511 ^ n498 ;
  assign n518 = n502 & ~n512 ;
  assign n525 = n518 ^ n512 ;
  assign n503 = n502 ^ n501 ;
  assign n504 = n503 ^ n500 ;
  assign n505 = n504 ^ n501 ;
  assign n523 = n505 & ~n512 ;
  assign n522 = n503 & ~n512 ;
  assign n524 = n523 ^ n522 ;
  assign n526 = n525 ^ n524 ;
  assign n507 = x96 ^ x32 ;
  assign n508 = x105 ^ x58 ;
  assign n509 = ~n507 & n508 ;
  assign n561 = n509 ^ n507 ;
  assign n577 = n561 ^ n508 ;
  assign n578 = n577 ^ n507 ;
  assign n596 = ~n526 & n578 ;
  assign n588 = n499 & n503 ;
  assign n540 = n524 ^ n505 ;
  assign n537 = n505 & ~n511 ;
  assign n538 = n537 ^ n522 ;
  assign n506 = n499 & n505 ;
  assign n539 = n538 ^ n506 ;
  assign n541 = n540 ^ n539 ;
  assign n589 = n588 ^ n541 ;
  assign n517 = n499 & n502 ;
  assign n519 = n518 ^ n517 ;
  assign n515 = n502 & ~n511 ;
  assign n516 = n515 ^ n502 ;
  assign n520 = n519 ^ n516 ;
  assign n513 = n512 ^ n497 ;
  assign n514 = ~n504 & ~n513 ;
  assign n521 = n520 ^ n514 ;
  assign n542 = n541 ^ n521 ;
  assign n543 = n542 ^ n513 ;
  assign n536 = n499 & ~n504 ;
  assign n544 = n543 ^ n536 ;
  assign n590 = n589 ^ n544 ;
  assign n593 = n508 & ~n590 ;
  assign n594 = n593 ^ n589 ;
  assign n595 = ~n507 & n594 ;
  assign n597 = n596 ^ n595 ;
  assign n585 = n524 & n577 ;
  assign n564 = n542 ^ n517 ;
  assign n565 = n564 ^ n561 ;
  assign n527 = n503 & ~n511 ;
  assign n528 = n527 ^ n526 ;
  assign n1185 = n538 ^ n528 ;
  assign n1186 = n1185 ^ n526 ;
  assign n566 = n565 & ~n1186 ;
  assign n567 = n566 ^ n561 ;
  assign n569 = n1186 ^ n511 ;
  assign n568 = n522 ^ n515 ;
  assign n570 = n569 ^ n568 ;
  assign n571 = n570 ^ n523 ;
  assign n574 = n507 & ~n571 ;
  assign n575 = n574 ^ n523 ;
  assign n576 = ~n508 & n575 ;
  assign n580 = n1186 ^ n576 ;
  assign n579 = n578 ^ n576 ;
  assign n581 = n580 ^ n579 ;
  assign n582 = ~n567 & n581 ;
  assign n583 = n582 ^ n579 ;
  assign n535 = n508 ^ n507 ;
  assign n552 = n520 ^ n506 ;
  assign n553 = n552 ^ n515 ;
  assign n551 = n537 ^ n517 ;
  assign n554 = n553 ^ n551 ;
  assign n557 = n507 & n554 ;
  assign n558 = n557 ^ n551 ;
  assign n559 = n535 & n558 ;
  assign n584 = n583 ^ n559 ;
  assign n586 = n585 ^ n584 ;
  assign n545 = n544 ^ n518 ;
  assign n548 = n507 & ~n545 ;
  assign n549 = n548 ^ n518 ;
  assign n550 = n535 & n549 ;
  assign n587 = n586 ^ n550 ;
  assign n598 = n597 ^ n587 ;
  assign n529 = n528 ^ n521 ;
  assign n532 = ~n508 & ~n529 ;
  assign n533 = n532 ^ n528 ;
  assign n534 = ~n507 & ~n533 ;
  assign n599 = n598 ^ n534 ;
  assign n510 = n506 & n509 ;
  assign n600 = n599 ^ n510 ;
  assign n601 = n600 ^ x27 ;
  assign n602 = n601 ^ x121 ;
  assign n751 = n406 ^ n403 ;
  assign n720 = ~n710 & n751 ;
  assign n721 = n720 ^ n405 ;
  assign n722 = ~n602 & ~n721 ;
  assign n723 = n722 ^ n405 ;
  assign n724 = n496 & ~n723 ;
  assign n725 = n232 & n724 ;
  assign n2572 = n2571 ^ n725 ;
  assign n2573 = n2572 ^ x56 ;
  assign n732 = n406 & ~n602 ;
  assign n711 = n602 & n710 ;
  assign n756 = ~n404 & ~n711 ;
  assign n712 = n710 ^ n602 ;
  assign n757 = n756 ^ n712 ;
  assign n758 = ~n732 & ~n757 ;
  assign n759 = n758 ^ n757 ;
  assign n754 = n406 & n711 ;
  assign n755 = n754 ^ n711 ;
  assign n729 = n404 & ~n602 ;
  assign n2562 = n755 ^ n729 ;
  assign n728 = ~n321 & n711 ;
  assign n2555 = n758 ^ n728 ;
  assign n2556 = n2555 ^ n403 ;
  assign n735 = ~n405 & ~n602 ;
  assign n713 = n712 ^ n711 ;
  assign n736 = n735 ^ n713 ;
  assign n2557 = n2556 ^ n736 ;
  assign n2558 = n2557 ^ n728 ;
  assign n2559 = n496 & n2558 ;
  assign n2560 = n2559 ^ n2555 ;
  assign n744 = n321 & n712 ;
  assign n2561 = n2560 ^ n744 ;
  assign n2563 = n2562 ^ n2561 ;
  assign n2564 = n2563 ^ n2560 ;
  assign n2565 = ~n496 & n2564 ;
  assign n2566 = n2565 ^ n2561 ;
  assign n2567 = n232 & ~n2566 ;
  assign n2568 = n2567 ^ n2560 ;
  assign n2569 = n759 & n2568 ;
  assign n2574 = n2573 ^ n2569 ;
  assign n3444 = n2574 ^ x70 ;
  assign n3445 = n3443 & ~n3444 ;
  assign n3475 = n3445 ^ n3444 ;
  assign n4454 = n3475 ^ n3443 ;
  assign n4476 = n4454 ^ n3444 ;
  assign n2610 = n433 & n475 ;
  assign n2604 = n479 ^ n463 ;
  assign n2605 = n487 & ~n2604 ;
  assign n2598 = n432 ^ n426 ;
  assign n2599 = n2598 ^ n461 ;
  assign n2600 = n409 & ~n2599 ;
  assign n1319 = n487 ^ n409 ;
  assign n2593 = ~n461 & ~n1319 ;
  assign n2591 = n446 & n475 ;
  assign n2589 = n452 ^ n444 ;
  assign n2590 = n2589 ^ n457 ;
  assign n2592 = n2591 ^ n2590 ;
  assign n2594 = n2593 ^ n2592 ;
  assign n2601 = n2600 ^ n2594 ;
  assign n2602 = n411 & ~n2601 ;
  assign n1325 = ~n410 & n450 ;
  assign n1326 = n1325 ^ n432 ;
  assign n1327 = n409 & n1326 ;
  assign n2595 = n2594 ^ n1327 ;
  assign n2588 = n481 ^ x21 ;
  assign n2596 = n2595 ^ n2588 ;
  assign n2603 = n2602 ^ n2596 ;
  assign n2606 = n2605 ^ n2603 ;
  assign n2586 = n436 ^ n426 ;
  assign n2587 = ~n1319 & n2586 ;
  assign n2607 = n2606 ^ n2587 ;
  assign n2580 = n477 ^ n444 ;
  assign n2583 = n410 & n2580 ;
  assign n2584 = n2583 ^ n444 ;
  assign n2585 = n409 & n2584 ;
  assign n2608 = n2607 ^ n2585 ;
  assign n2578 = n438 ^ n433 ;
  assign n2579 = n410 & ~n2578 ;
  assign n2609 = n2608 ^ n2579 ;
  assign n2611 = n2610 ^ n2609 ;
  assign n2612 = n2611 ^ x91 ;
  assign n810 = n809 ^ n354 ;
  assign n811 = ~n399 & n810 ;
  assign n804 = n353 ^ n329 ;
  assign n805 = n804 ^ n350 ;
  assign n806 = n805 ^ n359 ;
  assign n807 = ~n322 & n806 ;
  assign n802 = n359 ^ n346 ;
  assign n803 = n802 ^ n331 ;
  assign n808 = n807 ^ n803 ;
  assign n812 = n811 ^ n808 ;
  assign n795 = n778 ^ n391 ;
  assign n796 = n795 ^ n346 ;
  assign n799 = n322 & n796 ;
  assign n800 = n799 ^ n346 ;
  assign n801 = ~n323 & n800 ;
  assign n813 = n812 ^ n801 ;
  assign n785 = n374 ^ n349 ;
  assign n814 = n813 ^ n785 ;
  assign n793 = n362 ^ n346 ;
  assign n794 = ~n370 & n793 ;
  assign n815 = n814 ^ n794 ;
  assign n786 = n785 ^ n399 ;
  assign n787 = n370 ^ n334 ;
  assign n790 = ~n785 & ~n787 ;
  assign n791 = n790 ^ n370 ;
  assign n792 = ~n786 & ~n791 ;
  assign n816 = n815 ^ n792 ;
  assign n817 = n816 ^ n393 ;
  assign n818 = n817 ^ x29 ;
  assign n784 = n324 & n783 ;
  assign n819 = n818 ^ n784 ;
  assign n2577 = n819 ^ x85 ;
  assign n1621 = n233 & ~n244 ;
  assign n1653 = n246 & ~n252 ;
  assign n1654 = n1621 & n1653 ;
  assign n1631 = n244 ^ n233 ;
  assign n1286 = n291 ^ n276 ;
  assign n1289 = ~n252 & n1286 ;
  assign n1290 = n1289 ^ n276 ;
  assign n1291 = n233 & n1290 ;
  assign n1632 = n1631 ^ n1291 ;
  assign n1296 = ~n233 & n291 ;
  assign n1297 = n1296 ^ n271 ;
  assign n1298 = n258 & n1297 ;
  assign n1299 = n1298 ^ n271 ;
  assign n1633 = n1632 ^ n1299 ;
  assign n1634 = n1633 ^ n287 ;
  assign n1635 = n1634 ^ n1268 ;
  assign n1282 = n233 & n274 ;
  assign n1283 = n1282 ^ n280 ;
  assign n1284 = n258 & n1283 ;
  assign n1285 = n1284 ^ n280 ;
  assign n1636 = n1635 ^ n1285 ;
  assign n1648 = n1647 ^ n1636 ;
  assign n1649 = n1648 ^ x5 ;
  assign n1624 = n1623 ^ n287 ;
  assign n1625 = n1624 ^ n288 ;
  assign n1628 = ~n233 & n1625 ;
  assign n1629 = n1628 ^ n288 ;
  assign n1630 = n258 & n1629 ;
  assign n1650 = n1649 ^ n1630 ;
  assign n1651 = n1650 ^ n1621 ;
  assign n1655 = n1654 ^ n1651 ;
  assign n2615 = n1655 ^ x78 ;
  assign n2634 = n165 & ~n1812 ;
  assign n2631 = n1832 ^ n175 ;
  assign n2626 = n164 ^ n134 ;
  assign n2627 = n2626 ^ n172 ;
  assign n2628 = n129 & n2627 ;
  assign n2632 = n2631 ^ n2628 ;
  assign n2624 = n1816 ^ n162 ;
  assign n2622 = n150 ^ n146 ;
  assign n2623 = ~n129 & n2622 ;
  assign n2625 = n2624 ^ n2623 ;
  assign n2629 = n2628 ^ n2625 ;
  assign n2630 = n130 & n2629 ;
  assign n2633 = n2632 ^ n2630 ;
  assign n2635 = n2634 ^ n2633 ;
  assign n2619 = ~n129 & n179 ;
  assign n2620 = n2619 ^ n175 ;
  assign n2621 = ~n130 & n2620 ;
  assign n2636 = n2635 ^ n2621 ;
  assign n2637 = n2636 ^ n1369 ;
  assign n2638 = n2637 ^ n1368 ;
  assign n2639 = n2638 ^ n195 ;
  assign n2640 = n2639 ^ x13 ;
  assign n2641 = n2640 ^ x108 ;
  assign n2642 = ~n2615 & ~n2641 ;
  assign n2643 = ~n2577 & n2642 ;
  assign n2644 = n2643 ^ n2642 ;
  assign n2645 = n2612 & n2644 ;
  assign n2646 = n2645 ^ n2644 ;
  assign n970 = x104 ^ x60 ;
  assign n969 = x122 ^ x34 ;
  assign n975 = x81 ^ x2 ;
  assign n977 = x64 ^ x26 ;
  assign n978 = n975 & n977 ;
  assign n979 = n978 ^ n975 ;
  assign n972 = x99 ^ x18 ;
  assign n973 = x90 ^ x10 ;
  assign n983 = n972 & ~n973 ;
  assign n984 = n983 ^ n972 ;
  assign n988 = n984 ^ n973 ;
  assign n989 = n979 & n988 ;
  assign n990 = n989 ^ n978 ;
  assign n987 = ~n973 & n978 ;
  assign n991 = n990 ^ n987 ;
  assign n976 = n973 & n975 ;
  assign n992 = n991 ^ n976 ;
  assign n982 = n972 & n977 ;
  assign n985 = n984 ^ n982 ;
  assign n993 = n992 ^ n985 ;
  assign n986 = ~n975 & n985 ;
  assign n994 = n993 ^ n986 ;
  assign n974 = n973 ^ n972 ;
  assign n980 = n979 ^ n976 ;
  assign n981 = ~n974 & n980 ;
  assign n995 = n994 ^ n981 ;
  assign n1007 = n995 ^ n989 ;
  assign n1001 = n988 ^ n972 ;
  assign n1005 = n975 & ~n1001 ;
  assign n1006 = n1005 ^ n990 ;
  assign n1008 = n1007 ^ n1006 ;
  assign n1061 = n1008 ^ n992 ;
  assign n1064 = n969 & n1061 ;
  assign n1065 = n1064 ^ n992 ;
  assign n1066 = n970 & n1065 ;
  assign n1044 = n977 ^ n975 ;
  assign n1045 = n1044 ^ n972 ;
  assign n1021 = n1045 ^ n975 ;
  assign n1024 = ~n973 & ~n1021 ;
  assign n1025 = n1024 ^ n975 ;
  assign n1026 = n974 & ~n1025 ;
  assign n1018 = n977 ^ n973 ;
  assign n1027 = n1026 ^ n1018 ;
  assign n1028 = ~n969 & n1027 ;
  assign n1068 = n1066 ^ n1028 ;
  assign n997 = n978 ^ n977 ;
  assign n1002 = n997 & ~n1001 ;
  assign n1049 = n1002 ^ n1001 ;
  assign n1050 = n1049 ^ n1005 ;
  assign n998 = n997 ^ n975 ;
  assign n999 = n983 & ~n998 ;
  assign n1046 = n999 ^ n991 ;
  assign n1047 = n1046 ^ n1045 ;
  assign n1051 = n1050 ^ n1047 ;
  assign n1009 = n1008 ^ n981 ;
  assign n1033 = n1009 ^ n980 ;
  assign n1052 = n1051 ^ n1033 ;
  assign n1035 = n984 & n997 ;
  assign n1043 = n1035 ^ n999 ;
  assign n1048 = n1047 ^ n1043 ;
  assign n1053 = n1052 ^ n1048 ;
  assign n1042 = n1018 ^ n1009 ;
  assign n1054 = n1053 ^ n1042 ;
  assign n1055 = n1054 ^ n1050 ;
  assign n1058 = ~n969 & ~n1055 ;
  assign n1059 = n1058 ^ n1050 ;
  assign n1060 = n970 & ~n1059 ;
  assign n1069 = n1068 ^ n1060 ;
  assign n1070 = n1069 ^ x37 ;
  assign n1000 = n999 ^ n992 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n1034 = n1033 ^ n1003 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1039 = n969 & n1036 ;
  assign n1029 = n988 & ~n998 ;
  assign n1030 = n1029 ^ n1028 ;
  assign n1040 = n1039 ^ n1030 ;
  assign n1041 = n970 & n1040 ;
  assign n1071 = n1070 ^ n1041 ;
  assign n971 = n970 ^ n969 ;
  assign n1004 = n1003 ^ n986 ;
  assign n1010 = n1009 ^ n1004 ;
  assign n996 = n995 ^ n986 ;
  assign n1011 = n1010 ^ n996 ;
  assign n1014 = ~n969 & ~n1011 ;
  assign n1015 = n1014 ^ n1010 ;
  assign n1016 = n971 & ~n1015 ;
  assign n1072 = n1071 ^ n1016 ;
  assign n2576 = n1072 ^ x102 ;
  assign n1552 = n637 ^ n618 ;
  assign n1555 = n1554 ^ n1552 ;
  assign n1556 = n1555 ^ n647 ;
  assign n1557 = n603 & ~n1556 ;
  assign n1558 = n1557 ^ n637 ;
  assign n1559 = ~n604 & n1558 ;
  assign n1548 = n679 ^ n657 ;
  assign n1549 = n1520 & n1548 ;
  assign n1538 = n645 ^ n641 ;
  assign n1539 = n1538 ^ n1521 ;
  assign n1540 = ~n656 & n1539 ;
  assign n1541 = n1540 ^ n698 ;
  assign n1543 = n699 ^ n632 ;
  assign n1544 = n1543 ^ n644 ;
  assign n1542 = ~n656 & n1521 ;
  assign n1545 = n1544 ^ n1542 ;
  assign n1546 = n1541 & n1545 ;
  assign n1525 = n643 & n1520 ;
  assign n1536 = n1535 ^ n1525 ;
  assign n1524 = n1523 ^ x63 ;
  assign n1537 = n1536 ^ n1524 ;
  assign n1547 = n1546 ^ n1537 ;
  assign n1550 = n1549 ^ n1547 ;
  assign n1519 = ~n605 & n636 ;
  assign n1551 = n1550 ^ n1519 ;
  assign n1560 = n1559 ^ n1551 ;
  assign n2685 = n1560 ^ x84 ;
  assign n2686 = ~n2576 & n2685 ;
  assign n2687 = n2686 ^ n2576 ;
  assign n3126 = n2646 & ~n2687 ;
  assign n2663 = n2577 & n2615 ;
  assign n2657 = n2577 & n2641 ;
  assign n2658 = n2657 ^ n2577 ;
  assign n2659 = n2658 ^ n2644 ;
  assign n2688 = n2663 ^ n2659 ;
  assign n2648 = n2641 ^ n2615 ;
  assign n2649 = n2641 ^ n2612 ;
  assign n2650 = n2648 & ~n2649 ;
  assign n2651 = n2650 ^ n2641 ;
  assign n2652 = n2577 & n2651 ;
  assign n2613 = ~n2577 & ~n2612 ;
  assign n2614 = n2613 ^ n2612 ;
  assign n2647 = n2646 ^ n2614 ;
  assign n2653 = n2652 ^ n2647 ;
  assign n2689 = n2688 ^ n2653 ;
  assign n2705 = n2685 ^ n2576 ;
  assign n2992 = ~n2689 & ~n2705 ;
  assign n2690 = n2689 ^ n2646 ;
  assign n2660 = n2612 & n2659 ;
  assign n2661 = n2660 ^ n2659 ;
  assign n2691 = n2690 ^ n2661 ;
  assign n2692 = n2691 ^ n2614 ;
  assign n2693 = n2692 ^ n2653 ;
  assign n3149 = n2686 & ~n2693 ;
  assign n3142 = n2661 ^ n2613 ;
  assign n2654 = n2612 & n2641 ;
  assign n2655 = n2577 & n2654 ;
  assign n2667 = n2655 ^ n2654 ;
  assign n2665 = n2657 ^ n2641 ;
  assign n2670 = n2667 ^ n2665 ;
  assign n2671 = n2670 ^ n2613 ;
  assign n2672 = ~n2615 & n2671 ;
  assign n2675 = n2672 ^ n2613 ;
  assign n2676 = n2675 ^ n2670 ;
  assign n2673 = n2672 ^ n2643 ;
  assign n2668 = n2667 ^ n2613 ;
  assign n2669 = n2668 ^ n2577 ;
  assign n2674 = n2673 ^ n2669 ;
  assign n2677 = n2676 ^ n2674 ;
  assign n2664 = n2663 ^ n2615 ;
  assign n2666 = n2665 ^ n2664 ;
  assign n2678 = n2677 ^ n2666 ;
  assign n2679 = n2678 ^ n2672 ;
  assign n2680 = n2679 ^ n2613 ;
  assign n2681 = n2680 ^ n2650 ;
  assign n2656 = n2655 ^ n2653 ;
  assign n2662 = n2661 ^ n2656 ;
  assign n2682 = n2681 ^ n2662 ;
  assign n2700 = n2682 ^ n2670 ;
  assign n2701 = n2700 ^ n2678 ;
  assign n2715 = n2701 ^ n2645 ;
  assign n3143 = n3142 ^ n2715 ;
  assign n2702 = n2701 ^ n2667 ;
  assign n3139 = n2702 ^ n2646 ;
  assign n3144 = n3143 ^ n3139 ;
  assign n3145 = ~n2685 & n3144 ;
  assign n3136 = n2680 ^ n2673 ;
  assign n3134 = n2671 ^ n2577 ;
  assign n3135 = ~n2685 & ~n3134 ;
  assign n3137 = n3136 ^ n3135 ;
  assign n3140 = n3139 ^ n3137 ;
  assign n3146 = n3145 ^ n3140 ;
  assign n3147 = n2576 & n3146 ;
  assign n3127 = n2669 ^ n2643 ;
  assign n3128 = n3127 ^ n2653 ;
  assign n3131 = n2685 & n3128 ;
  assign n3132 = n3131 ^ n2653 ;
  assign n3133 = n2576 & ~n3132 ;
  assign n3138 = n3137 ^ n3133 ;
  assign n3148 = n3147 ^ n3138 ;
  assign n3150 = n3149 ^ n3148 ;
  assign n3151 = ~n2992 & n3150 ;
  assign n3152 = ~n3126 & n3151 ;
  assign n2694 = n2660 ^ n2656 ;
  assign n3153 = n2694 ^ n2690 ;
  assign n3156 = ~n2685 & n3153 ;
  assign n3157 = n3156 ^ n2690 ;
  assign n3158 = ~n2576 & ~n3157 ;
  assign n3159 = n3152 & ~n3158 ;
  assign n3162 = n3159 ^ x30 ;
  assign n3125 = n2694 ^ n2692 ;
  assign n2697 = n2687 ^ n2685 ;
  assign n2698 = n2697 ^ n2576 ;
  assign n3160 = n2698 & n3159 ;
  assign n3161 = ~n3125 & n3160 ;
  assign n3163 = n3162 ^ n3161 ;
  assign n3360 = n3163 ^ x116 ;
  assign n1413 = n872 ^ n846 ;
  assign n1386 = n857 ^ n824 ;
  assign n1387 = n1386 ^ n880 ;
  assign n1388 = n1387 ^ n875 ;
  assign n1389 = n1388 ^ n841 ;
  assign n882 = n834 ^ n823 ;
  assign n883 = n882 ^ n842 ;
  assign n901 = n883 ^ n837 ;
  assign n1383 = n1382 ^ n901 ;
  assign n1384 = n1383 ^ n858 ;
  assign n1385 = n1384 ^ n853 ;
  assign n1390 = n1389 ^ n1385 ;
  assign n1391 = ~n861 & ~n1390 ;
  assign n1392 = n1391 ^ n1389 ;
  assign n1414 = n1413 ^ n1392 ;
  assign n919 = n918 ^ n872 ;
  assign n1412 = n861 & n919 ;
  assign n1415 = n1414 ^ n1412 ;
  assign n1416 = ~n893 & ~n1415 ;
  assign n881 = n880 ^ n836 ;
  assign n884 = n883 ^ n881 ;
  assign n867 = n837 ^ n832 ;
  assign n878 = n877 ^ n867 ;
  assign n885 = n884 ^ n878 ;
  assign n1404 = n885 ^ n856 ;
  assign n1405 = n1404 ^ n1386 ;
  assign n1406 = n822 & n1405 ;
  assign n1407 = n1406 ^ n874 ;
  assign n1408 = ~n861 & n1407 ;
  assign n1393 = n1386 ^ n878 ;
  assign n1394 = n1393 ^ n875 ;
  assign n1395 = n872 ^ n861 ;
  assign n1396 = n1395 ^ n917 ;
  assign n1397 = ~n1394 & n1396 ;
  assign n1398 = n1397 ^ n872 ;
  assign n1399 = n1394 ^ n917 ;
  assign n1400 = n1399 ^ n822 ;
  assign n1401 = n1398 & ~n1400 ;
  assign n1402 = n1401 ^ n1394 ;
  assign n1403 = n1402 ^ n1392 ;
  assign n1409 = n1408 ^ n1403 ;
  assign n898 = n854 & ~n861 ;
  assign n899 = n898 ^ n878 ;
  assign n900 = ~n893 & n899 ;
  assign n1410 = n1409 ^ n900 ;
  assign n1411 = n1410 ^ x31 ;
  assign n1417 = n1416 ^ n1411 ;
  assign n1657 = n1417 ^ x75 ;
  assign n1656 = n1655 ^ x116 ;
  assign n1210 = n597 ^ n585 ;
  assign n1204 = n536 ^ n521 ;
  assign n1201 = n588 ^ n506 ;
  assign n1202 = n1201 ^ n536 ;
  assign n1203 = n508 & n1202 ;
  assign n1205 = n1204 ^ n1203 ;
  assign n1206 = n507 & n1205 ;
  assign n1207 = n1206 ^ n561 ;
  assign n1193 = n570 ^ n518 ;
  assign n1194 = n1193 ^ n561 ;
  assign n1195 = n578 ^ n543 ;
  assign n1198 = ~n1193 & n1195 ;
  assign n1199 = n1198 ^ n543 ;
  assign n1200 = n1194 & n1199 ;
  assign n1208 = n1207 ^ n1200 ;
  assign n1209 = n1208 ^ n517 ;
  assign n1211 = n1210 ^ n1209 ;
  assign n928 = ~n508 & n540 ;
  assign n929 = n928 ^ n541 ;
  assign n930 = ~n507 & n929 ;
  assign n1212 = n1211 ^ n930 ;
  assign n1187 = n1186 ^ n528 ;
  assign n1190 = ~n507 & ~n1187 ;
  assign n1191 = n1190 ^ n528 ;
  assign n1192 = n535 & ~n1191 ;
  assign n1213 = n1212 ^ n1192 ;
  assign n1214 = n1213 ^ x39 ;
  assign n940 = n523 ^ n515 ;
  assign n1182 = n508 & n940 ;
  assign n1183 = n1182 ^ n517 ;
  assign n1184 = ~n507 & n1183 ;
  assign n1215 = n1214 ^ n1184 ;
  assign n1599 = n1215 ^ x70 ;
  assign n1231 = n1054 ^ n992 ;
  assign n1232 = n1231 ^ n1050 ;
  assign n1233 = n1232 ^ n1029 ;
  assign n1234 = ~n969 & ~n1233 ;
  assign n1235 = n1234 ^ n1050 ;
  assign n1236 = ~n970 & ~n1235 ;
  assign n1610 = n1236 ^ x55 ;
  assign n1604 = n1027 ^ n996 ;
  assign n1605 = n970 & ~n1604 ;
  assign n1606 = n1605 ^ n996 ;
  assign n1611 = n1610 ^ n1606 ;
  assign n1607 = n1606 ^ n1010 ;
  assign n1600 = n1029 ^ n1008 ;
  assign n1601 = n1600 ^ n1010 ;
  assign n1602 = n1601 ^ n1036 ;
  assign n1603 = ~n970 & n1602 ;
  assign n1608 = n1607 ^ n1603 ;
  assign n1609 = n969 & n1608 ;
  assign n1612 = n1611 ^ n1609 ;
  assign n1613 = n1612 ^ x93 ;
  assign n1614 = ~n1599 & ~n1613 ;
  assign n1561 = n1560 ^ x76 ;
  assign n1578 = n343 ^ n326 ;
  assign n1579 = n1578 ^ n350 ;
  assign n1586 = n1579 ^ n336 ;
  assign n1580 = n1579 ^ n322 ;
  assign n1581 = n324 & n1580 ;
  assign n1582 = n1581 ^ n322 ;
  assign n1583 = n1579 ^ n378 ;
  assign n1584 = n1583 ^ n354 ;
  assign n1585 = n1582 & n1584 ;
  assign n1587 = n1586 ^ n1585 ;
  assign n1569 = n1568 ^ n778 ;
  assign n1570 = n322 & n1569 ;
  assign n1590 = n1587 ^ n1570 ;
  assign n1591 = n324 & n1590 ;
  assign n1588 = n1587 ^ n1577 ;
  assign n1592 = n1591 ^ n1588 ;
  assign n1562 = n780 ^ n343 ;
  assign n1565 = n323 & n1562 ;
  assign n1566 = n1565 ^ n780 ;
  assign n1567 = ~n322 & n1566 ;
  assign n1593 = n1592 ^ n1567 ;
  assign n1594 = n1593 ^ n393 ;
  assign n1595 = n1594 ^ x47 ;
  assign n1596 = n1595 ^ x118 ;
  assign n1597 = ~n1561 & n1596 ;
  assign n1663 = n1597 ^ n1596 ;
  assign n1681 = n1614 & n1663 ;
  assign n1617 = n1614 ^ n1599 ;
  assign n1660 = n1617 ^ n1613 ;
  assign n1664 = ~n1660 & n1663 ;
  assign n1682 = n1681 ^ n1664 ;
  assign n1615 = n1614 ^ n1613 ;
  assign n1679 = ~n1615 & n1663 ;
  assign n1680 = n1679 ^ n1663 ;
  assign n1683 = n1682 ^ n1680 ;
  assign n1598 = n1597 ^ n1561 ;
  assign n1665 = n1598 ^ n1596 ;
  assign n1671 = ~n1660 & n1665 ;
  assign n1670 = ~n1615 & n1665 ;
  assign n1672 = n1671 ^ n1670 ;
  assign n1666 = n1614 & n1665 ;
  assign n1669 = n1666 ^ n1665 ;
  assign n1673 = n1672 ^ n1669 ;
  assign n1684 = n1683 ^ n1673 ;
  assign n2296 = ~n1656 & n1684 ;
  assign n2297 = n2296 ^ n1673 ;
  assign n2298 = n1657 & n2297 ;
  assign n1618 = ~n1598 & ~n1617 ;
  assign n1678 = n1618 ^ n1617 ;
  assign n1685 = n1684 ^ n1678 ;
  assign n1668 = n1597 & ~n1615 ;
  assign n1686 = n1685 ^ n1668 ;
  assign n1676 = n1597 & n1614 ;
  assign n1677 = n1676 ^ n1597 ;
  assign n1687 = n1686 ^ n1677 ;
  assign n1716 = n1687 ^ n1618 ;
  assign n1717 = n1716 ^ n1686 ;
  assign n1720 = ~n1656 & n1717 ;
  assign n1721 = n1720 ^ n1686 ;
  assign n1722 = n1657 & ~n1721 ;
  assign n2299 = n2298 ^ n1722 ;
  assign n1731 = n1683 ^ n1679 ;
  assign n1616 = ~n1598 & ~n1615 ;
  assign n1619 = n1618 ^ n1616 ;
  assign n1620 = n1619 ^ n1598 ;
  assign n2271 = n1731 ^ n1620 ;
  assign n2262 = ~n1598 & n1614 ;
  assign n2263 = n2262 ^ n1668 ;
  assign n2268 = n1657 & n2263 ;
  assign n2269 = n2268 ^ n1682 ;
  assign n2270 = ~n1656 & n2269 ;
  assign n2272 = n2271 ^ n2270 ;
  assign n2259 = n1687 ^ n1679 ;
  assign n2258 = n1673 ^ n1620 ;
  assign n2260 = n2259 ^ n2258 ;
  assign n2261 = n2260 ^ n1685 ;
  assign n2273 = n2272 ^ n2261 ;
  assign n2274 = n2273 ^ n2270 ;
  assign n2275 = ~n1656 & n2274 ;
  assign n2276 = n2275 ^ n2272 ;
  assign n2300 = n2299 ^ n2276 ;
  assign n1699 = n1656 & n1672 ;
  assign n1700 = n1699 ^ n1671 ;
  assign n1701 = n1657 & n1700 ;
  assign n2301 = n2300 ^ n1701 ;
  assign n2302 = n2301 ^ x6 ;
  assign n1658 = n1657 ^ n1656 ;
  assign n2284 = n1615 ^ n1598 ;
  assign n2281 = n1671 ^ n1618 ;
  assign n2282 = n2281 ^ n1679 ;
  assign n2279 = n1676 ^ n1670 ;
  assign n2280 = n2279 ^ n2262 ;
  assign n2283 = n2282 ^ n2280 ;
  assign n2285 = n2284 ^ n2283 ;
  assign n2277 = n1613 ^ n1599 ;
  assign n2278 = n2277 ^ n1561 ;
  assign n2286 = n2285 ^ n2278 ;
  assign n2287 = ~n1656 & n2286 ;
  assign n2288 = n2287 ^ n2286 ;
  assign n2289 = n2288 ^ n2270 ;
  assign n2290 = n2289 ^ n2276 ;
  assign n2291 = n1658 & ~n2290 ;
  assign n2303 = n2302 ^ n2291 ;
  assign n3361 = n2303 ^ x94 ;
  assign n3362 = n3360 & ~n3361 ;
  assign n3363 = n3362 ^ n3360 ;
  assign n3364 = n3363 ^ n3361 ;
  assign n1335 = n1334 ^ n439 ;
  assign n1336 = n487 & ~n1335 ;
  assign n1331 = n444 ^ n423 ;
  assign n1332 = n410 & n1331 ;
  assign n1328 = n1327 ^ n481 ;
  assign n1329 = n1328 ^ n474 ;
  assign n1330 = n1329 ^ x7 ;
  assign n1333 = n1332 ^ n1330 ;
  assign n1337 = n1336 ^ n1333 ;
  assign n1320 = n493 & ~n1319 ;
  assign n1338 = n1337 ^ n1320 ;
  assign n1312 = n490 ^ n458 ;
  assign n1311 = n1310 ^ n458 ;
  assign n1313 = n1312 ^ n1311 ;
  assign n1316 = n410 & ~n1313 ;
  assign n1317 = n1316 ^ n1312 ;
  assign n1318 = n409 & n1317 ;
  assign n1339 = n1338 ^ n1318 ;
  assign n1950 = n1339 ^ x65 ;
  assign n2095 = n2094 ^ x72 ;
  assign n2140 = n1950 & n2095 ;
  assign n2141 = n2140 ^ n2095 ;
  assign n2147 = n2141 ^ n1950 ;
  assign n1237 = n1236 ^ x57 ;
  assign n1217 = n1033 ^ n987 ;
  assign n1218 = n1217 ^ n1052 ;
  assign n1219 = ~n969 & n1218 ;
  assign n1220 = n1219 ^ n1052 ;
  assign n1222 = n1220 ^ n1047 ;
  assign n1221 = n1220 ^ n1006 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1226 = n969 & n1223 ;
  assign n1227 = n1226 ^ n1222 ;
  assign n1228 = n971 & n1227 ;
  assign n1229 = n1228 ^ n1220 ;
  assign n1230 = ~n1043 & ~n1229 ;
  assign n1238 = n1237 ^ n1230 ;
  assign n2009 = n1238 ^ x106 ;
  assign n2018 = n570 ^ n552 ;
  assign n2021 = n589 ^ n536 ;
  assign n2022 = n2021 ^ n517 ;
  assign n2019 = n588 ^ n552 ;
  assign n2020 = n2019 ^ n570 ;
  assign n2023 = n2022 ^ n2020 ;
  assign n2024 = n2023 ^ n508 ;
  assign n2025 = n2024 ^ n2020 ;
  assign n2026 = ~n535 & n2025 ;
  assign n2027 = n2026 ^ n535 ;
  assign n2028 = n2018 & ~n2027 ;
  assign n2029 = n2028 ^ n2020 ;
  assign n2030 = n2025 ^ n507 ;
  assign n2031 = n2030 ^ n2026 ;
  assign n2032 = ~n2029 & n2031 ;
  assign n2033 = n2032 ^ n2020 ;
  assign n2042 = n2033 ^ n507 ;
  assign n931 = n537 ^ n526 ;
  assign n934 = n507 & ~n931 ;
  assign n935 = n934 ^ n526 ;
  assign n936 = ~n508 & ~n935 ;
  assign n2043 = n2042 ^ n936 ;
  assign n2044 = n2043 ^ n576 ;
  assign n952 = n509 & ~n570 ;
  assign n953 = n952 ^ n596 ;
  assign n2045 = n2044 ^ n953 ;
  assign n2046 = n2045 ^ n550 ;
  assign n2047 = n2046 ^ n1192 ;
  assign n2034 = n2033 ^ n520 ;
  assign n2035 = n2034 ^ n541 ;
  assign n2036 = n2035 ^ n2033 ;
  assign n2039 = ~n508 & ~n2036 ;
  assign n2040 = n2039 ^ n2033 ;
  assign n2041 = n535 & ~n2040 ;
  assign n2048 = n2047 ^ n2041 ;
  assign n2017 = n509 & n589 ;
  assign n2049 = n2048 ^ n2017 ;
  assign n2010 = n578 ^ n568 ;
  assign n2011 = n561 ^ n518 ;
  assign n2014 = ~n568 & n2011 ;
  assign n2015 = n2014 ^ n561 ;
  assign n2016 = n2010 & ~n2015 ;
  assign n2050 = n2049 ^ n2016 ;
  assign n2051 = n2050 ^ n510 ;
  assign n2052 = n2051 ^ x49 ;
  assign n2053 = n2052 ^ x89 ;
  assign n2054 = n2009 & n2053 ;
  assign n2055 = n2054 ^ n2009 ;
  assign n2056 = n2055 ^ n2053 ;
  assign n2058 = n2056 ^ n2009 ;
  assign n1959 = n701 ^ n662 ;
  assign n1958 = n1743 ^ n636 ;
  assign n1960 = n1959 ^ n1958 ;
  assign n1961 = ~n603 & ~n1960 ;
  assign n1962 = n1961 ^ n1959 ;
  assign n1965 = n1962 ^ n1536 ;
  assign n1966 = n1965 ^ n1764 ;
  assign n1967 = n1966 ^ n688 ;
  assign n1954 = n678 ^ n647 ;
  assign n1955 = n1954 ^ n1752 ;
  assign n1956 = n1955 ^ n1760 ;
  assign n1957 = n603 & n1956 ;
  assign n1963 = n1962 ^ n1957 ;
  assign n1964 = ~n604 & ~n1963 ;
  assign n1968 = n1967 ^ n1964 ;
  assign n1952 = n699 ^ n637 ;
  assign n1953 = ~n605 & n1952 ;
  assign n1969 = n1968 ^ n1953 ;
  assign n1970 = n1969 ^ n707 ;
  assign n1971 = n1970 ^ x41 ;
  assign n1951 = ~n656 & n679 ;
  assign n1972 = n1971 ^ n1951 ;
  assign n1973 = n1972 ^ x115 ;
  assign n2007 = n2006 ^ x104 ;
  assign n2008 = ~n1973 & ~n2007 ;
  assign n2064 = n2008 ^ n2007 ;
  assign n2097 = n2064 ^ n1973 ;
  assign n2098 = n2097 ^ n2007 ;
  assign n2100 = n2058 & ~n2098 ;
  assign n2099 = n2055 & ~n2098 ;
  assign n2907 = n2100 ^ n2099 ;
  assign n2908 = ~n2147 & n2907 ;
  assign n2122 = ~n2056 & ~n2098 ;
  assign n2123 = n2122 ^ n2056 ;
  assign n2117 = n2058 & ~n2097 ;
  assign n2118 = n2117 ^ n2058 ;
  assign n2059 = n2008 & n2058 ;
  assign n2101 = n2100 ^ n2059 ;
  assign n2119 = n2118 ^ n2101 ;
  assign n2114 = n2055 & ~n2064 ;
  assign n2065 = n2054 & ~n2064 ;
  assign n2115 = n2114 ^ n2065 ;
  assign n2116 = n2115 ^ n2064 ;
  assign n2120 = n2119 ^ n2116 ;
  assign n2057 = n2008 & ~n2056 ;
  assign n2121 = n2120 ^ n2057 ;
  assign n2124 = n2123 ^ n2121 ;
  assign n3389 = ~n2095 & n2124 ;
  assign n2881 = n2122 ^ n2057 ;
  assign n3382 = n2881 ^ n2119 ;
  assign n3379 = n2114 ^ n2057 ;
  assign n3380 = n3379 ^ n2064 ;
  assign n3381 = ~n2095 & ~n3380 ;
  assign n3383 = n3382 ^ n3381 ;
  assign n2096 = n2095 ^ n1950 ;
  assign n2061 = n2008 & n2055 ;
  assign n2062 = n2061 ^ n2008 ;
  assign n2060 = n2059 ^ n2057 ;
  assign n2063 = n2062 ^ n2060 ;
  assign n3368 = n2114 ^ n2063 ;
  assign n3366 = n1973 & n2009 ;
  assign n3367 = n2095 & n3366 ;
  assign n3369 = n3368 ^ n3367 ;
  assign n2105 = n2055 & ~n2097 ;
  assign n2125 = n2117 ^ n2105 ;
  assign n3370 = n3369 ^ n2125 ;
  assign n2129 = n2065 ^ n2054 ;
  assign n2126 = n2125 ^ n2097 ;
  assign n2127 = n2126 ^ n2124 ;
  assign n2128 = n2127 ^ n2063 ;
  assign n2130 = n2129 ^ n2128 ;
  assign n2131 = n2130 ^ n2061 ;
  assign n2132 = n2131 ^ n2127 ;
  assign n3371 = n3370 ^ n2132 ;
  assign n3372 = n3371 ^ n3369 ;
  assign n3375 = n2095 & n3372 ;
  assign n3376 = n3375 ^ n3369 ;
  assign n3377 = n2096 & n3376 ;
  assign n3378 = n3377 ^ n3369 ;
  assign n3384 = n3383 ^ n3378 ;
  assign n3387 = n3384 ^ n2059 ;
  assign n3388 = n3387 ^ n3378 ;
  assign n3390 = n3389 ^ n3388 ;
  assign n3391 = ~n1950 & n3390 ;
  assign n2875 = n2131 ^ n2100 ;
  assign n2878 = ~n2095 & ~n2875 ;
  assign n2879 = n2878 ^ n2100 ;
  assign n2880 = n1950 & n2879 ;
  assign n3385 = n3384 ^ n2880 ;
  assign n2110 = ~n2095 & n2105 ;
  assign n2102 = n2101 ^ n2099 ;
  assign n2103 = n2095 & n2102 ;
  assign n2104 = n2103 ^ n2101 ;
  assign n2111 = n2110 ^ n2104 ;
  assign n2112 = ~n2096 & n2111 ;
  assign n2113 = n2112 ^ n2104 ;
  assign n3386 = n3385 ^ n2113 ;
  assign n3392 = n3391 ^ n3386 ;
  assign n2153 = n2119 & ~n2147 ;
  assign n3393 = n3392 ^ n2153 ;
  assign n2161 = ~n2120 & n2141 ;
  assign n3394 = n3393 ^ n2161 ;
  assign n2158 = n2140 ^ n1950 ;
  assign n3365 = ~n2127 & n2158 ;
  assign n3395 = n3394 ^ n3365 ;
  assign n3396 = ~n2908 & ~n3395 ;
  assign n3397 = n3396 ^ x14 ;
  assign n3398 = n3397 ^ x101 ;
  assign n1741 = n601 ^ x113 ;
  assign n1772 = n1771 ^ x123 ;
  assign n1856 = n1741 & n1772 ;
  assign n1789 = n852 ^ n825 ;
  assign n1790 = n1789 ^ n841 ;
  assign n1791 = ~n822 & n1790 ;
  assign n1792 = n1791 ^ n858 ;
  assign n1793 = n893 & n1792 ;
  assign n890 = ~n822 & ~n885 ;
  assign n891 = n890 ^ n878 ;
  assign n892 = ~n861 & n891 ;
  assign n1783 = n892 ^ n858 ;
  assign n1784 = n1783 ^ n1402 ;
  assign n1785 = n1784 ^ n1408 ;
  assign n1786 = n1785 ^ x43 ;
  assign n1776 = n1383 ^ n880 ;
  assign n1774 = n854 ^ n851 ;
  assign n1775 = n1774 ^ n1382 ;
  assign n1777 = n1776 ^ n1775 ;
  assign n1780 = n861 & ~n1777 ;
  assign n1781 = n1780 ^ n1775 ;
  assign n1782 = ~n893 & n1781 ;
  assign n1787 = n1786 ^ n1782 ;
  assign n1773 = n822 & ~n847 ;
  assign n1788 = n1787 ^ n1773 ;
  assign n1794 = n1793 ^ n1788 ;
  assign n1795 = n1794 ^ x80 ;
  assign n1796 = n495 ^ x99 ;
  assign n1797 = n1795 & n1796 ;
  assign n1858 = n1797 ^ n1796 ;
  assign n1859 = n1858 ^ n1795 ;
  assign n1860 = n1859 ^ n1796 ;
  assign n1802 = ~n969 & n1053 ;
  assign n1803 = n1802 ^ n1052 ;
  assign n1807 = n1803 ^ n1066 ;
  assign n1808 = n1807 ^ n1060 ;
  assign n1809 = n1808 ^ x51 ;
  assign n1801 = n1043 ^ n1007 ;
  assign n1804 = n1803 ^ n1801 ;
  assign n1798 = n1029 ^ n1007 ;
  assign n1799 = n1798 ^ n1217 ;
  assign n1800 = ~n969 & n1799 ;
  assign n1805 = n1804 ^ n1800 ;
  assign n1806 = n970 & ~n1805 ;
  assign n1810 = n1809 ^ n1806 ;
  assign n1811 = n1810 ^ x81 ;
  assign n1842 = n1841 ^ x90 ;
  assign n1843 = ~n1811 & n1842 ;
  assign n1864 = n1843 ^ n1811 ;
  assign n1885 = n1860 & ~n1864 ;
  assign n1847 = n1843 ^ n1842 ;
  assign n1848 = n1847 ^ n1811 ;
  assign n1868 = n1848 & n1858 ;
  assign n1908 = n1885 ^ n1868 ;
  assign n3422 = n1856 & n1908 ;
  assign n1878 = n1848 & ~n1859 ;
  assign n1865 = n1797 & ~n1864 ;
  assign n1890 = n1878 ^ n1865 ;
  assign n1849 = n1797 & n1848 ;
  assign n1891 = n1890 ^ n1849 ;
  assign n1892 = n1891 ^ n1848 ;
  assign n1869 = n1868 ^ n1865 ;
  assign n1893 = n1892 ^ n1869 ;
  assign n1886 = n1885 ^ n1865 ;
  assign n1875 = ~n1859 & ~n1864 ;
  assign n1884 = n1875 ^ n1864 ;
  assign n1887 = n1886 ^ n1884 ;
  assign n1922 = n1893 ^ n1887 ;
  assign n2869 = ~n1772 & ~n1922 ;
  assign n2870 = n2869 ^ n1893 ;
  assign n2871 = n1741 & n2870 ;
  assign n1944 = n1856 ^ n1741 ;
  assign n1945 = n1849 & n1944 ;
  assign n1910 = n1772 ^ n1741 ;
  assign n1861 = n1847 & n1860 ;
  assign n1894 = n1893 ^ n1861 ;
  assign n1941 = n1772 & n1894 ;
  assign n1942 = n1941 ^ n1861 ;
  assign n1943 = n1910 & n1942 ;
  assign n1946 = n1945 ^ n1943 ;
  assign n1857 = n1856 ^ n1772 ;
  assign n3416 = n1857 & n1869 ;
  assign n2848 = n1857 ^ n1741 ;
  assign n1889 = n1885 ^ n1860 ;
  assign n1895 = n1894 ^ n1889 ;
  assign n1877 = n1875 ^ n1849 ;
  assign n1879 = n1878 ^ n1877 ;
  assign n1876 = n1875 ^ n1861 ;
  assign n1880 = n1879 ^ n1876 ;
  assign n1871 = n1796 ^ n1795 ;
  assign n1872 = n1871 ^ n1811 ;
  assign n1873 = n1872 ^ n1842 ;
  assign n1874 = n1811 & n1873 ;
  assign n1881 = n1880 ^ n1874 ;
  assign n1882 = n1881 ^ n1868 ;
  assign n1883 = n1882 ^ n1858 ;
  assign n1888 = n1887 ^ n1883 ;
  assign n1896 = n1895 ^ n1888 ;
  assign n1897 = n1896 ^ n1876 ;
  assign n1866 = n1865 ^ n1797 ;
  assign n1844 = n1797 & n1843 ;
  assign n1850 = n1849 ^ n1844 ;
  assign n1867 = n1866 ^ n1850 ;
  assign n1870 = n1869 ^ n1867 ;
  assign n1898 = n1897 ^ n1870 ;
  assign n1899 = n1898 ^ n1873 ;
  assign n1900 = n1899 ^ n1894 ;
  assign n1901 = n1900 ^ n1867 ;
  assign n3413 = n1901 ^ n1896 ;
  assign n3414 = ~n2848 & ~n3413 ;
  assign n3409 = n1857 & n1876 ;
  assign n3406 = n1888 ^ n1844 ;
  assign n2856 = n1901 & n1944 ;
  assign n3407 = n3406 ^ n2856 ;
  assign n2831 = n1895 ^ n1881 ;
  assign n3400 = n2831 ^ n1867 ;
  assign n1911 = n1890 ^ n1887 ;
  assign n1912 = n1772 & ~n1911 ;
  assign n1913 = n1912 ^ n1890 ;
  assign n3399 = n1913 ^ n1868 ;
  assign n3401 = n3400 ^ n3399 ;
  assign n3402 = n3401 ^ n1913 ;
  assign n3403 = n1772 & n3402 ;
  assign n3404 = n3403 ^ n3399 ;
  assign n3408 = n3407 ^ n3404 ;
  assign n3410 = n3409 ^ n3408 ;
  assign n3411 = n1910 & ~n3410 ;
  assign n2849 = n1893 & ~n2848 ;
  assign n3405 = n3404 ^ n2849 ;
  assign n3412 = n3411 ^ n3405 ;
  assign n3415 = n3414 ^ n3412 ;
  assign n3417 = n3416 ^ n3415 ;
  assign n3418 = ~n1946 & ~n3417 ;
  assign n3419 = ~n2871 & n3418 ;
  assign n3420 = ~n1878 & n3419 ;
  assign n3421 = n3420 ^ x22 ;
  assign n3424 = n3422 ^ n3421 ;
  assign n3425 = n3424 ^ x83 ;
  assign n3426 = ~n3398 & ~n3425 ;
  assign n3435 = n3426 ^ n3425 ;
  assign n3436 = n3364 & ~n3435 ;
  assign n3429 = n3362 ^ n3361 ;
  assign n3427 = n3426 ^ n3398 ;
  assign n3430 = n3427 ^ n3425 ;
  assign n3431 = ~n3429 & ~n3430 ;
  assign n3457 = n3436 ^ n3431 ;
  assign n3434 = ~n3427 & ~n3429 ;
  assign n3437 = n3436 ^ n3434 ;
  assign n3433 = ~n3360 & n3425 ;
  assign n3438 = n3437 ^ n3433 ;
  assign n3432 = n3431 ^ n3364 ;
  assign n3439 = n3438 ^ n3432 ;
  assign n3428 = n3364 & ~n3427 ;
  assign n3440 = n3439 ^ n3428 ;
  assign n3458 = n3457 ^ n3440 ;
  assign n3459 = n3458 ^ n3432 ;
  assign n3496 = n3459 ^ n3434 ;
  assign n3497 = n3496 ^ n3457 ;
  assign n3441 = n3426 & ~n3429 ;
  assign n3442 = n3441 ^ n3440 ;
  assign n3468 = n3442 ^ n3360 ;
  assign n3498 = n3497 ^ n3468 ;
  assign n4477 = n3498 ^ n3459 ;
  assign n4478 = n4476 & ~n4477 ;
  assign n3499 = n3445 & ~n3498 ;
  assign n3469 = n3468 ^ n3427 ;
  assign n3465 = n3398 ^ n3360 ;
  assign n3466 = n3465 ^ n3458 ;
  assign n3447 = n3361 ^ n3360 ;
  assign n3448 = n3447 ^ n3425 ;
  assign n3454 = ~n3360 & n3398 ;
  assign n3455 = n3454 ^ n3435 ;
  assign n3463 = n3455 ^ n3425 ;
  assign n3464 = n3448 & n3463 ;
  assign n3467 = n3466 ^ n3464 ;
  assign n3470 = n3469 ^ n3467 ;
  assign n3471 = n3470 ^ n3363 ;
  assign n3461 = n3363 & ~n3430 ;
  assign n3452 = n3362 & ~n3435 ;
  assign n3453 = n3452 ^ n3431 ;
  assign n3456 = n3455 ^ n3453 ;
  assign n3460 = n3459 ^ n3456 ;
  assign n3462 = n3461 ^ n3460 ;
  assign n3472 = n3471 ^ n3462 ;
  assign n3473 = n3472 ^ n3440 ;
  assign n3449 = n3448 ^ n3433 ;
  assign n3450 = ~n3398 & ~n3449 ;
  assign n3451 = n3450 ^ n3398 ;
  assign n3474 = n3473 ^ n3451 ;
  assign n3489 = n3474 ^ n3472 ;
  assign n3490 = n3489 ^ n3457 ;
  assign n3491 = n3457 ^ n3444 ;
  assign n3492 = n3491 ^ n3457 ;
  assign n3493 = ~n3490 & n3492 ;
  assign n3494 = n3493 ^ n3457 ;
  assign n3495 = ~n3443 & n3494 ;
  assign n3500 = n3499 ^ n3495 ;
  assign n4479 = n4478 ^ n3500 ;
  assign n3507 = n3470 ^ n3461 ;
  assign n3508 = n3507 ^ n3496 ;
  assign n4461 = n3444 & n3508 ;
  assign n4462 = n4461 ^ n3496 ;
  assign n4480 = n4479 ^ n4462 ;
  assign n3517 = n3472 ^ n3452 ;
  assign n4481 = n4480 ^ n3517 ;
  assign n3486 = n3445 & ~n3462 ;
  assign n4482 = n4481 ^ n3486 ;
  assign n4483 = n4482 ^ n402 ;
  assign n4484 = n4483 ^ n3517 ;
  assign n3485 = n3362 & ~n3430 ;
  assign n4468 = n3517 ^ n3485 ;
  assign n3518 = n3517 ^ n3362 ;
  assign n3516 = n3489 ^ n3485 ;
  assign n3519 = n3518 ^ n3516 ;
  assign n4469 = n4468 ^ n3519 ;
  assign n4470 = n4469 ^ n4468 ;
  assign n4471 = n4468 ^ n3444 ;
  assign n4472 = n4471 ^ n4468 ;
  assign n4473 = n4470 & n4472 ;
  assign n4474 = n4473 ^ n4468 ;
  assign n4475 = n3443 & ~n4474 ;
  assign n4485 = n4484 ^ n4475 ;
  assign n4466 = n3517 ^ n3474 ;
  assign n4467 = ~n3444 & ~n4466 ;
  assign n4486 = n4485 ^ n4467 ;
  assign n4460 = n3441 ^ n3439 ;
  assign n4463 = n4462 ^ n4460 ;
  assign n4456 = n3441 ^ n3433 ;
  assign n4457 = n4456 ^ n3432 ;
  assign n4458 = n4457 ^ n3428 ;
  assign n4459 = ~n3444 & n4458 ;
  assign n4464 = n4463 ^ n4459 ;
  assign n4465 = n3443 & n4464 ;
  assign n4487 = n4486 ^ n4465 ;
  assign n4455 = n3497 & n4454 ;
  assign n4488 = n4487 ^ n4455 ;
  assign n4453 = n3470 & ~n3475 ;
  assign n4489 = n4488 ^ n4453 ;
  assign n4490 = n4489 ^ x115 ;
  assign n3643 = n2881 ^ n2115 ;
  assign n3644 = n3643 ^ n2061 ;
  assign n3647 = ~n2095 & n3644 ;
  assign n3648 = n3647 ^ n2061 ;
  assign n3649 = n2096 & n3648 ;
  assign n2899 = n2125 ^ n2059 ;
  assign n2900 = ~n2095 & n2899 ;
  assign n2901 = n2900 ^ n2125 ;
  assign n3641 = n2908 ^ n2901 ;
  assign n2909 = n2124 ^ n2119 ;
  assign n2910 = n2909 ^ n2100 ;
  assign n2911 = ~n2095 & n2910 ;
  assign n2912 = n2911 ^ n2100 ;
  assign n2913 = n2096 & n2912 ;
  assign n2914 = n2913 ^ n2161 ;
  assign n3642 = n3641 ^ n2914 ;
  assign n3650 = n3649 ^ n3642 ;
  assign n3638 = n1950 & n2099 ;
  assign n3639 = n3638 ^ n2128 ;
  assign n3640 = n2095 & ~n3639 ;
  assign n3651 = n3650 ^ n3640 ;
  assign n3628 = n2125 ^ n2060 ;
  assign n3629 = n3628 ^ n2065 ;
  assign n3630 = n3629 ^ n2909 ;
  assign n3631 = ~n2095 & n3630 ;
  assign n3626 = n2909 ^ n2901 ;
  assign n3632 = n3631 ^ n3626 ;
  assign n3633 = ~n1950 & n3632 ;
  assign n3652 = n3651 ^ n3633 ;
  assign n3653 = n3652 ^ n2130 ;
  assign n3654 = n3653 ^ x58 ;
  assign n3625 = ~n2121 & n2140 ;
  assign n3655 = n3654 ^ n3625 ;
  assign n3961 = n3655 ^ x81 ;
  assign n2729 = n2672 & n2686 ;
  assign n2706 = n2698 & n2700 ;
  assign n2730 = n2729 ^ n2706 ;
  assign n2727 = ~n2677 & n2698 ;
  assign n2722 = n2660 ^ n2645 ;
  assign n2723 = n2722 ^ n2680 ;
  assign n2724 = n2697 & ~n2723 ;
  assign n2718 = n2685 & ~n2715 ;
  assign n2719 = n2718 ^ n2702 ;
  assign n2720 = n2705 & ~n2719 ;
  assign n2707 = n2706 ^ n2690 ;
  assign n2708 = n2707 ^ n2700 ;
  assign n2709 = n2708 ^ n2673 ;
  assign n2710 = n2709 ^ n2706 ;
  assign n2711 = ~n2705 & ~n2710 ;
  assign n2712 = n2711 ^ n2707 ;
  assign n2721 = n2720 ^ n2712 ;
  assign n2725 = n2724 ^ n2721 ;
  assign n2699 = n2692 ^ n2662 ;
  assign n2703 = n2702 ^ n2699 ;
  assign n2704 = n2698 & n2703 ;
  assign n2726 = n2725 ^ n2704 ;
  assign n2728 = n2727 ^ n2726 ;
  assign n2731 = n2730 ^ n2728 ;
  assign n2732 = n2731 ^ x32 ;
  assign n2695 = n2694 ^ n2693 ;
  assign n2696 = ~n2687 & n2695 ;
  assign n2733 = n2732 ^ n2696 ;
  assign n2683 = n2682 ^ n2674 ;
  assign n2684 = ~n2576 & ~n2683 ;
  assign n2734 = n2733 ^ n2684 ;
  assign n3962 = n2734 ^ x72 ;
  assign n3963 = ~n3961 & ~n3962 ;
  assign n3964 = n3963 ^ n3961 ;
  assign n3965 = n3964 ^ n3962 ;
  assign n4111 = n3965 ^ n3963 ;
  assign n777 = n320 ^ x77 ;
  assign n820 = n819 ^ x126 ;
  assign n1108 = n777 & ~n820 ;
  assign n1124 = n1108 ^ n777 ;
  assign n1125 = n1124 ^ n820 ;
  assign n920 = n917 & n919 ;
  assign n910 = n869 ^ n857 ;
  assign n911 = n910 ^ n832 ;
  assign n906 = n874 ^ n854 ;
  assign n907 = n906 ^ n847 ;
  assign n912 = n911 ^ n907 ;
  assign n913 = ~n822 & ~n912 ;
  assign n908 = n907 ^ n901 ;
  assign n914 = n913 ^ n908 ;
  assign n915 = n861 & n914 ;
  assign n902 = n901 ^ n858 ;
  assign n903 = n902 ^ n900 ;
  assign n904 = n903 ^ n892 ;
  assign n905 = n904 ^ x45 ;
  assign n916 = n915 ^ n905 ;
  assign n921 = n920 ^ n916 ;
  assign n864 = n856 & ~n861 ;
  assign n865 = n864 ^ n858 ;
  assign n866 = ~n822 & n865 ;
  assign n922 = n921 ^ n866 ;
  assign n923 = n922 ^ x109 ;
  assign n938 = n588 ^ n514 ;
  assign n939 = n938 ^ n544 ;
  assign n943 = n939 ^ n508 ;
  assign n944 = ~n507 & ~n943 ;
  assign n945 = n944 ^ n508 ;
  assign n946 = n940 ^ n552 ;
  assign n941 = n940 ^ n939 ;
  assign n947 = n946 ^ n941 ;
  assign n948 = n947 ^ n589 ;
  assign n949 = n945 & ~n948 ;
  assign n950 = n949 ^ n941 ;
  assign n951 = n950 ^ n527 ;
  assign n962 = n951 ^ n519 ;
  assign n960 = n543 ^ n502 ;
  assign n961 = n508 & ~n960 ;
  assign n963 = n962 ^ n961 ;
  assign n964 = ~n507 & ~n963 ;
  assign n954 = n953 ^ n951 ;
  assign n955 = n954 ^ n936 ;
  assign n956 = n955 ^ n534 ;
  assign n957 = n956 ^ n930 ;
  assign n958 = n957 ^ n510 ;
  assign n959 = n958 ^ x53 ;
  assign n965 = n964 ^ n959 ;
  assign n966 = n965 ^ x94 ;
  assign n967 = n923 & ~n966 ;
  assign n968 = n967 ^ n966 ;
  assign n1073 = n1072 ^ x92 ;
  assign n1074 = n231 ^ x83 ;
  assign n1075 = n1073 & n1074 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1110 = n1076 ^ n1073 ;
  assign n1117 = ~n968 & ~n1110 ;
  assign n1113 = n967 & ~n1110 ;
  assign n1118 = n1117 ^ n1113 ;
  assign n1082 = n967 ^ n923 ;
  assign n1111 = n1082 & ~n1110 ;
  assign n1116 = n1111 ^ n1110 ;
  assign n1119 = n1118 ^ n1116 ;
  assign n1094 = n968 ^ n923 ;
  assign n1120 = n1119 ^ n1094 ;
  assign n1095 = n1075 & n1094 ;
  assign n1086 = n967 & n1076 ;
  assign n1081 = ~n968 & n1075 ;
  assign n1087 = n1086 ^ n1081 ;
  assign n1088 = n1087 ^ n1076 ;
  assign n1083 = n1076 & n1082 ;
  assign n1084 = n1083 ^ n1081 ;
  assign n1077 = ~n968 & n1076 ;
  assign n1085 = n1084 ^ n1077 ;
  assign n1089 = n1088 ^ n1085 ;
  assign n1115 = n1095 ^ n1089 ;
  assign n1121 = n1120 ^ n1115 ;
  assign n1078 = n1075 ^ n1073 ;
  assign n1079 = n967 & n1078 ;
  assign n1090 = n1079 ^ n1078 ;
  assign n3557 = n1121 ^ n1090 ;
  assign n1096 = n1095 ^ n1079 ;
  assign n1097 = n1096 ^ n1083 ;
  assign n1146 = n1119 ^ n1097 ;
  assign n3574 = n1097 ^ n1086 ;
  assign n1092 = n967 & n1075 ;
  assign n1093 = n1092 ^ n1084 ;
  assign n3575 = n3574 ^ n1093 ;
  assign n3576 = n3575 ^ n1086 ;
  assign n1091 = n1090 ^ n1073 ;
  assign n1099 = n3576 ^ n1091 ;
  assign n1144 = n1099 ^ n1077 ;
  assign n1145 = n1144 ^ n1095 ;
  assign n1147 = n1146 ^ n1145 ;
  assign n1112 = n1111 ^ n1079 ;
  assign n1141 = n1112 ^ n1086 ;
  assign n1142 = n1141 ^ n1097 ;
  assign n1139 = n1074 ^ n1073 ;
  assign n1140 = n1139 ^ n966 ;
  assign n1143 = n1142 ^ n1140 ;
  assign n1148 = n1147 ^ n1143 ;
  assign n3558 = n3557 ^ n1148 ;
  assign n1151 = n3558 ^ n1119 ;
  assign n1152 = n1125 & ~n1151 ;
  assign n3587 = n1152 ^ x0 ;
  assign n1109 = n1108 ^ n820 ;
  assign n3555 = n1092 & ~n1109 ;
  assign n2514 = n777 & n1115 ;
  assign n2515 = n2514 ^ n1095 ;
  assign n2516 = ~n820 & n2515 ;
  assign n3556 = n3555 ^ n2516 ;
  assign n821 = n820 ^ n777 ;
  assign n3571 = n1093 ^ n777 ;
  assign n3572 = ~n821 & ~n3571 ;
  assign n3573 = n3572 ^ n777 ;
  assign n3577 = n3573 & n3576 ;
  assign n3578 = n3577 ^ n3574 ;
  assign n1149 = n1148 ^ n1121 ;
  assign n1157 = n1149 ^ n1111 ;
  assign n3568 = n1157 ^ n1117 ;
  assign n3569 = n3568 ^ n1077 ;
  assign n3570 = ~n820 & n3569 ;
  assign n3581 = n3578 ^ n3570 ;
  assign n3582 = ~n821 & n3581 ;
  assign n2524 = ~n820 & n1118 ;
  assign n2517 = n1117 ^ n1086 ;
  assign n2518 = ~n820 & n2517 ;
  assign n2519 = n2518 ^ n1117 ;
  assign n2525 = n2524 ^ n2519 ;
  assign n2526 = n777 & n2525 ;
  assign n2527 = n2526 ^ n2519 ;
  assign n3579 = n3578 ^ n2527 ;
  assign n3583 = n3582 ^ n3579 ;
  assign n3565 = n1143 ^ n1113 ;
  assign n3566 = n3565 ^ n1089 ;
  assign n3567 = n1124 & n3566 ;
  assign n3584 = n3583 ^ n3567 ;
  assign n3559 = n3558 ^ n1121 ;
  assign n3562 = n777 & ~n3559 ;
  assign n3563 = n3562 ^ n1121 ;
  assign n3564 = n821 & ~n3563 ;
  assign n3585 = n3584 ^ n3564 ;
  assign n3586 = ~n3556 & ~n3585 ;
  assign n3588 = n3587 ^ n3586 ;
  assign n3966 = n3588 ^ x123 ;
  assign n1914 = n1896 ^ n1844 ;
  assign n1915 = n1914 ^ n1843 ;
  assign n2859 = n1915 ^ n1900 ;
  assign n2860 = ~n2848 & ~n2859 ;
  assign n1853 = ~n1772 & n1850 ;
  assign n1854 = n1853 ^ n1844 ;
  assign n1855 = ~n1741 & n1854 ;
  assign n3972 = n1908 ^ n1898 ;
  assign n3973 = n3972 ^ n3406 ;
  assign n3974 = ~n1772 & n3973 ;
  assign n3967 = n3400 ^ n1890 ;
  assign n3970 = n3967 ^ n1898 ;
  assign n3975 = n3974 ^ n3970 ;
  assign n3976 = ~n1910 & ~n3975 ;
  assign n2850 = n1887 ^ n1875 ;
  assign n2853 = n1772 & ~n2850 ;
  assign n2854 = n2853 ^ n1875 ;
  assign n2855 = n1910 & n2854 ;
  assign n3968 = n3967 ^ n2855 ;
  assign n3969 = n3968 ^ n1943 ;
  assign n3977 = n3976 ^ n3969 ;
  assign n3978 = ~n1855 & ~n3977 ;
  assign n3979 = ~n2860 & n3978 ;
  assign n3980 = ~n2849 & n3979 ;
  assign n3981 = ~n2871 & n3980 ;
  assign n3982 = n3981 ^ x16 ;
  assign n3983 = n3982 ^ x106 ;
  assign n3984 = ~n3966 & n3983 ;
  assign n3985 = n3984 ^ n3966 ;
  assign n1300 = n1299 ^ n241 ;
  assign n1301 = n1300 ^ n1291 ;
  assign n1302 = n1301 ^ n1285 ;
  assign n1303 = n1302 ^ n1277 ;
  assign n1304 = n1303 ^ n1269 ;
  assign n1305 = n1304 ^ x23 ;
  assign n1251 = n1250 ^ n286 ;
  assign n1248 = n269 ^ n243 ;
  assign n1252 = n1251 ^ n1248 ;
  assign n1253 = n233 & n1252 ;
  assign n1249 = n1248 ^ n241 ;
  assign n1254 = n1253 ^ n1249 ;
  assign n1255 = ~n252 & n1254 ;
  assign n1306 = n1305 ^ n1255 ;
  assign n1247 = n246 & ~n258 ;
  assign n1307 = n1306 ^ n1247 ;
  assign n1244 = n233 & n1241 ;
  assign n1245 = n1244 ^ n1240 ;
  assign n1246 = n252 & n1245 ;
  assign n1308 = n1307 ^ n1246 ;
  assign n1309 = n1308 ^ x68 ;
  assign n1340 = n1339 ^ x110 ;
  assign n1341 = n1309 & ~n1340 ;
  assign n1342 = n1341 ^ n1340 ;
  assign n1376 = n178 ^ n155 ;
  assign n1377 = n130 & n1376 ;
  assign n1356 = n136 & ~n205 ;
  assign n1355 = n226 ^ n175 ;
  assign n1357 = n1356 ^ n1355 ;
  assign n1370 = n1369 ^ n1357 ;
  assign n1371 = n1370 ^ n203 ;
  assign n1372 = n1371 ^ n1368 ;
  assign n1373 = n1372 ^ x15 ;
  assign n1354 = n165 ^ n155 ;
  assign n1358 = n1357 ^ n1354 ;
  assign n1352 = n188 ^ n137 ;
  assign n1353 = ~n129 & n1352 ;
  assign n1359 = n1358 ^ n1353 ;
  assign n1360 = n1359 & n1812 ;
  assign n1374 = n1373 ^ n1360 ;
  assign n1350 = n189 ^ n181 ;
  assign n1351 = n132 & ~n1350 ;
  assign n1375 = n1374 ^ n1351 ;
  assign n1378 = n1377 ^ n1375 ;
  assign n1349 = ~n129 & n155 ;
  assign n1379 = n1378 ^ n1349 ;
  assign n1343 = n182 ^ n172 ;
  assign n1346 = ~n129 & n1343 ;
  assign n1347 = n1346 ^ n172 ;
  assign n1348 = ~n130 & n1347 ;
  assign n1380 = n1379 ^ n1348 ;
  assign n1381 = n1380 ^ x117 ;
  assign n1418 = n1417 ^ x69 ;
  assign n1419 = n1381 & n1418 ;
  assign n1420 = n1419 ^ n1418 ;
  assign n1421 = n1420 ^ n1381 ;
  assign n1422 = ~n1342 & ~n1421 ;
  assign n1440 = n1422 ^ n1421 ;
  assign n1425 = n1342 ^ n1309 ;
  assign n1434 = ~n1421 & n1425 ;
  assign n1431 = n1341 & ~n1421 ;
  assign n1439 = n1434 ^ n1431 ;
  assign n1441 = n1440 ^ n1439 ;
  assign n1442 = n1441 ^ n1418 ;
  assign n1424 = n1421 ^ n1418 ;
  assign n1430 = n1424 & n1425 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1433 = n1432 ^ n1422 ;
  assign n1435 = n1434 ^ n1433 ;
  assign n1428 = n1341 & n1424 ;
  assign n1426 = n1425 ^ n1340 ;
  assign n1427 = n1424 & n1426 ;
  assign n1429 = n1428 ^ n1427 ;
  assign n1436 = n1435 ^ n1429 ;
  assign n1443 = n1442 ^ n1436 ;
  assign n2324 = n1443 ^ n1441 ;
  assign n1216 = n1215 ^ x100 ;
  assign n1464 = n1341 & n1419 ;
  assign n2311 = n1464 ^ n1429 ;
  assign n1446 = n1341 & n1420 ;
  assign n1496 = n1446 ^ n1430 ;
  assign n1465 = n1419 & n1426 ;
  assign n2309 = n1496 ^ n1465 ;
  assign n2307 = ~n1216 & n1419 ;
  assign n1462 = n1419 & n1425 ;
  assign n1495 = n1464 ^ n1462 ;
  assign n2308 = n2307 ^ n1495 ;
  assign n2310 = n2309 ^ n2308 ;
  assign n2312 = n2311 ^ n2310 ;
  assign n2313 = n1216 & n2312 ;
  assign n2314 = n2313 ^ n2310 ;
  assign n2323 = n2314 ^ n2308 ;
  assign n2325 = n2324 ^ n2323 ;
  assign n1239 = n1238 ^ x86 ;
  assign n1458 = n1216 & n1239 ;
  assign n1459 = n1458 ^ n1216 ;
  assign n1449 = ~n1342 & n1420 ;
  assign n1448 = n1420 & n1425 ;
  assign n1450 = n1449 ^ n1448 ;
  assign n1447 = n1446 ^ n1420 ;
  assign n1451 = n1450 ^ n1447 ;
  assign n2321 = n1451 ^ n1449 ;
  assign n2322 = n1459 & n2321 ;
  assign n2326 = n2325 ^ n2322 ;
  assign n1494 = n1239 ^ n1216 ;
  assign n2318 = n1239 & ~n2324 ;
  assign n2315 = n2314 ^ n1450 ;
  assign n1471 = n1439 ^ n1428 ;
  assign n2306 = n1471 ^ n1441 ;
  assign n2316 = n2315 ^ n2306 ;
  assign n2319 = n2318 ^ n2316 ;
  assign n2320 = ~n1494 & ~n2319 ;
  assign n2327 = n2326 ^ n2320 ;
  assign n1460 = n1459 ^ n1239 ;
  assign n1461 = n1460 ^ n1216 ;
  assign n2305 = n1422 & n1461 ;
  assign n2328 = n2327 ^ n2305 ;
  assign n1470 = n1446 & n1459 ;
  assign n2329 = n2328 ^ n1470 ;
  assign n1466 = n1465 ^ n1464 ;
  assign n1463 = n1462 ^ n1419 ;
  assign n1467 = n1466 ^ n1463 ;
  assign n1468 = n1467 ^ n1448 ;
  assign n1469 = n1461 & n1468 ;
  assign n2330 = n2329 ^ n1469 ;
  assign n2331 = n2330 ^ x24 ;
  assign n3986 = n2331 ^ x96 ;
  assign n4012 = n2271 ^ n1672 ;
  assign n1689 = n1685 ^ n1616 ;
  assign n4013 = n4012 ^ n1689 ;
  assign n4014 = n1656 & n4013 ;
  assign n1702 = n1679 ^ n1666 ;
  assign n1703 = ~n1656 & n1702 ;
  assign n1704 = n1703 ^ n1666 ;
  assign n4011 = n1704 ^ n1670 ;
  assign n4015 = n4014 ^ n4011 ;
  assign n4016 = ~n1657 & n4015 ;
  assign n1723 = n1656 & ~n1657 ;
  assign n3603 = n1676 & n1723 ;
  assign n3604 = n3603 ^ n2298 ;
  assign n4005 = n3604 ^ n1704 ;
  assign n1674 = n1673 ^ n1668 ;
  assign n3989 = n1716 ^ n1674 ;
  assign n3995 = n3989 ^ n1682 ;
  assign n3988 = n2263 ^ n1687 ;
  assign n3990 = n3989 ^ n3988 ;
  assign n3991 = n3988 ^ n1656 ;
  assign n3992 = n1658 & n3991 ;
  assign n3993 = n3992 ^ n1656 ;
  assign n3994 = n3990 & n3993 ;
  assign n3996 = n3995 ^ n3994 ;
  assign n4006 = n4005 ^ n3996 ;
  assign n4007 = n4006 ^ n1701 ;
  assign n4008 = n4007 ^ x8 ;
  assign n1733 = n1676 ^ n1619 ;
  assign n3997 = n3996 ^ n1733 ;
  assign n3998 = n3997 ^ n1668 ;
  assign n3999 = n3998 ^ n3996 ;
  assign n4000 = n3996 ^ n1657 ;
  assign n4001 = n4000 ^ n3996 ;
  assign n4002 = n3999 & n4001 ;
  assign n4003 = n4002 ^ n3996 ;
  assign n4004 = n1658 & ~n4003 ;
  assign n4009 = n4008 ^ n4004 ;
  assign n3987 = ~n1656 & n1666 ;
  assign n4010 = n4009 ^ n3987 ;
  assign n4017 = n4016 ^ n4010 ;
  assign n4018 = n4017 ^ x113 ;
  assign n4019 = n3986 & ~n4018 ;
  assign n4020 = n4019 ^ n3986 ;
  assign n4021 = n4020 ^ n4018 ;
  assign n4026 = n4021 ^ n3986 ;
  assign n4039 = ~n3985 & ~n4026 ;
  assign n4036 = n3984 & n4019 ;
  assign n4024 = n3985 ^ n3983 ;
  assign n4028 = n4021 & n4024 ;
  assign n4027 = n3984 & ~n4026 ;
  assign n4029 = n4028 ^ n4027 ;
  assign n4037 = n4036 ^ n4029 ;
  assign n4032 = n4018 ^ n3966 ;
  assign n4033 = n3966 & ~n3986 ;
  assign n4034 = n4033 ^ n3983 ;
  assign n4035 = ~n4032 & n4034 ;
  assign n4038 = n4037 ^ n4035 ;
  assign n4040 = n4039 ^ n4038 ;
  assign n4041 = n4040 ^ n4036 ;
  assign n4025 = n4020 & n4024 ;
  assign n4030 = n4029 ^ n4025 ;
  assign n4023 = ~n3985 & n4019 ;
  assign n4031 = n4030 ^ n4023 ;
  assign n4042 = n4041 ^ n4031 ;
  assign n4043 = n4042 ^ n4032 ;
  assign n4047 = n4043 ^ n4027 ;
  assign n4046 = n4024 & ~n4026 ;
  assign n4048 = n4047 ^ n4046 ;
  assign n4044 = n4043 ^ n4039 ;
  assign n4045 = n4044 ^ n4026 ;
  assign n4049 = n4048 ^ n4045 ;
  assign n4074 = n4049 ^ n4030 ;
  assign n4066 = n4019 & n4024 ;
  assign n4067 = n4066 ^ n4036 ;
  assign n4022 = ~n3985 & n4021 ;
  assign n4073 = n4067 ^ n4022 ;
  assign n4075 = n4074 ^ n4073 ;
  assign n4071 = n3983 ^ n3966 ;
  assign n4052 = n4033 ^ n4021 ;
  assign n4072 = n4071 ^ n4052 ;
  assign n4076 = n4075 ^ n4072 ;
  assign n4077 = n4076 ^ n4025 ;
  assign n4070 = n4038 ^ n4020 ;
  assign n4078 = n4077 ^ n4070 ;
  assign n4068 = n4067 ^ n4019 ;
  assign n4069 = n4068 ^ n4023 ;
  assign n4079 = n4078 ^ n4069 ;
  assign n4361 = n4079 ^ n4039 ;
  assign n4362 = n4039 ^ n3961 ;
  assign n4363 = n4362 ^ n4039 ;
  assign n4364 = ~n4361 & ~n4363 ;
  assign n4365 = n4364 ^ n4039 ;
  assign n4366 = ~n4111 & n4365 ;
  assign n4367 = n3963 & n4039 ;
  assign n4368 = ~n4366 & n4367 ;
  assign n4369 = n4368 ^ n4366 ;
  assign n4380 = n4076 ^ n4066 ;
  assign n4381 = n3963 & n4380 ;
  assign n4393 = n4381 ^ n3963 ;
  assign n4382 = n4052 ^ n4028 ;
  assign n4050 = n4049 ^ n4022 ;
  assign n4383 = n4382 ^ n4050 ;
  assign n4384 = n3963 & ~n4383 ;
  assign n4385 = n4384 ^ n3965 ;
  assign n4394 = n4393 ^ n4385 ;
  assign n4387 = n4077 ^ n4050 ;
  assign n4388 = n4077 ^ n3962 ;
  assign n4389 = n4388 ^ n4077 ;
  assign n4390 = n4387 & ~n4389 ;
  assign n4391 = n4390 ^ n4077 ;
  assign n4392 = n3961 & ~n4391 ;
  assign n4395 = n4394 ^ n4392 ;
  assign n4062 = n3963 ^ n3962 ;
  assign n4063 = n4023 & ~n4062 ;
  assign n4061 = ~n3964 & ~n4044 ;
  assign n4064 = n4063 ^ n4061 ;
  assign n4411 = n4395 ^ n4064 ;
  assign n4405 = n4078 ^ n4043 ;
  assign n4406 = n4043 ^ n3961 ;
  assign n4407 = n4406 ^ n4043 ;
  assign n4408 = n4405 & ~n4407 ;
  assign n4409 = n4408 ^ n4043 ;
  assign n4410 = n4111 & ~n4409 ;
  assign n4412 = n4411 ^ n4410 ;
  assign n4399 = n4077 ^ n4067 ;
  assign n4400 = n4067 ^ n3961 ;
  assign n4401 = n4400 ^ n4067 ;
  assign n4402 = ~n4399 & n4401 ;
  assign n4403 = n4402 ^ n4067 ;
  assign n4404 = n4111 & n4403 ;
  assign n4413 = n4412 ^ n4404 ;
  assign n4386 = ~n4381 & ~n4385 ;
  assign n4396 = n4395 ^ n4029 ;
  assign n4397 = n4396 ^ n4392 ;
  assign n4398 = n4386 & ~n4397 ;
  assign n4414 = n4413 ^ n4398 ;
  assign n4378 = n4079 ^ n4046 ;
  assign n4379 = ~n3965 & ~n4378 ;
  assign n4415 = n4414 ^ n4379 ;
  assign n4371 = n4050 ^ n4038 ;
  assign n4370 = n4069 ^ n4027 ;
  assign n4372 = n4371 ^ n4370 ;
  assign n4373 = n4370 ^ n3961 ;
  assign n4374 = n4373 ^ n4370 ;
  assign n4375 = ~n4372 & ~n4374 ;
  assign n4376 = n4375 ^ n4370 ;
  assign n4377 = n4111 & n4376 ;
  assign n4416 = n4415 ^ n4377 ;
  assign n4417 = ~n4369 & n4416 ;
  assign n4418 = n4417 ^ n601 ;
  assign n4419 = n4418 ^ x89 ;
  assign n4539 = n4490 ^ n4419 ;
  assign n3589 = n3588 ^ x107 ;
  assign n2454 = n2419 ^ n2404 ;
  assign n2457 = n2334 & ~n2454 ;
  assign n2458 = n2457 ^ n2419 ;
  assign n2459 = ~n2335 & ~n2458 ;
  assign n3552 = n2459 ^ x26 ;
  assign n3541 = n2414 ^ n2401 ;
  assign n3542 = n3541 ^ n2412 ;
  assign n3543 = n3542 ^ n3215 ;
  assign n3544 = n2335 & n3543 ;
  assign n3545 = n3544 ^ n2414 ;
  assign n3546 = ~n2336 & n3545 ;
  assign n2466 = n2465 ^ n2416 ;
  assign n3539 = n2466 & ~n2494 ;
  assign n3530 = n2401 & n2493 ;
  assign n3529 = n2479 ^ n2421 ;
  assign n3531 = n3530 ^ n3529 ;
  assign n3532 = n3531 ^ n2927 ;
  assign n3535 = n2403 & n2493 ;
  assign n3533 = n3531 ^ n2466 ;
  assign n3534 = n3533 ^ n3227 ;
  assign n3536 = n3535 ^ n3534 ;
  assign n3537 = n3532 & n3536 ;
  assign n3538 = n3537 ^ n2927 ;
  assign n3540 = n3539 ^ n3538 ;
  assign n3547 = n3546 ^ n3540 ;
  assign n3548 = n3547 ^ n2944 ;
  assign n2487 = n2463 ^ n2410 ;
  assign n2490 = n2334 & n2487 ;
  assign n2491 = n2490 ^ n2410 ;
  assign n2492 = ~n2335 & n2491 ;
  assign n3549 = n3548 ^ n2492 ;
  assign n3550 = n3549 ^ n3229 ;
  assign n3551 = ~n3233 & n3550 ;
  assign n3553 = n3552 ^ n3551 ;
  assign n3554 = n3553 ^ x97 ;
  assign n3590 = n3589 ^ n3554 ;
  assign n733 = n732 ^ n406 ;
  assign n3595 = n733 ^ n711 ;
  assign n3596 = n3595 ^ n729 ;
  assign n3597 = n3596 ^ n744 ;
  assign n3598 = ~n496 & n3597 ;
  assign n3593 = n759 ^ n744 ;
  assign n3594 = n3593 ^ n2560 ;
  assign n3599 = n3598 ^ n3594 ;
  assign n3600 = ~n232 & ~n3599 ;
  assign n726 = n725 ^ n724 ;
  assign n408 = n407 ^ n406 ;
  assign n714 = ~n496 & ~n713 ;
  assign n715 = n408 & n714 ;
  assign n727 = n726 ^ n715 ;
  assign n3591 = n727 ^ x50 ;
  assign n3592 = n3591 ^ n2560 ;
  assign n3601 = n3600 ^ n3592 ;
  assign n3602 = n3601 ^ x65 ;
  assign n3614 = n1656 & n2283 ;
  assign n3610 = ~n1657 & n2260 ;
  assign n3611 = n3610 ^ n1664 ;
  assign n3612 = n1656 & n3611 ;
  assign n3613 = n3612 ^ n2280 ;
  assign n3615 = n3614 ^ n3613 ;
  assign n3619 = n3615 ^ n2287 ;
  assign n3620 = n3619 ^ n3612 ;
  assign n3621 = ~n1657 & n3620 ;
  assign n1709 = ~n1656 & n1673 ;
  assign n1710 = n1709 ^ n1704 ;
  assign n1711 = n1657 & n1710 ;
  assign n3605 = n3604 ^ n1711 ;
  assign n3616 = n3615 ^ n3605 ;
  assign n1724 = n1666 & n1723 ;
  assign n1725 = n1724 ^ n1722 ;
  assign n3617 = n3616 ^ n1725 ;
  assign n3618 = n3617 ^ x34 ;
  assign n3622 = n3621 ^ n3618 ;
  assign n3623 = n3622 ^ x112 ;
  assign n3624 = ~n3602 & n3623 ;
  assign n3687 = n3624 ^ n3623 ;
  assign n3690 = n3687 ^ n3602 ;
  assign n3691 = n3690 ^ n3623 ;
  assign n3656 = n3655 ^ x74 ;
  assign n3678 = n2686 & ~n2701 ;
  assign n2982 = ~n2646 & ~n2698 ;
  assign n3670 = n2692 & ~n2982 ;
  assign n2983 = n2653 & n2982 ;
  assign n3668 = n2983 ^ n2722 ;
  assign n2984 = ~n2722 & n2983 ;
  assign n3669 = n3668 ^ n2984 ;
  assign n3671 = n3670 ^ n3669 ;
  assign n3667 = n3126 ^ n2661 ;
  assign n3672 = n3671 ^ n3667 ;
  assign n3673 = n3672 ^ n2682 ;
  assign n3659 = n2694 ^ n2676 ;
  assign n3660 = ~n2576 & ~n3659 ;
  assign n3674 = n3673 ^ n3660 ;
  assign n3675 = ~n2705 & n3674 ;
  assign n3663 = n2648 ^ n2612 ;
  assign n3664 = n3663 ^ n2652 ;
  assign n3665 = n2697 & n3664 ;
  assign n2964 = ~n2656 & ~n2685 ;
  assign n2965 = n2964 ^ n2702 ;
  assign n2966 = n2576 & ~n2965 ;
  assign n2967 = n2966 ^ n2702 ;
  assign n3661 = n3660 ^ n2967 ;
  assign n3662 = n3661 ^ n3158 ;
  assign n3666 = n3665 ^ n3662 ;
  assign n3676 = n3675 ^ n3666 ;
  assign n3657 = n2701 ^ n2673 ;
  assign n3658 = ~n2576 & ~n3657 ;
  assign n3677 = n3676 ^ n3658 ;
  assign n3679 = n3678 ^ n3677 ;
  assign n3680 = ~n2730 & n3679 ;
  assign n3681 = ~n3133 & n3680 ;
  assign n3682 = n3681 ^ x42 ;
  assign n3683 = n3682 ^ x64 ;
  assign n3684 = ~n3656 & ~n3683 ;
  assign n3701 = n3684 ^ n3683 ;
  assign n3723 = ~n3691 & ~n3701 ;
  assign n3722 = n3687 & ~n3701 ;
  assign n3724 = n3723 ^ n3722 ;
  assign n3685 = n3684 ^ n3656 ;
  assign n3695 = ~n3685 & n3690 ;
  assign n3719 = n3695 ^ n3624 ;
  assign n3702 = n3701 ^ n3656 ;
  assign n3712 = n3624 & ~n3702 ;
  assign n3697 = n3623 ^ n3602 ;
  assign n3698 = n3697 ^ n3683 ;
  assign n3699 = n3698 ^ n3624 ;
  assign n3700 = n3656 & n3699 ;
  assign n3703 = n3702 ^ n3700 ;
  assign n3696 = n3695 ^ n3690 ;
  assign n3704 = n3703 ^ n3696 ;
  assign n3694 = n3684 & n3687 ;
  assign n3705 = n3704 ^ n3694 ;
  assign n3692 = n3684 & ~n3691 ;
  assign n3688 = ~n3685 & n3687 ;
  assign n3693 = n3692 ^ n3688 ;
  assign n3706 = n3705 ^ n3693 ;
  assign n3689 = n3688 ^ n3684 ;
  assign n3707 = n3706 ^ n3689 ;
  assign n3708 = n3707 ^ n3695 ;
  assign n3686 = n3624 & ~n3685 ;
  assign n3709 = n3708 ^ n3686 ;
  assign n3713 = n3712 ^ n3709 ;
  assign n3720 = n3719 ^ n3713 ;
  assign n3721 = n3720 ^ n3701 ;
  assign n3725 = n3724 ^ n3721 ;
  assign n3737 = n3725 ^ n3703 ;
  assign n3727 = ~n3691 & ~n3702 ;
  assign n3738 = n3737 ^ n3727 ;
  assign n4444 = n3738 ^ n3706 ;
  assign n3742 = n3708 ^ n3705 ;
  assign n3743 = n3742 ^ n3656 ;
  assign n3741 = n3693 ^ n3686 ;
  assign n3744 = n3743 ^ n3741 ;
  assign n4435 = n3744 ^ n3709 ;
  assign n3736 = n3712 ^ n3702 ;
  assign n3739 = n3738 ^ n3736 ;
  assign n4433 = n3739 ^ n3724 ;
  assign n4434 = n4433 ^ n3720 ;
  assign n4436 = n4435 ^ n4434 ;
  assign n4437 = ~n3589 & ~n4436 ;
  assign n4438 = n4437 ^ n4434 ;
  assign n4445 = n4444 ^ n4438 ;
  assign n4441 = n3704 ^ n3684 ;
  assign n4442 = n4441 ^ n3712 ;
  assign n4443 = ~n3589 & ~n4442 ;
  assign n4446 = n4445 ^ n4443 ;
  assign n4447 = n3590 & ~n4446 ;
  assign n4421 = n3723 ^ n3720 ;
  assign n4420 = n3695 ^ n3694 ;
  assign n4422 = n4421 ^ n4420 ;
  assign n4423 = ~n3554 & ~n4422 ;
  assign n4424 = n4423 ^ n4420 ;
  assign n4439 = n4438 ^ n4424 ;
  assign n3740 = n3739 ^ n3725 ;
  assign n3745 = n3744 ^ n3740 ;
  assign n3746 = n3744 ^ n3589 ;
  assign n3747 = n3746 ^ n3744 ;
  assign n3748 = ~n3745 & ~n3747 ;
  assign n3749 = n3748 ^ n3744 ;
  assign n3750 = ~n3590 & ~n3749 ;
  assign n4440 = n4439 ^ n3750 ;
  assign n4448 = n4447 ^ n4440 ;
  assign n4425 = n4424 ^ n3724 ;
  assign n4428 = n4425 ^ n3701 ;
  assign n4429 = n4428 ^ n4425 ;
  assign n4430 = n3554 & ~n4429 ;
  assign n4431 = n4430 ^ n4425 ;
  assign n4432 = ~n3589 & n4431 ;
  assign n4449 = n4448 ^ n4432 ;
  assign n3774 = ~n3554 & ~n3589 ;
  assign n3775 = n3774 ^ n3554 ;
  assign n3776 = n3775 ^ n3589 ;
  assign n3777 = n3686 & ~n3776 ;
  assign n4450 = n4449 ^ n3777 ;
  assign n4451 = n4450 ^ n320 ;
  assign n4452 = n4451 ^ x106 ;
  assign n2959 = ~n2335 & n2431 ;
  assign n2953 = n2430 ^ n2414 ;
  assign n2954 = n2953 ^ n2952 ;
  assign n2955 = ~n2495 & ~n2954 ;
  assign n2467 = n2466 ^ n2464 ;
  assign n2470 = ~n2335 & ~n2467 ;
  assign n2471 = n2470 ^ n2464 ;
  assign n2472 = ~n2334 & ~n2471 ;
  assign n2947 = n2946 ^ n2472 ;
  assign n2948 = n2947 ^ n2943 ;
  assign n2949 = n2948 ^ n2936 ;
  assign n2950 = n2949 ^ n2459 ;
  assign n2951 = n2950 ^ x52 ;
  assign n2956 = n2955 ^ n2951 ;
  assign n2928 = n2412 ^ n2403 ;
  assign n2929 = n2928 ^ n2444 ;
  assign n2930 = ~n2927 & ~n2929 ;
  assign n2957 = n2956 ^ n2930 ;
  assign n2925 = n2465 ^ n2401 ;
  assign n2926 = ~n2494 & n2925 ;
  assign n2958 = n2957 ^ n2926 ;
  assign n2960 = n2959 ^ n2958 ;
  assign n2961 = n2960 ^ x78 ;
  assign n3000 = n2727 ^ x44 ;
  assign n2976 = n2666 ^ n2656 ;
  assign n2977 = n2976 ^ n2715 ;
  assign n2978 = n2685 & n2977 ;
  assign n2979 = n2978 ^ n2666 ;
  assign n2993 = n2992 ^ n2979 ;
  assign n2985 = n2984 ^ n2979 ;
  assign n2980 = n2979 ^ n2699 ;
  assign n2986 = n2985 ^ n2980 ;
  assign n2989 = n2685 & n2986 ;
  assign n2990 = n2989 ^ n2980 ;
  assign n2991 = ~n2576 & ~n2990 ;
  assign n2994 = n2993 ^ n2991 ;
  assign n2975 = ~n2691 & n2697 ;
  assign n2995 = n2994 ^ n2975 ;
  assign n2974 = n2672 & ~n2705 ;
  assign n2996 = n2995 ^ n2974 ;
  assign n2968 = n2675 ^ n2669 ;
  assign n2971 = ~n2685 & ~n2968 ;
  assign n2972 = n2971 ^ n2675 ;
  assign n2973 = ~n2576 & n2972 ;
  assign n2997 = n2996 ^ n2973 ;
  assign n2998 = n2997 ^ n2706 ;
  assign n2999 = n2967 & ~n2998 ;
  assign n3001 = n3000 ^ n2999 ;
  assign n3002 = n3001 ^ x93 ;
  assign n3003 = ~n2961 & ~n3002 ;
  assign n3004 = n3003 ^ n2961 ;
  assign n2159 = ~n2128 & n2158 ;
  assign n2915 = n2159 ^ n2153 ;
  assign n2916 = n2915 ^ n2914 ;
  assign n2917 = n2916 ^ n2908 ;
  assign n2918 = n2917 ^ x60 ;
  assign n2893 = n2115 ^ n2060 ;
  assign n2894 = n2095 & n2893 ;
  assign n2888 = n2881 ^ n2127 ;
  assign n2885 = n2130 ^ n2105 ;
  assign n2886 = n2095 & ~n2885 ;
  assign n2887 = n2886 ^ n2105 ;
  assign n2889 = n2888 ^ n2887 ;
  assign n2882 = n2881 ^ n2063 ;
  assign n2133 = n2099 ^ n2065 ;
  assign n2883 = n2882 ^ n2133 ;
  assign n2884 = n2095 & n2883 ;
  assign n2890 = n2889 ^ n2884 ;
  assign n2891 = n2890 ^ n2115 ;
  assign n2892 = n2891 ^ n2887 ;
  assign n2895 = n2894 ^ n2892 ;
  assign n2898 = n2895 ^ n2891 ;
  assign n2902 = ~n2898 & ~n2901 ;
  assign n2903 = n2902 ^ n2895 ;
  assign n2904 = n1950 & n2903 ;
  assign n2905 = n2904 ^ n2895 ;
  assign n2906 = ~n2880 & n2905 ;
  assign n2919 = n2918 ^ n2906 ;
  assign n2920 = n2919 ^ x67 ;
  assign n752 = n751 ^ n405 ;
  assign n749 = n711 ^ n602 ;
  assign n750 = n749 ^ n733 ;
  assign n753 = n752 ^ n750 ;
  assign n767 = n753 ^ n232 ;
  assign n760 = n759 ^ n754 ;
  assign n761 = n760 ^ n733 ;
  assign n762 = n761 ^ n755 ;
  assign n738 = n710 ^ n403 ;
  assign n739 = n735 & ~n738 ;
  assign n763 = n762 ^ n739 ;
  assign n764 = n763 ^ n753 ;
  assign n765 = ~n232 & n764 ;
  assign n766 = n765 ^ n763 ;
  assign n768 = n767 ^ n766 ;
  assign n769 = n768 ^ n763 ;
  assign n737 = n736 ^ n722 ;
  assign n740 = n739 ^ n737 ;
  assign n730 = n602 ^ n403 ;
  assign n731 = n730 ^ n729 ;
  assign n734 = n733 ^ n731 ;
  assign n741 = n740 ^ n734 ;
  assign n742 = n741 ^ n728 ;
  assign n770 = n769 ^ n742 ;
  assign n745 = n744 ^ n734 ;
  assign n746 = n745 ^ n739 ;
  assign n743 = n742 ^ n733 ;
  assign n747 = n746 ^ n743 ;
  assign n748 = ~n232 & ~n747 ;
  assign n771 = n770 ^ n748 ;
  assign n772 = ~n496 & ~n771 ;
  assign n773 = n772 ^ n769 ;
  assign n774 = ~n727 & n773 ;
  assign n775 = n774 ^ x36 ;
  assign n2921 = n775 ^ x76 ;
  assign n2922 = n2920 & n2921 ;
  assign n3008 = n2922 ^ n2921 ;
  assign n3017 = ~n3004 & n3008 ;
  assign n2923 = n2922 ^ n2920 ;
  assign n2924 = n2923 ^ n2921 ;
  assign n3026 = n3017 ^ n2924 ;
  assign n3005 = n3004 ^ n3002 ;
  assign n3019 = n3005 ^ n2961 ;
  assign n3021 = n2923 & ~n3019 ;
  assign n3020 = n2922 & ~n3019 ;
  assign n3022 = n3021 ^ n3020 ;
  assign n3014 = n3002 ^ n2961 ;
  assign n3015 = n2961 ^ n2920 ;
  assign n3016 = n3014 & ~n3015 ;
  assign n3018 = n3017 ^ n3016 ;
  assign n3023 = n3022 ^ n3018 ;
  assign n3009 = n3003 & n3008 ;
  assign n3024 = n3023 ^ n3009 ;
  assign n3012 = n2961 ^ n2921 ;
  assign n3013 = ~n2920 & n3012 ;
  assign n3025 = n3024 ^ n3013 ;
  assign n3027 = n3026 ^ n3025 ;
  assign n3011 = n2922 & n3003 ;
  assign n3028 = n3027 ^ n3011 ;
  assign n3010 = n3009 ^ n3003 ;
  assign n3029 = n3028 ^ n3010 ;
  assign n1506 = n1465 ^ n1449 ;
  assign n1507 = n1506 ^ n1443 ;
  assign n1504 = n1430 ^ n1422 ;
  assign n1505 = n1504 ^ n1427 ;
  assign n1508 = n1507 ^ n1505 ;
  assign n1509 = n1216 & n1508 ;
  assign n1510 = n1509 ^ n1507 ;
  assign n1511 = n1494 & n1510 ;
  assign n1497 = n1434 ^ n1427 ;
  assign n1498 = n1497 ^ n1496 ;
  assign n1499 = n1239 & ~n1498 ;
  assign n1500 = n1499 ^ n1495 ;
  assign n1501 = ~n1494 & n1500 ;
  assign n3874 = n1464 ^ n1463 ;
  assign n1476 = n3874 ^ n1494 ;
  assign n1479 = n1451 & ~n1476 ;
  assign n1480 = n3874 ^ n1479 ;
  assign n1486 = ~n1239 & n1429 ;
  assign n1487 = n1486 ^ n1428 ;
  assign n1488 = ~n1216 & n1487 ;
  assign n1490 = n1488 ^ n1216 ;
  assign n1481 = n1458 ^ n1451 ;
  assign n1489 = n1488 ^ n1481 ;
  assign n1491 = n1490 ^ n1489 ;
  assign n1492 = ~n1480 & n1491 ;
  assign n1493 = n1492 ^ n1490 ;
  assign n1502 = n1501 ^ n1493 ;
  assign n1472 = n1471 ^ n1449 ;
  assign n1473 = ~n1460 & n1472 ;
  assign n1503 = n1502 ^ n1473 ;
  assign n1512 = n1511 ^ n1503 ;
  assign n1513 = n1512 ^ n1470 ;
  assign n1514 = n1513 ^ n1469 ;
  assign n1452 = n1451 ^ n1434 ;
  assign n1455 = n1239 & n1452 ;
  assign n1456 = n1455 ^ n1451 ;
  assign n1457 = ~n1216 & n1456 ;
  assign n1515 = n1514 ^ n1457 ;
  assign n1423 = n1422 ^ n1418 ;
  assign n1437 = n1436 ^ n1423 ;
  assign n1438 = n1239 & ~n1437 ;
  assign n1444 = n1443 ^ n1438 ;
  assign n1445 = n1216 & n1444 ;
  assign n1516 = n1515 ^ n1445 ;
  assign n1517 = n1516 ^ x28 ;
  assign n2828 = n1517 ^ x110 ;
  assign n1862 = n1857 & n1861 ;
  assign n1863 = n1862 ^ n1855 ;
  assign n2832 = n2831 ^ n1865 ;
  assign n2833 = n2832 ^ n1875 ;
  assign n2829 = n1888 ^ n1878 ;
  assign n2830 = n2829 ^ n1901 ;
  assign n2840 = n2833 ^ n2830 ;
  assign n2841 = n1772 & ~n2840 ;
  assign n2834 = n1891 ^ n1868 ;
  assign n2835 = n2834 ^ n1915 ;
  assign n2836 = n1772 & ~n2835 ;
  assign n2837 = n2836 ^ n1882 ;
  assign n2838 = n2837 ^ n2833 ;
  assign n2842 = n2841 ^ n2838 ;
  assign n2843 = ~n1741 & n2842 ;
  assign n2844 = n2843 ^ n2837 ;
  assign n2845 = ~n1863 & ~n2844 ;
  assign n2861 = n2860 ^ n2845 ;
  assign n2857 = n2856 ^ n2855 ;
  assign n1929 = n1772 & ~n1914 ;
  assign n1930 = n1929 ^ n1844 ;
  assign n1931 = n1741 & n1930 ;
  assign n2858 = n2857 ^ n1931 ;
  assign n2862 = n2861 ^ n2858 ;
  assign n2863 = n2862 ^ n2849 ;
  assign n2847 = n1885 & n1910 ;
  assign n2864 = n2863 ^ n2847 ;
  assign n2872 = n2864 & ~n2871 ;
  assign n2873 = n2872 ^ x2 ;
  assign n2874 = n2873 ^ x124 ;
  assign n3058 = n2828 & ~n2874 ;
  assign n3059 = n3058 ^ n2874 ;
  assign n4161 = ~n3029 & ~n3059 ;
  assign n4529 = n4161 ^ n709 ;
  assign n3063 = n3058 ^ n2828 ;
  assign n3094 = n3063 ^ n3059 ;
  assign n3114 = n3027 ^ n3019 ;
  assign n3006 = ~n2924 & ~n3005 ;
  assign n3037 = n3024 ^ n3006 ;
  assign n3035 = ~n2920 & n3002 ;
  assign n3036 = n3035 ^ n3008 ;
  assign n3038 = n3037 ^ n3036 ;
  assign n3071 = n3038 ^ n3027 ;
  assign n3072 = n3071 ^ n3022 ;
  assign n3115 = n3114 ^ n3072 ;
  assign n3039 = n3038 ^ n3017 ;
  assign n3040 = n3039 ^ n3009 ;
  assign n3041 = n3040 ^ n3008 ;
  assign n3116 = n3115 ^ n3041 ;
  assign n3117 = n3115 ^ n2828 ;
  assign n3118 = n3117 ^ n3115 ;
  assign n3119 = ~n3116 & n3118 ;
  assign n3120 = n3119 ^ n3115 ;
  assign n3121 = ~n3094 & ~n3120 ;
  assign n4530 = n4529 ^ n3121 ;
  assign n3088 = n3029 ^ n3006 ;
  assign n3089 = n3006 ^ n2828 ;
  assign n3090 = n3089 ^ n3006 ;
  assign n3091 = ~n3088 & n3090 ;
  assign n3092 = n3091 ^ n3006 ;
  assign n3093 = n2874 & n3092 ;
  assign n3032 = n2923 & ~n3004 ;
  assign n3033 = n3032 ^ n3020 ;
  assign n4526 = n3033 & n3063 ;
  assign n4501 = n3032 ^ n3011 ;
  assign n4502 = n4501 ^ n3022 ;
  assign n3074 = n3027 ^ n3006 ;
  assign n3075 = n3074 ^ n3017 ;
  assign n3077 = n3028 ^ n3021 ;
  assign n4498 = n3075 & n3077 ;
  assign n3030 = n3029 ^ n3022 ;
  assign n3031 = n3030 ^ n2923 ;
  assign n3034 = n3033 ^ n3031 ;
  assign n4499 = n4498 ^ n3034 ;
  assign n4500 = n3094 & n4499 ;
  assign n4503 = n3058 & ~n4500 ;
  assign n4504 = n4502 & n4503 ;
  assign n4505 = n4504 ^ n4500 ;
  assign n3103 = n3011 ^ n2922 ;
  assign n3042 = n3041 ^ n3034 ;
  assign n3007 = n3006 ^ n3005 ;
  assign n3043 = n3042 ^ n3007 ;
  assign n3044 = n3043 ^ n3020 ;
  assign n3104 = n3103 ^ n3044 ;
  assign n4129 = n3104 ^ n3034 ;
  assign n4493 = ~n3059 & ~n4129 ;
  assign n4506 = n4505 ^ n4493 ;
  assign n3070 = n2874 ^ n2828 ;
  assign n4507 = n3115 ^ n3024 ;
  assign n4508 = n4507 ^ n2828 ;
  assign n4509 = n3070 & n4508 ;
  assign n4510 = n4509 ^ n2828 ;
  assign n4513 = n4507 ^ n3040 ;
  assign n4514 = n4510 & ~n4513 ;
  assign n4511 = n3043 ^ n3040 ;
  assign n4515 = n4514 ^ n4511 ;
  assign n4516 = n4515 ^ n3039 ;
  assign n4517 = n4516 ^ n3023 ;
  assign n4518 = n4517 ^ n4515 ;
  assign n4521 = ~n2828 & n4518 ;
  assign n4522 = n4521 ^ n4515 ;
  assign n4523 = n3070 & n4522 ;
  assign n4524 = n4523 ^ n4515 ;
  assign n4525 = ~n4506 & ~n4524 ;
  assign n4527 = n4526 ^ n4525 ;
  assign n4528 = ~n3093 & n4527 ;
  assign n4531 = n4530 ^ n4528 ;
  assign n4532 = n4531 ^ x88 ;
  assign n4548 = n4452 & ~n4532 ;
  assign n4563 = n4539 & n4548 ;
  assign n3190 = n1464 ^ n1448 ;
  assign n3191 = n3190 ^ n1441 ;
  assign n3192 = n3191 ^ n1464 ;
  assign n3193 = n3192 ^ n1462 ;
  assign n3194 = ~n1216 & ~n3193 ;
  assign n3195 = n3194 ^ n3190 ;
  assign n3196 = n1239 & n3195 ;
  assign n3181 = n3874 ^ n1507 ;
  assign n3182 = n3181 ^ n1446 ;
  assign n3183 = n3874 ^ n3182 ;
  assign n3186 = ~n1239 & n3183 ;
  assign n3187 = n3874 ^ n3186 ;
  assign n3188 = ~n1216 & n3187 ;
  assign n3189 = n3874 ^ n3188 ;
  assign n3197 = n3196 ^ n3189 ;
  assign n3198 = n3197 ^ n1471 ;
  assign n3178 = n1432 & n1461 ;
  assign n3177 = n1471 ^ n1432 ;
  assign n3179 = n3178 ^ n3177 ;
  assign n3180 = ~n1459 & n3179 ;
  assign n3199 = n3198 ^ n3180 ;
  assign n3200 = n3199 ^ n2322 ;
  assign n3201 = n3200 ^ n1488 ;
  assign n3202 = n3201 ^ n2305 ;
  assign n3203 = n3202 ^ n1469 ;
  assign n3204 = n3203 ^ n1457 ;
  assign n3205 = n3204 ^ n1445 ;
  assign n3206 = n3205 ^ x46 ;
  assign n3207 = n3206 ^ x102 ;
  assign n1171 = n1089 ^ n1084 ;
  assign n1172 = n1124 & n1171 ;
  assign n1167 = n1145 ^ n1111 ;
  assign n1168 = ~n820 & n1167 ;
  assign n1158 = n1157 ^ n1145 ;
  assign n1159 = n1158 ^ n1117 ;
  assign n1160 = n1159 ^ n1157 ;
  assign n1163 = ~n820 & n1160 ;
  assign n1164 = n1163 ^ n1157 ;
  assign n1165 = n777 & n1164 ;
  assign n1153 = n1152 ^ n1111 ;
  assign n1133 = n1118 ^ n1089 ;
  assign n1136 = ~n777 & n1133 ;
  assign n1137 = n1136 ^ n1118 ;
  assign n1138 = ~n821 & n1137 ;
  assign n1154 = n1153 ^ n1138 ;
  assign n1127 = n1092 ^ n1087 ;
  assign n1130 = ~n777 & n1127 ;
  assign n1131 = n1130 ^ n1092 ;
  assign n1132 = n820 & n1131 ;
  assign n1155 = n1154 ^ n1132 ;
  assign n1156 = n1155 ^ x62 ;
  assign n1166 = n1165 ^ n1156 ;
  assign n1169 = n1168 ^ n1166 ;
  assign n1126 = n1113 & n1125 ;
  assign n1170 = n1169 ^ n1126 ;
  assign n1173 = n1172 ^ n1170 ;
  assign n1114 = n1113 ^ n1112 ;
  assign n1122 = n1121 ^ n1114 ;
  assign n1123 = ~n1109 & ~n1122 ;
  assign n1174 = n1173 ^ n1123 ;
  assign n1100 = n1099 ^ n1089 ;
  assign n1101 = n1100 ^ n1087 ;
  assign n1080 = n1079 ^ n1077 ;
  assign n1102 = n1101 ^ n1080 ;
  assign n1105 = n777 & n1102 ;
  assign n1106 = n1105 ^ n1080 ;
  assign n1107 = n821 & n1106 ;
  assign n1175 = n1174 ^ n1107 ;
  assign n3238 = n1175 ^ x91 ;
  assign n3252 = ~n3207 & n3238 ;
  assign n3165 = n754 ^ n742 ;
  assign n3166 = n3165 ^ n746 ;
  assign n3167 = n232 & n3166 ;
  assign n3168 = n3167 ^ n742 ;
  assign n3169 = n3168 ^ n766 ;
  assign n3172 = n496 & n3169 ;
  assign n3173 = n3172 ^ n3168 ;
  assign n3174 = ~n2572 & n3173 ;
  assign n3175 = n3174 ^ x54 ;
  assign n3176 = n3175 ^ x77 ;
  assign n3237 = n3236 ^ x117 ;
  assign n3253 = n3176 & ~n3237 ;
  assign n3254 = n3253 ^ n3176 ;
  assign n3271 = n3252 & n3254 ;
  assign n3259 = n3252 ^ n3238 ;
  assign n3263 = n3259 ^ n3207 ;
  assign n3265 = n3263 ^ n3238 ;
  assign n3266 = n3253 & ~n3265 ;
  assign n3264 = n3253 & n3263 ;
  assign n3267 = n3266 ^ n3264 ;
  assign n3261 = n3253 & n3259 ;
  assign n3262 = n3261 ^ n3253 ;
  assign n3268 = n3267 ^ n3262 ;
  assign n3272 = n3271 ^ n3268 ;
  assign n3255 = n3254 ^ n3237 ;
  assign n3256 = n3252 & n3255 ;
  assign n3270 = n3256 ^ n3252 ;
  assign n3273 = n3272 ^ n3270 ;
  assign n3260 = n3255 & n3259 ;
  assign n3269 = n3268 ^ n3260 ;
  assign n3274 = n3273 ^ n3269 ;
  assign n3239 = n3237 & n3238 ;
  assign n3258 = n3252 ^ n3239 ;
  assign n3275 = n3274 ^ n3258 ;
  assign n3276 = n3275 ^ n3273 ;
  assign n4356 = n3276 ^ n495 ;
  assign n3164 = n3163 ^ x126 ;
  assign n3277 = n3276 ^ n3261 ;
  assign n3249 = n3237 ^ n3207 ;
  assign n3250 = n3249 ^ n3176 ;
  assign n3251 = n3250 ^ n3237 ;
  assign n3257 = n3256 ^ n3251 ;
  assign n3278 = n3277 ^ n3257 ;
  assign n3279 = n3278 ^ n3249 ;
  assign n3242 = n3237 ^ n3176 ;
  assign n3243 = n3242 ^ n3238 ;
  assign n3245 = n3238 ^ n3207 ;
  assign n3246 = n3176 & ~n3245 ;
  assign n3247 = ~n3243 & n3246 ;
  assign n3248 = n3247 ^ n3243 ;
  assign n3280 = n3279 ^ n3248 ;
  assign n4347 = ~n3164 & ~n3280 ;
  assign n4348 = n4347 ^ n3248 ;
  assign n4357 = n4356 ^ n4348 ;
  assign n1947 = n1946 ^ x4 ;
  assign n1916 = n1915 ^ n1881 ;
  assign n1917 = n1916 ^ n1887 ;
  assign n1932 = n1931 ^ n1917 ;
  assign n1920 = n1889 ^ n1872 ;
  assign n1921 = n1920 ^ n1867 ;
  assign n1923 = n1922 ^ n1921 ;
  assign n1924 = ~n1772 & ~n1923 ;
  assign n1918 = n1917 ^ n1879 ;
  assign n1919 = n1918 ^ n1913 ;
  assign n1925 = n1924 ^ n1919 ;
  assign n1926 = ~n1910 & n1925 ;
  assign n1933 = n1932 ^ n1926 ;
  assign n1909 = n1857 & n1908 ;
  assign n1934 = n1933 ^ n1909 ;
  assign n1902 = n1901 ^ n1886 ;
  assign n1905 = n1772 & n1902 ;
  assign n1906 = n1905 ^ n1886 ;
  assign n1907 = n1741 & n1906 ;
  assign n1935 = n1934 ^ n1907 ;
  assign n1936 = ~n1863 & ~n1935 ;
  assign n1948 = n1947 ^ n1936 ;
  assign n3308 = n1948 ^ x100 ;
  assign n3208 = n3207 ^ n3176 ;
  assign n3240 = n3239 ^ n3176 ;
  assign n3241 = ~n3208 & ~n3240 ;
  assign n3244 = n3243 ^ n3241 ;
  assign n4349 = n4348 ^ n3244 ;
  assign n4350 = n4349 ^ n4348 ;
  assign n4353 = n3164 & n4350 ;
  assign n4354 = n4353 ^ n4348 ;
  assign n4355 = n3308 & ~n4354 ;
  assign n4358 = n4357 ^ n4355 ;
  assign n3282 = n3245 ^ n3176 ;
  assign n3283 = n3282 ^ n3245 ;
  assign n3284 = n3245 ^ n3237 ;
  assign n3287 = ~n3283 & n3284 ;
  assign n3288 = n3287 ^ n3245 ;
  assign n3289 = ~n3208 & ~n3288 ;
  assign n3290 = n3289 ^ n3284 ;
  assign n4344 = n3290 & n3308 ;
  assign n4345 = n4344 ^ n3276 ;
  assign n4346 = ~n3164 & n4345 ;
  assign n4359 = n4358 ^ n4346 ;
  assign n4360 = n4359 ^ x82 ;
  assign n4491 = n4490 ^ n4452 ;
  assign n4545 = n4532 ^ n4419 ;
  assign n4535 = n4532 ^ n4490 ;
  assign n6441 = n4535 ^ n4532 ;
  assign n6442 = ~n4545 & ~n6441 ;
  assign n6443 = n6442 ^ n4532 ;
  assign n6444 = ~n4491 & n6443 ;
  assign n4561 = n4548 ^ n4532 ;
  assign n4562 = n4419 & ~n4561 ;
  assign n4564 = n4563 ^ n4562 ;
  assign n6455 = n6444 ^ n4564 ;
  assign n6456 = n6455 ^ n4539 ;
  assign n4556 = n4452 ^ n4419 ;
  assign n4557 = n4556 ^ n4452 ;
  assign n4558 = n4490 & ~n4557 ;
  assign n4559 = n4558 ^ n4452 ;
  assign n4560 = n4532 & n4559 ;
  assign n4565 = n4564 ^ n4560 ;
  assign n4553 = n4539 ^ n4532 ;
  assign n4546 = n4545 ^ n4452 ;
  assign n4547 = n4546 ^ n4532 ;
  assign n4549 = n4548 ^ n4452 ;
  assign n4550 = n4549 ^ n4490 ;
  assign n4492 = n4452 & ~n4491 ;
  assign n4551 = n4550 ^ n4492 ;
  assign n4552 = ~n4547 & n4551 ;
  assign n4554 = n4553 ^ n4552 ;
  assign n4566 = n4565 ^ n4554 ;
  assign n6457 = n6456 ^ n4566 ;
  assign n2304 = n2303 ^ x114 ;
  assign n2332 = n2331 ^ x121 ;
  assign n2784 = ~n2304 & ~n2332 ;
  assign n2785 = n2784 ^ n2332 ;
  assign n2497 = n2496 ^ n2492 ;
  assign n2427 = ~n2334 & n2404 ;
  assign n2428 = n2427 ^ n2422 ;
  assign n2429 = ~n2335 & ~n2428 ;
  assign n2433 = n2432 ^ n2429 ;
  assign n2434 = n2433 ^ n2414 ;
  assign n2436 = n2435 ^ n2434 ;
  assign n2437 = n2436 ^ n2429 ;
  assign n2438 = n2334 & ~n2437 ;
  assign n2439 = n2438 ^ n2433 ;
  assign n2498 = n2497 ^ n2439 ;
  assign n2499 = n2498 ^ n2486 ;
  assign n2500 = n2499 ^ n2478 ;
  assign n2501 = n2500 ^ n2472 ;
  assign n2502 = n2501 ^ n2459 ;
  assign n2503 = n2502 ^ x48 ;
  assign n2451 = n2334 & n2448 ;
  assign n2440 = n2439 ^ n2429 ;
  assign n2452 = n2451 ^ n2440 ;
  assign n2453 = ~n2336 & n2452 ;
  assign n2504 = n2503 ^ n2453 ;
  assign n2505 = n2504 ^ x73 ;
  assign n2544 = n1094 ^ n1092 ;
  assign n2545 = n2544 ^ n1112 ;
  assign n2546 = n2545 ^ n1115 ;
  assign n2547 = ~n820 & n2546 ;
  assign n2548 = n2547 ^ n1112 ;
  assign n2549 = n777 & n2548 ;
  assign n2535 = n3557 ^ n1112 ;
  assign n2538 = n2535 ^ n1144 ;
  assign n2533 = n1095 ^ n1085 ;
  assign n2536 = n2535 ^ n2533 ;
  assign n2537 = n777 & ~n2536 ;
  assign n2539 = n2538 ^ n2537 ;
  assign n2540 = ~n821 & ~n2539 ;
  assign n2528 = n2527 ^ n1144 ;
  assign n2529 = n2528 ^ n2516 ;
  assign n2530 = n2529 ^ n1138 ;
  assign n2531 = n2530 ^ n1152 ;
  assign n2532 = n2531 ^ x40 ;
  assign n2541 = n2540 ^ n2532 ;
  assign n2507 = n1113 ^ n1095 ;
  assign n2508 = n2507 ^ n1148 ;
  assign n2509 = n1125 & ~n2508 ;
  assign n2542 = n2541 ^ n2509 ;
  assign n2506 = n1083 & ~n1109 ;
  assign n2543 = n2542 ^ n2506 ;
  assign n2550 = n2549 ^ n2543 ;
  assign n2551 = n2550 ^ x99 ;
  assign n2552 = ~n2505 & ~n2551 ;
  assign n2575 = n2574 ^ x90 ;
  assign n2735 = n2734 ^ x88 ;
  assign n2736 = ~n2575 & ~n2735 ;
  assign n2741 = n2552 & n2736 ;
  assign n2788 = n2741 ^ n2552 ;
  assign n2553 = n2552 ^ n2551 ;
  assign n2554 = n2553 ^ n2505 ;
  assign n2737 = n2736 ^ n2575 ;
  assign n2752 = n2737 ^ n2735 ;
  assign n2764 = ~n2554 & ~n2752 ;
  assign n2757 = ~n2551 & ~n2752 ;
  assign n2763 = n2757 ^ n2752 ;
  assign n2765 = n2764 ^ n2763 ;
  assign n2753 = n2752 ^ n2575 ;
  assign n2754 = ~n2553 & ~n2753 ;
  assign n2766 = n2765 ^ n2754 ;
  assign n2740 = ~n2553 & n2736 ;
  assign n2742 = n2741 ^ n2740 ;
  assign n2743 = n2742 ^ n2736 ;
  assign n2739 = ~n2554 & n2736 ;
  assign n2744 = n2743 ^ n2739 ;
  assign n2767 = n2766 ^ n2744 ;
  assign n2747 = n2552 ^ n2505 ;
  assign n2748 = ~n2737 & ~n2747 ;
  assign n2761 = n2754 ^ n2748 ;
  assign n2762 = n2761 ^ n2747 ;
  assign n2768 = n2767 ^ n2762 ;
  assign n2769 = n2768 ^ n2753 ;
  assign n2759 = ~n2554 & ~n2753 ;
  assign n2760 = n2759 ^ n2754 ;
  assign n2770 = n2769 ^ n2760 ;
  assign n2756 = ~n2553 & ~n2752 ;
  assign n2758 = n2757 ^ n2756 ;
  assign n2771 = n2770 ^ n2758 ;
  assign n2789 = n2788 ^ n2771 ;
  assign n2821 = n2789 ^ n2737 ;
  assign n2738 = ~n2554 & ~n2737 ;
  assign n2782 = n2748 ^ n2738 ;
  assign n2822 = n2821 ^ n2782 ;
  assign n2823 = ~n2785 & n2822 ;
  assign n2819 = ~n2765 & ~n2785 ;
  assign n2745 = n2744 ^ n2738 ;
  assign n2772 = n2771 ^ n2745 ;
  assign n4328 = n2304 & ~n2772 ;
  assign n2786 = n2785 ^ n2304 ;
  assign n2800 = n2786 ^ n2332 ;
  assign n2795 = n2768 ^ n2764 ;
  assign n2796 = n2795 ^ n2770 ;
  assign n4325 = n2796 ^ n2765 ;
  assign n4326 = ~n2800 & n4325 ;
  assign n2790 = n2789 ^ n2739 ;
  assign n2791 = n2790 ^ n2756 ;
  assign n4322 = n2791 ^ n2759 ;
  assign n4323 = ~n2786 & ~n4322 ;
  assign n2814 = n2789 ^ n2740 ;
  assign n4315 = n2814 ^ n2754 ;
  assign n4312 = n2768 ^ n2757 ;
  assign n4313 = n4312 ^ n2814 ;
  assign n4314 = ~n2332 & ~n4313 ;
  assign n4316 = n4315 ^ n4314 ;
  assign n4318 = n2784 ^ n2304 ;
  assign n4317 = n2784 ^ n2754 ;
  assign n4319 = n4318 ^ n4317 ;
  assign n4320 = n4316 & ~n4319 ;
  assign n4321 = n4320 ^ n4318 ;
  assign n4324 = n4323 ^ n4321 ;
  assign n4327 = n4326 ^ n4324 ;
  assign n4329 = n4328 ^ n4327 ;
  assign n4305 = n2784 ^ n2748 ;
  assign n2746 = n2745 ^ n2741 ;
  assign n4306 = n2746 ^ n2332 ;
  assign n4309 = ~n2748 & n4306 ;
  assign n4310 = n4309 ^ n2332 ;
  assign n4311 = n4305 & ~n4310 ;
  assign n4330 = n4329 ^ n4311 ;
  assign n4331 = ~n2819 & n4330 ;
  assign n2333 = n2332 ^ n2304 ;
  assign n4332 = n2759 ^ n2748 ;
  assign n4307 = n2748 ^ n2332 ;
  assign n4333 = n4307 ^ n2748 ;
  assign n4334 = n4332 & ~n4333 ;
  assign n4335 = n4334 ^ n2748 ;
  assign n4336 = n2333 & n4335 ;
  assign n4337 = n4331 & ~n4336 ;
  assign n4338 = ~n2823 & n4337 ;
  assign n4339 = n4338 ^ n231 ;
  assign n4340 = n4339 ^ x64 ;
  assign n6445 = n4549 ^ n4532 ;
  assign n4536 = ~n4419 & ~n4532 ;
  assign n4537 = n4536 ^ n4452 ;
  assign n6446 = n6445 ^ n4537 ;
  assign n6447 = n6446 ^ n4452 ;
  assign n6448 = n4490 & n6447 ;
  assign n6449 = n6448 ^ n4546 ;
  assign n6450 = n6449 ^ n4562 ;
  assign n6451 = n6450 ^ n6444 ;
  assign n6452 = n4340 & ~n6451 ;
  assign n6453 = n6452 ^ n6449 ;
  assign n6458 = n6457 ^ n6453 ;
  assign n4538 = ~n4535 & n4537 ;
  assign n4540 = n4539 ^ n4538 ;
  assign n6435 = n4554 ^ n4540 ;
  assign n6436 = n6435 ^ n4492 ;
  assign n6437 = n6436 ^ n4560 ;
  assign n6438 = n6437 ^ n4553 ;
  assign n6454 = n6453 ^ n6438 ;
  assign n6459 = n6458 ^ n6454 ;
  assign n6460 = n6458 ^ n4340 ;
  assign n6461 = n6460 ^ n6458 ;
  assign n6462 = ~n6459 & ~n6461 ;
  assign n6463 = n6462 ^ n6458 ;
  assign n6464 = n4360 & ~n6463 ;
  assign n6465 = n6464 ^ n6453 ;
  assign n6466 = ~n4563 & n6465 ;
  assign n6467 = n6466 ^ n2574 ;
  assign n6468 = n6467 ^ x123 ;
  assign n3122 = n3121 ^ n1771 ;
  assign n3045 = n3044 ^ n3041 ;
  assign n3046 = ~n2874 & n3045 ;
  assign n3047 = n3046 ^ n3041 ;
  assign n3050 = n3047 ^ n3033 ;
  assign n3048 = n3043 ^ n3034 ;
  assign n3049 = n3048 ^ n3047 ;
  assign n3051 = n3050 ^ n3049 ;
  assign n3054 = ~n2874 & ~n3051 ;
  assign n3055 = n3054 ^ n3050 ;
  assign n3056 = n2828 & n3055 ;
  assign n3057 = n3056 ^ n3047 ;
  assign n3102 = n3059 ^ n2828 ;
  assign n3105 = n3104 ^ n3029 ;
  assign n3106 = n3102 & ~n3105 ;
  assign n3107 = n3106 ^ n3017 ;
  assign n3073 = n3072 ^ n3036 ;
  assign n3076 = n3075 ^ n3073 ;
  assign n3078 = n3077 ^ n3076 ;
  assign n3079 = n2828 & ~n3078 ;
  assign n3080 = n3079 ^ n3072 ;
  assign n3108 = n3107 ^ n3080 ;
  assign n3097 = n3041 ^ n2874 ;
  assign n3098 = n3097 ^ n3041 ;
  assign n3099 = ~n3042 & n3098 ;
  assign n3100 = n3099 ^ n3041 ;
  assign n3101 = ~n3094 & n3100 ;
  assign n3109 = n3108 ^ n3101 ;
  assign n3110 = n3109 ^ n3093 ;
  assign n3085 = n2828 & ~n3028 ;
  assign n3086 = n3085 ^ n3080 ;
  assign n3087 = ~n3070 & ~n3086 ;
  assign n3111 = n3110 ^ n3087 ;
  assign n3060 = n3059 ^ n3017 ;
  assign n3061 = n3032 ^ n3009 ;
  assign n3062 = n3061 ^ n3006 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3065 = n3063 ^ n3017 ;
  assign n3066 = n3065 ^ n3063 ;
  assign n3067 = ~n3064 & ~n3066 ;
  assign n3068 = n3067 ^ n3063 ;
  assign n3069 = ~n3060 & ~n3068 ;
  assign n3112 = n3111 ^ n3069 ;
  assign n3113 = ~n3057 & n3112 ;
  assign n3123 = n3122 ^ n3113 ;
  assign n3124 = n3123 ^ x107 ;
  assign n3326 = n3164 & ~n3308 ;
  assign n3327 = n3326 ^ n3308 ;
  assign n3328 = n3327 ^ n3164 ;
  assign n3329 = n3328 ^ n3308 ;
  assign n3330 = n3329 ^ n3327 ;
  assign n3336 = n3261 ^ n3260 ;
  assign n3337 = n3336 ^ n3259 ;
  assign n3291 = n3290 ^ n3276 ;
  assign n3281 = n3280 ^ n3244 ;
  assign n3292 = n3291 ^ n3281 ;
  assign n3297 = n3292 ^ n3256 ;
  assign n3296 = n3249 ^ n3248 ;
  assign n3298 = n3297 ^ n3296 ;
  assign n3299 = n3298 ^ n3266 ;
  assign n3316 = n3299 ^ n3265 ;
  assign n3350 = n3337 ^ n3316 ;
  assign n3351 = n3316 ^ n3164 ;
  assign n3352 = n3351 ^ n3316 ;
  assign n3353 = ~n3350 & ~n3352 ;
  assign n3354 = n3353 ^ n3316 ;
  assign n3355 = ~n3330 & ~n3354 ;
  assign n3356 = n3355 ^ n2363 ;
  assign n3315 = n3261 ^ n3247 ;
  assign n3334 = n3315 & ~n3327 ;
  assign n3335 = n3334 ^ n3329 ;
  assign n3338 = n3268 ^ n3256 ;
  assign n3339 = n3338 ^ n3334 ;
  assign n3340 = n3339 ^ n3337 ;
  assign n3341 = n3335 & n3340 ;
  assign n3331 = n3269 ^ n3261 ;
  assign n3332 = n3331 ^ n3271 ;
  assign n3333 = n3330 & n3332 ;
  assign n3342 = n3341 ^ n3333 ;
  assign n3317 = n3316 ^ n3315 ;
  assign n3294 = n3255 ^ n3176 ;
  assign n3295 = n3263 & ~n3294 ;
  assign n3300 = n3299 ^ n3295 ;
  assign n3293 = n3292 ^ n3276 ;
  assign n3301 = n3300 ^ n3293 ;
  assign n3304 = n3301 ^ n3295 ;
  assign n3303 = n3264 ^ n3263 ;
  assign n3305 = n3304 ^ n3303 ;
  assign n3318 = n3317 ^ n3305 ;
  assign n3319 = n3318 ^ n3301 ;
  assign n3314 = n3300 ^ n3256 ;
  assign n3320 = n3319 ^ n3314 ;
  assign n3321 = n3319 ^ n3308 ;
  assign n3322 = n3321 ^ n3319 ;
  assign n3323 = ~n3320 & ~n3322 ;
  assign n3324 = n3323 ^ n3319 ;
  assign n3325 = ~n3164 & ~n3324 ;
  assign n3343 = n3342 ^ n3325 ;
  assign n3344 = n3273 ^ n3264 ;
  assign n3347 = ~n3330 & n3344 ;
  assign n3348 = n3347 ^ n3273 ;
  assign n3349 = ~n3343 & ~n3348 ;
  assign n3357 = n3356 ^ n3349 ;
  assign n3302 = n3301 ^ n3266 ;
  assign n3306 = n3305 ^ n3302 ;
  assign n3307 = n3306 ^ n3305 ;
  assign n3311 = n3307 & ~n3308 ;
  assign n3312 = n3311 ^ n3305 ;
  assign n3313 = n3164 & n3312 ;
  assign n3358 = n3357 ^ n3313 ;
  assign n3359 = n3358 ^ x97 ;
  assign n3524 = ~n3473 & ~n3475 ;
  assign n3520 = n3519 ^ n3485 ;
  assign n3521 = n3443 & n3520 ;
  assign n3506 = n3468 ^ n3439 ;
  assign n3509 = n3508 ^ n3506 ;
  assign n3510 = n3509 ^ n3485 ;
  assign n3504 = n3450 ^ n3448 ;
  assign n3505 = n3504 ^ n3485 ;
  assign n3511 = n3510 ^ n3505 ;
  assign n3512 = ~n3443 & n3511 ;
  assign n3513 = n3512 ^ n3510 ;
  assign n3514 = n3444 & ~n3513 ;
  assign n3487 = n3486 ^ n3485 ;
  assign n3477 = n3461 ^ n3452 ;
  assign n3480 = n3461 ^ n3443 ;
  assign n3481 = n3480 ^ n3461 ;
  assign n3482 = n3477 & n3481 ;
  assign n3483 = n3482 ^ n3461 ;
  assign n3484 = ~n3444 & n3483 ;
  assign n3488 = n3487 ^ n3484 ;
  assign n3501 = n3500 ^ n3488 ;
  assign n3476 = n3474 & ~n3475 ;
  assign n3502 = n3501 ^ n3476 ;
  assign n3503 = n3502 ^ n2094 ;
  assign n3515 = n3514 ^ n3503 ;
  assign n3522 = n3521 ^ n3515 ;
  assign n3446 = n3442 & n3445 ;
  assign n3523 = n3522 ^ n3446 ;
  assign n3525 = n3524 ^ n3523 ;
  assign n3526 = n3525 ^ x80 ;
  assign n3766 = n3737 ^ n3693 ;
  assign n3767 = n3766 ^ n3722 ;
  assign n3763 = n3695 ^ n3686 ;
  assign n3761 = n3712 ^ n3692 ;
  assign n3762 = n3761 ^ n3694 ;
  assign n3764 = n3763 ^ n3762 ;
  assign n3755 = n3708 ^ n3694 ;
  assign n3756 = n3755 ^ n3737 ;
  assign n3757 = ~n3589 & n3756 ;
  assign n3752 = n3739 ^ n3723 ;
  assign n3753 = n3752 ^ n3727 ;
  assign n3754 = n3753 ^ n3742 ;
  assign n3758 = n3757 ^ n3754 ;
  assign n3765 = n3764 ^ n3758 ;
  assign n3768 = n3767 ^ n3765 ;
  assign n3769 = n3768 ^ n3758 ;
  assign n3770 = n3589 & ~n3769 ;
  assign n3771 = n3770 ^ n3765 ;
  assign n3772 = ~n3590 & n3771 ;
  assign n3726 = n3725 ^ n3720 ;
  assign n3728 = n3727 ^ n3726 ;
  assign n3731 = n3727 ^ n3554 ;
  assign n3732 = n3731 ^ n3727 ;
  assign n3733 = ~n3728 & n3732 ;
  assign n3734 = n3733 ^ n3727 ;
  assign n3735 = ~n3590 & n3734 ;
  assign n3751 = n3750 ^ n3735 ;
  assign n3759 = n3758 ^ n3751 ;
  assign n3710 = n3709 ^ n3589 ;
  assign n3711 = n3710 ^ n3709 ;
  assign n3716 = n3711 & ~n3713 ;
  assign n3717 = n3716 ^ n3709 ;
  assign n3718 = n3590 & ~n3717 ;
  assign n3760 = n3759 ^ n3718 ;
  assign n3773 = n3772 ^ n3760 ;
  assign n3778 = n3777 ^ n3773 ;
  assign n3779 = n3778 ^ n2390 ;
  assign n3780 = n3779 ^ x90 ;
  assign n3781 = n3526 & ~n3780 ;
  assign n3782 = n3359 & n3781 ;
  assign n3792 = n3124 & n3782 ;
  assign n3793 = n3792 ^ n3782 ;
  assign n1176 = n1175 ^ x68 ;
  assign n776 = n775 ^ x86 ;
  assign n2228 = n1176 ^ n776 ;
  assign n1949 = n1948 ^ x125 ;
  assign n2170 = n2065 & n2095 ;
  assign n2167 = n2100 & ~n2147 ;
  assign n2144 = n2124 ^ n2057 ;
  assign n2165 = n2144 & n2158 ;
  assign n2148 = n2122 ^ n2120 ;
  assign n2151 = n2148 ^ n2060 ;
  assign n2152 = n2140 & ~n2151 ;
  assign n2154 = n2153 ^ n2152 ;
  assign n2149 = n2148 ^ n2117 ;
  assign n2150 = ~n2147 & ~n2149 ;
  assign n2155 = n2154 ^ n2150 ;
  assign n2142 = n2130 ^ n2114 ;
  assign n2143 = n2142 ^ n2117 ;
  assign n2145 = n2144 ^ n2143 ;
  assign n2146 = n2141 & ~n2145 ;
  assign n2156 = n2155 ^ n2146 ;
  assign n2134 = n2133 ^ n2132 ;
  assign n2137 = n2095 & n2134 ;
  assign n2138 = n2137 ^ n2133 ;
  assign n2139 = n1950 & n2138 ;
  assign n2157 = n2156 ^ n2139 ;
  assign n2160 = n2159 ^ n2157 ;
  assign n2162 = n2161 ^ n2160 ;
  assign n2163 = n2162 ^ n2113 ;
  assign n2164 = n2163 ^ x12 ;
  assign n2166 = n2165 ^ n2164 ;
  assign n2168 = n2167 ^ n2166 ;
  assign n2066 = n2065 ^ n2063 ;
  assign n2067 = ~n1950 & n2066 ;
  assign n2169 = n2168 ^ n2067 ;
  assign n2171 = n2170 ^ n2169 ;
  assign n2172 = n2171 ^ x92 ;
  assign n2173 = n1949 & ~n2172 ;
  assign n2174 = n2173 ^ n2172 ;
  assign n2199 = n2174 ^ n1949 ;
  assign n1518 = n1517 ^ x69 ;
  assign n1732 = n1731 ^ n1670 ;
  assign n1734 = n1733 ^ n1732 ;
  assign n1735 = n1656 & n1734 ;
  assign n1713 = n1676 ^ n1671 ;
  assign n1736 = n1735 ^ n1713 ;
  assign n1737 = n1658 & n1736 ;
  assign n1659 = ~n1620 & ~n1658 ;
  assign n1712 = n1687 ^ n1659 ;
  assign n1714 = n1713 ^ n1712 ;
  assign n1715 = n1714 ^ n1711 ;
  assign n1726 = n1725 ^ n1715 ;
  assign n1727 = n1726 ^ n1701 ;
  assign n1728 = n1727 ^ x20 ;
  assign n1690 = n1689 ^ n1681 ;
  assign n1667 = n1666 ^ n1664 ;
  assign n1675 = n1674 ^ n1667 ;
  assign n1691 = n1690 ^ n1675 ;
  assign n1692 = n1657 & ~n1691 ;
  assign n1688 = n1687 ^ n1675 ;
  assign n1693 = n1692 ^ n1688 ;
  assign n1694 = ~n1656 & ~n1693 ;
  assign n1729 = n1728 ^ n1694 ;
  assign n1661 = n1657 & n1660 ;
  assign n1662 = n1659 & n1661 ;
  assign n1730 = n1729 ^ n1662 ;
  assign n1738 = n1737 ^ n1730 ;
  assign n1739 = n1738 ^ x75 ;
  assign n1740 = n1518 & n1739 ;
  assign n2176 = n1740 ^ n1518 ;
  assign n2211 = n2176 ^ n1739 ;
  assign n2212 = n2199 & ~n2211 ;
  assign n2180 = n1740 ^ n1739 ;
  assign n2192 = n2173 & n2180 ;
  assign n2193 = n2192 ^ n2173 ;
  assign n2184 = n2172 ^ n1949 ;
  assign n2185 = n1739 ^ n1518 ;
  assign n2187 = n2185 ^ n1949 ;
  assign n2188 = n2187 ^ n2172 ;
  assign n2189 = n1518 & ~n2188 ;
  assign n2186 = n2185 ^ n2172 ;
  assign n2190 = n2189 ^ n2186 ;
  assign n2191 = n2184 & ~n2190 ;
  assign n2194 = n2193 ^ n2191 ;
  assign n2195 = n2194 ^ n2192 ;
  assign n2181 = n2173 ^ n1949 ;
  assign n2182 = n2180 & n2181 ;
  assign n2183 = n2182 ^ n2180 ;
  assign n2196 = n2195 ^ n2183 ;
  assign n2177 = ~n2174 & n2176 ;
  assign n2175 = n1740 & ~n2174 ;
  assign n2178 = n2177 ^ n2175 ;
  assign n2179 = n2178 ^ n2174 ;
  assign n2197 = n2196 ^ n2179 ;
  assign n2230 = n2212 ^ n2197 ;
  assign n2253 = n1176 & ~n2230 ;
  assign n2219 = n2173 & ~n2211 ;
  assign n2220 = n2219 ^ n2196 ;
  assign n2213 = n2212 ^ n2182 ;
  assign n2221 = n2220 ^ n2213 ;
  assign n2222 = n2221 ^ n2175 ;
  assign n2206 = n1740 & n2173 ;
  assign n2201 = n1740 & n2181 ;
  assign n2202 = n2201 ^ n2175 ;
  assign n2200 = n2176 & n2199 ;
  assign n2203 = n2202 ^ n2200 ;
  assign n2204 = n2203 ^ n2189 ;
  assign n2205 = n2204 ^ n2200 ;
  assign n2207 = n2206 ^ n2205 ;
  assign n2223 = n2222 ^ n2207 ;
  assign n2224 = ~n1176 & n2223 ;
  assign n2225 = n2224 ^ n2221 ;
  assign n2251 = n2225 ^ n2212 ;
  assign n1177 = ~n776 & ~n1176 ;
  assign n2214 = n1177 ^ n776 ;
  assign n2215 = n2214 ^ n1176 ;
  assign n2243 = n2215 ^ n776 ;
  assign n2245 = n2201 ^ n2194 ;
  assign n2239 = n2177 ^ n2176 ;
  assign n2240 = n2239 ^ n2205 ;
  assign n2244 = n2240 ^ n2177 ;
  assign n2246 = n2245 ^ n2244 ;
  assign n2247 = n2243 & ~n2246 ;
  assign n2236 = n2206 ^ n1740 ;
  assign n2237 = n2236 ^ n2202 ;
  assign n2238 = n2214 & ~n2237 ;
  assign n2241 = ~n2202 & ~n2240 ;
  assign n2242 = n2238 & n2241 ;
  assign n2248 = n2247 ^ n2242 ;
  assign n2229 = n2219 ^ n2211 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2232 = n2231 ^ n2196 ;
  assign n2233 = n2232 ^ n2192 ;
  assign n2249 = n2248 ^ n2233 ;
  assign n2198 = n2197 ^ n2194 ;
  assign n2216 = ~n2213 & n2215 ;
  assign n2217 = n2198 & n2216 ;
  assign n2208 = n2207 ^ n2198 ;
  assign n2209 = n2208 ^ n2197 ;
  assign n2210 = ~n1177 & ~n2209 ;
  assign n2218 = n2217 ^ n2210 ;
  assign n2250 = n2249 ^ n2218 ;
  assign n2252 = n2251 ^ n2250 ;
  assign n2254 = n2253 ^ n2252 ;
  assign n2255 = n2228 & n2254 ;
  assign n2226 = n2225 ^ n2006 ;
  assign n2227 = n2226 ^ n2218 ;
  assign n2256 = n2255 ^ n2227 ;
  assign n2257 = n2256 ^ x121 ;
  assign n2815 = n2814 ^ n2744 ;
  assign n2816 = ~n2785 & ~n2815 ;
  assign n2806 = n2796 ^ n2768 ;
  assign n2807 = n2806 ^ n2760 ;
  assign n2808 = n2760 ^ n2332 ;
  assign n2809 = n2808 ^ n2760 ;
  assign n2810 = ~n2807 & ~n2809 ;
  assign n2811 = n2810 ^ n2760 ;
  assign n2812 = n2304 & n2811 ;
  assign n2783 = n2782 ^ n2740 ;
  assign n2787 = n2786 ^ n2783 ;
  assign n2792 = n2791 ^ n2787 ;
  assign n2793 = ~n2758 & ~n2792 ;
  assign n2794 = n2793 ^ n2786 ;
  assign n2802 = n2768 ^ n2758 ;
  assign n2801 = n2800 ^ n2768 ;
  assign n2803 = n2802 ^ n2801 ;
  assign n2804 = n2794 & ~n2803 ;
  assign n2805 = n2804 ^ n2802 ;
  assign n2813 = n2812 ^ n2805 ;
  assign n2817 = n2816 ^ n2813 ;
  assign n2755 = n2754 ^ n2738 ;
  assign n2773 = n2772 ^ n2755 ;
  assign n2750 = n2735 ^ n2575 ;
  assign n2751 = n2750 ^ n2505 ;
  assign n2774 = n2773 ^ n2751 ;
  assign n2775 = n2774 ^ n2754 ;
  assign n2749 = n2748 ^ n2746 ;
  assign n2776 = n2775 ^ n2749 ;
  assign n2777 = n2775 ^ n2332 ;
  assign n2778 = n2777 ^ n2775 ;
  assign n2779 = n2776 & n2778 ;
  assign n2780 = n2779 ^ n2775 ;
  assign n2781 = ~n2333 & n2780 ;
  assign n2818 = n2817 ^ n2781 ;
  assign n2820 = n2819 ^ n2818 ;
  assign n2824 = n2823 ^ n2820 ;
  assign n2825 = n2824 ^ n1841 ;
  assign n2826 = n2825 ^ x65 ;
  assign n2827 = ~n2257 & ~n2826 ;
  assign n3800 = n2827 ^ n2826 ;
  assign n6398 = n3793 & ~n3800 ;
  assign n3828 = n3782 ^ n3781 ;
  assign n3787 = ~n3124 & ~n3359 ;
  assign n3796 = ~n3526 & n3787 ;
  assign n3788 = n3781 ^ n3526 ;
  assign n3789 = n3787 & n3788 ;
  assign n3795 = n3789 ^ n3787 ;
  assign n3797 = n3796 ^ n3795 ;
  assign n3829 = n3828 ^ n3797 ;
  assign n3527 = n3359 & ~n3526 ;
  assign n3528 = n3527 ^ n3359 ;
  assign n3783 = n3782 ^ n3528 ;
  assign n3830 = n3829 ^ n3783 ;
  assign n3831 = n3783 ^ n2257 ;
  assign n3832 = n3831 ^ n3783 ;
  assign n3833 = n3830 & ~n3832 ;
  assign n3834 = n3833 ^ n3783 ;
  assign n3835 = n2826 & n3834 ;
  assign n6023 = n2827 & n3783 ;
  assign n3801 = n3800 ^ n2257 ;
  assign n3802 = n3801 ^ n2826 ;
  assign n3784 = ~n3124 & n3783 ;
  assign n3785 = n3784 ^ n3783 ;
  assign n3836 = n3793 ^ n3785 ;
  assign n6426 = ~n3802 & n3836 ;
  assign n3805 = ~n3124 & n3527 ;
  assign n3814 = n3780 & n3805 ;
  assign n3815 = n3814 ^ n3805 ;
  assign n3810 = n3527 ^ n3526 ;
  assign n3811 = n3810 ^ n3796 ;
  assign n6420 = n3815 ^ n3811 ;
  assign n3790 = n3788 ^ n3783 ;
  assign n3791 = n3790 ^ n3789 ;
  assign n6032 = n3791 ^ n3784 ;
  assign n6421 = n6420 ^ n6032 ;
  assign n6422 = ~n2826 & ~n6421 ;
  assign n3812 = ~n3780 & ~n3811 ;
  assign n3813 = n3812 ^ n3811 ;
  assign n6399 = n3814 ^ n3813 ;
  assign n6400 = n6399 ^ n3789 ;
  assign n6401 = n2826 & ~n6400 ;
  assign n6402 = n6401 ^ n3789 ;
  assign n6419 = n6402 ^ n3791 ;
  assign n6423 = n6422 ^ n6419 ;
  assign n6424 = n2257 & n6423 ;
  assign n3803 = n3802 ^ n3800 ;
  assign n6408 = n3815 ^ n3812 ;
  assign n3808 = ~n3780 & n3796 ;
  assign n3809 = n3808 ^ n3796 ;
  assign n6404 = n3809 ^ n3792 ;
  assign n6405 = n6404 ^ n3797 ;
  assign n6406 = n6405 ^ n3809 ;
  assign n6407 = n6406 ^ n3797 ;
  assign n6409 = n6408 ^ n6407 ;
  assign n6410 = ~n2827 & ~n6409 ;
  assign n6411 = n6410 ^ n6405 ;
  assign n3804 = n3797 ^ n3792 ;
  assign n6412 = n6411 ^ n3804 ;
  assign n3821 = n3780 ^ n3124 ;
  assign n3822 = ~n3526 & ~n3821 ;
  assign n3806 = n3805 ^ n3527 ;
  assign n6413 = n3822 ^ n3806 ;
  assign n6414 = n3801 & ~n6413 ;
  assign n6415 = ~n6412 & n6414 ;
  assign n6416 = n6415 ^ n6411 ;
  assign n6417 = ~n3803 & ~n6416 ;
  assign n6403 = n6402 ^ n3792 ;
  assign n6418 = n6417 ^ n6403 ;
  assign n6425 = n6424 ^ n6418 ;
  assign n6427 = n6426 ^ n6425 ;
  assign n6428 = ~n6023 & ~n6427 ;
  assign n6429 = ~n3835 & n6428 ;
  assign n6040 = n3822 ^ n3796 ;
  assign n3816 = n3815 ^ n3813 ;
  assign n3817 = n3816 ^ n3809 ;
  assign n6041 = n6040 ^ n3817 ;
  assign n6055 = n6041 ^ n3806 ;
  assign n6063 = n6055 ^ n3809 ;
  assign n6064 = ~n3802 & ~n6063 ;
  assign n3842 = n3829 ^ n3789 ;
  assign n6062 = ~n3800 & n3842 ;
  assign n6065 = n6064 ^ n6062 ;
  assign n6430 = n6429 ^ n6065 ;
  assign n6431 = ~n6398 & n6430 ;
  assign n6432 = n6431 ^ n2504 ;
  assign n6433 = n6432 ^ x106 ;
  assign n4602 = n3022 ^ n3019 ;
  assign n4603 = n3063 & ~n4602 ;
  assign n4597 = n3043 ^ n3030 ;
  assign n4141 = ~n3043 & n3059 ;
  assign n4585 = n4501 ^ n4141 ;
  assign n4586 = n3063 & ~n4585 ;
  assign n4584 = n3022 & ~n4141 ;
  assign n4587 = n4586 ^ n4584 ;
  assign n4588 = n4587 ^ n3104 ;
  assign n4598 = n4597 ^ n4588 ;
  assign n4593 = n3071 ^ n3024 ;
  assign n4594 = n4593 ^ n3030 ;
  assign n4595 = n4594 ^ n3043 ;
  assign n4596 = ~n2828 & n4595 ;
  assign n4599 = n4598 ^ n4596 ;
  assign n4600 = n3094 & ~n4599 ;
  assign n4583 = n4161 ^ n3106 ;
  assign n4589 = n4588 ^ n4583 ;
  assign n4590 = n4589 ^ n3101 ;
  assign n4591 = n4590 ^ n3121 ;
  assign n4592 = n4591 ^ n1560 ;
  assign n4601 = n4600 ^ n4592 ;
  assign n4604 = n4603 ^ n4601 ;
  assign n4582 = ~n3048 & n3102 ;
  assign n4605 = n4604 ^ n4582 ;
  assign n4577 = n3024 ^ n2828 ;
  assign n4578 = n4577 ^ n3024 ;
  assign n4579 = n3025 & n4578 ;
  assign n4580 = n4579 ^ n3024 ;
  assign n4581 = ~n2874 & n4580 ;
  assign n4606 = n4605 ^ n4581 ;
  assign n4607 = n4606 ^ x83 ;
  assign n3857 = n1146 ^ n1117 ;
  assign n3858 = n3857 ^ n3557 ;
  assign n3859 = n777 & n3858 ;
  assign n3863 = n3859 ^ n3556 ;
  assign n3864 = n3863 ^ n1132 ;
  assign n3865 = n3864 ^ x18 ;
  assign n3860 = n3859 ^ n1122 ;
  assign n3855 = n3568 ^ n1078 ;
  assign n3856 = ~n777 & n3855 ;
  assign n3861 = n3860 ^ n3856 ;
  assign n3862 = n821 & ~n3861 ;
  assign n3866 = n3865 ^ n3862 ;
  assign n3854 = n1085 & n1108 ;
  assign n3867 = n3866 ^ n3854 ;
  assign n3848 = n1143 ^ n1100 ;
  assign n3851 = n820 & n3848 ;
  assign n3852 = n3851 ^ n1143 ;
  assign n3853 = ~n777 & n3852 ;
  assign n3868 = n3867 ^ n3853 ;
  assign n3869 = n3868 ^ x104 ;
  assign n3870 = n3553 ^ x105 ;
  assign n3913 = n3869 & ~n3870 ;
  assign n3915 = n3913 ^ n3870 ;
  assign n3916 = n3915 ^ n3869 ;
  assign n3911 = n2919 ^ x80 ;
  assign n3895 = n1462 ^ n1451 ;
  assign n3896 = n1458 & n3895 ;
  assign n3888 = n1441 ^ n1432 ;
  assign n3883 = ~n1216 & n1436 ;
  assign n3884 = n3883 ^ n1429 ;
  assign n3889 = n3888 ^ n3884 ;
  assign n3886 = n1463 ^ n1449 ;
  assign n3887 = n3886 ^ n3884 ;
  assign n3890 = n3889 ^ n3887 ;
  assign n3891 = ~n1216 & ~n3890 ;
  assign n3892 = n3891 ^ n3889 ;
  assign n3893 = n1494 & ~n3892 ;
  assign n3882 = n3178 ^ n1445 ;
  assign n3885 = n3884 ^ n3882 ;
  assign n3894 = n3893 ^ n3885 ;
  assign n3897 = n3896 ^ n3894 ;
  assign n3875 = n3874 ^ n1449 ;
  assign n3876 = n3875 ^ n1463 ;
  assign n3879 = n1216 & n3876 ;
  assign n3880 = n3879 ^ n1463 ;
  assign n3881 = ~n1239 & n3880 ;
  assign n3898 = n3897 ^ n3881 ;
  assign n3899 = n3898 ^ n2305 ;
  assign n3900 = n3899 ^ n1470 ;
  assign n3873 = n1216 & n1468 ;
  assign n3901 = n3900 ^ n3873 ;
  assign n3902 = ~n1457 & ~n3901 ;
  assign n3903 = n3902 ^ x10 ;
  assign n3904 = n3903 ^ x66 ;
  assign n3910 = n3622 ^ x98 ;
  assign n3952 = ~n3904 & n3910 ;
  assign n3871 = n2873 ^ x122 ;
  assign n3905 = ~n3871 & ~n3904 ;
  assign n3953 = n3952 ^ n3905 ;
  assign n3954 = ~n3911 & n3953 ;
  assign n4831 = n3954 ^ n3953 ;
  assign n4832 = n3916 & n4831 ;
  assign n3918 = n3870 ^ n3869 ;
  assign n3917 = ~n3871 & ~n3916 ;
  assign n3919 = n3918 ^ n3917 ;
  assign n3872 = n3870 & n3871 ;
  assign n3912 = n3872 ^ n3871 ;
  assign n3914 = n3913 ^ n3912 ;
  assign n3920 = n3919 ^ n3914 ;
  assign n3906 = n3905 ^ n3871 ;
  assign n3907 = n3906 ^ n3904 ;
  assign n4823 = n3920 ^ n3907 ;
  assign n4818 = n3904 ^ n3870 ;
  assign n3938 = n3870 & ~n3906 ;
  assign n4819 = n4818 ^ n3938 ;
  assign n4820 = n3869 & ~n4819 ;
  assign n3930 = ~n3869 & n3905 ;
  assign n3931 = n3930 ^ n3871 ;
  assign n3932 = ~n3918 & ~n3931 ;
  assign n4821 = n4820 ^ n3932 ;
  assign n3933 = n3904 ^ n3871 ;
  assign n3934 = ~n3915 & ~n3933 ;
  assign n3935 = n3934 ^ n3932 ;
  assign n3926 = n3920 ^ n3918 ;
  assign n3936 = n3935 ^ n3926 ;
  assign n4822 = n4821 ^ n3936 ;
  assign n4824 = n4823 ^ n4822 ;
  assign n3925 = ~n3871 & n3913 ;
  assign n3937 = n3936 ^ n3925 ;
  assign n4825 = n4824 ^ n3937 ;
  assign n4826 = ~n3910 & n4825 ;
  assign n4827 = n4826 ^ n4822 ;
  assign n3921 = n3920 ^ n3871 ;
  assign n3922 = n3904 & n3921 ;
  assign n3923 = n3922 ^ n3917 ;
  assign n3943 = n3936 ^ n3923 ;
  assign n3908 = n3907 ^ n3872 ;
  assign n3909 = n3869 & ~n3908 ;
  assign n4814 = n3943 ^ n3909 ;
  assign n4812 = n3904 ^ n3869 ;
  assign n4813 = n4812 ^ n3872 ;
  assign n4815 = n4814 ^ n4813 ;
  assign n4810 = n3925 ^ n3913 ;
  assign n4811 = n4810 ^ n3906 ;
  assign n4816 = n4815 ^ n4811 ;
  assign n3927 = n3871 ^ n3869 ;
  assign n4805 = n3870 & ~n3904 ;
  assign n4806 = n4805 ^ n3869 ;
  assign n4807 = n3927 & ~n4806 ;
  assign n4808 = n4807 ^ n3869 ;
  assign n4809 = n3910 & n4808 ;
  assign n4817 = n4816 ^ n4809 ;
  assign n4828 = n4827 ^ n4817 ;
  assign n4829 = ~n3911 & ~n4828 ;
  assign n4830 = n4829 ^ n4827 ;
  assign n4833 = n4832 ^ n4830 ;
  assign n4834 = n4833 ^ n1072 ;
  assign n4835 = n4834 ^ x70 ;
  assign n5834 = n4607 & n4835 ;
  assign n5835 = n5834 ^ n4835 ;
  assign n5836 = n5835 ^ n4607 ;
  assign n4755 = n3301 ^ n3264 ;
  assign n4756 = n4755 ^ n3316 ;
  assign n4757 = ~n3327 & ~n4756 ;
  assign n4752 = n3339 ^ n3271 ;
  assign n4753 = n4752 ^ n3264 ;
  assign n4758 = n4757 ^ n4753 ;
  assign n4759 = ~n3326 & n4758 ;
  assign n4751 = n3304 ^ n3256 ;
  assign n4754 = n4753 ^ n4751 ;
  assign n4760 = n4759 ^ n4754 ;
  assign n4745 = n3308 ^ n3256 ;
  assign n4746 = n4745 ^ n3328 ;
  assign n4747 = n3308 ^ n3277 ;
  assign n4748 = n3329 & ~n4747 ;
  assign n4749 = n4748 ^ n3308 ;
  assign n4750 = n4746 & ~n4749 ;
  assign n4761 = n4760 ^ n4750 ;
  assign n4744 = n3274 & n3328 ;
  assign n4762 = n4761 ^ n4744 ;
  assign n4742 = n3305 ^ n3298 ;
  assign n4743 = n3330 & n4742 ;
  assign n4763 = n4762 ^ n4743 ;
  assign n4735 = n3304 ^ n3267 ;
  assign n4734 = n3304 ^ n3272 ;
  assign n4736 = n4735 ^ n4734 ;
  assign n4737 = n4735 ^ n3308 ;
  assign n4738 = n4737 ^ n4735 ;
  assign n4739 = n4736 & ~n4738 ;
  assign n4740 = n4739 ^ n4735 ;
  assign n4741 = ~n3164 & n4740 ;
  assign n4764 = n4763 ^ n4741 ;
  assign n4765 = ~n3355 & ~n4764 ;
  assign n4766 = n4765 ^ n2611 ;
  assign n4767 = n4766 ^ x126 ;
  assign n4626 = n3737 ^ n3708 ;
  assign n4627 = n4626 ^ n3737 ;
  assign n4628 = n3737 ^ n3554 ;
  assign n4629 = n4628 ^ n3737 ;
  assign n4630 = ~n4627 & n4629 ;
  assign n4631 = n4630 ^ n3737 ;
  assign n4632 = ~n3590 & ~n4631 ;
  assign n4633 = n4632 ^ n3737 ;
  assign n4617 = ~n3741 & n3775 ;
  assign n4611 = n3776 ^ n3554 ;
  assign n4613 = n3695 ^ n3688 ;
  assign n4612 = n3744 ^ n3704 ;
  assign n4614 = n4613 ^ n4612 ;
  assign n4615 = n4611 & ~n4614 ;
  assign n4618 = n3704 & ~n4615 ;
  assign n4619 = n4617 & n4618 ;
  assign n4610 = n3724 ^ n3712 ;
  assign n4616 = n4615 ^ n4610 ;
  assign n4620 = n4619 ^ n4616 ;
  assign n4634 = n4633 ^ n4620 ;
  assign n4635 = n4634 ^ n3751 ;
  assign n4636 = n4635 ^ n1655 ;
  assign n4621 = n3712 ^ n3688 ;
  assign n4622 = n4621 ^ n3694 ;
  assign n4623 = n4622 ^ n4620 ;
  assign n4608 = n3700 ^ n3698 ;
  assign n4609 = ~n3589 & n4608 ;
  assign n4624 = n4623 ^ n4609 ;
  assign n4625 = ~n3590 & ~n4624 ;
  assign n4637 = n4636 ^ n4625 ;
  assign n4638 = n4637 ^ x109 ;
  assign n4797 = n4767 ^ n4638 ;
  assign n4714 = n2742 ^ n2738 ;
  assign n4710 = n2740 ^ n2738 ;
  assign n4711 = n4710 ^ n2822 ;
  assign n4712 = n4711 ^ n2790 ;
  assign n4713 = n2332 & ~n4712 ;
  assign n4715 = n4714 ^ n4713 ;
  assign n4725 = n4715 ^ n2823 ;
  assign n4717 = n2765 ^ n2759 ;
  assign n4716 = n4715 ^ n2771 ;
  assign n4718 = n4717 ^ n4716 ;
  assign n4719 = n4718 ^ n4715 ;
  assign n4720 = n4715 ^ n2332 ;
  assign n4721 = n4720 ^ n4715 ;
  assign n4722 = n4719 & n4721 ;
  assign n4723 = n4722 ^ n4715 ;
  assign n4724 = ~n2304 & n4723 ;
  assign n4726 = n4725 ^ n4724 ;
  assign n4702 = n2822 ^ n2739 ;
  assign n4703 = n4702 ^ n2782 ;
  assign n4701 = n2768 ^ n2756 ;
  assign n4704 = n4703 ^ n4701 ;
  assign n4705 = n4701 ^ n2304 ;
  assign n4706 = n4705 ^ n4701 ;
  assign n4707 = n4704 & ~n4706 ;
  assign n4708 = n4707 ^ n4701 ;
  assign n4709 = ~n2332 & n4708 ;
  assign n4727 = n4726 ^ n4709 ;
  assign n4699 = n2745 ^ n2740 ;
  assign n4700 = ~n2800 & n4699 ;
  assign n4728 = n4727 ^ n4700 ;
  assign n4692 = n2767 ^ n2758 ;
  assign n4693 = n4692 ^ n2770 ;
  assign n4694 = n4693 ^ n2758 ;
  assign n4695 = n4694 ^ n2795 ;
  assign n4696 = ~n2332 & n4695 ;
  assign n4697 = n4696 ^ n4692 ;
  assign n4698 = ~n2333 & ~n4697 ;
  assign n4729 = n4728 ^ n4698 ;
  assign n4730 = n4729 ^ n2819 ;
  assign n4731 = n4730 ^ n4336 ;
  assign n4732 = n4731 ^ n2640 ;
  assign n4733 = n4732 ^ x76 ;
  assign n4798 = n4797 ^ n4733 ;
  assign n4639 = n3445 & ~n3489 ;
  assign n4640 = n4639 ^ n3484 ;
  assign n4662 = n3444 ^ n3443 ;
  assign n4663 = n3519 ^ n3470 ;
  assign n4664 = ~n4662 & n4663 ;
  assign n4651 = n3443 ^ n3441 ;
  assign n4652 = n3441 ^ n3431 ;
  assign n4653 = n4652 ^ n3433 ;
  assign n4654 = n4653 ^ n4652 ;
  assign n4655 = n4652 ^ n3444 ;
  assign n4656 = n4655 ^ n4652 ;
  assign n4657 = n4654 & ~n4656 ;
  assign n4658 = n4657 ^ n4652 ;
  assign n4659 = n4651 & ~n4658 ;
  assign n4660 = n4659 ^ n3443 ;
  assign n4649 = n3477 ^ n3440 ;
  assign n4650 = n4454 & n4649 ;
  assign n4661 = n4660 ^ n4650 ;
  assign n4665 = n4664 ^ n4661 ;
  assign n4648 = n3439 & ~n3475 ;
  assign n4666 = n4665 ^ n4648 ;
  assign n4641 = n3460 ^ n3444 ;
  assign n4642 = n4641 ^ n3460 ;
  assign n4643 = n3460 ^ n3434 ;
  assign n4644 = n4643 ^ n3460 ;
  assign n4645 = n4642 & n4644 ;
  assign n4646 = n4645 ^ n3460 ;
  assign n4647 = n3443 & ~n4646 ;
  assign n4667 = n4666 ^ n4647 ;
  assign n4668 = ~n4640 & ~n4667 ;
  assign n4669 = ~n3495 & n4668 ;
  assign n4674 = ~n3444 & n3453 ;
  assign n4675 = n4674 ^ n3431 ;
  assign n4676 = ~n3443 & n4675 ;
  assign n4677 = n4669 & ~n4676 ;
  assign n4678 = n3485 ^ n3441 ;
  assign n4679 = n3444 & n4678 ;
  assign n4680 = n4679 ^ n3441 ;
  assign n4685 = ~n3443 & n4680 ;
  assign n4686 = n4685 ^ n4478 ;
  assign n4687 = n4677 & ~n4686 ;
  assign n4688 = n4687 ^ n819 ;
  assign n4689 = n4688 ^ x116 ;
  assign n4690 = n4638 & n4689 ;
  assign n4768 = ~n4733 & n4767 ;
  assign n4769 = n4768 ^ n4733 ;
  assign n4775 = n4769 ^ n4767 ;
  assign n4782 = n4690 & n4775 ;
  assign n4771 = n4690 ^ n4689 ;
  assign n4781 = n4771 & n4775 ;
  assign n4783 = n4782 ^ n4781 ;
  assign n4777 = ~n4689 & n4768 ;
  assign n4691 = n4690 ^ n4638 ;
  assign n4779 = n4777 ^ n4691 ;
  assign n4780 = n4779 ^ n4775 ;
  assign n4784 = n4783 ^ n4780 ;
  assign n4799 = n4798 ^ n4784 ;
  assign n4793 = n4690 & n4768 ;
  assign n4792 = n4777 ^ n4768 ;
  assign n4794 = n4793 ^ n4792 ;
  assign n4791 = n4690 & ~n4769 ;
  assign n4795 = n4794 ^ n4791 ;
  assign n4796 = n4795 ^ n4781 ;
  assign n4800 = n4799 ^ n4796 ;
  assign n5841 = n4800 ^ n4794 ;
  assign n4844 = n4779 ^ n4689 ;
  assign n4772 = n4771 ^ n4638 ;
  assign n4773 = n4768 & ~n4772 ;
  assign n4841 = n4777 ^ n4773 ;
  assign n4789 = n4768 ^ n4767 ;
  assign n4801 = n4771 & n4789 ;
  assign n4802 = n4801 ^ n4800 ;
  assign n4785 = n4784 ^ n4691 ;
  assign n4776 = ~n4772 & n4775 ;
  assign n4778 = n4777 ^ n4776 ;
  assign n4786 = n4785 ^ n4778 ;
  assign n4770 = n4691 & ~n4769 ;
  assign n4774 = n4773 ^ n4770 ;
  assign n4787 = n4786 ^ n4774 ;
  assign n4788 = n4787 ^ n4779 ;
  assign n4790 = n4789 ^ n4788 ;
  assign n4803 = n4802 ^ n4790 ;
  assign n4842 = n4841 ^ n4803 ;
  assign n4843 = n4842 ^ n4776 ;
  assign n4845 = n4844 ^ n4843 ;
  assign n5842 = n5841 ^ n4845 ;
  assign n5843 = n5842 ^ n4782 ;
  assign n5838 = n5834 ^ n4607 ;
  assign n5839 = n4803 ^ n4774 ;
  assign n5840 = n5838 & n5839 ;
  assign n5844 = n5843 ^ n5840 ;
  assign n5847 = n5836 & ~n5844 ;
  assign n5848 = n5847 ^ n4778 ;
  assign n5849 = ~n5834 & n5848 ;
  assign n5850 = n5849 ^ n4778 ;
  assign n5837 = n4843 & ~n5836 ;
  assign n5851 = n5850 ^ n5837 ;
  assign n5872 = n4784 & n5835 ;
  assign n5865 = n4791 ^ n4781 ;
  assign n4868 = ~n4769 & n4771 ;
  assign n5859 = n4868 ^ n4793 ;
  assign n5860 = n5834 & ~n5859 ;
  assign n4853 = n4835 ^ n4607 ;
  assign n5861 = n5860 ^ n4853 ;
  assign n5862 = n4845 ^ n4781 ;
  assign n4874 = n4801 ^ n4793 ;
  assign n5863 = n5862 ^ n4874 ;
  assign n5864 = ~n5861 & n5863 ;
  assign n5866 = n5865 ^ n5864 ;
  assign n5868 = n5834 ^ n4786 ;
  assign n5867 = n5861 ^ n4786 ;
  assign n5869 = n5868 ^ n5867 ;
  assign n5870 = ~n5866 & ~n5869 ;
  assign n5871 = n5870 ^ n5868 ;
  assign n5873 = n5872 ^ n5871 ;
  assign n5856 = n4783 & ~n4835 ;
  assign n5857 = n5856 ^ n4786 ;
  assign n5858 = n4853 & n5857 ;
  assign n5874 = n5873 ^ n5858 ;
  assign n5875 = ~n5851 & ~n5874 ;
  assign n5876 = n5875 ^ n2734 ;
  assign n6434 = n5876 ^ x121 ;
  assign n6546 = n6433 & n6434 ;
  assign n6550 = ~n6468 & n6546 ;
  assign n5759 = n4451 ^ x108 ;
  assign n5760 = n4688 ^ x94 ;
  assign n5761 = n5759 & ~n5760 ;
  assign n5764 = n5761 ^ n5759 ;
  assign n5762 = n5761 ^ n5760 ;
  assign n5990 = n5764 ^ n5762 ;
  assign n5144 = n2201 ^ n2200 ;
  assign n5673 = n2228 & n5144 ;
  assign n5665 = n2206 ^ n2185 ;
  assign n5666 = n5665 ^ n2201 ;
  assign n5667 = n5666 ^ n2191 ;
  assign n5668 = n1176 & ~n5667 ;
  assign n5669 = n5668 ^ n2182 ;
  assign n5670 = n776 & n5669 ;
  assign n5152 = n2206 ^ n2197 ;
  assign n5153 = n2197 ^ n1176 ;
  assign n5154 = n5153 ^ n2197 ;
  assign n5155 = ~n5152 & n5154 ;
  assign n5156 = n5155 ^ n2197 ;
  assign n5157 = ~n776 & ~n5156 ;
  assign n5661 = n5157 ^ n2182 ;
  assign n5647 = n2220 ^ n2195 ;
  assign n5648 = n5647 ^ n2197 ;
  assign n5649 = n5648 ^ n2220 ;
  assign n5650 = n5649 ^ n2231 ;
  assign n5651 = n1176 & ~n5650 ;
  assign n5652 = n5651 ^ n5647 ;
  assign n5662 = n5661 ^ n5652 ;
  assign n5663 = n5662 ^ n922 ;
  assign n5653 = n5652 ^ n2191 ;
  assign n5654 = n5653 ^ n2187 ;
  assign n5655 = n5654 ^ n5652 ;
  assign n5656 = n5652 ^ n776 ;
  assign n5657 = n5656 ^ n5652 ;
  assign n5658 = n5655 & ~n5657 ;
  assign n5659 = n5658 ^ n5652 ;
  assign n5660 = ~n2228 & n5659 ;
  assign n5664 = n5663 ^ n5660 ;
  assign n5671 = n5670 ^ n5664 ;
  assign n5646 = ~n2243 & n2244 ;
  assign n5672 = n5671 ^ n5646 ;
  assign n5674 = n5673 ^ n5672 ;
  assign n5675 = n5674 ^ x77 ;
  assign n4109 = n4046 & ~n4062 ;
  assign n5698 = ~n3961 & n4042 ;
  assign n5692 = n4049 ^ n4041 ;
  assign n4055 = n4046 ^ n4022 ;
  assign n4056 = n4046 ^ n3961 ;
  assign n4057 = n4056 ^ n4046 ;
  assign n4058 = n4055 & ~n4057 ;
  assign n4059 = n4058 ^ n4046 ;
  assign n4060 = n3962 & n4059 ;
  assign n5693 = n5692 ^ n4060 ;
  assign n5694 = n5693 ^ n4392 ;
  assign n5695 = n5694 ^ n4404 ;
  assign n5696 = n5695 ^ n4369 ;
  assign n4102 = n3962 ^ n3961 ;
  assign n5685 = n4035 ^ n3983 ;
  assign n5686 = n5685 ^ n4049 ;
  assign n5687 = n4049 ^ n3962 ;
  assign n5688 = n5687 ^ n4049 ;
  assign n5689 = ~n5686 & n5688 ;
  assign n5690 = n5689 ^ n4049 ;
  assign n5691 = n4102 & ~n5690 ;
  assign n5697 = n5696 ^ n5691 ;
  assign n5699 = n5698 ^ n5697 ;
  assign n5678 = n4067 ^ n4041 ;
  assign n5676 = n4042 ^ n4041 ;
  assign n5679 = n5678 ^ n5676 ;
  assign n5680 = n5676 ^ n3961 ;
  assign n5681 = n5680 ^ n5676 ;
  assign n5682 = n5679 & n5681 ;
  assign n5683 = n5682 ^ n5676 ;
  assign n5684 = n3962 & n5683 ;
  assign n5700 = n5699 ^ n5684 ;
  assign n4051 = n4050 ^ n4046 ;
  assign n4053 = n4052 ^ n4051 ;
  assign n4054 = ~n3965 & ~n4053 ;
  assign n5701 = n5700 ^ n4054 ;
  assign n5702 = ~n4109 & n5701 ;
  assign n5703 = n5702 ^ n965 ;
  assign n5704 = n5703 ^ x125 ;
  assign n5705 = ~n5675 & n5704 ;
  assign n5706 = n4339 ^ x118 ;
  assign n5707 = n4834 ^ x91 ;
  assign n5708 = ~n5706 & n5707 ;
  assign n5712 = n5708 ^ n5706 ;
  assign n5733 = n5705 & ~n5712 ;
  assign n5714 = n5705 & ~n5706 ;
  assign n5771 = n5733 ^ n5714 ;
  assign n5717 = n5705 ^ n5704 ;
  assign n5718 = n5717 ^ n5675 ;
  assign n5719 = n5718 ^ n5704 ;
  assign n5723 = ~n5712 & ~n5719 ;
  assign n5722 = n5708 & ~n5719 ;
  assign n5724 = n5723 ^ n5722 ;
  assign n5734 = n5733 ^ n5724 ;
  assign n5735 = n5734 ^ n5712 ;
  assign n5729 = ~n5712 & n5717 ;
  assign n5730 = n5729 ^ n5722 ;
  assign n5736 = n5735 ^ n5730 ;
  assign n5731 = n5730 ^ n5723 ;
  assign n5726 = n5704 ^ n5675 ;
  assign n5727 = n5706 & ~n5726 ;
  assign n5728 = n5727 ^ n5726 ;
  assign n5732 = n5731 ^ n5728 ;
  assign n5737 = n5736 ^ n5732 ;
  assign n6469 = n5771 ^ n5737 ;
  assign n5715 = n5714 ^ n5705 ;
  assign n6470 = n6469 ^ n5715 ;
  assign n5738 = n5707 ^ n5704 ;
  assign n5739 = n5738 ^ n5675 ;
  assign n5740 = n5706 ^ n5675 ;
  assign n5741 = n5706 ^ n5704 ;
  assign n5742 = n5741 ^ n5706 ;
  assign n5743 = ~n5740 & ~n5742 ;
  assign n5744 = n5743 ^ n5706 ;
  assign n5745 = n5739 & ~n5744 ;
  assign n5746 = n5745 ^ n5733 ;
  assign n5747 = n5746 ^ n5737 ;
  assign n5709 = n5708 ^ n5707 ;
  assign n5720 = n5709 & ~n5719 ;
  assign n5721 = n5720 ^ n5719 ;
  assign n5725 = n5724 ^ n5721 ;
  assign n5748 = n5747 ^ n5725 ;
  assign n5710 = n5705 & n5709 ;
  assign n5749 = n5748 ^ n5710 ;
  assign n5713 = n5712 ^ n5707 ;
  assign n5716 = n5715 ^ n5713 ;
  assign n5750 = n5749 ^ n5716 ;
  assign n5751 = n5750 ^ n5710 ;
  assign n5752 = n5751 ^ n5720 ;
  assign n5753 = n5752 ^ n5747 ;
  assign n5754 = n5753 ^ n5727 ;
  assign n5755 = n5754 ^ n5749 ;
  assign n5756 = n5755 ^ n5720 ;
  assign n5711 = n5710 ^ n5709 ;
  assign n5757 = n5756 ^ n5711 ;
  assign n5758 = n5757 ^ n5755 ;
  assign n6471 = n6470 ^ n5758 ;
  assign n6472 = n6471 ^ n5771 ;
  assign n6473 = n5759 & n6472 ;
  assign n6474 = n6473 ^ n6469 ;
  assign n6475 = n5990 & n6474 ;
  assign n6476 = n6475 ^ n5771 ;
  assign n6481 = n5747 ^ n5715 ;
  assign n5773 = n5714 ^ n5706 ;
  assign n5774 = n5773 ^ n5731 ;
  assign n5775 = n5774 ^ n5737 ;
  assign n6482 = n6481 ^ n5775 ;
  assign n6483 = n5760 & ~n6482 ;
  assign n6484 = n6483 ^ n5753 ;
  assign n6485 = ~n5990 & ~n6484 ;
  assign n6480 = n5775 ^ n5722 ;
  assign n6486 = n6485 ^ n6480 ;
  assign n6493 = n6486 ^ n5773 ;
  assign n5802 = n5715 ^ n5710 ;
  assign n6187 = n5802 ^ n5720 ;
  assign n6487 = n6187 ^ n5733 ;
  assign n6488 = n6487 ^ n5725 ;
  assign n6489 = n6488 ^ n5755 ;
  assign n6490 = n5760 & ~n6489 ;
  assign n6491 = n6490 ^ n5733 ;
  assign n6492 = n6486 & ~n6491 ;
  assign n6494 = n6493 ^ n6492 ;
  assign n6477 = n5733 ^ n5712 ;
  assign n6478 = n6477 ^ n5732 ;
  assign n6479 = n5760 & n6478 ;
  assign n6495 = n6494 ^ n6479 ;
  assign n6496 = n5759 & ~n6495 ;
  assign n6497 = n6496 ^ n6492 ;
  assign n6498 = ~n6476 & n6497 ;
  assign n6500 = n5731 & n5764 ;
  assign n6501 = n6498 & n6500 ;
  assign n6499 = n6498 ^ n2550 ;
  assign n6502 = n6501 ^ n6499 ;
  assign n6503 = n6502 ^ x96 ;
  assign n6504 = n6468 & ~n6503 ;
  assign n6547 = n6504 ^ n6468 ;
  assign n6548 = n6546 & n6547 ;
  assign n6549 = n6548 ^ n6546 ;
  assign n6551 = n6550 ^ n6549 ;
  assign n6505 = ~n6434 & n6504 ;
  assign n6506 = n6433 & n6505 ;
  assign n6507 = n6506 ^ n6505 ;
  assign n6552 = n6551 ^ n6507 ;
  assign n4984 = n2220 ^ n2204 ;
  assign n4982 = n2237 ^ n2206 ;
  assign n4981 = n2182 ^ n2177 ;
  assign n4983 = n4982 ^ n4981 ;
  assign n4985 = n4984 ^ n4983 ;
  assign n4986 = ~n1176 & n4985 ;
  assign n4987 = n4986 ^ n4984 ;
  assign n4988 = ~n776 & n4987 ;
  assign n4977 = n2232 ^ n2197 ;
  assign n4978 = ~n2243 & ~n4977 ;
  assign n4960 = ~n2205 & n2238 ;
  assign n4963 = ~n2203 & n2215 ;
  assign n4964 = ~n4960 & n4963 ;
  assign n4961 = n4960 ^ n2240 ;
  assign n4965 = n4964 ^ n4961 ;
  assign n4974 = n4965 ^ n1417 ;
  assign n4967 = n4965 ^ n2189 ;
  assign n4966 = n4965 ^ n2211 ;
  assign n4968 = n4967 ^ n4966 ;
  assign n4969 = n4967 ^ n776 ;
  assign n4970 = n4969 ^ n4967 ;
  assign n4971 = ~n4968 & ~n4970 ;
  assign n4972 = n4971 ^ n4967 ;
  assign n4973 = ~n1176 & ~n4972 ;
  assign n4975 = n4974 ^ n4973 ;
  assign n4957 = n1949 ^ n1739 ;
  assign n4958 = ~n1518 & ~n2215 ;
  assign n4959 = ~n4957 & n4958 ;
  assign n4976 = n4975 ^ n4959 ;
  assign n4979 = n4978 ^ n4976 ;
  assign n4956 = n2194 & n2228 ;
  assign n4980 = n4979 ^ n4956 ;
  assign n4989 = n4988 ^ n4980 ;
  assign n5513 = n4989 ^ x110 ;
  assign n5512 = n4637 ^ x84 ;
  assign n5515 = n4827 ^ n3911 ;
  assign n5516 = n5515 ^ n4830 ;
  assign n5517 = n5516 ^ n4817 ;
  assign n3955 = n3916 & n3954 ;
  assign n5518 = n5517 ^ n3955 ;
  assign n5519 = n5518 ^ n1612 ;
  assign n5520 = n5519 ^ x124 ;
  assign n4913 = n4038 ^ n4023 ;
  assign n4914 = n4913 ^ n3963 ;
  assign n4915 = n4051 ^ n3965 ;
  assign n4918 = ~n4913 & ~n4915 ;
  assign n4919 = n4918 ^ n3965 ;
  assign n4920 = n4914 & ~n4919 ;
  assign n4906 = n4066 ^ n4029 ;
  assign n4907 = n4906 ^ n4077 ;
  assign n4911 = ~n3964 & n4907 ;
  assign n4908 = n4410 ^ n3961 ;
  assign n4912 = n4911 ^ n4908 ;
  assign n4921 = n4920 ^ n4912 ;
  assign n4901 = n4073 ^ n3962 ;
  assign n4902 = n4901 ^ n4073 ;
  assign n4903 = ~n4075 & n4902 ;
  assign n4904 = n4903 ^ n4073 ;
  assign n4905 = n3961 & n4904 ;
  assign n4922 = n4921 ^ n4905 ;
  assign n4923 = n4922 ^ n4061 ;
  assign n4080 = n4079 ^ n4076 ;
  assign n4081 = n4080 ^ n4053 ;
  assign n4082 = n4053 ^ n3961 ;
  assign n4083 = n4082 ^ n4053 ;
  assign n4084 = ~n4081 & n4083 ;
  assign n4085 = n4084 ^ n4053 ;
  assign n4086 = ~n3962 & ~n4085 ;
  assign n4924 = n4923 ^ n4086 ;
  assign n4925 = n4924 ^ n4366 ;
  assign n4926 = n4925 ^ n4054 ;
  assign n4927 = n4926 ^ n4109 ;
  assign n4928 = n4927 ^ n1215 ;
  assign n5521 = n4928 ^ x101 ;
  assign n5522 = n5520 & ~n5521 ;
  assign n5523 = n5522 ^ n5520 ;
  assign n5524 = n5523 ^ n5521 ;
  assign n5543 = n4680 ^ n3461 ;
  assign n5544 = n5543 ^ n3470 ;
  assign n5545 = n5544 ^ n3516 ;
  assign n5546 = n5545 ^ n4680 ;
  assign n5547 = n3444 & ~n5546 ;
  assign n5548 = n5547 ^ n5543 ;
  assign n5549 = n3443 & n5548 ;
  assign n5540 = n3460 ^ n3428 ;
  assign n5541 = ~n3475 & ~n5540 ;
  assign n5533 = n4676 ^ n3437 ;
  assign n5534 = n5533 ^ n4680 ;
  assign n5535 = n5534 ^ n4640 ;
  assign n5536 = n5535 ^ n3476 ;
  assign n5537 = n5536 ^ n4478 ;
  assign n5538 = n5537 ^ n1595 ;
  assign n5525 = n3458 ^ n3437 ;
  assign n5526 = n5525 ^ n3467 ;
  assign n5527 = n5526 ^ n5525 ;
  assign n5528 = n5525 ^ n3444 ;
  assign n5529 = n5528 ^ n5525 ;
  assign n5530 = n5527 & n5529 ;
  assign n5531 = n5530 ^ n5525 ;
  assign n5532 = n4662 & n5531 ;
  assign n5539 = n5538 ^ n5532 ;
  assign n5542 = n5541 ^ n5539 ;
  assign n5550 = n5549 ^ n5542 ;
  assign n5551 = n5550 ^ x86 ;
  assign n5552 = n4606 ^ x75 ;
  assign n5553 = n5551 & ~n5552 ;
  assign n5562 = n5553 ^ n5551 ;
  assign n5575 = n5524 & n5562 ;
  assign n5563 = n5562 ^ n5552 ;
  assign n5564 = n5524 & n5563 ;
  assign n5576 = n5575 ^ n5564 ;
  assign n5554 = n5553 ^ n5552 ;
  assign n5555 = n5524 & ~n5554 ;
  assign n5574 = n5555 ^ n5524 ;
  assign n5577 = n5576 ^ n5574 ;
  assign n5557 = n5522 & n5553 ;
  assign n5556 = n5523 & n5553 ;
  assign n5558 = n5557 ^ n5556 ;
  assign n5580 = n5577 ^ n5558 ;
  assign n5581 = n5580 ^ n5553 ;
  assign n5579 = n5523 & ~n5554 ;
  assign n5582 = n5581 ^ n5579 ;
  assign n5571 = n5521 ^ n5520 ;
  assign n5583 = n5582 ^ n5571 ;
  assign n5560 = n5522 & ~n5554 ;
  assign n5578 = n5577 ^ n5560 ;
  assign n5584 = n5583 ^ n5578 ;
  assign n5572 = n5571 ^ n5552 ;
  assign n5559 = n5558 ^ n5555 ;
  assign n5573 = n5572 ^ n5559 ;
  assign n5585 = n5584 ^ n5573 ;
  assign n6122 = n5585 ^ n5582 ;
  assign n6123 = n5512 & ~n6122 ;
  assign n6124 = n6123 ^ n5582 ;
  assign n6534 = n5513 & n6124 ;
  assign n5614 = n5512 & ~n5513 ;
  assign n5615 = n5614 ^ n5513 ;
  assign n5616 = n5615 ^ n5512 ;
  assign n5617 = n5616 ^ n5513 ;
  assign n6258 = n5578 & n5617 ;
  assign n5590 = n5585 ^ n5556 ;
  assign n5591 = n5590 ^ n5523 ;
  assign n5588 = n5585 ^ n5579 ;
  assign n5587 = n5523 & n5562 ;
  assign n5589 = n5588 ^ n5587 ;
  assign n5592 = n5591 ^ n5589 ;
  assign n5593 = n5592 ^ n5581 ;
  assign n5566 = n5552 ^ n5520 ;
  assign n5567 = n5551 ^ n5521 ;
  assign n5568 = n5552 & n5567 ;
  assign n5569 = n5568 ^ n5521 ;
  assign n5570 = ~n5566 & ~n5569 ;
  assign n5586 = n5585 ^ n5570 ;
  assign n5594 = n5593 ^ n5586 ;
  assign n6138 = n5594 ^ n5563 ;
  assign n5598 = n5522 & n5562 ;
  assign n5619 = n5598 ^ n5592 ;
  assign n5620 = n5619 ^ n5564 ;
  assign n5621 = n5620 ^ n5568 ;
  assign n6139 = n6138 ^ n5621 ;
  assign n6140 = ~n5512 & ~n6139 ;
  assign n5622 = n5621 ^ n5564 ;
  assign n6141 = n6140 ^ n5622 ;
  assign n6142 = n5513 & n6141 ;
  assign n6530 = n6258 ^ n6142 ;
  assign n6517 = n5570 ^ n5551 ;
  assign n6515 = n5619 ^ n5555 ;
  assign n5599 = n5598 ^ n5575 ;
  assign n6508 = n5616 ^ n5599 ;
  assign n6509 = n5614 ^ n5590 ;
  assign n6510 = n5614 ^ n5599 ;
  assign n6511 = n6510 ^ n5614 ;
  assign n6512 = n6509 & ~n6511 ;
  assign n6513 = n6512 ^ n5614 ;
  assign n6514 = n6508 & n6513 ;
  assign n6516 = n6515 ^ n6514 ;
  assign n6518 = n6517 ^ n6516 ;
  assign n6519 = n6518 ^ n6514 ;
  assign n6520 = ~n5513 & ~n6519 ;
  assign n6521 = n6520 ^ n6516 ;
  assign n6531 = n6530 ^ n6521 ;
  assign n6532 = n6531 ^ n2303 ;
  assign n6522 = n6521 ^ n6514 ;
  assign n6127 = n5599 ^ n5592 ;
  assign n6128 = n6127 ^ n5594 ;
  assign n6126 = n5598 ^ n5577 ;
  assign n6129 = n6128 ^ n6126 ;
  assign n6130 = n6129 ^ n5572 ;
  assign n6523 = n6522 ^ n6130 ;
  assign n6524 = n6523 ^ n6522 ;
  assign n6527 = ~n5513 & n6524 ;
  assign n6528 = n6527 ^ n6522 ;
  assign n6529 = ~n5512 & ~n6528 ;
  assign n6533 = n6532 ^ n6529 ;
  assign n6535 = n6534 ^ n6533 ;
  assign n6536 = n6535 ^ x82 ;
  assign n3939 = n3938 ^ n3937 ;
  assign n3924 = ~n3914 & ~n3923 ;
  assign n3940 = n3939 ^ n3924 ;
  assign n3941 = n3911 & n3940 ;
  assign n3942 = n3941 ^ n3939 ;
  assign n3956 = n3955 ^ n3942 ;
  assign n3945 = n3942 ^ n3935 ;
  assign n3944 = n3943 ^ n3942 ;
  assign n3946 = n3945 ^ n3944 ;
  assign n3949 = n3911 & n3946 ;
  assign n3950 = n3949 ^ n3945 ;
  assign n3951 = ~n3910 & n3950 ;
  assign n3957 = n3956 ^ n3951 ;
  assign n3958 = ~n3909 & ~n3957 ;
  assign n3959 = n3958 ^ n1238 ;
  assign n4898 = n3959 ^ x117 ;
  assign n4929 = n4928 ^ x68 ;
  assign n4930 = ~n4898 & n4929 ;
  assign n4931 = n4930 ^ n4929 ;
  assign n4932 = n4931 ^ n4898 ;
  assign n4953 = n3777 ^ n1308 ;
  assign n4947 = n3753 ^ n3704 ;
  assign n4948 = n3774 & ~n4947 ;
  assign n4943 = n3762 ^ n3725 ;
  assign n4944 = ~n4611 & n4943 ;
  assign n4941 = n4612 ^ n3774 ;
  assign n4942 = ~n4617 & n4941 ;
  assign n4945 = n4944 ^ n4942 ;
  assign n4946 = n4945 ^ n3707 ;
  assign n4949 = n4948 ^ n4946 ;
  assign n4933 = n3739 ^ n3728 ;
  assign n4934 = n4933 ^ n3692 ;
  assign n4935 = n4934 ^ n3728 ;
  assign n4936 = n3728 ^ n3554 ;
  assign n4937 = n4936 ^ n3728 ;
  assign n4938 = n4935 & n4937 ;
  assign n4939 = n4938 ^ n3728 ;
  assign n4940 = n3589 & ~n4939 ;
  assign n4950 = n4949 ^ n4940 ;
  assign n4951 = n4633 & n4950 ;
  assign n4952 = ~n3718 & n4951 ;
  assign n4954 = n4953 ^ n4952 ;
  assign n4955 = n4954 ^ x67 ;
  assign n4990 = n4989 ^ x100 ;
  assign n4991 = ~n4955 & n4990 ;
  assign n4992 = n4991 ^ n4955 ;
  assign n4197 = n3336 ^ n1339 ;
  assign n4178 = n3337 ^ n3275 ;
  assign n4183 = n4178 ^ n3302 ;
  assign n4184 = n4183 ^ n3318 ;
  assign n4179 = n3295 ^ n3265 ;
  assign n4180 = n4179 ^ n3315 ;
  assign n4181 = n4180 ^ n3302 ;
  assign n4182 = ~n3308 & ~n4181 ;
  assign n4185 = n4184 ^ n4182 ;
  assign n4186 = ~n4178 & n4185 ;
  assign n4187 = n3164 & ~n4186 ;
  assign n4198 = n4197 ^ n4187 ;
  assign n4192 = n3256 ^ n3164 ;
  assign n4193 = n4192 ^ n3256 ;
  assign n4194 = n3297 & ~n4193 ;
  assign n4195 = n4194 ^ n3256 ;
  assign n4196 = n3308 & n4195 ;
  assign n4199 = n4198 ^ n4196 ;
  assign n4177 = n3276 ^ n3271 ;
  assign n4188 = n3326 & ~n4187 ;
  assign n4189 = n4177 & n4188 ;
  assign n4200 = n4199 ^ n4189 ;
  assign n4170 = n3336 ^ n3290 ;
  assign n4171 = n4170 ^ n3336 ;
  assign n4172 = n3336 ^ n3164 ;
  assign n4173 = n4172 ^ n3336 ;
  assign n4174 = n4171 & ~n4173 ;
  assign n4175 = n4174 ^ n3336 ;
  assign n4176 = ~n3308 & n4175 ;
  assign n4201 = n4200 ^ n4176 ;
  assign n4995 = n4201 ^ x78 ;
  assign n5015 = n2823 ^ n2761 ;
  assign n5016 = n5015 ^ n4336 ;
  assign n5017 = n5016 ^ n1380 ;
  assign n5010 = n2790 ^ n2766 ;
  assign n5011 = n5010 ^ n2772 ;
  assign n5012 = ~n2332 & ~n5011 ;
  assign n5013 = n5012 ^ n2761 ;
  assign n5014 = ~n2304 & ~n5013 ;
  assign n5018 = n5017 ^ n5014 ;
  assign n5003 = n2796 ^ n2741 ;
  assign n5004 = n5003 ^ n2758 ;
  assign n5005 = n5004 ^ n2796 ;
  assign n5006 = n5005 ^ n4702 ;
  assign n5007 = n2332 & ~n5006 ;
  assign n5008 = n5007 ^ n5003 ;
  assign n5009 = n2333 & n5008 ;
  assign n5019 = n5018 ^ n5009 ;
  assign n4996 = n2814 ^ n2756 ;
  assign n4997 = n4996 ^ n2800 ;
  assign n4998 = n4997 ^ n4717 ;
  assign n4999 = ~n2744 & n4998 ;
  assign n5000 = n4999 ^ n2800 ;
  assign n5001 = n2786 ^ n2744 ;
  assign n5002 = ~n5000 & ~n5001 ;
  assign n5020 = n5019 ^ n5002 ;
  assign n5021 = n5020 ^ x85 ;
  assign n5022 = ~n4995 & ~n5021 ;
  assign n5034 = n5022 ^ n4995 ;
  assign n5043 = n5034 ^ n5021 ;
  assign n5044 = ~n4992 & ~n5043 ;
  assign n5469 = n4932 & n5044 ;
  assign n5030 = n4995 ^ n4955 ;
  assign n5031 = n4995 ^ n4990 ;
  assign n5032 = n5030 & n5031 ;
  assign n5037 = n5032 ^ n4995 ;
  assign n5038 = n5030 ^ n5021 ;
  assign n5039 = ~n5037 & ~n5038 ;
  assign n5028 = n4991 & n5022 ;
  assign n5046 = n5039 ^ n5028 ;
  assign n5042 = ~n4992 & n5022 ;
  assign n5045 = n5044 ^ n5042 ;
  assign n5047 = n5046 ^ n5045 ;
  assign n4993 = n4992 ^ n4990 ;
  assign n5041 = n4993 & n5022 ;
  assign n5048 = n5047 ^ n5041 ;
  assign n5049 = n5048 ^ n5044 ;
  assign n5040 = n5039 ^ n5022 ;
  assign n5050 = n5049 ^ n5040 ;
  assign n5023 = n5022 ^ n5021 ;
  assign n5024 = n4990 & ~n5023 ;
  assign n5027 = n4955 & n5024 ;
  assign n5036 = n5027 ^ n5024 ;
  assign n5051 = n5050 ^ n5036 ;
  assign n4994 = n4993 ^ n4955 ;
  assign n5035 = n4994 & ~n5034 ;
  assign n5052 = n5051 ^ n5035 ;
  assign n5053 = n5052 ^ n5027 ;
  assign n5054 = n5053 ^ n5044 ;
  assign n5033 = n5032 ^ n5023 ;
  assign n5055 = n5054 ^ n5033 ;
  assign n5056 = n5055 ^ n5023 ;
  assign n5057 = n5056 ^ n5024 ;
  assign n5058 = n5057 ^ n5049 ;
  assign n5059 = n5058 ^ n5030 ;
  assign n5060 = n5059 ^ n5052 ;
  assign n5458 = n5060 ^ n4929 ;
  assign n5459 = n5458 ^ n5060 ;
  assign n5462 = n5047 & ~n5459 ;
  assign n5463 = n5462 ^ n5060 ;
  assign n5464 = n4898 & n5463 ;
  assign n5465 = n5464 ^ n5060 ;
  assign n5442 = n4990 ^ n4955 ;
  assign n5443 = n5021 & n5442 ;
  assign n5029 = n5028 ^ n5027 ;
  assign n5061 = n5060 ^ n5029 ;
  assign n5025 = n5024 ^ n4994 ;
  assign n5026 = n5025 ^ n4990 ;
  assign n5062 = n5061 ^ n5026 ;
  assign n5439 = n5062 ^ n5051 ;
  assign n5430 = n5035 ^ n5028 ;
  assign n5089 = n5057 ^ n5055 ;
  assign n5429 = n5089 ^ n5048 ;
  assign n5431 = n5430 ^ n5429 ;
  assign n5432 = n5431 ^ n5089 ;
  assign n5433 = n5089 ^ n4929 ;
  assign n5434 = n5433 ^ n5089 ;
  assign n5435 = n5432 & n5434 ;
  assign n5436 = n5435 ^ n5089 ;
  assign n5437 = ~n4898 & ~n5436 ;
  assign n5440 = n5439 ^ n5437 ;
  assign n5087 = n5057 ^ n4992 ;
  assign n5088 = n5087 ^ n5045 ;
  assign n5099 = n5088 ^ n5029 ;
  assign n5438 = n5099 ^ n5055 ;
  assign n5441 = n5440 ^ n5438 ;
  assign n5444 = n5443 ^ n5441 ;
  assign n5445 = n5444 ^ n5437 ;
  assign n5446 = n4929 & n5445 ;
  assign n5447 = n5446 ^ n5440 ;
  assign n5466 = n5465 ^ n5447 ;
  assign n5428 = n4929 ^ n4898 ;
  assign n5100 = n5052 ^ n5025 ;
  assign n5101 = n5100 ^ n5042 ;
  assign n5451 = n5101 ^ n5057 ;
  assign n5452 = n5451 ^ n5050 ;
  assign n5455 = ~n4929 & n5452 ;
  assign n5448 = n5447 ^ n5437 ;
  assign n5456 = n5455 ^ n5448 ;
  assign n5457 = n5428 & n5456 ;
  assign n5467 = n5466 ^ n5457 ;
  assign n5063 = n5062 ^ n5036 ;
  assign n5064 = n4932 & n5063 ;
  assign n5468 = n5467 ^ n5064 ;
  assign n5470 = n5469 ^ n5468 ;
  assign n5111 = n5055 ^ n4993 ;
  assign n5112 = n5111 ^ n5048 ;
  assign n5113 = n5112 ^ n5088 ;
  assign n5114 = n5113 ^ n5100 ;
  assign n5115 = n5100 ^ n4929 ;
  assign n5116 = n5115 ^ n5100 ;
  assign n5117 = n5114 & ~n5116 ;
  assign n5118 = n5117 ^ n5100 ;
  assign n5119 = ~n4898 & n5118 ;
  assign n5471 = n5470 ^ n5119 ;
  assign n5472 = n5471 ^ n2331 ;
  assign n6537 = n5472 ^ x89 ;
  assign n6538 = ~n6536 & n6537 ;
  assign n6539 = n6538 ^ n6536 ;
  assign n6563 = n6539 ^ n6537 ;
  assign n7440 = n6552 & n6563 ;
  assign n6557 = n6505 ^ n6504 ;
  assign n6558 = n6557 ^ n6551 ;
  assign n6554 = n6546 ^ n6434 ;
  assign n6555 = n6503 & n6554 ;
  assign n6556 = n6555 ^ n6554 ;
  assign n6559 = n6558 ^ n6556 ;
  assign n6543 = n6434 ^ n6433 ;
  assign n6544 = n6543 ^ n6468 ;
  assign n6545 = ~n6503 & n6544 ;
  assign n6553 = n6552 ^ n6545 ;
  assign n6560 = n6559 ^ n6553 ;
  assign n6540 = ~n6434 & ~n6468 ;
  assign n6541 = n6503 & n6540 ;
  assign n6542 = n6541 ^ n6540 ;
  assign n6561 = n6560 ^ n6542 ;
  assign n6562 = ~n6539 & n6561 ;
  assign n7441 = n7440 ^ n6562 ;
  assign n7954 = n7441 ^ n4339 ;
  assign n6579 = n6505 ^ n6434 ;
  assign n6580 = n6579 ^ n6540 ;
  assign n6581 = ~n6433 & ~n6580 ;
  assign n6609 = n6581 ^ n6580 ;
  assign n6616 = n6609 ^ n6559 ;
  assign n6617 = n6559 ^ n6537 ;
  assign n6618 = n6617 ^ n6559 ;
  assign n6619 = ~n6616 & n6618 ;
  assign n6620 = n6619 ^ n6559 ;
  assign n6621 = n6536 & n6620 ;
  assign n7955 = n7954 ^ n6621 ;
  assign n6587 = n6580 ^ n6547 ;
  assign n6588 = n6587 ^ n6556 ;
  assign n6589 = n6588 ^ n6434 ;
  assign n6590 = n6589 ^ n6549 ;
  assign n6601 = n6590 ^ n6555 ;
  assign n6611 = n6601 ^ n6506 ;
  assign n6612 = ~n6539 & ~n6611 ;
  assign n6570 = n6560 ^ n6555 ;
  assign n7452 = n6581 ^ n6570 ;
  assign n7945 = n6581 ^ n6536 ;
  assign n7946 = n7945 ^ n6581 ;
  assign n7947 = n7452 & ~n7946 ;
  assign n7948 = n7947 ^ n6581 ;
  assign n7949 = ~n6537 & n7948 ;
  assign n6565 = n6537 ^ n6536 ;
  assign n6566 = n6503 & n6550 ;
  assign n7938 = n6548 ^ n6537 ;
  assign n7939 = n7938 ^ n6548 ;
  assign n7940 = n6566 & n7939 ;
  assign n7941 = n7940 ^ n6548 ;
  assign n7942 = n6565 & n7941 ;
  assign n7950 = n7949 ^ n7942 ;
  assign n6568 = ~n6433 & n6541 ;
  assign n7923 = n6601 ^ n6568 ;
  assign n7924 = n7923 ^ n6507 ;
  assign n6567 = n6566 ^ n6550 ;
  assign n7451 = n6567 ^ n6561 ;
  assign n7922 = n7451 ^ n6559 ;
  assign n7925 = n7924 ^ n7922 ;
  assign n7918 = n6558 ^ n6505 ;
  assign n7919 = n7918 ^ n6581 ;
  assign n7920 = n7919 ^ n6568 ;
  assign n7921 = ~n6536 & n7920 ;
  assign n7926 = n7925 ^ n7921 ;
  assign n7935 = n7926 ^ n6548 ;
  assign n7951 = n7950 ^ n7935 ;
  assign n6586 = n6568 ^ n6541 ;
  assign n6591 = n6590 ^ n6586 ;
  assign n7928 = n6591 ^ n6558 ;
  assign n7929 = n7928 ^ n6609 ;
  assign n7930 = n7929 ^ n7926 ;
  assign n7917 = n6581 ^ n6567 ;
  assign n7927 = n7926 ^ n7917 ;
  assign n7931 = n7930 ^ n7927 ;
  assign n7932 = ~n6536 & n7931 ;
  assign n7933 = n7932 ^ n7930 ;
  assign n7934 = ~n6537 & ~n7933 ;
  assign n7952 = n7951 ^ n7934 ;
  assign n7953 = ~n6612 & n7952 ;
  assign n7956 = n7955 ^ n7953 ;
  assign n8185 = n7956 ^ x86 ;
  assign n4127 = n2256 ^ x72 ;
  assign n4162 = n4161 ^ n1972 ;
  assign n4135 = n3104 ^ n3020 ;
  assign n4136 = n3072 ^ n3019 ;
  assign n4137 = n4136 ^ n3039 ;
  assign n4138 = n3058 & ~n4137 ;
  assign n4139 = ~n4135 & n4138 ;
  assign n4140 = n4139 ^ n3058 ;
  assign n4147 = n4140 ^ n3021 ;
  assign n4142 = n3071 & n4141 ;
  assign n4143 = ~n3023 & n4142 ;
  assign n4144 = n4143 ^ n3094 ;
  assign n4145 = ~n3094 & ~n4144 ;
  assign n4146 = ~n4140 & n4145 ;
  assign n4148 = n4147 ^ n4146 ;
  assign n4149 = n4148 ^ n4140 ;
  assign n4150 = n4149 ^ n4146 ;
  assign n4151 = n4150 ^ n4149 ;
  assign n4152 = n4149 ^ n3036 ;
  assign n4153 = n4152 ^ n4149 ;
  assign n4154 = n4151 & n4153 ;
  assign n4155 = n4154 ^ n4149 ;
  assign n4156 = ~n3063 & n4155 ;
  assign n4157 = n4156 ^ n4148 ;
  assign n4158 = n4157 ^ n3011 ;
  assign n4128 = n3075 ^ n3021 ;
  assign n4130 = n4129 ^ n4128 ;
  assign n4131 = n4130 ^ n3062 ;
  assign n4132 = n2874 & n4131 ;
  assign n4133 = n4132 ^ n3011 ;
  assign n4134 = n3094 & n4133 ;
  assign n4159 = n4158 ^ n4134 ;
  assign n4160 = ~n3057 & ~n4159 ;
  assign n4163 = n4162 ^ n4160 ;
  assign n4164 = n4163 ^ x112 ;
  assign n4165 = n4127 & ~n4164 ;
  assign n3960 = n3959 ^ x74 ;
  assign n4088 = n3961 & ~n4048 ;
  assign n4089 = n4088 ^ n4046 ;
  assign n4090 = n4089 ^ n4049 ;
  assign n4091 = n4090 ^ n4040 ;
  assign n4092 = n4091 ^ n4089 ;
  assign n4095 = ~n3961 & ~n4092 ;
  assign n4096 = n4095 ^ n4089 ;
  assign n4097 = ~n3962 & n4096 ;
  assign n4098 = n4097 ^ n4089 ;
  assign n4117 = ~n3965 & n4023 ;
  assign n4115 = n3963 & n4066 ;
  assign n4112 = n4036 ^ n4025 ;
  assign n4113 = n4112 ^ n4078 ;
  assign n4100 = n4077 ^ n4069 ;
  assign n4107 = n4100 ^ n4038 ;
  assign n4099 = n4053 ^ n4049 ;
  assign n4101 = n4100 ^ n4099 ;
  assign n4103 = n4099 ^ n3962 ;
  assign n4104 = ~n4102 & n4103 ;
  assign n4105 = n4104 ^ n3962 ;
  assign n4106 = ~n4101 & ~n4105 ;
  assign n4108 = n4107 ^ n4106 ;
  assign n4114 = n4113 ^ n4108 ;
  assign n4116 = n4115 ^ n4114 ;
  assign n4118 = n4117 ^ n4116 ;
  assign n4119 = ~n4111 & n4118 ;
  assign n4110 = n4109 ^ n4108 ;
  assign n4120 = n4119 ^ n4110 ;
  assign n4121 = ~n4098 & n4120 ;
  assign n4065 = n4064 ^ n4060 ;
  assign n4087 = n4086 ^ n4065 ;
  assign n4122 = n4121 ^ n4087 ;
  assign n4123 = ~n4054 & n4122 ;
  assign n4124 = n4123 ^ n2052 ;
  assign n4125 = n4124 ^ x122 ;
  assign n4126 = ~n3960 & n4125 ;
  assign n4206 = n4126 ^ n3960 ;
  assign n4207 = n4206 ^ n4125 ;
  assign n4219 = n4207 ^ n3960 ;
  assign n4225 = n4165 & n4219 ;
  assign n4269 = n4225 ^ n4219 ;
  assign n4166 = n4165 ^ n4164 ;
  assign n4167 = n4166 ^ n4127 ;
  assign n4215 = n4126 & n4167 ;
  assign n4168 = n4167 ^ n4164 ;
  assign n4169 = n4126 & n4168 ;
  assign n4226 = n4215 ^ n4169 ;
  assign n4227 = n4226 ^ n4225 ;
  assign n4223 = n4164 ^ n3960 ;
  assign n4224 = n4125 & n4223 ;
  assign n4228 = n4227 ^ n4224 ;
  assign n4220 = n4167 & n4219 ;
  assign n4248 = n4228 ^ n4220 ;
  assign n4270 = n4269 ^ n4248 ;
  assign n4202 = n4201 ^ x98 ;
  assign n4203 = n3525 ^ x105 ;
  assign n4204 = n4202 & n4203 ;
  assign n4253 = n4167 & n4207 ;
  assign n4273 = n4253 ^ n4207 ;
  assign n4232 = n4126 & ~n4166 ;
  assign n4233 = n4232 ^ n4126 ;
  assign n4234 = n4233 ^ n4226 ;
  assign n4231 = ~n4166 & ~n4206 ;
  assign n4235 = n4234 ^ n4231 ;
  assign n4236 = n4235 ^ n4169 ;
  assign n4229 = n4228 ^ n4215 ;
  assign n4222 = n4166 ^ n4126 ;
  assign n4230 = n4229 ^ n4222 ;
  assign n4237 = n4236 ^ n4230 ;
  assign n4208 = n4168 & n4207 ;
  assign n4239 = n4237 ^ n4208 ;
  assign n4274 = n4273 ^ n4239 ;
  assign n5418 = n4204 & ~n4274 ;
  assign n4205 = n4169 & n4204 ;
  assign n5419 = n5418 ^ n4205 ;
  assign n4289 = n4204 ^ n4202 ;
  assign n4291 = n4231 & n4289 ;
  assign n4290 = n4169 & n4289 ;
  assign n4292 = n4291 ^ n4290 ;
  assign n5420 = n5419 ^ n4292 ;
  assign n4251 = n4168 & ~n4206 ;
  assign n4258 = n4251 ^ n4167 ;
  assign n4256 = n4248 ^ n4231 ;
  assign n4252 = n4251 ^ n4231 ;
  assign n4254 = n4253 ^ n4252 ;
  assign n4255 = n4254 ^ n4229 ;
  assign n4257 = n4256 ^ n4255 ;
  assign n4259 = n4258 ^ n4257 ;
  assign n4262 = n4259 ^ n4229 ;
  assign n4263 = n4262 ^ n4234 ;
  assign n5401 = n4263 ^ n4208 ;
  assign n4271 = n4253 ^ n4225 ;
  assign n4265 = n4252 ^ n4206 ;
  assign n4266 = n4265 ^ n4259 ;
  assign n4267 = n4266 ^ n4232 ;
  assign n4268 = n4267 ^ n4220 ;
  assign n5400 = n4271 ^ n4268 ;
  assign n5402 = n5401 ^ n5400 ;
  assign n5403 = ~n4203 & ~n5402 ;
  assign n5404 = n5403 ^ n5401 ;
  assign n5421 = n5420 ^ n5404 ;
  assign n4297 = n4204 ^ n4203 ;
  assign n4298 = n4297 ^ n4202 ;
  assign n4299 = ~n4274 & ~n4298 ;
  assign n5422 = n5421 ^ n4299 ;
  assign n5412 = n4259 ^ n4225 ;
  assign n5413 = n5412 ^ n4228 ;
  assign n4241 = n4228 ^ n4203 ;
  assign n5414 = n4241 ^ n4228 ;
  assign n5415 = n5413 & ~n5414 ;
  assign n5416 = n5415 ^ n4228 ;
  assign n5417 = ~n4202 & n5416 ;
  assign n5423 = n5422 ^ n5417 ;
  assign n5406 = n4230 ^ n3960 ;
  assign n5407 = n5406 ^ n5404 ;
  assign n4221 = n4220 ^ n4208 ;
  assign n5399 = n4235 ^ n4221 ;
  assign n5405 = n5404 ^ n5399 ;
  assign n5408 = n5407 ^ n5405 ;
  assign n5409 = ~n4203 & n5408 ;
  assign n5410 = n5409 ^ n5407 ;
  assign n5411 = ~n4202 & n5410 ;
  assign n5424 = n5423 ^ n5411 ;
  assign n5425 = ~n4270 & ~n5424 ;
  assign n5426 = n5425 ^ n3655 ;
  assign n5427 = n5426 ^ x114 ;
  assign n5473 = n5472 ^ x64 ;
  assign n5125 = n4359 ^ x96 ;
  assign n5126 = n2825 ^ x123 ;
  assign n5127 = n5125 & ~n5126 ;
  assign n5128 = n5127 ^ n5126 ;
  assign n5129 = n5128 ^ n5125 ;
  assign n5191 = n5129 ^ n5126 ;
  assign n5162 = n2231 ^ n2195 ;
  assign n5163 = n1177 & n5162 ;
  assign n5145 = n5144 ^ n4982 ;
  assign n5142 = n2232 ^ n2212 ;
  assign n5143 = n5142 ^ n2219 ;
  assign n5146 = n5145 ^ n5143 ;
  assign n5147 = ~n1176 & n5146 ;
  assign n5148 = n5147 ^ n5143 ;
  assign n5158 = n5148 ^ n1794 ;
  assign n5159 = n5158 ^ n5157 ;
  assign n5149 = n5148 ^ n2195 ;
  assign n5139 = n2243 ^ n2219 ;
  assign n5140 = n5139 ^ n2197 ;
  assign n5141 = ~n2216 & n5140 ;
  assign n5150 = n5149 ^ n5141 ;
  assign n5151 = n776 & n5150 ;
  assign n5160 = n5159 ^ n5151 ;
  assign n5138 = n2178 & n2228 ;
  assign n5161 = n5160 ^ n5138 ;
  assign n5164 = n5163 ^ n5161 ;
  assign n5137 = n2189 & ~n2215 ;
  assign n5165 = n5164 ^ n5137 ;
  assign n5130 = n2204 ^ n2201 ;
  assign n5131 = n5130 ^ n2240 ;
  assign n5132 = n2240 ^ n1176 ;
  assign n5133 = n5132 ^ n2240 ;
  assign n5134 = n5131 & ~n5133 ;
  assign n5135 = n5134 ^ n2240 ;
  assign n5136 = n2228 & n5135 ;
  assign n5166 = n5165 ^ n5136 ;
  assign n5167 = n5166 ^ x113 ;
  assign n5181 = ~n3909 & n3911 ;
  assign n5185 = n3910 & n3939 ;
  assign n5186 = n5181 & n5185 ;
  assign n5182 = n5181 ^ n1810 ;
  assign n5179 = n4832 ^ n3911 ;
  assign n5169 = n3935 ^ n3924 ;
  assign n5170 = ~n3911 & ~n5169 ;
  assign n5171 = n5170 ^ n3935 ;
  assign n5180 = n5179 ^ n5171 ;
  assign n5183 = n5182 ^ n5180 ;
  assign n5168 = n3911 ^ n3910 ;
  assign n5172 = n5171 ^ n3910 ;
  assign n5173 = n5172 ^ n5171 ;
  assign n5174 = n5171 ^ n4814 ;
  assign n5175 = n5174 ^ n5171 ;
  assign n5176 = ~n5173 & ~n5175 ;
  assign n5177 = n5176 ^ n5171 ;
  assign n5178 = ~n5168 & n5177 ;
  assign n5184 = n5183 ^ n5178 ;
  assign n5187 = n5186 ^ n5184 ;
  assign n5188 = n5187 ^ x114 ;
  assign n5189 = n5167 & n5188 ;
  assign n5196 = n5189 ^ n5167 ;
  assign n5197 = n5191 & n5196 ;
  assign n5194 = n5189 ^ n5188 ;
  assign n5195 = n5191 & n5194 ;
  assign n5198 = n5197 ^ n5195 ;
  assign n5192 = n5189 & n5191 ;
  assign n5193 = n5192 ^ n5191 ;
  assign n5199 = n5198 ^ n5193 ;
  assign n5123 = n4418 ^ x81 ;
  assign n5124 = n3123 ^ x120 ;
  assign n5237 = ~n5123 & n5124 ;
  assign n5266 = n5237 ^ n5124 ;
  assign n5267 = n5266 ^ n5123 ;
  assign n5268 = n5267 ^ n5124 ;
  assign n5282 = n5199 & ~n5268 ;
  assign n5505 = n5282 ^ n3982 ;
  assign n5212 = n5196 ^ n5188 ;
  assign n5213 = n5129 & ~n5212 ;
  assign n5203 = n5129 & n5194 ;
  assign n5214 = n5213 ^ n5203 ;
  assign n5190 = n5129 & n5189 ;
  assign n5211 = n5190 ^ n5129 ;
  assign n5215 = n5214 ^ n5211 ;
  assign n5243 = n5215 ^ n5197 ;
  assign n5240 = n5127 & n5189 ;
  assign n5227 = n5127 & ~n5167 ;
  assign n5228 = n5227 ^ n5127 ;
  assign n5241 = n5240 ^ n5228 ;
  assign n5242 = n5241 ^ n5196 ;
  assign n5244 = n5243 ^ n5242 ;
  assign n5225 = n5127 & ~n5212 ;
  assign n5239 = n5227 ^ n5225 ;
  assign n5245 = n5244 ^ n5239 ;
  assign n5493 = n5245 ^ n5228 ;
  assign n5494 = ~n5268 & n5493 ;
  assign n5210 = n5124 ^ n5123 ;
  assign n5480 = n5244 ^ n5240 ;
  assign n5481 = n5480 ^ n5195 ;
  assign n5482 = n5481 ^ n5190 ;
  assign n5489 = n5482 ^ n5203 ;
  assign n5484 = n5215 ^ n5195 ;
  assign n5238 = ~n5128 & ~n5212 ;
  assign n5485 = n5484 ^ n5238 ;
  assign n5486 = n5485 ^ n5241 ;
  assign n5483 = n5482 ^ n5197 ;
  assign n5487 = n5486 ^ n5483 ;
  assign n5488 = ~n5123 & n5487 ;
  assign n5490 = n5489 ^ n5488 ;
  assign n5491 = n5210 & n5490 ;
  assign n5249 = n5192 ^ n5190 ;
  assign n5250 = n5249 ^ n5225 ;
  assign n5251 = n5249 ^ n5123 ;
  assign n5252 = n5251 ^ n5249 ;
  assign n5253 = n5250 & n5252 ;
  assign n5254 = n5253 ^ n5249 ;
  assign n5255 = n5210 & n5254 ;
  assign n5204 = n5203 ^ n5197 ;
  assign n5479 = n5255 ^ n5204 ;
  assign n5492 = n5491 ^ n5479 ;
  assign n5495 = n5494 ^ n5492 ;
  assign n5269 = n5240 ^ n5189 ;
  assign n5270 = n5269 ^ n5249 ;
  assign n5477 = n5270 ^ n5213 ;
  assign n5478 = n5123 & n5477 ;
  assign n5496 = n5495 ^ n5478 ;
  assign n5474 = n5245 ^ n5199 ;
  assign n5475 = n5474 ^ n5240 ;
  assign n5476 = n5266 & n5475 ;
  assign n5497 = n5496 ^ n5476 ;
  assign n5224 = ~n5128 & n5194 ;
  assign n5226 = n5225 ^ n5224 ;
  assign n5498 = n5226 ^ n5190 ;
  assign n5499 = n5190 ^ n5124 ;
  assign n5500 = n5499 ^ n5190 ;
  assign n5501 = n5498 & n5500 ;
  assign n5502 = n5501 ^ n5190 ;
  assign n5503 = ~n5123 & n5502 ;
  assign n5504 = ~n5497 & ~n5503 ;
  assign n5506 = n5505 ^ n5504 ;
  assign n5507 = n5506 ^ x74 ;
  assign n5508 = ~n5473 & n5507 ;
  assign n5509 = n5508 ^ n5507 ;
  assign n5510 = n5509 ^ n5473 ;
  assign n5511 = n5510 ^ n5507 ;
  assign n5642 = n5587 & ~n5615 ;
  assign n5637 = n5577 ^ n5557 ;
  assign n5638 = n5637 ^ n5588 ;
  assign n5639 = n5617 & ~n5638 ;
  assign n5633 = n5620 ^ n5581 ;
  assign n5634 = n5616 & n5633 ;
  assign n5630 = n5594 ^ n5577 ;
  assign n5631 = ~n5615 & ~n5630 ;
  assign n5618 = ~n5594 & n5617 ;
  assign n5623 = n5622 ^ n5618 ;
  assign n5624 = n5623 ^ n5593 ;
  assign n5595 = n5594 ^ n5592 ;
  assign n5625 = n5621 ^ n5595 ;
  assign n5626 = n5617 & ~n5625 ;
  assign n5627 = n5626 ^ n5614 ;
  assign n5628 = n5624 & n5627 ;
  assign n5514 = n5513 ^ n5512 ;
  assign n5607 = n5588 ^ n5513 ;
  assign n5608 = n5607 ^ n5588 ;
  assign n5611 = ~n5589 & n5608 ;
  assign n5612 = n5611 ^ n5588 ;
  assign n5613 = ~n5514 & ~n5612 ;
  assign n5629 = n5628 ^ n5613 ;
  assign n5632 = n5631 ^ n5629 ;
  assign n5635 = n5634 ^ n5632 ;
  assign n5561 = n5560 ^ n5559 ;
  assign n5636 = n5635 ^ n5561 ;
  assign n5640 = n5639 ^ n5636 ;
  assign n5565 = n5564 ^ n5563 ;
  assign n5596 = n5595 ^ n5565 ;
  assign n5597 = n5596 ^ n5561 ;
  assign n5600 = n5599 ^ n5597 ;
  assign n5601 = n5600 ^ n5561 ;
  assign n5602 = n5561 ^ n5512 ;
  assign n5603 = n5602 ^ n5561 ;
  assign n5604 = ~n5601 & ~n5603 ;
  assign n5605 = n5604 ^ n5561 ;
  assign n5606 = ~n5514 & n5605 ;
  assign n5641 = n5640 ^ n5606 ;
  assign n5643 = n5642 ^ n5641 ;
  assign n5644 = n5643 ^ n4017 ;
  assign n5645 = n5644 ^ x81 ;
  assign n5803 = n5802 ^ n5736 ;
  assign n5804 = n5803 ^ n5752 ;
  assign n5805 = n5759 ^ n5752 ;
  assign n5806 = n5805 ^ n5752 ;
  assign n5807 = ~n5804 & n5806 ;
  assign n5808 = n5807 ^ n5752 ;
  assign n5809 = n5760 & n5808 ;
  assign n5781 = ~n5764 & n5775 ;
  assign n5785 = n5781 ^ n5737 ;
  assign n5786 = ~n5733 & n5785 ;
  assign n5787 = n5786 ^ n5733 ;
  assign n5788 = n5787 ^ n5785 ;
  assign n5783 = n5781 ^ n5710 ;
  assign n5784 = ~n5762 & ~n5783 ;
  assign n5789 = n5788 ^ n5784 ;
  assign n5790 = n5789 ^ n5730 ;
  assign n5782 = n5771 & ~n5781 ;
  assign n5791 = n5790 ^ n5782 ;
  assign n5778 = n5736 ^ n5723 ;
  assign n5779 = n5778 ^ n5758 ;
  assign n5780 = n5779 ^ n5739 ;
  assign n5792 = n5791 ^ n5780 ;
  assign n5772 = n5771 ^ n5723 ;
  assign n5776 = n5775 ^ n5772 ;
  assign n5777 = n5776 ^ n5736 ;
  assign n5793 = n5792 ^ n5777 ;
  assign n5794 = n5793 ^ n5791 ;
  assign n5795 = ~n5759 & ~n5794 ;
  assign n5796 = n5795 ^ n5792 ;
  assign n5798 = n5791 ^ n5759 ;
  assign n5797 = n5791 ^ n5760 ;
  assign n5799 = n5798 ^ n5797 ;
  assign n5800 = ~n5796 & n5799 ;
  assign n5801 = n5800 ^ n5798 ;
  assign n5810 = n5809 ^ n5801 ;
  assign n5763 = n5762 ^ n5758 ;
  assign n5765 = n5764 ^ n5747 ;
  assign n5766 = n5764 ^ n5758 ;
  assign n5767 = n5766 ^ n5764 ;
  assign n5768 = ~n5765 & ~n5767 ;
  assign n5769 = n5768 ^ n5764 ;
  assign n5770 = ~n5763 & n5769 ;
  assign n5811 = n5810 ^ n5770 ;
  assign n5812 = n5755 ^ n5725 ;
  assign n5815 = n5760 & ~n5812 ;
  assign n5816 = n5815 ^ n5725 ;
  assign n5817 = ~n5759 & ~n5816 ;
  assign n5818 = n5811 & ~n5817 ;
  assign n5819 = n5818 ^ n3588 ;
  assign n5820 = n5819 ^ x120 ;
  assign n5821 = ~n5645 & ~n5820 ;
  assign n5826 = n5821 ^ n5820 ;
  assign n5892 = ~n5511 & ~n5826 ;
  assign n5822 = n5821 ^ n5645 ;
  assign n5823 = ~n5511 & ~n5822 ;
  assign n5922 = n5892 ^ n5823 ;
  assign n5894 = ~n5511 & n5821 ;
  assign n5921 = n5894 ^ n5511 ;
  assign n5923 = n5922 ^ n5921 ;
  assign n5883 = n5509 & ~n5822 ;
  assign n5958 = n5923 ^ n5883 ;
  assign n5877 = n5876 ^ x105 ;
  assign n5959 = n5883 ^ n5877 ;
  assign n5960 = n5959 ^ n5883 ;
  assign n5961 = ~n5958 & ~n5960 ;
  assign n5962 = n5961 ^ n5883 ;
  assign n5963 = n5427 & n5962 ;
  assign n5830 = n5826 ^ n5645 ;
  assign n5884 = n5509 & ~n5830 ;
  assign n5885 = n5884 ^ n5883 ;
  assign n5886 = n5884 ^ n5877 ;
  assign n5887 = n5886 ^ n5884 ;
  assign n5888 = n5885 & ~n5887 ;
  assign n5889 = n5888 ^ n5884 ;
  assign n5890 = ~n5427 & n5889 ;
  assign n5897 = n5508 & ~n5830 ;
  assign n5898 = n5897 ^ n5894 ;
  assign n5896 = n5508 & ~n5822 ;
  assign n5899 = n5898 ^ n5896 ;
  assign n5900 = n5899 ^ n5508 ;
  assign n5828 = n5473 & ~n5826 ;
  assign n5891 = n5828 ^ n5826 ;
  assign n5893 = n5892 ^ n5891 ;
  assign n5895 = n5894 ^ n5893 ;
  assign n5901 = n5900 ^ n5895 ;
  assign n6917 = n5901 ^ n5823 ;
  assign n8206 = n6917 ^ n5894 ;
  assign n6895 = n5899 ^ n5884 ;
  assign n6896 = n5427 & n6895 ;
  assign n6897 = n6896 ^ n5899 ;
  assign n8207 = n8206 ^ n6897 ;
  assign n8204 = n5922 ^ n5511 ;
  assign n8205 = n5427 & ~n8204 ;
  assign n8208 = n8207 ^ n8205 ;
  assign n8209 = n5877 & ~n8208 ;
  assign n5948 = n5877 ^ n5427 ;
  assign n8199 = n6897 ^ n5893 ;
  assign n5824 = n5510 & n5821 ;
  assign n8196 = n5883 ^ n5824 ;
  assign n5935 = n5894 ^ n5821 ;
  assign n5915 = n5901 ^ n5824 ;
  assign n5936 = n5935 ^ n5915 ;
  assign n8197 = n8196 ^ n5936 ;
  assign n8198 = ~n5877 & ~n8197 ;
  assign n8200 = n8199 ^ n8198 ;
  assign n8201 = n8200 ^ n6897 ;
  assign n8202 = n5948 & ~n8201 ;
  assign n8203 = n8202 ^ n8199 ;
  assign n8210 = n8209 ^ n8203 ;
  assign n5937 = n5427 & ~n5877 ;
  assign n5938 = n5937 ^ n5427 ;
  assign n5939 = n5938 ^ n5877 ;
  assign n6927 = ~n5923 & n5939 ;
  assign n8211 = n8210 ^ n6927 ;
  assign n5904 = n5828 ^ n5824 ;
  assign n5831 = n5510 & ~n5830 ;
  assign n5827 = n5510 & ~n5826 ;
  assign n5829 = n5828 ^ n5827 ;
  assign n5832 = n5831 ^ n5829 ;
  assign n5903 = n5832 ^ n5510 ;
  assign n5905 = n5904 ^ n5903 ;
  assign n5906 = n5905 ^ n5829 ;
  assign n8214 = ~n5427 & n5906 ;
  assign n8215 = n8214 ^ n5831 ;
  assign n8216 = ~n5877 & n8215 ;
  assign n8217 = n8216 ^ n5831 ;
  assign n8218 = n8211 & n8217 ;
  assign n8219 = n8218 ^ n8211 ;
  assign n8222 = n8219 ^ n5824 ;
  assign n8195 = n5922 ^ n5893 ;
  assign n8220 = n5937 & n8219 ;
  assign n8221 = ~n8195 & n8220 ;
  assign n8223 = n8222 ^ n8221 ;
  assign n5913 = n5824 ^ n5427 ;
  assign n5914 = n5913 ^ n5824 ;
  assign n8192 = n5828 & ~n5914 ;
  assign n8193 = n8192 ^ n5824 ;
  assign n8194 = n5948 & n8193 ;
  assign n8224 = n8223 ^ n8194 ;
  assign n5945 = ~n5936 & n5938 ;
  assign n8225 = n8224 ^ n5945 ;
  assign n8226 = ~n5890 & n8225 ;
  assign n8227 = ~n5963 & n8226 ;
  assign n8228 = n8227 ^ n5703 ;
  assign n8229 = n8228 ^ x93 ;
  assign n4216 = n4203 ^ n4202 ;
  assign n4217 = n4215 & n4216 ;
  assign n4209 = n4208 ^ n4169 ;
  assign n4212 = n4202 & n4209 ;
  assign n4213 = n4212 ^ n4169 ;
  assign n4214 = ~n4203 & n4213 ;
  assign n4218 = n4217 ^ n4214 ;
  assign n4249 = n4248 ^ n4225 ;
  assign n4238 = n4237 ^ n4221 ;
  assign n4240 = n4239 ^ n4203 ;
  assign n4242 = n4241 ^ n4240 ;
  assign n4243 = n4242 ^ n4203 ;
  assign n4244 = n4216 ^ n4203 ;
  assign n4245 = n4243 & ~n4244 ;
  assign n4246 = n4245 ^ n4203 ;
  assign n4247 = ~n4238 & n4246 ;
  assign n4250 = n4249 ^ n4247 ;
  assign n4260 = n4259 ^ n4250 ;
  assign n4293 = n4292 ^ n4260 ;
  assign n4282 = n4251 ^ n4232 ;
  assign n4283 = n4282 ^ n4270 ;
  assign n4284 = n4270 ^ n4203 ;
  assign n4285 = n4284 ^ n4270 ;
  assign n4286 = n4283 & n4285 ;
  assign n4287 = n4286 ^ n4270 ;
  assign n4288 = ~n4216 & n4287 ;
  assign n4294 = n4293 ^ n4288 ;
  assign n4272 = n4271 ^ n4270 ;
  assign n4275 = n4274 ^ n4272 ;
  assign n4276 = n4275 ^ n4268 ;
  assign n4277 = n4276 ^ n4260 ;
  assign n4261 = n4260 ^ n4237 ;
  assign n4264 = n4263 ^ n4261 ;
  assign n4278 = n4277 ^ n4264 ;
  assign n4279 = ~n4203 & ~n4278 ;
  assign n4280 = n4279 ^ n4277 ;
  assign n4281 = ~n4202 & n4280 ;
  assign n4295 = n4294 ^ n4281 ;
  assign n4296 = ~n4218 & ~n4295 ;
  assign n4300 = n4299 ^ n4296 ;
  assign n4301 = ~n4205 & n4300 ;
  assign n4302 = n4301 ^ n2919 ;
  assign n5968 = n4302 ^ x113 ;
  assign n5283 = n5282 ^ n2873 ;
  assign n5271 = n5270 ^ n5203 ;
  assign n5272 = ~n5268 & n5271 ;
  assign n5256 = n5213 ^ n5197 ;
  assign n5246 = n5245 ^ n5238 ;
  assign n5257 = n5256 ^ n5246 ;
  assign n5258 = n5246 ^ n5123 ;
  assign n5259 = n5258 ^ n5246 ;
  assign n5260 = n5257 & ~n5259 ;
  assign n5261 = n5260 ^ n5246 ;
  assign n5262 = n5210 & n5261 ;
  assign n5263 = n5262 ^ n5255 ;
  assign n5247 = n5246 ^ n5224 ;
  assign n5248 = n5237 & n5247 ;
  assign n5264 = n5263 ^ n5248 ;
  assign n5229 = n5228 ^ n5226 ;
  assign n5232 = n5229 ^ n5123 ;
  assign n5233 = n5232 ^ n5229 ;
  assign n5234 = n5227 & n5233 ;
  assign n5235 = n5234 ^ n5229 ;
  assign n5236 = ~n5210 & n5235 ;
  assign n5265 = n5264 ^ n5236 ;
  assign n5273 = n5272 ^ n5265 ;
  assign n5216 = n5215 ^ n5213 ;
  assign n5217 = n5216 ^ n5195 ;
  assign n5218 = n5217 ^ n5215 ;
  assign n5219 = n5215 ^ n5123 ;
  assign n5220 = n5219 ^ n5215 ;
  assign n5221 = n5218 & n5220 ;
  assign n5222 = n5221 ^ n5215 ;
  assign n5223 = ~n5210 & n5222 ;
  assign n5274 = n5273 ^ n5223 ;
  assign n5284 = n5283 ^ n5274 ;
  assign n5205 = n5204 ^ n5192 ;
  assign n5277 = ~n5124 & ~n5274 ;
  assign n5278 = n5205 & n5277 ;
  assign n5279 = n5278 ^ n5205 ;
  assign n5200 = n5199 ^ n5190 ;
  assign n5201 = ~n5124 & n5200 ;
  assign n5202 = n5201 ^ n5199 ;
  assign n5206 = n5205 ^ n5202 ;
  assign n5280 = n5279 ^ n5206 ;
  assign n5281 = n5123 & n5280 ;
  assign n5285 = n5284 ^ n5281 ;
  assign n6071 = n5285 ^ x90 ;
  assign n3837 = ~n3800 & n3836 ;
  assign n6066 = n6065 ^ n3837 ;
  assign n6056 = n6055 ^ n6032 ;
  assign n6057 = n6055 ^ n2257 ;
  assign n6058 = n6057 ^ n6055 ;
  assign n6059 = ~n6056 & ~n6058 ;
  assign n6060 = n6059 ^ n6055 ;
  assign n6061 = n3803 & ~n6060 ;
  assign n6067 = n6066 ^ n6061 ;
  assign n6068 = n6067 ^ n3553 ;
  assign n6046 = n3813 ^ n3809 ;
  assign n6044 = n2827 & n3808 ;
  assign n6042 = n6041 ^ n3793 ;
  assign n6043 = n6042 ^ n3829 ;
  assign n6045 = n6044 ^ n6043 ;
  assign n6047 = n6046 ^ n6045 ;
  assign n6039 = ~n3801 & n3815 ;
  assign n6048 = n6047 ^ n6039 ;
  assign n6049 = n2826 ^ n2257 ;
  assign n6050 = ~n6048 & ~n6049 ;
  assign n6051 = n6050 ^ n2257 ;
  assign n6033 = n6032 ^ n3808 ;
  assign n6034 = n3808 ^ n2826 ;
  assign n6035 = n6034 ^ n3808 ;
  assign n6036 = ~n6033 & n6035 ;
  assign n6037 = n6036 ^ n3808 ;
  assign n6038 = n2257 & n6037 ;
  assign n6052 = n6051 ^ n6038 ;
  assign n6024 = n3814 ^ n3812 ;
  assign n6025 = n6024 ^ n3802 ;
  assign n6026 = n3804 ^ n3800 ;
  assign n6029 = ~n6024 & n6026 ;
  assign n6030 = n6029 ^ n3800 ;
  assign n6031 = ~n6025 & ~n6030 ;
  assign n6053 = n6052 ^ n6031 ;
  assign n6054 = ~n6023 & n6053 ;
  assign n6069 = n6068 ^ n6054 ;
  assign n6070 = n6069 ^ x73 ;
  assign n6072 = n6071 ^ n6070 ;
  assign n5066 = ~n4898 & n5058 ;
  assign n5067 = n5066 ^ n5049 ;
  assign n5070 = n5067 ^ n5060 ;
  assign n5071 = n5070 ^ n5067 ;
  assign n5072 = n4898 & n5071 ;
  assign n5073 = n5072 ^ n5067 ;
  assign n5074 = ~n4929 & n5073 ;
  assign n5075 = n5074 ^ n5067 ;
  assign n5983 = n5469 ^ n5075 ;
  assign n5972 = n5021 ^ n4990 ;
  assign n5973 = n5972 ^ n5039 ;
  assign n5970 = n5430 ^ n5055 ;
  assign n5971 = n5970 ^ n5063 ;
  assign n5974 = n5973 ^ n5971 ;
  assign n5975 = ~n4929 & ~n5974 ;
  assign n5976 = n5975 ^ n5971 ;
  assign n5984 = n5983 ^ n5976 ;
  assign n5978 = n5054 ^ n5050 ;
  assign n5979 = n5978 ^ n5443 ;
  assign n5980 = n4929 & n5979 ;
  assign n5969 = n5054 ^ n5042 ;
  assign n5977 = n5976 ^ n5969 ;
  assign n5981 = n5980 ^ n5977 ;
  assign n5982 = ~n4898 & ~n5981 ;
  assign n5985 = n5984 ^ n5982 ;
  assign n5986 = ~n5119 & n5985 ;
  assign n5987 = n5986 ^ n3903 ;
  assign n5988 = n5987 ^ x99 ;
  assign n6083 = n6071 ^ n5988 ;
  assign n5989 = n5775 ^ n5733 ;
  assign n5993 = n5803 ^ n5772 ;
  assign n5994 = n5993 ^ n5761 ;
  assign n5995 = n5750 ^ n5747 ;
  assign n5996 = n5995 ^ n5993 ;
  assign n5997 = ~n5994 & ~n5996 ;
  assign n5998 = n5997 ^ n5761 ;
  assign n5992 = n5817 ^ n5764 ;
  assign n6004 = n5998 ^ n5992 ;
  assign n6000 = n5817 ^ n5751 ;
  assign n6001 = n6000 ^ n5757 ;
  assign n6002 = n5725 & n6001 ;
  assign n6003 = n5992 & n6002 ;
  assign n6005 = n6004 ^ n6003 ;
  assign n5991 = n5756 & ~n5760 ;
  assign n6006 = n6005 ^ n5991 ;
  assign n6007 = ~n5759 & ~n6006 ;
  assign n6009 = n5737 ^ n5710 ;
  assign n6008 = n5993 ^ n5747 ;
  assign n6010 = n6009 ^ n6008 ;
  assign n6011 = ~n5760 & ~n6010 ;
  assign n6012 = n6011 ^ n6008 ;
  assign n6013 = n6007 & ~n6012 ;
  assign n6014 = n6013 ^ n6006 ;
  assign n6015 = ~n5990 & ~n6014 ;
  assign n6016 = ~n5989 & n6015 ;
  assign n6017 = n6016 ^ n6014 ;
  assign n6019 = n5730 & n5760 ;
  assign n6020 = ~n6017 & n6019 ;
  assign n6018 = n6017 ^ n3868 ;
  assign n6021 = n6020 ^ n6018 ;
  assign n6022 = n6021 ^ x72 ;
  assign n6092 = n6083 ^ n6022 ;
  assign n6093 = n6070 & n6092 ;
  assign n6094 = n6093 ^ n6022 ;
  assign n6095 = ~n6072 & ~n6094 ;
  assign n6096 = n6095 ^ n6094 ;
  assign n6079 = n6022 ^ n5988 ;
  assign n6073 = n6022 & ~n6072 ;
  assign n6074 = n6073 ^ n6071 ;
  assign n6088 = n6074 ^ n6022 ;
  assign n6085 = n6022 & n6071 ;
  assign n6089 = n6088 ^ n6085 ;
  assign n6090 = n6079 & n6089 ;
  assign n6091 = ~n6083 & n6090 ;
  assign n6097 = n6096 ^ n6091 ;
  assign n6086 = n6085 ^ n6071 ;
  assign n6076 = n6070 ^ n6022 ;
  assign n6080 = n6071 & ~n6076 ;
  assign n6087 = n6086 ^ n6080 ;
  assign n6098 = n6097 ^ n6087 ;
  assign n6099 = n6098 ^ n6022 ;
  assign n6109 = n6099 ^ n5988 ;
  assign n6110 = n6109 ^ n6091 ;
  assign n6103 = n6070 ^ n5988 ;
  assign n6106 = n6103 ^ n6090 ;
  assign n6081 = n6080 ^ n6070 ;
  assign n6082 = ~n6079 & ~n6081 ;
  assign n6105 = n6095 ^ n6082 ;
  assign n6107 = n6106 ^ n6105 ;
  assign n6077 = n6076 ^ n6071 ;
  assign n6108 = n6107 ^ n6077 ;
  assign n6111 = n6110 ^ n6108 ;
  assign n6131 = n6130 ^ n5584 ;
  assign n6132 = n5512 & ~n6131 ;
  assign n6133 = n6132 ^ n5584 ;
  assign n6137 = n6133 ^ n5618 ;
  assign n6143 = n6142 ^ n6137 ;
  assign n6144 = n6143 ^ n3622 ;
  assign n6120 = n5637 ^ n5555 ;
  assign n6121 = n6120 ^ n5621 ;
  assign n6125 = n6124 ^ n6121 ;
  assign n6134 = n6133 ^ n6125 ;
  assign n6115 = n5552 ^ n5551 ;
  assign n6116 = n5567 ^ n5551 ;
  assign n6117 = ~n6115 & n6116 ;
  assign n6118 = n6117 ^ n5551 ;
  assign n6119 = n5512 & n6118 ;
  assign n6135 = n6134 ^ n6119 ;
  assign n6136 = n5513 & n6135 ;
  assign n6145 = n6144 ^ n6136 ;
  assign n6146 = n6145 ^ x66 ;
  assign n7138 = n6111 & ~n6146 ;
  assign n7139 = n7138 ^ n6108 ;
  assign n7131 = n6071 ^ n6022 ;
  assign n7132 = n5988 & n6070 ;
  assign n7133 = n7132 ^ n6022 ;
  assign n7134 = n7131 & ~n7133 ;
  assign n7135 = n7134 ^ n6022 ;
  assign n7136 = n6146 & n7135 ;
  assign n7137 = n7136 ^ n6106 ;
  assign n7141 = n7139 ^ n7137 ;
  assign n7142 = ~n5968 & n7141 ;
  assign n7143 = n7142 ^ n7139 ;
  assign n8189 = n7143 ^ n4834 ;
  assign n8190 = n8189 ^ x126 ;
  assign n8277 = n8229 ^ n8190 ;
  assign n8278 = n8185 & n8277 ;
  assign n8279 = n8278 ^ n8185 ;
  assign n6188 = n6187 ^ n5751 ;
  assign n6189 = n6188 ^ n5786 ;
  assign n6190 = n5761 & ~n6189 ;
  assign n6178 = n5764 ^ n5732 ;
  assign n6179 = n5745 ^ n5741 ;
  assign n6180 = n6179 ^ n5762 ;
  assign n6182 = n5764 & n6180 ;
  assign n6183 = n6182 ^ n5762 ;
  assign n6184 = ~n6178 & ~n6183 ;
  assign n6185 = n6184 ^ n1175 ;
  assign n6175 = n6001 ^ n5734 ;
  assign n6168 = n6001 ^ n5749 ;
  assign n6169 = n6168 ^ n6001 ;
  assign n6170 = n6001 ^ n5755 ;
  assign n6171 = n6170 ^ n6001 ;
  assign n6172 = n6169 & ~n6171 ;
  assign n6173 = n6172 ^ n6001 ;
  assign n6174 = n5760 & n6173 ;
  assign n6176 = n6175 ^ n6174 ;
  assign n6177 = ~n5759 & n6176 ;
  assign n6186 = n6185 ^ n6177 ;
  assign n6191 = n6190 ^ n6186 ;
  assign n6167 = n5760 & ~n5775 ;
  assign n6192 = n6191 ^ n6167 ;
  assign n6193 = n6192 ^ x67 ;
  assign n6216 = n5477 ^ n5215 ;
  assign n6217 = n6216 ^ n5205 ;
  assign n6218 = ~n5123 & n6217 ;
  assign n6207 = n5480 ^ n5226 ;
  assign n6213 = n6207 ^ n5126 ;
  assign n6219 = n6218 ^ n6213 ;
  assign n6220 = n5210 & ~n6219 ;
  assign n6210 = n5195 ^ n5191 ;
  assign n6211 = n6210 ^ n5215 ;
  assign n6206 = n5211 ^ n5197 ;
  assign n6208 = n6207 ^ n6206 ;
  assign n6209 = n5267 & n6208 ;
  assign n6212 = n6211 ^ n6209 ;
  assign n6214 = n6213 ^ n6212 ;
  assign n6201 = n5191 ^ n5124 ;
  assign n6202 = n6201 ^ n5191 ;
  assign n6203 = n5484 & n6202 ;
  assign n6204 = n6203 ^ n5191 ;
  assign n6205 = ~n5123 & n6204 ;
  assign n6215 = n6214 ^ n6205 ;
  assign n6221 = n6220 ^ n6215 ;
  assign n6222 = n6221 ^ n5282 ;
  assign n6223 = ~n5503 & n6222 ;
  assign n6224 = n6223 ^ n1948 ;
  assign n6225 = n6224 ^ x93 ;
  assign n6249 = n4202 & n4234 ;
  assign n6233 = n4265 ^ n4226 ;
  assign n6234 = n6233 ^ n4265 ;
  assign n6235 = n6234 ^ n4238 ;
  assign n6236 = n6235 ^ n4270 ;
  assign n6237 = ~n4203 & ~n6236 ;
  assign n6238 = n6237 ^ n6233 ;
  assign n6242 = n4225 ^ n4204 ;
  assign n6243 = n6242 ^ n4221 ;
  assign n6244 = n4297 & n6243 ;
  assign n6239 = n5419 ^ n4216 ;
  assign n6240 = n6239 ^ n4288 ;
  assign n6241 = n6240 ^ n5419 ;
  assign n6245 = n6244 ^ n6241 ;
  assign n6246 = n6245 ^ n4288 ;
  assign n6247 = n6238 & n6246 ;
  assign n6248 = n6247 ^ n6240 ;
  assign n6250 = n6249 ^ n6248 ;
  assign n6226 = n4256 ^ n4203 ;
  assign n6227 = n6226 ^ n4256 ;
  assign n6230 = n4257 & ~n6227 ;
  assign n6231 = n6230 ^ n4256 ;
  assign n6232 = ~n4216 & n6231 ;
  assign n6251 = n6250 ^ n6232 ;
  assign n6252 = ~n4291 & ~n6251 ;
  assign n6253 = ~n5417 & n6252 ;
  assign n6254 = n6253 ^ n2171 ;
  assign n6255 = n6254 ^ x91 ;
  assign n6256 = n6225 & n6255 ;
  assign n6267 = n5594 ^ n5512 ;
  assign n6269 = n5594 ^ n5580 ;
  assign n6268 = n5622 ^ n5594 ;
  assign n6270 = n6269 ^ n6268 ;
  assign n6271 = n6269 ^ n5513 ;
  assign n6272 = n6271 ^ n6269 ;
  assign n6273 = n6270 & ~n6272 ;
  assign n6274 = n6273 ^ n6269 ;
  assign n6275 = n6267 & n6274 ;
  assign n6276 = n6275 ^ n5512 ;
  assign n6266 = n5582 & n5617 ;
  assign n6277 = n6276 ^ n6266 ;
  assign n6259 = n6120 ^ n5581 ;
  assign n6260 = n6259 ^ n5576 ;
  assign n6261 = n5576 ^ n5513 ;
  assign n6262 = n6261 ^ n5576 ;
  assign n6263 = n6260 & ~n6262 ;
  assign n6264 = n6263 ^ n5576 ;
  assign n6265 = n5514 & n6264 ;
  assign n6278 = n6277 ^ n6265 ;
  assign n6279 = ~n5642 & n6278 ;
  assign n6280 = ~n6258 & n6279 ;
  assign n6281 = n5596 ^ n5558 ;
  assign n6282 = n5512 & ~n6281 ;
  assign n6283 = n6282 ^ n5558 ;
  assign n6284 = n6283 ^ n5514 ;
  assign n6285 = n6284 ^ n6283 ;
  assign n6286 = n5512 & ~n6128 ;
  assign n6287 = n6286 ^ n6283 ;
  assign n6288 = n6285 & n6287 ;
  assign n6289 = n6288 ^ n6283 ;
  assign n6290 = n6280 & n6289 ;
  assign n6291 = n6290 ^ n6280 ;
  assign n6292 = ~n5613 & n6291 ;
  assign n6293 = ~n6142 & n6292 ;
  assign n6294 = n6293 ^ n1738 ;
  assign n6295 = n6294 ^ x110 ;
  assign n5065 = n4930 & n5052 ;
  assign n5105 = n4932 & n5050 ;
  assign n5102 = n5101 ^ n5099 ;
  assign n5103 = n4931 & ~n5102 ;
  assign n5097 = n4930 & n5045 ;
  assign n5083 = n5035 ^ n4929 ;
  assign n5084 = n5061 ^ n5035 ;
  assign n5085 = n5084 ^ n4898 ;
  assign n5086 = n5085 ^ n5084 ;
  assign n5090 = n5089 ^ n5088 ;
  assign n5091 = n5090 ^ n5035 ;
  assign n5092 = n5091 ^ n5084 ;
  assign n5093 = n5086 & n5092 ;
  assign n5094 = n5093 ^ n5084 ;
  assign n5095 = ~n5083 & ~n5094 ;
  assign n5096 = n5095 ^ n4929 ;
  assign n5098 = n5097 ^ n5096 ;
  assign n5104 = n5103 ^ n5098 ;
  assign n5106 = n5105 ^ n5104 ;
  assign n5078 = n5041 ^ n4929 ;
  assign n5079 = n5078 ^ n5041 ;
  assign n5080 = ~n5055 & ~n5079 ;
  assign n5081 = n5080 ^ n5041 ;
  assign n5082 = ~n4898 & n5081 ;
  assign n5107 = n5106 ^ n5082 ;
  assign n5108 = ~n5075 & n5107 ;
  assign n5109 = ~n5065 & n5108 ;
  assign n5110 = ~n5064 & n5109 ;
  assign n5120 = n5110 & ~n5119 ;
  assign n5121 = n5120 ^ n1517 ;
  assign n6296 = n5121 ^ x100 ;
  assign n6297 = ~n6295 & n6296 ;
  assign n6302 = n6297 ^ n6295 ;
  assign n6356 = n6256 & ~n6302 ;
  assign n4567 = n4360 & ~n4566 ;
  assign n4568 = n4567 ^ n4554 ;
  assign n4571 = n4568 ^ n4340 ;
  assign n4541 = n4540 ^ n4491 ;
  assign n4533 = n4532 ^ n4492 ;
  assign n4534 = n4419 & n4533 ;
  assign n4542 = n4541 ^ n4534 ;
  assign n4543 = n4360 & n4542 ;
  assign n4544 = n4543 ^ n4540 ;
  assign n4569 = n4568 ^ n4544 ;
  assign n4570 = n4340 & ~n4569 ;
  assign n4572 = n4571 ^ n4570 ;
  assign n4573 = n4572 ^ n775 ;
  assign n6194 = n4573 ^ x117 ;
  assign n7189 = n6356 ^ n6194 ;
  assign n7190 = n7189 ^ n6356 ;
  assign n6306 = n6256 ^ n6255 ;
  assign n6307 = n6306 ^ n6225 ;
  assign n6308 = ~n6302 & ~n6307 ;
  assign n7191 = n6356 ^ n6308 ;
  assign n7194 = n7190 & n7191 ;
  assign n7195 = n7194 ^ n6356 ;
  assign n7196 = ~n6193 & n7195 ;
  assign n6331 = n6302 ^ n6296 ;
  assign n6365 = n6256 & n6331 ;
  assign n6355 = ~n6307 & n6331 ;
  assign n6380 = n6365 ^ n6355 ;
  assign n6257 = n6256 ^ n6225 ;
  assign n6300 = n6257 & n6297 ;
  assign n6381 = n6380 ^ n6300 ;
  assign n6351 = n6256 & n6297 ;
  assign n6332 = n6306 & n6331 ;
  assign n6330 = ~n6302 & n6306 ;
  assign n6333 = n6332 ^ n6330 ;
  assign n6321 = n6297 & n6306 ;
  assign n6329 = n6321 ^ n6306 ;
  assign n6334 = n6333 ^ n6329 ;
  assign n6379 = n6351 ^ n6334 ;
  assign n6382 = n6381 ^ n6379 ;
  assign n6383 = ~n6193 & n6382 ;
  assign n6384 = n6383 ^ n6300 ;
  assign n6311 = n6297 & ~n6307 ;
  assign n6385 = n6384 ^ n6311 ;
  assign n6386 = n6385 ^ n6384 ;
  assign n6387 = n6384 ^ n6193 ;
  assign n6388 = n6387 ^ n6384 ;
  assign n6389 = n6386 & n6388 ;
  assign n6390 = n6389 ^ n6384 ;
  assign n6391 = n6194 & n6390 ;
  assign n6392 = n6391 ^ n6384 ;
  assign n8178 = n7196 ^ n6392 ;
  assign n6320 = n6194 ^ n6193 ;
  assign n7181 = n6379 ^ n6321 ;
  assign n6298 = n6297 ^ n6296 ;
  assign n6350 = n6298 & ~n6307 ;
  assign n7180 = n6379 ^ n6350 ;
  assign n7182 = n7181 ^ n7180 ;
  assign n7183 = n7181 ^ n6194 ;
  assign n7184 = n7183 ^ n7181 ;
  assign n7185 = n7182 & ~n7184 ;
  assign n7186 = n7185 ^ n7181 ;
  assign n7187 = ~n6320 & n7186 ;
  assign n7188 = n7187 ^ n6379 ;
  assign n8179 = n8178 ^ n7188 ;
  assign n6195 = n6193 & n6194 ;
  assign n6196 = n6195 ^ n6194 ;
  assign n6197 = n6196 ^ n6193 ;
  assign n6198 = n6197 ^ n6194 ;
  assign n7702 = n6198 & n6380 ;
  assign n6374 = n6195 & n6330 ;
  assign n7703 = n7702 ^ n6374 ;
  assign n8180 = n8179 ^ n7703 ;
  assign n6303 = n6257 & ~n6302 ;
  assign n6304 = n6303 ^ n6257 ;
  assign n6299 = n6257 & n6298 ;
  assign n6301 = n6300 ^ n6299 ;
  assign n6305 = n6304 ^ n6301 ;
  assign n6309 = n6308 ^ n6305 ;
  assign n6310 = n6198 & n6309 ;
  assign n8181 = n8180 ^ n6310 ;
  assign n8182 = n8181 ^ n5674 ;
  assign n7730 = n6195 & n6301 ;
  assign n6314 = n6198 ^ n6196 ;
  assign n8161 = n6309 ^ n6299 ;
  assign n8162 = n8161 ^ n6334 ;
  assign n8160 = n6296 ^ n6295 ;
  assign n8163 = n8162 ^ n8160 ;
  assign n8164 = ~n6193 & ~n8163 ;
  assign n8165 = n8164 ^ n6356 ;
  assign n8166 = n8165 ^ n6308 ;
  assign n7721 = n6332 ^ n6299 ;
  assign n7722 = ~n6193 & n7721 ;
  assign n7723 = n7722 ^ n6332 ;
  assign n8167 = n8166 ^ n7723 ;
  assign n8168 = n8167 ^ n6380 ;
  assign n8169 = n8168 ^ n6308 ;
  assign n8170 = n8169 ^ n8167 ;
  assign n8173 = n6193 & n8170 ;
  assign n8174 = n8173 ^ n8167 ;
  assign n8175 = ~n6314 & n8174 ;
  assign n8176 = n8175 ^ n8165 ;
  assign n8177 = ~n7730 & ~n8176 ;
  assign n8183 = n8182 ^ n8177 ;
  assign n8184 = n8183 ^ x108 ;
  assign n8186 = n8184 & ~n8185 ;
  assign n8230 = ~n8190 & n8229 ;
  assign n8236 = n8230 ^ n8190 ;
  assign n8256 = n8186 & ~n8236 ;
  assign n8245 = n8185 ^ n8184 ;
  assign n8246 = n8229 ^ n8184 ;
  assign n8247 = ~n8190 & n8246 ;
  assign n8248 = n8247 ^ n8184 ;
  assign n8249 = ~n8245 & n8248 ;
  assign n8250 = n8249 ^ n8185 ;
  assign n8187 = n8186 ^ n8184 ;
  assign n8237 = n8187 & ~n8236 ;
  assign n8188 = n8187 ^ n8185 ;
  assign n8244 = n8237 ^ n8188 ;
  assign n8251 = n8250 ^ n8244 ;
  assign n8239 = n8186 ^ n8185 ;
  assign n8231 = n8230 ^ n8229 ;
  assign n8242 = n8231 ^ n8190 ;
  assign n8243 = ~n8239 & n8242 ;
  assign n8252 = n8251 ^ n8243 ;
  assign n8240 = n8231 & ~n8239 ;
  assign n8241 = n8240 ^ n8239 ;
  assign n8253 = n8252 ^ n8241 ;
  assign n8262 = n8256 ^ n8253 ;
  assign n8263 = n8262 ^ n8240 ;
  assign n8233 = n8187 & n8230 ;
  assign n8264 = n8263 ^ n8233 ;
  assign n8258 = n8186 & n8230 ;
  assign n8259 = n8258 ^ n8186 ;
  assign n8255 = n8186 & n8242 ;
  assign n8257 = n8256 ^ n8255 ;
  assign n8260 = n8259 ^ n8257 ;
  assign n8261 = n8260 ^ n8256 ;
  assign n8265 = n8264 ^ n8261 ;
  assign n8254 = n8253 ^ n8231 ;
  assign n8266 = n8265 ^ n8254 ;
  assign n8232 = n8188 & n8231 ;
  assign n8234 = n8233 ^ n8232 ;
  assign n8267 = n8266 ^ n8234 ;
  assign n8238 = n8237 ^ n8232 ;
  assign n8268 = n8267 ^ n8238 ;
  assign n8280 = n8279 ^ n8268 ;
  assign n7212 = n6069 ^ x65 ;
  assign n7213 = n5819 ^ x104 ;
  assign n7214 = ~n7212 & n7213 ;
  assign n7215 = n7214 ^ n7212 ;
  assign n7216 = n7215 ^ n7213 ;
  assign n7239 = n4783 ^ n4777 ;
  assign n4875 = n4874 ^ n4776 ;
  assign n7240 = n7239 ^ n4875 ;
  assign n7241 = ~n5836 & n7240 ;
  assign n6649 = n5865 ^ n4803 ;
  assign n6650 = n4835 ^ n4803 ;
  assign n6651 = n6650 ^ n4803 ;
  assign n6652 = n6649 & n6651 ;
  assign n6653 = n6652 ^ n4803 ;
  assign n6654 = n4607 & n6653 ;
  assign n6629 = n4868 ^ n4782 ;
  assign n6630 = n5838 & n6629 ;
  assign n7232 = n6654 ^ n6630 ;
  assign n4846 = n4845 ^ n4786 ;
  assign n4847 = n4846 ^ n4795 ;
  assign n4850 = n4835 & ~n4847 ;
  assign n4851 = n4850 ^ n4795 ;
  assign n4852 = n4607 & n4851 ;
  assign n7233 = n7232 ^ n4852 ;
  assign n4804 = n4803 ^ n4788 ;
  assign n4838 = n4804 & n4835 ;
  assign n4839 = n4838 ^ n4788 ;
  assign n4840 = ~n4607 & n4839 ;
  assign n7234 = n7233 ^ n4840 ;
  assign n7235 = n7234 ^ n3682 ;
  assign n7225 = n4846 ^ n4835 ;
  assign n7226 = n7225 ^ n4846 ;
  assign n7227 = n4846 ^ n4788 ;
  assign n7228 = n7227 ^ n4846 ;
  assign n7229 = n7226 & n7228 ;
  assign n7230 = n7229 ^ n4846 ;
  assign n7231 = n4853 & ~n7230 ;
  assign n7236 = n7235 ^ n7231 ;
  assign n7218 = n4802 ^ n4774 ;
  assign n7219 = n7218 ^ n4841 ;
  assign n7220 = n4841 ^ n4835 ;
  assign n7221 = n7220 ^ n4841 ;
  assign n7222 = n7219 & n7221 ;
  assign n7223 = n7222 ^ n4841 ;
  assign n7224 = n4607 & n7223 ;
  assign n7237 = n7236 ^ n7224 ;
  assign n7217 = n4799 & n5835 ;
  assign n7238 = n7237 ^ n7217 ;
  assign n7242 = n7241 ^ n7238 ;
  assign n7243 = n7242 ^ x97 ;
  assign n7244 = n5426 ^ x107 ;
  assign n7245 = n6145 ^ x80 ;
  assign n7246 = ~n7244 & n7245 ;
  assign n7247 = n6449 ^ n6438 ;
  assign n7248 = n4360 & n7247 ;
  assign n7249 = n7248 ^ n6449 ;
  assign n7257 = n7249 ^ n3601 ;
  assign n7250 = n7249 ^ n6455 ;
  assign n7251 = n7250 ^ n4563 ;
  assign n7252 = n7251 ^ n6457 ;
  assign n7253 = n7252 ^ n7249 ;
  assign n7254 = n4360 & n7253 ;
  assign n7255 = n7254 ^ n7250 ;
  assign n7256 = ~n4340 & n7255 ;
  assign n7258 = n7257 ^ n7256 ;
  assign n7259 = n7258 ^ x98 ;
  assign n7260 = n7246 & n7259 ;
  assign n7261 = n7260 ^ n7246 ;
  assign n7262 = ~n7243 & n7261 ;
  assign n7263 = n7262 ^ n7261 ;
  assign n7264 = n7216 & n7263 ;
  assign n7270 = ~n7244 & ~n7259 ;
  assign n7269 = n7259 ^ n7244 ;
  assign n7271 = n7270 ^ n7269 ;
  assign n7276 = n7271 ^ n7244 ;
  assign n7324 = n7243 & ~n7276 ;
  assign n7335 = n7324 ^ n7276 ;
  assign n7336 = n7245 & ~n7335 ;
  assign n7337 = n7336 ^ n7335 ;
  assign n7277 = n7243 & ~n7245 ;
  assign n7293 = n7259 & n7277 ;
  assign n7294 = n7293 ^ n7277 ;
  assign n7278 = ~n7276 & n7277 ;
  assign n7295 = n7294 ^ n7278 ;
  assign n7292 = n7270 ^ n7261 ;
  assign n7296 = n7295 ^ n7292 ;
  assign n7265 = ~n7243 & n7259 ;
  assign n7279 = n7271 ^ n7265 ;
  assign n7272 = n7243 & ~n7271 ;
  assign n7280 = n7279 ^ n7272 ;
  assign n7266 = n7246 & n7265 ;
  assign n7281 = n7280 ^ n7266 ;
  assign n7297 = n7296 ^ n7281 ;
  assign n7291 = n7277 ^ n7245 ;
  assign n7298 = n7297 ^ n7291 ;
  assign n7290 = n7280 ^ n7265 ;
  assign n7299 = n7298 ^ n7290 ;
  assign n7338 = n7337 ^ n7299 ;
  assign n8031 = n7214 & n7338 ;
  assign n7268 = n7214 ^ n7213 ;
  assign n7273 = n7245 & n7272 ;
  assign n7274 = n7268 & n7273 ;
  assign n8032 = n8031 ^ n7274 ;
  assign n7323 = n7213 ^ n7212 ;
  assign n7325 = n7324 ^ n7278 ;
  assign n7492 = n7325 ^ n7299 ;
  assign n8066 = n7492 ^ n7325 ;
  assign n8067 = n7325 ^ n7213 ;
  assign n8068 = n8067 ^ n7325 ;
  assign n8069 = ~n8066 & n8068 ;
  assign n8070 = n8069 ^ n7325 ;
  assign n8071 = ~n7323 & n8070 ;
  assign n8063 = n7214 & n7245 ;
  assign n8064 = n8063 ^ n7215 ;
  assign n8065 = ~n7335 & ~n8064 ;
  assign n8072 = n8071 ^ n8065 ;
  assign n7306 = n7293 ^ n7272 ;
  assign n7307 = n7306 ^ n7273 ;
  assign n8038 = n7307 ^ n7278 ;
  assign n8037 = n7281 ^ n7262 ;
  assign n8039 = n8038 ^ n8037 ;
  assign n8040 = n8039 ^ n7307 ;
  assign n8041 = ~n7212 & ~n8040 ;
  assign n8042 = n8041 ^ n8038 ;
  assign n8052 = n8042 ^ n7266 ;
  assign n7478 = n7296 ^ n7295 ;
  assign n7479 = n7295 ^ n7212 ;
  assign n7480 = n7479 ^ n7295 ;
  assign n7481 = n7478 & n7480 ;
  assign n7482 = n7481 ^ n7295 ;
  assign n7483 = n7213 & n7482 ;
  assign n8053 = n8052 ^ n7483 ;
  assign n7328 = n7266 ^ n7260 ;
  assign n7329 = n7328 ^ n7296 ;
  assign n8044 = n7329 ^ n7263 ;
  assign n8045 = n8044 ^ n8042 ;
  assign n8049 = n8045 ^ n7266 ;
  assign n7339 = n7338 ^ n7290 ;
  assign n7326 = n7307 ^ n7293 ;
  assign n8033 = n7339 ^ n7326 ;
  assign n8043 = n8033 ^ n7335 ;
  assign n8046 = n8045 ^ n8043 ;
  assign n8047 = n8046 ^ n8042 ;
  assign n8048 = n7212 & n8047 ;
  assign n8050 = n8049 ^ n8048 ;
  assign n8051 = n7323 & n8050 ;
  assign n8054 = n8053 ^ n8051 ;
  assign n8073 = n8072 ^ n8054 ;
  assign n7507 = ~n7215 & n7273 ;
  assign n7506 = n7216 & n7295 ;
  assign n7508 = n7507 ^ n7506 ;
  assign n8074 = n8073 ^ n7508 ;
  assign n8034 = n8033 ^ n7213 ;
  assign n8035 = n8034 ^ n8033 ;
  assign n8036 = n7328 ^ n7281 ;
  assign n8055 = ~n8036 & ~n8054 ;
  assign n8056 = n8055 ^ n8033 ;
  assign n8057 = ~n8035 & ~n8056 ;
  assign n8058 = n8057 ^ n8033 ;
  assign n8059 = n7323 & ~n8058 ;
  assign n8075 = n8074 ^ n8059 ;
  assign n8076 = ~n8032 & ~n8075 ;
  assign n8077 = ~n7264 & n8076 ;
  assign n8078 = n8077 ^ n4451 ;
  assign n8271 = n8078 ^ x76 ;
  assign n6717 = n6398 ^ n3236 ;
  assign n3786 = n2827 & n3785 ;
  assign n6706 = n3811 ^ n3805 ;
  assign n6707 = ~n3801 & n6706 ;
  assign n6697 = n3822 ^ n3816 ;
  assign n6698 = n6697 ^ n6408 ;
  assign n6699 = n6698 ^ n6697 ;
  assign n6700 = n6697 ^ n2826 ;
  assign n6701 = n6700 ^ n6697 ;
  assign n6702 = ~n6699 & ~n6701 ;
  assign n6703 = n6702 ^ n6697 ;
  assign n6704 = ~n2257 & n6703 ;
  assign n6705 = n6704 ^ n2826 ;
  assign n6708 = n6707 ^ n6705 ;
  assign n6695 = n3792 ^ n3789 ;
  assign n6696 = ~n3803 & n6695 ;
  assign n6709 = n6708 ^ n6696 ;
  assign n6690 = n3797 ^ n3791 ;
  assign n6691 = n6690 ^ n6399 ;
  assign n6692 = ~n2826 & ~n6691 ;
  assign n6693 = n6692 ^ n3784 ;
  assign n6694 = n2257 & n6693 ;
  assign n6710 = n6709 ^ n6694 ;
  assign n6711 = n6710 ^ n3829 ;
  assign n6712 = n6711 ^ n6064 ;
  assign n6683 = n3829 ^ n2826 ;
  assign n6684 = n6683 ^ n3829 ;
  assign n6685 = n3829 ^ n3809 ;
  assign n6686 = n6685 ^ n3829 ;
  assign n6687 = ~n6684 & n6686 ;
  assign n6688 = n6687 ^ n3829 ;
  assign n6689 = ~n2257 & n6688 ;
  assign n6713 = n6712 ^ n6689 ;
  assign n6714 = n6713 ^ n6426 ;
  assign n6715 = n6714 ^ n6061 ;
  assign n6716 = ~n3786 & ~n6715 ;
  assign n6718 = n6717 ^ n6716 ;
  assign n7050 = n6718 ^ x83 ;
  assign n7051 = n6467 ^ x101 ;
  assign n7061 = n7050 & ~n7051 ;
  assign n7062 = n7061 ^ n7050 ;
  assign n7063 = n7062 ^ n7051 ;
  assign n7064 = n7063 ^ n7061 ;
  assign n6997 = n5203 ^ n5190 ;
  assign n6998 = n6997 ^ n5480 ;
  assign n6999 = n5124 & n6998 ;
  assign n6996 = n5202 ^ n5198 ;
  assign n7000 = n6999 ^ n6996 ;
  assign n7001 = ~n5123 & n7000 ;
  assign n7002 = n7001 ^ n5202 ;
  assign n7021 = n5270 ^ n5192 ;
  assign n7022 = n5266 & n7021 ;
  assign n7003 = n5270 ^ n5188 ;
  assign n7004 = ~n5266 & n7003 ;
  assign n7009 = ~n5268 & n5477 ;
  assign n7010 = n7009 ^ n5229 ;
  assign n7011 = ~n7004 & n7010 ;
  assign n7012 = n7011 ^ n5484 ;
  assign n7013 = n7012 ^ n5475 ;
  assign n7014 = n7013 ^ n7011 ;
  assign n7017 = n5123 & n7014 ;
  assign n7018 = n7017 ^ n7011 ;
  assign n7019 = n5210 & n7018 ;
  assign n7020 = n7019 ^ n7011 ;
  assign n7023 = n7022 ^ n7020 ;
  assign n7024 = ~n7002 & ~n7023 ;
  assign n7025 = ~n5503 & n7024 ;
  assign n7026 = ~n5203 & n7025 ;
  assign n7027 = n7026 ^ n3424 ;
  assign n7028 = n7027 ^ x118 ;
  assign n7029 = n6535 ^ x125 ;
  assign n7030 = ~n7028 & n7029 ;
  assign n7031 = n7030 ^ n7029 ;
  assign n6643 = n4801 ^ n4691 ;
  assign n6644 = n6643 ^ n4786 ;
  assign n6645 = n6644 ^ n4773 ;
  assign n6646 = n5838 & n6645 ;
  assign n6638 = n5859 ^ n4787 ;
  assign n6639 = n4835 & n6638 ;
  assign n6634 = n4842 & ~n5834 ;
  assign n6631 = n4844 ^ n4800 ;
  assign n6632 = n6631 ^ n6630 ;
  assign n6633 = n6632 ^ n4840 ;
  assign n6635 = n6634 ^ n6633 ;
  assign n6636 = n6635 ^ n6630 ;
  assign n6637 = n6636 ^ n4840 ;
  assign n6640 = n6639 ^ n6637 ;
  assign n6641 = n4853 & ~n6640 ;
  assign n6642 = n6641 ^ n6635 ;
  assign n6647 = n6646 ^ n6642 ;
  assign n6627 = n4796 ^ n4793 ;
  assign n6628 = ~n5836 & n6627 ;
  assign n6648 = n6647 ^ n6628 ;
  assign n6655 = n6648 & ~n6654 ;
  assign n6658 = n6655 ^ n3163 ;
  assign n6656 = n4835 & n6655 ;
  assign n6657 = n5841 & n6656 ;
  assign n6659 = n6658 ^ n6657 ;
  assign n6969 = n6659 ^ x84 ;
  assign n6975 = n4234 ^ n4215 ;
  assign n6976 = n6975 ^ n4267 ;
  assign n6977 = n6976 ^ n4238 ;
  assign n6978 = n4203 & n6977 ;
  assign n6979 = n6978 ^ n4234 ;
  assign n6986 = n6979 ^ n4274 ;
  assign n6985 = n4299 ^ n4218 ;
  assign n6987 = n6986 ^ n6985 ;
  assign n6984 = ~n4203 & n4272 ;
  assign n6988 = n6987 ^ n6984 ;
  assign n6974 = n4282 ^ n4248 ;
  assign n6980 = n6979 ^ n6974 ;
  assign n6981 = n6980 ^ n4275 ;
  assign n6970 = n4232 ^ n4169 ;
  assign n6971 = n6970 ^ n4231 ;
  assign n6972 = n6971 ^ n4248 ;
  assign n6973 = n4203 & n6972 ;
  assign n6982 = n6981 ^ n6973 ;
  assign n6983 = ~n4202 & ~n6982 ;
  assign n6989 = n6988 ^ n6983 ;
  assign n6990 = n6989 ^ n4291 ;
  assign n6991 = ~n4205 & n6990 ;
  assign n6992 = ~n5417 & n6991 ;
  assign n6993 = n6992 ^ n3397 ;
  assign n6994 = n6993 ^ x69 ;
  assign n6995 = ~n6969 & n6994 ;
  assign n7033 = n6995 ^ n6994 ;
  assign n7034 = n7033 ^ n6969 ;
  assign n7090 = n7031 & n7034 ;
  assign n7067 = n7028 & n7034 ;
  assign n7091 = n7090 ^ n7067 ;
  assign n7038 = n7030 ^ n7028 ;
  assign n7070 = n6995 & ~n7038 ;
  assign n7035 = n7034 ^ n6994 ;
  assign n7039 = ~n7035 & ~n7038 ;
  assign n7071 = n7070 ^ n7039 ;
  assign n7047 = n7033 & ~n7038 ;
  assign n7069 = n7047 ^ n7038 ;
  assign n7072 = n7071 ^ n7069 ;
  assign n7068 = n7067 ^ n7034 ;
  assign n7073 = n7072 ^ n7068 ;
  assign n7092 = n7091 ^ n7073 ;
  assign n7046 = n7031 & n7033 ;
  assign n7048 = n7047 ^ n7046 ;
  assign n8150 = n7092 ^ n7048 ;
  assign n7032 = n6995 & n7031 ;
  assign n8144 = n7072 ^ n7032 ;
  assign n8145 = n8144 ^ n7092 ;
  assign n7052 = n7051 ^ n7050 ;
  assign n8146 = n7092 ^ n7051 ;
  assign n8147 = n7052 & ~n8146 ;
  assign n8148 = n8147 ^ n7051 ;
  assign n8149 = n8145 & n8148 ;
  assign n8151 = n8150 ^ n8149 ;
  assign n7066 = n6995 & n7030 ;
  assign n7074 = n7073 ^ n7066 ;
  assign n7041 = n7031 ^ n7028 ;
  assign n7042 = ~n7035 & n7041 ;
  assign n7040 = n7039 ^ n7032 ;
  assign n7043 = n7042 ^ n7040 ;
  assign n7037 = n7031 & ~n7035 ;
  assign n7044 = n7043 ^ n7037 ;
  assign n7036 = n7035 ^ n7032 ;
  assign n7045 = n7044 ^ n7036 ;
  assign n7065 = n7045 ^ n7030 ;
  assign n7075 = n7074 ^ n7065 ;
  assign n7108 = n7075 ^ n7072 ;
  assign n7984 = n7108 ^ n7037 ;
  assign n7985 = n7050 & ~n7984 ;
  assign n7986 = n7985 ^ n7037 ;
  assign n8139 = n7986 ^ n7073 ;
  assign n8143 = n8139 ^ n7066 ;
  assign n8152 = n8151 ^ n8143 ;
  assign n8153 = ~n7064 & n8152 ;
  assign n7669 = n7066 ^ n7037 ;
  assign n7085 = n7070 ^ n7066 ;
  assign n7086 = n7085 ^ n6969 ;
  assign n7087 = n7086 ^ n7036 ;
  assign n7668 = n7087 ^ n7037 ;
  assign n7670 = n7669 ^ n7668 ;
  assign n7671 = n7669 ^ n7050 ;
  assign n7672 = n7671 ^ n7669 ;
  assign n7673 = n7670 & ~n7672 ;
  assign n7674 = n7673 ^ n7669 ;
  assign n7675 = n7052 & n7674 ;
  assign n7676 = n7675 ^ n7037 ;
  assign n8140 = n8139 ^ n7676 ;
  assign n7077 = n7046 ^ n7033 ;
  assign n7076 = n7075 ^ n7047 ;
  assign n7078 = n7077 ^ n7076 ;
  assign n7079 = n7078 ^ n7070 ;
  assign n7080 = n7070 ^ n7050 ;
  assign n7081 = n7080 ^ n7070 ;
  assign n7082 = n7079 & n7081 ;
  assign n7083 = n7082 ^ n7070 ;
  assign n7084 = n7064 & n7083 ;
  assign n8141 = n8140 ^ n7084 ;
  assign n7088 = n7087 ^ n7050 ;
  assign n7089 = n7088 ^ n7087 ;
  assign n7679 = n7091 ^ n7075 ;
  assign n8002 = n7679 ^ n7087 ;
  assign n8003 = ~n7089 & n8002 ;
  assign n8004 = n8003 ^ n7087 ;
  assign n8005 = n7064 & n8004 ;
  assign n8142 = n8141 ^ n8005 ;
  assign n8154 = n8153 ^ n8142 ;
  assign n7124 = n7045 ^ n7042 ;
  assign n7125 = n7062 & ~n7124 ;
  assign n8155 = n8154 ^ n7125 ;
  assign n8132 = n7071 ^ n7050 ;
  assign n8133 = n8132 ^ n7071 ;
  assign n8134 = n7042 ^ n7032 ;
  assign n8135 = n8134 ^ n7071 ;
  assign n8136 = n8133 & n8135 ;
  assign n8137 = n8136 ^ n7071 ;
  assign n8138 = ~n7051 & n8137 ;
  assign n8156 = n8155 ^ n8138 ;
  assign n7099 = n7090 ^ n7078 ;
  assign n7127 = n7063 & n7099 ;
  assign n8157 = n8156 ^ n7127 ;
  assign n8158 = n8157 ^ n4688 ;
  assign n8159 = n8158 ^ x125 ;
  assign n8281 = n8271 ^ n8159 ;
  assign n8282 = n8280 & n8281 ;
  assign n8235 = n8234 ^ n8187 ;
  assign n8269 = n8268 ^ n8235 ;
  assign n8270 = n8269 ^ n8267 ;
  assign n8274 = n8270 & n8271 ;
  assign n8275 = n8274 ^ n8267 ;
  assign n8276 = ~n8159 & n8275 ;
  assign n8283 = n8282 ^ n8276 ;
  assign n8284 = n8159 & ~n8271 ;
  assign n8285 = n8284 ^ n8271 ;
  assign n8890 = n8280 & ~n8285 ;
  assign n8318 = n8258 ^ n8240 ;
  assign n8319 = n8284 & n8318 ;
  assign n8891 = n8890 ^ n8319 ;
  assign n8871 = n8188 & n8230 ;
  assign n8298 = n8269 ^ n8237 ;
  assign n8870 = n8298 ^ n8233 ;
  assign n8872 = n8871 ^ n8870 ;
  assign n8869 = n8278 ^ n8188 ;
  assign n8873 = n8872 ^ n8869 ;
  assign n8874 = n8873 ^ n8244 ;
  assign n8306 = n8259 ^ n8251 ;
  assign n8868 = n8306 ^ n8237 ;
  assign n8875 = n8874 ^ n8868 ;
  assign n8864 = n8229 ^ n8185 ;
  assign n8865 = n8864 ^ n8248 ;
  assign n8866 = n8865 ^ n8278 ;
  assign n8867 = n8159 & ~n8866 ;
  assign n8876 = n8875 ^ n8867 ;
  assign n8892 = n8891 ^ n8876 ;
  assign n8286 = n8285 ^ n8159 ;
  assign n8888 = n8874 ^ n8871 ;
  assign n8889 = n8286 & n8888 ;
  assign n8893 = n8892 ^ n8889 ;
  assign n8885 = n8871 ^ n8267 ;
  assign n8886 = n8885 ^ n8243 ;
  assign n8887 = n8284 & n8886 ;
  assign n8894 = n8893 ^ n8887 ;
  assign n8877 = n8876 ^ n8261 ;
  assign n8878 = n8877 ^ n8265 ;
  assign n8879 = n8878 ^ n8877 ;
  assign n8880 = n8877 ^ n8271 ;
  assign n8881 = n8880 ^ n8877 ;
  assign n8882 = ~n8879 & n8881 ;
  assign n8883 = n8882 ^ n8877 ;
  assign n8884 = n8281 & n8883 ;
  assign n8895 = n8894 ^ n8884 ;
  assign n8896 = ~n8283 & ~n8895 ;
  assign n8897 = n8896 ^ n5819 ;
  assign n8898 = n8897 ^ x72 ;
  assign n6328 = n6256 & n6298 ;
  assign n6335 = n6334 ^ n6328 ;
  assign n6336 = n6334 ^ n6194 ;
  assign n6337 = n6336 ^ n6334 ;
  assign n6338 = n6335 & ~n6337 ;
  assign n6339 = n6338 ^ n6334 ;
  assign n6340 = n6193 & n6339 ;
  assign n6342 = n6305 ^ n6300 ;
  assign n6345 = n6300 ^ n6193 ;
  assign n6346 = n6345 ^ n6300 ;
  assign n6347 = n6342 & n6346 ;
  assign n6348 = n6347 ^ n6300 ;
  assign n6349 = ~n6314 & n6348 ;
  assign n7713 = n6308 ^ n6303 ;
  assign n7709 = n6321 ^ n6311 ;
  assign n7707 = n6350 ^ n6330 ;
  assign n7708 = n7707 ^ n6328 ;
  assign n7710 = n7709 ^ n7708 ;
  assign n7711 = ~n6193 & n7710 ;
  assign n7705 = n6351 ^ n6330 ;
  assign n7706 = n7705 ^ n6350 ;
  assign n7712 = n7711 ^ n7706 ;
  assign n7714 = n7713 ^ n7712 ;
  assign n7715 = n6314 & n7714 ;
  assign n6366 = n6365 ^ n6332 ;
  assign n7704 = n6196 & n6366 ;
  assign n7716 = n7715 ^ n7704 ;
  assign n7724 = n7723 ^ n7191 ;
  assign n7717 = n6308 ^ n6306 ;
  assign n7718 = n7717 ^ n6355 ;
  assign n7719 = n7718 ^ n7709 ;
  assign n7720 = ~n6193 & n7719 ;
  assign n7725 = n7724 ^ n7720 ;
  assign n7726 = ~n6314 & ~n7725 ;
  assign n7727 = ~n7723 & n7726 ;
  assign n7728 = n7727 ^ n6314 ;
  assign n7729 = ~n7716 & n7728 ;
  assign n7731 = n7730 ^ n7729 ;
  assign n7732 = ~n6349 & n7731 ;
  assign n7733 = ~n6340 & n7732 ;
  assign n7734 = ~n7703 & n7733 ;
  assign n7735 = n7734 ^ n2256 ;
  assign n8499 = n7735 ^ x89 ;
  assign n6610 = ~n6539 & ~n6609 ;
  assign n6613 = n6612 ^ n6610 ;
  assign n6571 = n6570 ^ n6541 ;
  assign n6569 = n6568 ^ n6567 ;
  assign n6572 = n6571 ^ n6569 ;
  assign n6573 = n6569 ^ n6537 ;
  assign n6574 = n6573 ^ n6569 ;
  assign n6575 = n6572 & ~n6574 ;
  assign n6576 = n6575 ^ n6569 ;
  assign n6577 = n6565 & n6576 ;
  assign n6578 = n6577 ^ n6569 ;
  assign n6582 = n6581 ^ n6566 ;
  assign n6583 = n6582 ^ n6537 ;
  assign n6594 = n6558 ^ n6506 ;
  assign n6595 = n6594 ^ n6537 ;
  assign n6584 = n6551 ^ n6506 ;
  assign n6585 = n6584 ^ n6561 ;
  assign n6592 = n6591 ^ n6585 ;
  assign n6593 = ~n6536 & ~n6592 ;
  assign n6596 = n6595 ^ n6593 ;
  assign n6597 = n6583 & n6596 ;
  assign n6598 = n6597 ^ n6537 ;
  assign n6599 = ~n6578 & ~n6598 ;
  assign n6564 = n6548 & n6563 ;
  assign n6600 = n6599 ^ n6564 ;
  assign n6602 = n6601 ^ n6559 ;
  assign n6603 = n6559 ^ n6536 ;
  assign n6604 = n6603 ^ n6559 ;
  assign n6605 = ~n6602 & n6604 ;
  assign n6606 = n6605 ^ n6559 ;
  assign n6607 = ~n6537 & n6606 ;
  assign n6608 = n6600 & ~n6607 ;
  assign n6614 = n6613 ^ n6608 ;
  assign n6615 = ~n6562 & n6614 ;
  assign n6622 = n6615 & ~n6621 ;
  assign n6623 = ~n6507 & n6622 ;
  assign n6624 = n6623 ^ n2825 ;
  assign n8498 = n6624 ^ x98 ;
  assign n8505 = n8499 ^ n8498 ;
  assign n6660 = n6659 ^ x94 ;
  assign n6626 = n6224 ^ x68 ;
  assign n6787 = n6660 ^ n6626 ;
  assign n6722 = n6192 ^ x126 ;
  assign n6723 = n4570 ^ n4544 ;
  assign n6724 = n6723 ^ n3175 ;
  assign n6725 = n6724 ^ x108 ;
  assign n6726 = n6722 & ~n6725 ;
  assign n6727 = n6726 ^ n6725 ;
  assign n6672 = n5452 ^ n5041 ;
  assign n6671 = n5112 ^ n5035 ;
  assign n6673 = n6672 ^ n6671 ;
  assign n6664 = n5112 ^ n5090 ;
  assign n6662 = n5058 ^ n5037 ;
  assign n6663 = n6662 ^ n5972 ;
  assign n6665 = n6664 ^ n6663 ;
  assign n6666 = n4898 & n6665 ;
  assign n6667 = n6666 ^ n6664 ;
  assign n6669 = n6667 ^ n5438 ;
  assign n6670 = n6669 ^ n6667 ;
  assign n6674 = n6673 ^ n6670 ;
  assign n6675 = ~n4898 & ~n6674 ;
  assign n6676 = n6675 ^ n6669 ;
  assign n6677 = ~n4929 & ~n6676 ;
  assign n6661 = n5465 ^ n5065 ;
  assign n6668 = n6667 ^ n6661 ;
  assign n6678 = n6677 ^ n6668 ;
  assign n6679 = n6678 ^ n5064 ;
  assign n6680 = ~n5469 & n6679 ;
  assign n6681 = n6680 ^ n3206 ;
  assign n6682 = n6681 ^ x70 ;
  assign n6719 = n6718 ^ x85 ;
  assign n6720 = ~n6682 & n6719 ;
  assign n6721 = n6720 ^ n6682 ;
  assign n6739 = n6721 ^ n6719 ;
  assign n6743 = n6739 ^ n6682 ;
  assign n6752 = ~n6727 & n6743 ;
  assign n6728 = n6727 ^ n6722 ;
  assign n6749 = n6720 & n6728 ;
  assign n6740 = n6728 & n6739 ;
  assign n6750 = n6749 ^ n6740 ;
  assign n6729 = ~n6721 & n6728 ;
  assign n6730 = n6729 ^ n6728 ;
  assign n6751 = n6750 ^ n6730 ;
  assign n6753 = n6752 ^ n6751 ;
  assign n8474 = ~n6660 & n6753 ;
  assign n8475 = n8474 ^ n6752 ;
  assign n6764 = n6726 & n6739 ;
  assign n8476 = n8475 ^ n6764 ;
  assign n6744 = n6726 & n6743 ;
  assign n6748 = n6744 ^ n6743 ;
  assign n6754 = n6753 ^ n6748 ;
  assign n8477 = n8476 ^ n6754 ;
  assign n8478 = n8477 ^ n8475 ;
  assign n8479 = n8475 ^ n6626 ;
  assign n8480 = n8479 ^ n8475 ;
  assign n8481 = n8478 & ~n8480 ;
  assign n8482 = n8481 ^ n8475 ;
  assign n8483 = ~n6787 & n8482 ;
  assign n8484 = n8483 ^ n8475 ;
  assign n8485 = n8484 ^ n3358 ;
  assign n6804 = n6626 & ~n6660 ;
  assign n6805 = n6804 ^ n6626 ;
  assign n6810 = n6764 & n6805 ;
  assign n6808 = n6804 ^ n6660 ;
  assign n6809 = n6740 & ~n6808 ;
  assign n6811 = n6810 ^ n6809 ;
  assign n8469 = ~n6626 & n6660 ;
  assign n6742 = ~n6721 & n6726 ;
  assign n7530 = n6751 ^ n6729 ;
  assign n8470 = ~n6742 & n7530 ;
  assign n8471 = n8469 & n8470 ;
  assign n6765 = n6764 ^ n6726 ;
  assign n6745 = n6744 ^ n6742 ;
  assign n6766 = n6765 ^ n6745 ;
  assign n6732 = n6722 ^ n6719 ;
  assign n6733 = ~n6682 & ~n6732 ;
  assign n6771 = n6766 ^ n6733 ;
  assign n6734 = n6733 ^ n6722 ;
  assign n6735 = n6725 ^ n6682 ;
  assign n6736 = ~n6734 & ~n6735 ;
  assign n6731 = n6730 ^ n6720 ;
  assign n6737 = n6736 ^ n6731 ;
  assign n6738 = n6737 ^ n6729 ;
  assign n6772 = n6771 ^ n6738 ;
  assign n6795 = n6772 ^ n6752 ;
  assign n8467 = n6795 & n6804 ;
  assign n6762 = n6728 ^ n6725 ;
  assign n6763 = n6739 & n6762 ;
  assign n6767 = n6766 ^ n6763 ;
  assign n6757 = n6725 ^ n6722 ;
  assign n6758 = n6757 ^ n6719 ;
  assign n6759 = n6743 ^ n6722 ;
  assign n6760 = ~n6758 & n6759 ;
  assign n6761 = n6760 ^ n6751 ;
  assign n6768 = n6767 ^ n6761 ;
  assign n6769 = n6768 ^ n6766 ;
  assign n6770 = n6769 ^ n6754 ;
  assign n6773 = n6772 ^ n6770 ;
  assign n8461 = n6773 ^ n6730 ;
  assign n8462 = n6660 & n8461 ;
  assign n6746 = n6720 & ~n6727 ;
  assign n6747 = n6746 ^ n6729 ;
  assign n8454 = n6766 ^ n6747 ;
  assign n6794 = n6746 ^ n6727 ;
  assign n6796 = n6795 ^ n6794 ;
  assign n8453 = n6796 ^ n6749 ;
  assign n8455 = n8454 ^ n8453 ;
  assign n8456 = ~n6808 & ~n8455 ;
  assign n8451 = n6762 ^ n6743 ;
  assign n8452 = n8451 ^ n6753 ;
  assign n8457 = n8456 ^ n8452 ;
  assign n8460 = n8457 ^ n8456 ;
  assign n8463 = n8462 ^ n8460 ;
  assign n8458 = n8457 ^ n6742 ;
  assign n8459 = n8458 ^ n8457 ;
  assign n8464 = n8463 ^ n8459 ;
  assign n8465 = ~n6787 & n8464 ;
  assign n8466 = n8465 ^ n8458 ;
  assign n8468 = n8467 ^ n8466 ;
  assign n8472 = n8471 ^ n8468 ;
  assign n8473 = ~n6811 & ~n8472 ;
  assign n8486 = n8485 ^ n8473 ;
  assign n8487 = n8486 ^ x65 ;
  assign n3843 = ~n3801 & n3842 ;
  assign n3823 = n2257 & n3822 ;
  assign n3818 = n3817 ^ n3812 ;
  assign n3824 = n3823 ^ n3818 ;
  assign n3838 = n3837 ^ n3824 ;
  assign n3839 = n3838 ^ n3835 ;
  assign n3825 = n3824 ^ n3527 ;
  assign n3807 = n3806 ^ n3804 ;
  assign n3819 = n3818 ^ n3807 ;
  assign n3820 = n2257 & ~n3819 ;
  assign n3826 = n3825 ^ n3820 ;
  assign n3827 = n3803 & ~n3826 ;
  assign n3840 = n3839 ^ n3827 ;
  assign n3794 = n3793 ^ n3791 ;
  assign n3798 = n3797 ^ n3794 ;
  assign n3799 = ~n2257 & n3798 ;
  assign n3841 = n3840 ^ n3799 ;
  assign n3844 = n3843 ^ n3841 ;
  assign n3845 = ~n3786 & n3844 ;
  assign n3846 = n3845 ^ n2960 ;
  assign n3847 = n3846 ^ x109 ;
  assign n4303 = n4302 ^ x102 ;
  assign n4304 = ~n3847 & n4303 ;
  assign n4574 = n4573 ^ x75 ;
  assign n4869 = n4868 ^ n4783 ;
  assign n4870 = n4869 ^ n4800 ;
  assign n4860 = n4843 ^ n4770 ;
  assign n4871 = n4870 ^ n4860 ;
  assign n4872 = ~n4607 & n4871 ;
  assign n4873 = n4872 ^ n4860 ;
  assign n4876 = n4875 ^ n4873 ;
  assign n4877 = n4876 ^ n4788 ;
  assign n4878 = n4877 ^ n4873 ;
  assign n4879 = n4873 ^ n4835 ;
  assign n4880 = n4879 ^ n4873 ;
  assign n4881 = n4878 & n4880 ;
  assign n4882 = n4881 ^ n4873 ;
  assign n4883 = ~n4853 & n4882 ;
  assign n4884 = n4883 ^ n4873 ;
  assign n4861 = n4860 ^ n4782 ;
  assign n4859 = n4845 ^ n4777 ;
  assign n4862 = n4861 ^ n4859 ;
  assign n4863 = n4859 ^ n4835 ;
  assign n4864 = n4863 ^ n4859 ;
  assign n4865 = ~n4862 & ~n4864 ;
  assign n4866 = n4865 ^ n4859 ;
  assign n4867 = ~n4607 & ~n4866 ;
  assign n4885 = n4884 ^ n4867 ;
  assign n4886 = n4885 ^ n4795 ;
  assign n4856 = n4802 & ~n4835 ;
  assign n4857 = n4856 ^ n4795 ;
  assign n4858 = n4853 & n4857 ;
  assign n4887 = n4886 ^ n4858 ;
  assign n4888 = n4887 ^ n4852 ;
  assign n4889 = n4888 ^ n4840 ;
  assign n4890 = n4889 ^ n3001 ;
  assign n4891 = n4890 ^ x124 ;
  assign n4892 = ~n4574 & n4891 ;
  assign n4896 = n4304 & n4892 ;
  assign n4893 = n4892 ^ n4574 ;
  assign n4894 = n4893 ^ n4891 ;
  assign n4895 = n4304 & n4894 ;
  assign n4897 = n4896 ^ n4895 ;
  assign n5122 = n5121 ^ x78 ;
  assign n5286 = n5285 ^ x92 ;
  assign n5287 = ~n5122 & ~n5286 ;
  assign n5288 = n5287 ^ n5286 ;
  assign n5289 = n5288 ^ n5122 ;
  assign n5290 = n4897 & ~n5289 ;
  assign n5292 = n4304 ^ n4303 ;
  assign n5293 = n5292 ^ n3847 ;
  assign n5319 = ~n4893 & n5293 ;
  assign n5318 = n4894 & n5293 ;
  assign n5320 = n5319 ^ n5318 ;
  assign n5321 = n5320 ^ n5293 ;
  assign n5294 = n4894 ^ n4574 ;
  assign n5295 = n5293 & n5294 ;
  assign n5322 = n5321 ^ n5295 ;
  assign n5323 = n5322 ^ n4892 ;
  assign n5304 = n4304 & n5294 ;
  assign n5305 = n5304 ^ n4304 ;
  assign n5306 = n5305 ^ n4897 ;
  assign n5303 = n4303 & ~n4891 ;
  assign n5307 = n5306 ^ n5303 ;
  assign n5298 = n4574 ^ n3847 ;
  assign n5299 = n5298 ^ n4891 ;
  assign n5300 = ~n4574 & ~n5299 ;
  assign n5301 = n5300 ^ n4891 ;
  assign n5302 = n4303 & ~n5301 ;
  assign n5308 = n5307 ^ n5302 ;
  assign n5317 = n5308 ^ n4896 ;
  assign n5324 = n5323 ^ n5317 ;
  assign n5336 = n5324 ^ n5318 ;
  assign n5329 = n5322 ^ n5306 ;
  assign n5328 = n5308 ^ n5300 ;
  assign n5330 = n5329 ^ n5328 ;
  assign n5331 = n5330 ^ n5308 ;
  assign n5327 = n5306 ^ n5304 ;
  assign n5332 = n5331 ^ n5327 ;
  assign n5326 = n5320 ^ n5304 ;
  assign n5333 = n5332 ^ n5326 ;
  assign n5334 = n5333 ^ n4891 ;
  assign n5335 = n5334 ^ n5302 ;
  assign n5337 = n5336 ^ n5335 ;
  assign n5338 = n5337 ^ n4895 ;
  assign n5325 = n5324 ^ n4894 ;
  assign n5339 = n5338 ^ n5325 ;
  assign n5384 = n5339 ^ n5330 ;
  assign n5385 = ~n5289 & ~n5384 ;
  assign n5315 = n5299 & n5303 ;
  assign n5316 = n5315 ^ n4895 ;
  assign n5340 = n5339 ^ n5316 ;
  assign n5314 = n5308 ^ n5292 ;
  assign n5341 = n5340 ^ n5314 ;
  assign n5378 = n5341 ^ n5339 ;
  assign n5379 = n5339 ^ n5122 ;
  assign n5380 = n5379 ^ n5339 ;
  assign n5381 = n5378 & n5380 ;
  assign n5382 = n5381 ^ n5339 ;
  assign n5383 = ~n5286 & ~n5382 ;
  assign n5386 = n5385 ^ n5383 ;
  assign n5291 = n5286 ^ n5122 ;
  assign n5349 = n4304 ^ n3847 ;
  assign n5350 = n5294 & ~n5349 ;
  assign n5351 = n5350 ^ n5318 ;
  assign n5346 = n5340 ^ n5327 ;
  assign n5352 = n5351 ^ n5346 ;
  assign n5344 = n5335 ^ n5324 ;
  assign n5345 = n5344 ^ n5315 ;
  assign n5347 = n5346 ^ n5345 ;
  assign n5348 = n5122 & n5347 ;
  assign n5353 = n5352 ^ n5348 ;
  assign n5354 = n5291 & ~n5353 ;
  assign n5355 = n5354 ^ n5350 ;
  assign n5342 = n5341 ^ n4896 ;
  assign n5343 = n5287 & ~n5342 ;
  assign n5356 = n5355 ^ n5343 ;
  assign n5359 = n5322 ^ n5122 ;
  assign n5360 = n5359 ^ n5322 ;
  assign n5361 = n5329 & n5360 ;
  assign n5362 = n5361 ^ n5322 ;
  assign n5363 = n5286 & n5362 ;
  assign n5364 = ~n5356 & ~n5363 ;
  assign n5296 = n5295 ^ n5122 ;
  assign n5297 = n5296 ^ n5295 ;
  assign n5311 = n5297 & n5308 ;
  assign n5312 = n5311 ^ n5295 ;
  assign n5313 = ~n5291 & n5312 ;
  assign n5365 = n5364 ^ n5313 ;
  assign n5309 = n5308 ^ n5295 ;
  assign n5366 = n5330 ^ n5309 ;
  assign n5367 = ~n5122 & n5366 ;
  assign n5368 = n5367 ^ n5308 ;
  assign n5369 = n5368 ^ n5322 ;
  assign n5370 = n5369 ^ n5368 ;
  assign n5371 = n5368 ^ n5286 ;
  assign n5372 = n5371 ^ n5368 ;
  assign n5373 = n5370 & ~n5372 ;
  assign n5374 = n5373 ^ n5368 ;
  assign n5375 = ~n5291 & n5374 ;
  assign n5376 = n5375 ^ n5368 ;
  assign n5377 = n5365 & ~n5376 ;
  assign n5387 = n5386 ^ n5377 ;
  assign n5388 = ~n5290 & n5387 ;
  assign n5389 = n5335 ^ n5319 ;
  assign n5390 = n5389 ^ n5350 ;
  assign n5391 = n5350 ^ n5122 ;
  assign n5392 = n5391 ^ n5350 ;
  assign n5393 = ~n5390 & ~n5392 ;
  assign n5394 = n5393 ^ n5350 ;
  assign n5395 = ~n5286 & n5394 ;
  assign n5396 = n5388 & ~n5395 ;
  assign n5397 = n5396 ^ n3123 ;
  assign n8488 = n5397 ^ x104 ;
  assign n8489 = n8487 & ~n8488 ;
  assign n7696 = n7127 ^ n3525 ;
  assign n7122 = n7042 & n7063 ;
  assign n7049 = n7048 ^ n7045 ;
  assign n7684 = n7067 ^ n7049 ;
  assign n7685 = n7050 & ~n7684 ;
  assign n7686 = n7685 ^ n7071 ;
  assign n7691 = n7686 ^ n7050 ;
  assign n7692 = n7051 & n7691 ;
  assign n7683 = n7679 ^ n7099 ;
  assign n7687 = n7686 ^ n7683 ;
  assign n7678 = n7108 ^ n7032 ;
  assign n7680 = n7679 ^ n7678 ;
  assign n7681 = n7680 ^ n7099 ;
  assign n7682 = n7051 & ~n7681 ;
  assign n7688 = n7687 ^ n7682 ;
  assign n7689 = ~n7050 & ~n7688 ;
  assign n7095 = n7089 & ~n7092 ;
  assign n7096 = n7095 ^ n7087 ;
  assign n7097 = ~n7051 & n7096 ;
  assign n7677 = n7676 ^ n7097 ;
  assign n7690 = n7689 ^ n7677 ;
  assign n7693 = n7692 ^ n7690 ;
  assign n7661 = n7070 ^ n7063 ;
  assign n7662 = n7661 ^ n7072 ;
  assign n7663 = n7662 ^ n7046 ;
  assign n7664 = n7061 & n7663 ;
  assign n7665 = n7664 ^ n7063 ;
  assign n7666 = n7061 ^ n7045 ;
  assign n7667 = n7665 & ~n7666 ;
  assign n7694 = n7693 ^ n7667 ;
  assign n7695 = ~n7122 & n7694 ;
  assign n7697 = n7696 ^ n7695 ;
  assign n8424 = n7697 ^ x113 ;
  assign n7353 = n7266 & ~n7323 ;
  assign n8446 = n7353 ^ n3779 ;
  assign n7484 = ~n7215 & n7278 ;
  assign n7485 = n7484 ^ n7483 ;
  assign n8443 = n8032 ^ n7485 ;
  assign n7486 = n7268 & n7328 ;
  assign n7300 = n7299 ^ n7295 ;
  assign n7301 = n7295 ^ n7213 ;
  assign n7302 = n7301 ^ n7295 ;
  assign n7303 = ~n7300 & ~n7302 ;
  assign n7304 = n7303 ^ n7295 ;
  assign n7305 = n7212 & n7304 ;
  assign n7487 = n7486 ^ n7305 ;
  assign n8439 = ~n7215 & n7296 ;
  assign n8437 = ~n7323 & n7336 ;
  assign n7327 = n7326 ^ n7325 ;
  assign n8435 = n7268 & n7327 ;
  assign n8432 = n7278 ^ n7262 ;
  assign n8433 = n7214 & n8432 ;
  assign n8426 = n7339 ^ n7273 ;
  assign n7308 = n7307 ^ n7262 ;
  assign n8427 = n8426 ^ n7308 ;
  assign n8428 = ~n7213 & ~n8427 ;
  assign n8425 = n8036 ^ n7327 ;
  assign n8429 = n8428 ^ n8425 ;
  assign n8430 = ~n7212 & ~n8429 ;
  assign n8431 = n8430 ^ n8428 ;
  assign n8434 = n8433 ^ n8431 ;
  assign n8436 = n8435 ^ n8434 ;
  assign n8438 = n8437 ^ n8436 ;
  assign n8440 = n8439 ^ n8438 ;
  assign n8441 = ~n7506 & ~n8440 ;
  assign n8442 = ~n7487 & n8441 ;
  assign n8444 = n8443 ^ n8442 ;
  assign n8445 = ~n7264 & n8444 ;
  assign n8447 = n8446 ^ n8445 ;
  assign n8448 = n8447 ^ x123 ;
  assign n8449 = n8424 & ~n8448 ;
  assign n8450 = n8449 ^ n8448 ;
  assign n8506 = n8450 ^ n8424 ;
  assign n8552 = n8489 & n8506 ;
  assign n8494 = n8489 ^ n8488 ;
  assign n8520 = n8494 ^ n8487 ;
  assign n8521 = n8449 & n8520 ;
  assign n8572 = n8552 ^ n8521 ;
  assign n8525 = n8449 & ~n8494 ;
  assign n8526 = n8525 ^ n8521 ;
  assign n8490 = n8489 ^ n8487 ;
  assign n8523 = n8449 & n8490 ;
  assign n8524 = n8523 ^ n8449 ;
  assign n8527 = n8526 ^ n8524 ;
  assign n8516 = n8449 ^ n8424 ;
  assign n8517 = n8490 & n8516 ;
  assign n8528 = n8527 ^ n8517 ;
  assign n8573 = n8572 ^ n8528 ;
  assign n8574 = ~n8499 & n8573 ;
  assign n8500 = n8498 & n8499 ;
  assign n8547 = n8500 & n8527 ;
  assign n8501 = n8500 ^ n8498 ;
  assign n8545 = n8516 & n8520 ;
  assign n8546 = ~n8501 & ~n8545 ;
  assign n8548 = n8547 ^ n8546 ;
  assign n8519 = n8489 & n8516 ;
  assign n8522 = n8521 ^ n8519 ;
  assign n8549 = n8548 ^ n8522 ;
  assign n8575 = n8574 ^ n8549 ;
  assign n8576 = n8505 & ~n8575 ;
  assign n8502 = n8501 ^ n8499 ;
  assign n8507 = n8490 & n8506 ;
  assign n8569 = n8525 ^ n8507 ;
  assign n8570 = ~n8502 & n8569 ;
  assign n8562 = n8528 ^ n8520 ;
  assign n8529 = n8528 ^ n8522 ;
  assign n8511 = n8488 ^ n8448 ;
  assign n8512 = n8424 & n8511 ;
  assign n8492 = ~n8450 & n8489 ;
  assign n8513 = n8512 ^ n8492 ;
  assign n8509 = n8448 ^ n8424 ;
  assign n8510 = n8509 ^ n8488 ;
  assign n8514 = n8513 ^ n8510 ;
  assign n8495 = ~n8450 & ~n8494 ;
  assign n8508 = n8507 ^ n8495 ;
  assign n8515 = n8514 ^ n8508 ;
  assign n8518 = n8517 ^ n8515 ;
  assign n8530 = n8529 ^ n8518 ;
  assign n8531 = n8530 ^ n8509 ;
  assign n8491 = ~n8450 & n8490 ;
  assign n8493 = n8492 ^ n8491 ;
  assign n8496 = n8495 ^ n8493 ;
  assign n8532 = n8531 ^ n8496 ;
  assign n8563 = n8562 ^ n8532 ;
  assign n8564 = n8501 & n8563 ;
  assign n8553 = n8552 ^ n8515 ;
  assign n8551 = n8507 ^ n8506 ;
  assign n8554 = n8553 ^ n8551 ;
  assign n8497 = n8496 ^ n8450 ;
  assign n8555 = n8554 ^ n8497 ;
  assign n8556 = n8555 ^ n8545 ;
  assign n8557 = n8545 ^ n8499 ;
  assign n8558 = n8557 ^ n8545 ;
  assign n8559 = n8556 & ~n8558 ;
  assign n8560 = n8559 ^ n8545 ;
  assign n8561 = n8505 & n8560 ;
  assign n8565 = n8564 ^ n8561 ;
  assign n8550 = n8549 ^ n8496 ;
  assign n8566 = n8565 ^ n8550 ;
  assign n8539 = n8515 ^ n8491 ;
  assign n8540 = n8515 ^ n8499 ;
  assign n8541 = n8540 ^ n8515 ;
  assign n8542 = ~n8539 & ~n8541 ;
  assign n8543 = n8542 ^ n8515 ;
  assign n8544 = n8498 & ~n8543 ;
  assign n8567 = n8566 ^ n8544 ;
  assign n8534 = n8499 ^ n8496 ;
  assign n8535 = n8534 ^ n8496 ;
  assign n8536 = ~n8531 & n8535 ;
  assign n8537 = n8536 ^ n8496 ;
  assign n8538 = n8505 & n8537 ;
  assign n8568 = n8567 ^ n8538 ;
  assign n8571 = n8570 ^ n8568 ;
  assign n8577 = n8576 ^ n8571 ;
  assign n8503 = n8502 ^ n8498 ;
  assign n8504 = ~n8497 & n8503 ;
  assign n8578 = n8577 ^ n8504 ;
  assign n8579 = n8578 ^ n6069 ;
  assign n8580 = n8579 ^ x98 ;
  assign n8899 = n8898 ^ n8580 ;
  assign n7698 = n7697 ^ x73 ;
  assign n7532 = n6796 ^ n6763 ;
  assign n6755 = n6754 ^ n6747 ;
  assign n6756 = n6755 ^ n6752 ;
  assign n7533 = n7532 ^ n6756 ;
  assign n6780 = n6758 ^ n6736 ;
  assign n7534 = n7533 ^ n6780 ;
  assign n7535 = n6626 & n7534 ;
  assign n7536 = n7535 ^ n6780 ;
  assign n7540 = n7536 ^ n6810 ;
  assign n6797 = n6796 ^ n6751 ;
  assign n6798 = n6797 ^ n6795 ;
  assign n6799 = n6795 ^ n6626 ;
  assign n6800 = n6799 ^ n6795 ;
  assign n6801 = ~n6798 & ~n6800 ;
  assign n6802 = n6801 ^ n6795 ;
  assign n6803 = n6660 & n6802 ;
  assign n7541 = n7540 ^ n6803 ;
  assign n7531 = n7530 ^ n6744 ;
  assign n7537 = n7536 ^ n7531 ;
  assign n7528 = n6760 ^ n6722 ;
  assign n7529 = ~n6626 & n7528 ;
  assign n7538 = n7537 ^ n7529 ;
  assign n7539 = n6660 & ~n7538 ;
  assign n7542 = n7541 ^ n7539 ;
  assign n7527 = n6767 & n6805 ;
  assign n7543 = n7542 ^ n7527 ;
  assign n7544 = n6746 ^ n6745 ;
  assign n7545 = n6745 ^ n6660 ;
  assign n7546 = n7545 ^ n6745 ;
  assign n7547 = n7544 & n7546 ;
  assign n7548 = n7547 ^ n6745 ;
  assign n7549 = n6787 & n7548 ;
  assign n7550 = n7543 & ~n7549 ;
  assign n7551 = n7550 ^ n4201 ;
  assign n7699 = n7551 ^ x66 ;
  assign n7700 = ~n7698 & n7699 ;
  assign n7862 = n7700 ^ n7698 ;
  assign n7872 = n7862 ^ n7699 ;
  assign n6100 = n6077 & ~n6099 ;
  assign n6101 = n6100 ^ n6071 ;
  assign n6084 = n6083 ^ n6082 ;
  assign n6102 = n6101 ^ n6084 ;
  assign n6104 = n6103 ^ n6102 ;
  assign n6112 = n6111 ^ n6104 ;
  assign n6075 = n5988 & ~n6074 ;
  assign n6078 = n6077 ^ n6075 ;
  assign n7583 = n6084 ^ n6078 ;
  assign n7584 = n5968 & n7583 ;
  assign n7585 = n7584 ^ n6084 ;
  assign n7587 = n7585 ^ n6101 ;
  assign n6156 = n6095 ^ n6092 ;
  assign n7586 = n7585 ^ n6156 ;
  assign n7588 = n7587 ^ n7586 ;
  assign n7591 = n5968 & n7588 ;
  assign n7592 = n7591 ^ n7587 ;
  assign n7593 = n6146 & n7592 ;
  assign n7594 = n7593 ^ n7585 ;
  assign n7595 = ~n6112 & n7594 ;
  assign n7596 = n7595 ^ n3959 ;
  assign n7701 = n7596 ^ x107 ;
  assign n7736 = n7735 ^ x105 ;
  assign n7737 = ~n7701 & ~n7736 ;
  assign n7754 = n5384 ^ n5320 ;
  assign n7755 = n7754 ^ n5350 ;
  assign n7756 = n5122 & ~n7755 ;
  assign n7757 = n7756 ^ n5316 ;
  assign n7758 = ~n5286 & n7757 ;
  assign n7759 = n7758 ^ n5316 ;
  assign n7747 = n5338 ^ n5306 ;
  assign n7748 = n7747 ^ n5317 ;
  assign n7749 = n5317 ^ n5286 ;
  assign n7750 = n7749 ^ n5317 ;
  assign n7751 = ~n7748 & ~n7750 ;
  assign n7752 = n7751 ^ n5317 ;
  assign n7753 = ~n5122 & n7752 ;
  assign n7760 = n7759 ^ n7753 ;
  assign n7761 = n7760 ^ n5304 ;
  assign n6939 = n5341 ^ n5335 ;
  assign n6940 = n5335 ^ n5122 ;
  assign n6941 = n6940 ^ n5335 ;
  assign n6942 = n6939 & n6941 ;
  assign n6943 = n6942 ^ n5335 ;
  assign n6944 = n5286 & ~n6943 ;
  assign n7762 = n7761 ^ n6944 ;
  assign n7763 = n7762 ^ n5376 ;
  assign n7764 = n7763 ^ n5383 ;
  assign n7740 = n5304 ^ n5286 ;
  assign n7741 = n7740 ^ n5304 ;
  assign n7742 = n5336 ^ n5304 ;
  assign n7743 = n7742 ^ n5304 ;
  assign n7744 = n7741 & n7743 ;
  assign n7745 = n7744 ^ n5304 ;
  assign n7746 = ~n5291 & n7745 ;
  assign n7765 = n7764 ^ n7746 ;
  assign n7766 = n5350 ^ n5341 ;
  assign n7767 = n5341 ^ n5286 ;
  assign n7768 = n7767 ^ n5341 ;
  assign n7769 = ~n7766 & n7768 ;
  assign n7770 = n7769 ^ n5341 ;
  assign n7771 = ~n5122 & ~n7770 ;
  assign n7772 = ~n7765 & ~n7771 ;
  assign n7738 = n5290 ^ n4163 ;
  assign n7739 = n7738 ^ n5385 ;
  assign n7773 = n7772 ^ n7739 ;
  assign n7774 = n7773 ^ x80 ;
  assign n7814 = n6927 ^ n4124 ;
  assign n5944 = n5892 & n5939 ;
  assign n5946 = n5945 ^ n5944 ;
  assign n5928 = n5883 ^ n5827 ;
  assign n5929 = n5928 ^ n5893 ;
  assign n5930 = n5893 ^ n5427 ;
  assign n5931 = n5930 ^ n5893 ;
  assign n5932 = ~n5929 & ~n5931 ;
  assign n5933 = n5932 ^ n5893 ;
  assign n5934 = n5877 & ~n5933 ;
  assign n5918 = ~n5914 & ~n5915 ;
  assign n5919 = n5918 ^ n5824 ;
  assign n5920 = ~n5877 & n5919 ;
  assign n6908 = n5936 ^ n5896 ;
  assign n6909 = n5896 ^ n5877 ;
  assign n6910 = n6909 ^ n5896 ;
  assign n6911 = ~n6908 & ~n6910 ;
  assign n6912 = n6911 ^ n5896 ;
  assign n6913 = n5427 & n6912 ;
  assign n6899 = n5892 ^ n5831 ;
  assign n6900 = n6899 ^ n5824 ;
  assign n7782 = n6900 ^ n5883 ;
  assign n5949 = n5905 ^ n5827 ;
  assign n7781 = n5949 ^ n5831 ;
  assign n7783 = n7782 ^ n7781 ;
  assign n7784 = n7781 ^ n5427 ;
  assign n7785 = n5948 & ~n7784 ;
  assign n7786 = n7785 ^ n5427 ;
  assign n7787 = n7783 & ~n7786 ;
  assign n7788 = n7787 ^ n7781 ;
  assign n7789 = n7788 ^ n5897 ;
  assign n7790 = n7789 ^ n5823 ;
  assign n5951 = n5895 ^ n5884 ;
  assign n7777 = n5951 ^ n5936 ;
  assign n7775 = n5923 ^ n5899 ;
  assign n7776 = n7775 ^ n6899 ;
  assign n7778 = n7777 ^ n7776 ;
  assign n7779 = ~n5877 & ~n7778 ;
  assign n7780 = n7779 ^ n7777 ;
  assign n7791 = n7790 ^ n7780 ;
  assign n7798 = n7791 ^ n5893 ;
  assign n7799 = n7798 ^ n7791 ;
  assign n7802 = n7791 ^ n5427 ;
  assign n7803 = n7802 ^ n7791 ;
  assign n7804 = ~n7790 & ~n7803 ;
  assign n7805 = ~n7799 & n7804 ;
  assign n7806 = n7805 ^ n7799 ;
  assign n7807 = n7806 ^ n7798 ;
  assign n7808 = ~n5948 & n7807 ;
  assign n7809 = n7808 ^ n7780 ;
  assign n7810 = ~n6913 & ~n7809 ;
  assign n7811 = ~n5920 & n7810 ;
  assign n7812 = ~n5934 & n7811 ;
  assign n7813 = ~n5946 & n7812 ;
  assign n7815 = n7814 ^ n7813 ;
  assign n7816 = n7815 ^ x90 ;
  assign n7817 = n7774 & n7816 ;
  assign n7829 = n7817 ^ n7816 ;
  assign n7833 = n7829 ^ n7774 ;
  assign n7835 = n7737 & ~n7833 ;
  assign n7819 = n7737 & ~n7774 ;
  assign n7838 = n7835 ^ n7819 ;
  assign n7822 = n7737 ^ n7701 ;
  assign n7823 = n7817 ^ n7774 ;
  assign n7824 = ~n7822 & n7823 ;
  assign n7905 = n7838 ^ n7824 ;
  assign n7906 = n7872 & n7905 ;
  assign n7827 = n7737 ^ n7736 ;
  assign n7830 = n7827 ^ n7701 ;
  assign n7831 = n7829 & ~n7830 ;
  assign n7820 = n7819 ^ n7737 ;
  assign n7818 = n7737 & n7817 ;
  assign n7821 = n7820 ^ n7818 ;
  assign n7825 = n7824 ^ n7821 ;
  assign n7826 = n7700 & n7825 ;
  assign n8610 = n7831 ^ n7826 ;
  assign n7870 = n7699 ^ n7698 ;
  assign n7854 = n7823 & ~n7830 ;
  assign n7850 = ~n7827 & ~n7833 ;
  assign n7851 = n7850 ^ n7833 ;
  assign n7834 = ~n7822 & ~n7833 ;
  assign n7836 = n7835 ^ n7834 ;
  assign n7852 = n7851 ^ n7836 ;
  assign n7866 = n7854 ^ n7852 ;
  assign n7865 = n7831 ^ n7830 ;
  assign n7867 = n7866 ^ n7865 ;
  assign n7879 = n7867 ^ n7852 ;
  assign n7840 = n7817 & ~n7822 ;
  assign n7839 = n7838 ^ n7821 ;
  assign n7841 = n7840 ^ n7839 ;
  assign n7837 = n7836 ^ n7818 ;
  assign n7842 = n7841 ^ n7837 ;
  assign n7832 = n7824 ^ n7701 ;
  assign n7843 = n7842 ^ n7832 ;
  assign n7844 = n7843 ^ n7838 ;
  assign n7845 = n7844 ^ n7829 ;
  assign n7846 = n7845 ^ n7831 ;
  assign n8603 = n7879 ^ n7846 ;
  assign n7828 = n7817 & ~n7827 ;
  assign n8602 = n7866 ^ n7828 ;
  assign n8604 = n8603 ^ n8602 ;
  assign n8605 = n8602 ^ n7699 ;
  assign n8606 = n8605 ^ n8602 ;
  assign n8607 = ~n8604 & ~n8606 ;
  assign n8608 = n8607 ^ n8602 ;
  assign n8609 = ~n7870 & ~n8608 ;
  assign n8611 = n8610 ^ n8609 ;
  assign n7847 = n7846 ^ n7828 ;
  assign n7855 = n7854 ^ n7847 ;
  assign n7881 = n7855 ^ n7701 ;
  assign n7863 = n7850 ^ n7831 ;
  assign n7880 = n7879 ^ n7863 ;
  assign n7882 = n7881 ^ n7880 ;
  assign n8599 = n7882 ^ n7828 ;
  assign n8600 = n8599 ^ n7837 ;
  assign n8601 = n7872 & ~n8600 ;
  assign n8612 = n8611 ^ n8601 ;
  assign n8590 = n7846 ^ n7818 ;
  assign n8591 = n8590 ^ n7843 ;
  assign n8589 = n7867 ^ n7850 ;
  assign n8592 = n8591 ^ n8589 ;
  assign n8588 = n7854 ^ n7821 ;
  assign n8593 = n8592 ^ n8588 ;
  assign n8594 = n8592 ^ n7699 ;
  assign n8595 = n8594 ^ n8592 ;
  assign n8596 = n8593 & ~n8595 ;
  assign n8597 = n8596 ^ n8592 ;
  assign n8598 = ~n7698 & ~n8597 ;
  assign n8613 = n8612 ^ n8598 ;
  assign n7886 = n7840 ^ n7835 ;
  assign n7873 = n7872 ^ n7698 ;
  assign n8581 = n7886 ^ n7873 ;
  assign n8582 = n7862 ^ n7844 ;
  assign n8583 = n7873 ^ n7862 ;
  assign n8584 = n8583 ^ n7862 ;
  assign n8585 = ~n8582 & n8584 ;
  assign n8586 = n8585 ^ n7862 ;
  assign n8587 = n8581 & ~n8586 ;
  assign n8614 = n8613 ^ n8587 ;
  assign n8615 = ~n7906 & n8614 ;
  assign n8616 = n8615 ^ n5426 ;
  assign n8617 = n8616 ^ x104 ;
  assign n7205 = n6380 ^ n6328 ;
  assign n7206 = n7205 ^ n6342 ;
  assign n7207 = ~n6193 & n7206 ;
  assign n7204 = n6332 ^ n6328 ;
  assign n7208 = n7207 ^ n7204 ;
  assign n7209 = ~n6314 & n7208 ;
  assign n7167 = n6380 ^ n6330 ;
  assign n7168 = n7167 ^ n6303 ;
  assign n6357 = n6356 ^ n6355 ;
  assign n7169 = n7168 ^ n6357 ;
  assign n7170 = n6193 & n7169 ;
  assign n7171 = n7170 ^ n7167 ;
  assign n6322 = n6321 ^ n6299 ;
  assign n6323 = n6321 ^ n6194 ;
  assign n6324 = n6323 ^ n6321 ;
  assign n6325 = n6322 & n6324 ;
  assign n6326 = n6325 ^ n6321 ;
  assign n6327 = ~n6320 & n6326 ;
  assign n6341 = n6340 ^ n6327 ;
  assign n7197 = n7171 ^ n6341 ;
  assign n6312 = n6311 ^ n6196 ;
  assign n6313 = n6299 ^ n6198 ;
  assign n6316 = n6196 & ~n6313 ;
  assign n6317 = n6316 ^ n6198 ;
  assign n6318 = n6312 & ~n6317 ;
  assign n6319 = n6318 ^ n6311 ;
  assign n7198 = n7197 ^ n6319 ;
  assign n7199 = n7198 ^ n7196 ;
  assign n7200 = n7199 ^ n7188 ;
  assign n7201 = n7200 ^ n6310 ;
  assign n7202 = n7201 ^ n4989 ;
  assign n7172 = n7171 ^ n6299 ;
  assign n7173 = n7172 ^ n6330 ;
  assign n7174 = n7173 ^ n7171 ;
  assign n7177 = n6193 & n7174 ;
  assign n7178 = n7177 ^ n7171 ;
  assign n7179 = ~n6194 & n7178 ;
  assign n7203 = n7202 ^ n7179 ;
  assign n7210 = n7209 ^ n7203 ;
  assign n7211 = n7210 ^ x78 ;
  assign n7354 = n7353 ^ n4637 ;
  assign n7267 = n7214 & n7266 ;
  assign n7275 = n7274 ^ n7267 ;
  assign n7330 = n7329 ^ n7327 ;
  assign n7331 = ~n7212 & n7330 ;
  assign n7332 = n7331 ^ n7329 ;
  assign n7342 = n7328 & ~n7332 ;
  assign n7340 = n7339 ^ n7336 ;
  assign n7333 = n7332 ^ n7307 ;
  assign n7334 = n7333 ^ n7278 ;
  assign n7341 = n7340 ^ n7334 ;
  assign n7343 = n7342 ^ n7341 ;
  assign n7344 = ~n7323 & ~n7343 ;
  assign n7345 = n7344 ^ n7333 ;
  assign n7315 = n7307 ^ n7299 ;
  assign n7317 = n7315 ^ n7306 ;
  assign n7318 = n7306 ^ n7213 ;
  assign n7319 = n7318 ^ n7306 ;
  assign n7320 = ~n7317 & n7319 ;
  assign n7321 = n7320 ^ n7306 ;
  assign n7322 = ~n7212 & n7321 ;
  assign n7346 = n7345 ^ n7322 ;
  assign n7309 = n7308 ^ n7297 ;
  assign n7310 = n7297 ^ n7212 ;
  assign n7311 = n7310 ^ n7297 ;
  assign n7312 = ~n7309 & n7311 ;
  assign n7313 = n7312 ^ n7297 ;
  assign n7314 = n7213 & ~n7313 ;
  assign n7347 = n7346 ^ n7314 ;
  assign n7348 = n7347 ^ n7263 ;
  assign n7349 = n7348 ^ n7305 ;
  assign n7282 = n7281 ^ n7278 ;
  assign n7285 = n7263 ^ n7213 ;
  assign n7286 = n7285 ^ n7263 ;
  assign n7287 = ~n7282 & ~n7286 ;
  assign n7288 = n7287 ^ n7263 ;
  assign n7289 = n7212 & n7288 ;
  assign n7350 = n7349 ^ n7289 ;
  assign n7351 = ~n7275 & ~n7350 ;
  assign n7352 = ~n7264 & n7351 ;
  assign n7355 = n7354 ^ n7352 ;
  assign n7356 = n7355 ^ x83 ;
  assign n7357 = n7211 & ~n7356 ;
  assign n8633 = n7357 ^ n7356 ;
  assign n6920 = n5906 ^ n5893 ;
  assign n6918 = n6917 ^ n5898 ;
  assign n6919 = n6918 ^ n5827 ;
  assign n6921 = n6920 ^ n6919 ;
  assign n6922 = ~n5877 & ~n6921 ;
  assign n6923 = n6922 ^ n6920 ;
  assign n6924 = n5948 & n6923 ;
  assign n5902 = n5901 ^ n5897 ;
  assign n5907 = n5906 ^ n5902 ;
  assign n5908 = n5906 ^ n5427 ;
  assign n5909 = n5908 ^ n5906 ;
  assign n5910 = ~n5907 & ~n5909 ;
  assign n5911 = n5910 ^ n5906 ;
  assign n5912 = n5877 & n5911 ;
  assign n6914 = n5912 ^ n5427 ;
  assign n6915 = n6914 ^ n6913 ;
  assign n5940 = n5939 ^ n5427 ;
  assign n5941 = ~n5936 & ~n5940 ;
  assign n5942 = n5941 ^ n5934 ;
  assign n6916 = n6915 ^ n5942 ;
  assign n6925 = n6924 ^ n6916 ;
  assign n6901 = n6900 ^ n5940 ;
  assign n6902 = n5938 ^ n5884 ;
  assign n6905 = ~n5940 & ~n6902 ;
  assign n6906 = n6905 ^ n5938 ;
  assign n6907 = ~n6901 & n6906 ;
  assign n6926 = n6925 ^ n6907 ;
  assign n6928 = n6927 ^ n6926 ;
  assign n6929 = n6928 ^ n5963 ;
  assign n6930 = n6929 ^ n4928 ;
  assign n6898 = ~n5877 & n6897 ;
  assign n6931 = n6930 ^ n6898 ;
  assign n6932 = n6931 ^ x69 ;
  assign n6959 = n5291 & ~n5341 ;
  assign n6954 = n5346 ^ n5324 ;
  assign n6945 = ~n5122 & n5333 ;
  assign n6946 = n6945 ^ n5326 ;
  assign n6955 = n6954 ^ n6946 ;
  assign n6950 = n5329 ^ n5324 ;
  assign n6951 = n6950 ^ n5346 ;
  assign n6952 = n6951 ^ n5389 ;
  assign n6953 = n5122 & n6952 ;
  assign n6956 = n6955 ^ n6953 ;
  assign n6957 = ~n5286 & ~n6956 ;
  assign n6947 = n6946 ^ n5313 ;
  assign n6948 = n6947 ^ n6944 ;
  assign n6933 = n5340 ^ n5336 ;
  assign n6934 = n5336 ^ n5122 ;
  assign n6935 = n6934 ^ n5336 ;
  assign n6936 = ~n6933 & n6935 ;
  assign n6937 = n6936 ^ n5336 ;
  assign n6938 = n5291 & n6937 ;
  assign n6949 = n6948 ^ n6938 ;
  assign n6958 = n6957 ^ n6949 ;
  assign n6960 = n6959 ^ n6958 ;
  assign n6961 = ~n5290 & ~n6960 ;
  assign n6962 = ~n5395 & n6961 ;
  assign n6963 = n6962 ^ n4606 ;
  assign n6964 = n6963 ^ x110 ;
  assign n6965 = n6932 & ~n6964 ;
  assign n6966 = n6965 ^ n6932 ;
  assign n6967 = n6966 ^ n6964 ;
  assign n7109 = n7108 ^ n7066 ;
  assign n7110 = n7109 ^ n7092 ;
  assign n7107 = n7075 ^ n7071 ;
  assign n7111 = n7110 ^ n7107 ;
  assign n7112 = n7110 ^ n7050 ;
  assign n7113 = n7112 ^ n7110 ;
  assign n7114 = n7111 & n7113 ;
  assign n7115 = n7114 ^ n7110 ;
  assign n7116 = ~n7051 & n7115 ;
  assign n7098 = n7076 ^ n7040 ;
  assign n7100 = n7099 ^ n7098 ;
  assign n7101 = n7100 ^ n7040 ;
  assign n7104 = n7050 & n7101 ;
  assign n7105 = n7104 ^ n7040 ;
  assign n7106 = ~n7052 & n7105 ;
  assign n7117 = n7116 ^ n7106 ;
  assign n7118 = n7117 ^ n7037 ;
  assign n7119 = n7118 ^ n7097 ;
  assign n7120 = n7119 ^ n7084 ;
  assign n7053 = n7052 ^ n7049 ;
  assign n7058 = ~n7049 & ~n7050 ;
  assign n7059 = n7058 ^ n7037 ;
  assign n7060 = n7053 & n7059 ;
  assign n7121 = n7120 ^ n7060 ;
  assign n7123 = n7122 ^ n7121 ;
  assign n7126 = n7125 ^ n7123 ;
  assign n7128 = n7127 ^ n7126 ;
  assign n7129 = n7128 ^ n5550 ;
  assign n7130 = n7129 ^ x117 ;
  assign n7140 = n7139 ^ n5968 ;
  assign n7144 = n7143 ^ n7140 ;
  assign n7145 = n7144 ^ n7137 ;
  assign n7146 = n7145 ^ n5519 ;
  assign n7147 = n7146 ^ x92 ;
  assign n7148 = n7130 & n7147 ;
  assign n7387 = n6967 & n7148 ;
  assign n7149 = n7148 ^ n7147 ;
  assign n7156 = n6965 & n7149 ;
  assign n7393 = n7387 ^ n7156 ;
  assign n7153 = n7148 ^ n7130 ;
  assign n7154 = n7153 ^ n7147 ;
  assign n7371 = n6967 & ~n7154 ;
  assign n8645 = n7393 ^ n7371 ;
  assign n8646 = ~n8633 & n8645 ;
  assign n6968 = n6967 ^ n6932 ;
  assign n7157 = ~n6968 & n7153 ;
  assign n8634 = n8633 ^ n7211 ;
  assign n8638 = n7157 & n8634 ;
  assign n7384 = n6966 & ~n7154 ;
  assign n7163 = n7130 ^ n6932 ;
  assign n7379 = n7154 ^ n6964 ;
  assign n7380 = ~n7163 & ~n7379 ;
  assign n7151 = n6965 & n7148 ;
  assign n7158 = n7157 ^ n7151 ;
  assign n7159 = n7158 ^ n7156 ;
  assign n7155 = n6965 & ~n7154 ;
  assign n7160 = n7159 ^ n7155 ;
  assign n7381 = n7380 ^ n7160 ;
  assign n7378 = n6966 & n7153 ;
  assign n7382 = n7381 ^ n7378 ;
  assign n7164 = ~n6964 & ~n7163 ;
  assign n7161 = n7160 ^ n6965 ;
  assign n7162 = n7161 ^ n7157 ;
  assign n7165 = n7164 ^ n7162 ;
  assign n7150 = ~n6968 & n7149 ;
  assign n7152 = n7151 ^ n7150 ;
  assign n7166 = n7165 ^ n7152 ;
  assign n7376 = n7166 ^ n7159 ;
  assign n7374 = n6966 & n7148 ;
  assign n7375 = n7374 ^ n7155 ;
  assign n7377 = n7376 ^ n7375 ;
  assign n7383 = n7382 ^ n7377 ;
  assign n7385 = n7384 ^ n7383 ;
  assign n8637 = n7357 & n7385 ;
  assign n8639 = n8638 ^ n8637 ;
  assign n8635 = n7383 & n8634 ;
  assign n7418 = n7378 ^ n7371 ;
  assign n7407 = n6967 & n7153 ;
  assign n7417 = n7407 ^ n7374 ;
  assign n7419 = n7418 ^ n7417 ;
  assign n7420 = n7418 ^ n7356 ;
  assign n7421 = n7420 ^ n7418 ;
  assign n7422 = n7419 & ~n7421 ;
  assign n7423 = n7422 ^ n7418 ;
  assign n7424 = ~n7211 & n7423 ;
  assign n8636 = n8635 ^ n7424 ;
  assign n8640 = n8639 ^ n8636 ;
  assign n8641 = n8640 ^ n7393 ;
  assign n7360 = n7356 ^ n7211 ;
  assign n7427 = n7165 ^ n7150 ;
  assign n7428 = n7427 ^ n7387 ;
  assign n7429 = n7387 ^ n7356 ;
  assign n7430 = n7429 ^ n7387 ;
  assign n7431 = n7428 & n7430 ;
  assign n7432 = n7431 ^ n7387 ;
  assign n7433 = n7360 & n7432 ;
  assign n8642 = n8641 ^ n7433 ;
  assign n8643 = n8642 ^ n6145 ;
  assign n8626 = n7164 ^ n7155 ;
  assign n8627 = n8626 ^ n7164 ;
  assign n8630 = ~n7211 & n8627 ;
  assign n8631 = n8630 ^ n7164 ;
  assign n8632 = ~n7356 & n8631 ;
  assign n8644 = n8643 ^ n8632 ;
  assign n8647 = n8646 ^ n8644 ;
  assign n8619 = n7393 ^ n7381 ;
  assign n8618 = n7393 ^ n7378 ;
  assign n8620 = n8619 ^ n8618 ;
  assign n8621 = n8619 ^ n7356 ;
  assign n8622 = n8621 ^ n8619 ;
  assign n8623 = ~n8620 & ~n8622 ;
  assign n8624 = n8623 ^ n8619 ;
  assign n8625 = n7211 & ~n8624 ;
  assign n8648 = n8647 ^ n8625 ;
  assign n8649 = n8648 ^ x113 ;
  assign n8650 = n8617 & n8649 ;
  assign n5950 = n5949 ^ n5896 ;
  assign n5952 = n5951 ^ n5950 ;
  assign n5953 = ~n5877 & ~n5952 ;
  assign n5924 = n5923 ^ n5898 ;
  assign n5954 = n5953 ^ n5924 ;
  assign n5955 = n5948 & ~n5954 ;
  assign n5925 = n5924 ^ n5920 ;
  assign n5926 = n5925 ^ n5912 ;
  assign n5927 = n5926 ^ n5890 ;
  assign n5943 = n5942 ^ n5927 ;
  assign n5947 = n5946 ^ n5943 ;
  assign n5956 = n5955 ^ n5947 ;
  assign n5825 = n5824 ^ n5823 ;
  assign n5833 = n5832 ^ n5825 ;
  assign n5880 = n5833 & n5877 ;
  assign n5881 = n5880 ^ n5832 ;
  assign n5882 = ~n5427 & n5881 ;
  assign n5957 = n5956 ^ n5882 ;
  assign n5964 = n5957 & ~n5963 ;
  assign n5965 = n5964 ^ n4418 ;
  assign n7982 = n5965 ^ x122 ;
  assign n7979 = n5395 ^ n4531 ;
  assign n7966 = n5302 ^ n5299 ;
  assign n7964 = n5331 ^ n5316 ;
  assign n7963 = n5322 ^ n4895 ;
  assign n7965 = n7964 ^ n7963 ;
  assign n7967 = n7966 ^ n7965 ;
  assign n7968 = n7965 ^ n5286 ;
  assign n7969 = n7968 ^ n7965 ;
  assign n7970 = ~n7967 & ~n7969 ;
  assign n7971 = n7970 ^ n7965 ;
  assign n7972 = ~n5291 & n7971 ;
  assign n7973 = n7972 ^ n7965 ;
  assign n7960 = n5339 ^ n5299 ;
  assign n7961 = n7960 ^ n5315 ;
  assign n7962 = ~n5289 & ~n7961 ;
  assign n7974 = n7973 ^ n7962 ;
  assign n7959 = n4896 & ~n5288 ;
  assign n7975 = n7974 ^ n7959 ;
  assign n7976 = ~n5363 & ~n7975 ;
  assign n7977 = n7976 ^ n7771 ;
  assign n7978 = ~n6938 & n7977 ;
  assign n7980 = n7979 ^ n7978 ;
  assign n7981 = n7980 ^ x121 ;
  assign n8029 = n7982 ^ n7981 ;
  assign n8079 = n8078 ^ x74 ;
  assign n8093 = n8079 ^ n7981 ;
  assign n8108 = ~n8029 & n8093 ;
  assign n8018 = n7078 ^ n7073 ;
  assign n8019 = ~n7064 & ~n8018 ;
  assign n8013 = n7039 ^ n7035 ;
  assign n8014 = n7050 & ~n8013 ;
  assign n8006 = n7085 ^ n7047 ;
  assign n8007 = n8006 ^ n7078 ;
  assign n8008 = ~n7050 & n8007 ;
  assign n8009 = n8008 ^ n7085 ;
  assign n8012 = n8009 ^ n7044 ;
  assign n8015 = n8014 ^ n8012 ;
  assign n8016 = ~n7051 & n8015 ;
  assign n8010 = n8009 ^ n7125 ;
  assign n8011 = n8010 ^ n8005 ;
  assign n8017 = n8016 ^ n8011 ;
  assign n8020 = n8019 ^ n8017 ;
  assign n7994 = n7034 & n7050 ;
  assign n7999 = n7041 & n7051 ;
  assign n8000 = n7999 ^ n7028 ;
  assign n8001 = n7994 & n8000 ;
  assign n8021 = n8020 ^ n8001 ;
  assign n7993 = n7046 & n7062 ;
  assign n8022 = n8021 ^ n7993 ;
  assign n7988 = n7051 ^ n7040 ;
  assign n7989 = n7988 ^ n7040 ;
  assign n7990 = n7098 & ~n7989 ;
  assign n7991 = n7990 ^ n7040 ;
  assign n7992 = ~n7050 & n7991 ;
  assign n8023 = n8022 ^ n7992 ;
  assign n8024 = n8023 ^ n7122 ;
  assign n8025 = n8024 ^ n4489 ;
  assign n7987 = n7064 & n7986 ;
  assign n8026 = n8025 ^ n7987 ;
  assign n8027 = n8026 ^ x112 ;
  assign n8109 = n8093 ^ n8027 ;
  assign n8110 = ~n8108 & n8109 ;
  assign n8085 = ~n7982 & n8079 ;
  assign n8086 = n8027 & n8085 ;
  assign n8111 = n8110 ^ n8086 ;
  assign n8083 = n8079 ^ n7982 ;
  assign n8084 = ~n8027 & ~n8083 ;
  assign n8087 = n8086 ^ n8084 ;
  assign n8028 = n8027 ^ n7981 ;
  assign n8030 = ~n8027 & n8029 ;
  assign n8080 = n8079 ^ n8030 ;
  assign n8081 = n8028 & n8080 ;
  assign n8082 = n8081 ^ n8029 ;
  assign n8088 = n8087 ^ n8082 ;
  assign n7983 = n7981 & n7982 ;
  assign n8089 = n8088 ^ n7983 ;
  assign n8112 = n8111 ^ n8089 ;
  assign n8103 = n8029 ^ n8027 ;
  assign n8104 = n8027 ^ n7982 ;
  assign n8105 = n8103 & ~n8104 ;
  assign n8106 = n8105 ^ n7981 ;
  assign n8107 = ~n8079 & n8106 ;
  assign n7957 = n7956 ^ x97 ;
  assign n8665 = n8107 ^ n7957 ;
  assign n6806 = n6742 & n6805 ;
  assign n6807 = n6806 ^ n6803 ;
  assign n6812 = n6811 ^ n6807 ;
  assign n6774 = n6773 ^ n6756 ;
  assign n6775 = n6773 ^ n6660 ;
  assign n6776 = n6775 ^ n6773 ;
  assign n6777 = n6774 & ~n6776 ;
  assign n6778 = n6777 ^ n6773 ;
  assign n6779 = ~n6745 & ~n6778 ;
  assign n6813 = n6812 ^ n6779 ;
  assign n6788 = n6768 ^ n6754 ;
  assign n6789 = n6754 ^ n6660 ;
  assign n6790 = n6789 ^ n6754 ;
  assign n6791 = n6788 & ~n6790 ;
  assign n6792 = n6791 ^ n6754 ;
  assign n6793 = ~n6787 & n6792 ;
  assign n6814 = n6813 ^ n6793 ;
  assign n6815 = n6814 ^ n4359 ;
  assign n6781 = n6780 ^ n6779 ;
  assign n6741 = n6740 ^ n6738 ;
  assign n6782 = n6781 ^ n6741 ;
  assign n6783 = n6782 ^ n6779 ;
  assign n6784 = n6660 & ~n6783 ;
  assign n6785 = n6784 ^ n6781 ;
  assign n6786 = n6626 & n6785 ;
  assign n6816 = n6815 ^ n6786 ;
  assign n7958 = n6816 ^ x115 ;
  assign n8666 = n8665 ^ n7958 ;
  assign n8667 = n8666 ^ n8665 ;
  assign n8668 = n8112 & n8667 ;
  assign n8669 = n8668 ^ n7957 ;
  assign n8655 = n8108 ^ n8103 ;
  assign n8656 = n8655 ^ n8030 ;
  assign n8095 = n8079 ^ n8027 ;
  assign n8657 = n8656 ^ n8095 ;
  assign n8670 = ~n8028 & n8657 ;
  assign n8671 = n8670 ^ n8095 ;
  assign n8674 = n8667 & n8671 ;
  assign n8672 = n8671 ^ n8665 ;
  assign n8675 = n8674 ^ n8672 ;
  assign n8676 = n7957 & n8675 ;
  assign n8677 = n8669 & n8676 ;
  assign n8678 = n8677 ^ n8674 ;
  assign n8679 = n8678 ^ n8672 ;
  assign n8680 = n8679 ^ n7258 ;
  assign n8653 = n7958 ^ n7957 ;
  assign n8654 = n8111 ^ n8084 ;
  assign n8658 = n8657 ^ n8654 ;
  assign n8094 = n8093 ^ n7982 ;
  assign n8098 = n8093 ^ n8029 ;
  assign n8099 = ~n8095 & n8098 ;
  assign n8100 = n8099 ^ n8029 ;
  assign n8101 = n8094 & n8100 ;
  assign n8102 = n8101 ^ n8029 ;
  assign n8659 = n8658 ^ n8102 ;
  assign n8660 = n8658 ^ n7957 ;
  assign n8661 = n8660 ^ n8658 ;
  assign n8662 = ~n8659 & ~n8661 ;
  assign n8663 = n8662 ^ n8658 ;
  assign n8664 = n8653 & ~n8663 ;
  assign n8681 = n8680 ^ n8664 ;
  assign n8682 = n8681 ^ x66 ;
  assign n8684 = n6963 ^ x118 ;
  assign n8687 = n8158 ^ x84 ;
  assign n8725 = n7355 ^ x77 ;
  assign n8726 = n8687 & ~n8725 ;
  assign n8719 = n6538 & n6586 ;
  assign n8709 = n6601 ^ n6581 ;
  assign n8710 = n8709 ^ n6556 ;
  assign n8711 = n8710 ^ n6506 ;
  assign n8712 = n8711 ^ n6601 ;
  assign n8713 = ~n6537 & n8712 ;
  assign n8714 = n8713 ^ n8709 ;
  assign n8715 = n6536 & ~n8714 ;
  assign n8691 = n6558 ^ n6545 ;
  assign n8692 = n8691 ^ n7923 ;
  assign n8693 = ~n6536 & ~n8692 ;
  assign n8694 = n8693 ^ n6545 ;
  assign n8716 = n8715 ^ n8694 ;
  assign n8703 = n6565 ^ n6537 ;
  assign n8704 = n6537 ^ n6503 ;
  assign n8705 = n8704 ^ n6537 ;
  assign n8706 = ~n8703 & n8705 ;
  assign n8707 = n8706 ^ n6537 ;
  assign n8708 = n6550 & n8707 ;
  assign n8717 = n8716 ^ n8708 ;
  assign n8697 = n7451 ^ n6507 ;
  assign n8698 = n8697 ^ n6586 ;
  assign n7458 = n6594 ^ n6548 ;
  assign n8699 = n8698 ^ n7458 ;
  assign n8700 = ~n6537 & n8699 ;
  assign n8695 = n8694 ^ n6507 ;
  assign n8696 = n8695 ^ n7458 ;
  assign n8701 = n8700 ^ n8696 ;
  assign n8702 = n6565 & n8701 ;
  assign n8718 = n8717 ^ n8702 ;
  assign n8720 = n8719 ^ n8718 ;
  assign n8721 = ~n7949 & ~n8720 ;
  assign n7460 = n6568 ^ n6566 ;
  assign n7461 = n6538 & n7460 ;
  assign n8688 = n7461 ^ n6610 ;
  assign n8689 = n8688 ^ n6562 ;
  assign n8690 = n8689 ^ n4732 ;
  assign n8722 = n8721 ^ n8690 ;
  assign n8723 = n8722 ^ x75 ;
  assign n8748 = n6747 & n6804 ;
  assign n8744 = n8484 ^ n6807 ;
  assign n8734 = n6769 ^ n6740 ;
  assign n8743 = n8734 ^ n6737 ;
  assign n8745 = n8744 ^ n8743 ;
  assign n8746 = n8745 ^ n6793 ;
  assign n8735 = n8734 ^ n6795 ;
  assign n8736 = n8735 ^ n6750 ;
  assign n8737 = n8736 ^ n8734 ;
  assign n8738 = n8734 ^ n6626 ;
  assign n8739 = n8738 ^ n8734 ;
  assign n8740 = n8737 & ~n8739 ;
  assign n8741 = n8740 ^ n8734 ;
  assign n8742 = ~n6787 & n8741 ;
  assign n8747 = n8746 ^ n8742 ;
  assign n8749 = n8748 ^ n8747 ;
  assign n8729 = n6737 ^ n6660 ;
  assign n8730 = n8729 ^ n6737 ;
  assign n8731 = ~n8453 & n8730 ;
  assign n8732 = n8731 ^ n6737 ;
  assign n8733 = n6626 & n8732 ;
  assign n8750 = n8749 ^ n8733 ;
  assign n8751 = n8750 ^ n7527 ;
  assign n8752 = ~n7549 & ~n8751 ;
  assign n8753 = n8752 ^ n4766 ;
  assign n8754 = n8753 ^ x94 ;
  assign n8755 = n8723 & ~n8754 ;
  assign n8756 = n8755 ^ n8723 ;
  assign n8798 = n8726 & n8756 ;
  assign n8683 = n8189 ^ x101 ;
  assign n8838 = n8798 ^ n8683 ;
  assign n8839 = ~n8684 & n8838 ;
  assign n8685 = n8683 & ~n8684 ;
  assign n8686 = n8685 ^ n8683 ;
  assign n8762 = n8726 ^ n8687 ;
  assign n8807 = n8756 & n8762 ;
  assign n8757 = n8756 ^ n8754 ;
  assign n8761 = n8726 & n8757 ;
  assign n8808 = n8807 ^ n8761 ;
  assign n8834 = n8686 & n8808 ;
  assign n8724 = n8687 & ~n8723 ;
  assign n8774 = n8724 ^ n8723 ;
  assign n8775 = n8774 ^ n8687 ;
  assign n8767 = n8726 ^ n8725 ;
  assign n8768 = n8756 & ~n8767 ;
  assign n8763 = n8762 ^ n8725 ;
  assign n8766 = n8755 & n8763 ;
  assign n8769 = n8768 ^ n8766 ;
  assign n8765 = n8756 & n8763 ;
  assign n8770 = n8769 ^ n8765 ;
  assign n8776 = n8775 ^ n8770 ;
  assign n8772 = n8757 & ~n8767 ;
  assign n8773 = n8772 ^ n8765 ;
  assign n8777 = n8776 ^ n8773 ;
  assign n8778 = n8777 ^ n8766 ;
  assign n8771 = n8770 ^ n8767 ;
  assign n8779 = n8778 ^ n8771 ;
  assign n8764 = n8757 & n8763 ;
  assign n8780 = n8779 ^ n8764 ;
  assign n8781 = n8780 ^ n8772 ;
  assign n8782 = n8781 ^ n8774 ;
  assign n8832 = n8782 ^ n8776 ;
  assign n8833 = n8686 & n8832 ;
  assign n8835 = n8834 ^ n8833 ;
  assign n8821 = n8778 ^ n8684 ;
  assign n8822 = n8821 ^ n8778 ;
  assign n8823 = ~n8765 & n8781 ;
  assign n8824 = n8823 ^ n8778 ;
  assign n8825 = n8822 & ~n8824 ;
  assign n8826 = n8825 ^ n8778 ;
  assign n8827 = ~n8683 & ~n8826 ;
  assign n8828 = n8827 ^ n8683 ;
  assign n8790 = n8685 ^ n8684 ;
  assign n8797 = n8790 ^ n8686 ;
  assign n8758 = n8757 ^ n8723 ;
  assign n8759 = n8726 & ~n8758 ;
  assign n8760 = n8759 ^ n8724 ;
  assign n8806 = n8762 ^ n8760 ;
  assign n8809 = n8808 ^ n8806 ;
  assign n8817 = n8809 ^ n8798 ;
  assign n8818 = n8817 ^ n8807 ;
  assign n8816 = n8775 ^ n8723 ;
  assign n8819 = n8818 ^ n8816 ;
  assign n8820 = n8797 & n8819 ;
  assign n8829 = n8828 ^ n8820 ;
  assign n8783 = n8782 ^ n8779 ;
  assign n8813 = n8783 ^ n8769 ;
  assign n8814 = n8813 ^ n8807 ;
  assign n8815 = n8685 & ~n8814 ;
  assign n8830 = n8829 ^ n8815 ;
  assign n8810 = ~n8683 & n8809 ;
  assign n8784 = n8759 ^ n8758 ;
  assign n8785 = n8784 ^ n8783 ;
  assign n8786 = n8785 ^ n8761 ;
  assign n8787 = n8786 ^ n8760 ;
  assign n8799 = n8798 ^ n8787 ;
  assign n8800 = n8799 ^ n8785 ;
  assign n8801 = n8785 ^ n8684 ;
  assign n8802 = n8801 ^ n8785 ;
  assign n8803 = n8800 & n8802 ;
  assign n8804 = n8803 ^ n8785 ;
  assign n8805 = n8797 & n8804 ;
  assign n8811 = n8810 ^ n8805 ;
  assign n8812 = n8811 ^ n8683 ;
  assign n8831 = n8830 ^ n8812 ;
  assign n8836 = n8835 ^ n8831 ;
  assign n8837 = n8836 ^ n7242 ;
  assign n8840 = n8839 ^ n8837 ;
  assign n8788 = n8787 ^ n8759 ;
  assign n8789 = n8788 ^ n8686 ;
  assign n8791 = n8790 ^ n8773 ;
  assign n8792 = n8773 ^ n8686 ;
  assign n8793 = n8792 ^ n8773 ;
  assign n8794 = n8791 & ~n8793 ;
  assign n8795 = n8794 ^ n8773 ;
  assign n8796 = n8789 & ~n8795 ;
  assign n8841 = n8840 ^ n8796 ;
  assign n8842 = n8841 ^ x65 ;
  assign n8843 = ~n8682 & ~n8842 ;
  assign n8849 = n8650 & n8843 ;
  assign n10570 = n8849 ^ n8843 ;
  assign n8651 = n8650 ^ n8617 ;
  assign n8652 = n8651 ^ n8649 ;
  assign n8856 = ~n8652 & n8843 ;
  assign n8846 = n8650 ^ n8649 ;
  assign n8847 = n8843 & n8846 ;
  assign n8857 = n8856 ^ n8847 ;
  assign n10571 = n10570 ^ n8857 ;
  assign n8844 = n8843 ^ n8682 ;
  assign n8921 = n8844 ^ n8842 ;
  assign n8922 = n8650 & ~n8921 ;
  assign n8923 = n8922 ^ n8921 ;
  assign n8909 = n8682 ^ n8649 ;
  assign n8910 = n8909 ^ n8842 ;
  assign n8911 = n8617 & n8910 ;
  assign n8912 = n8911 ^ n8910 ;
  assign n8858 = n8857 ^ n8652 ;
  assign n8850 = n8842 ^ n8649 ;
  assign n8851 = n8682 ^ n8617 ;
  assign n8852 = ~n8842 & n8851 ;
  assign n8853 = n8852 ^ n8617 ;
  assign n8854 = n8850 & ~n8853 ;
  assign n8855 = n8854 ^ n8849 ;
  assign n8859 = n8858 ^ n8855 ;
  assign n8845 = ~n8652 & ~n8844 ;
  assign n8848 = n8847 ^ n8845 ;
  assign n8860 = n8859 ^ n8848 ;
  assign n8913 = n8912 ^ n8860 ;
  assign n8861 = n8860 ^ n8858 ;
  assign n8914 = n8913 ^ n8861 ;
  assign n8924 = n8923 ^ n8914 ;
  assign n8920 = n8650 & ~n8844 ;
  assign n8925 = n8924 ^ n8920 ;
  assign n10831 = n10571 ^ n8925 ;
  assign n8949 = n8911 ^ n8617 ;
  assign n10845 = n10831 ^ n8949 ;
  assign n8915 = n8914 ^ n8845 ;
  assign n8916 = n8915 ^ n8617 ;
  assign n8908 = n8852 ^ n8843 ;
  assign n8917 = n8916 ^ n8908 ;
  assign n10547 = n8917 ^ n8849 ;
  assign n10548 = n10547 ^ n8915 ;
  assign n8926 = n8925 ^ n8911 ;
  assign n10546 = n8926 ^ n8842 ;
  assign n10549 = n10548 ^ n10546 ;
  assign n10572 = n10571 ^ n10549 ;
  assign n10569 = n8924 ^ n8651 ;
  assign n10573 = n10572 ^ n10569 ;
  assign n10846 = n10845 ^ n10573 ;
  assign n10847 = n10846 ^ n8922 ;
  assign n10848 = ~n8899 & ~n10847 ;
  assign n8905 = n8580 & n8898 ;
  assign n8906 = n8905 ^ n8580 ;
  assign n8907 = n8906 ^ n8898 ;
  assign n10839 = ~n8907 & n8924 ;
  assign n10832 = n10831 ^ n8651 ;
  assign n10833 = n10832 ^ n10831 ;
  assign n10834 = n10831 ^ n8580 ;
  assign n10835 = n10834 ^ n10831 ;
  assign n10836 = n10833 & ~n10835 ;
  assign n10837 = n10836 ^ n10831 ;
  assign n10838 = n8899 & n10837 ;
  assign n10840 = n10839 ^ n10838 ;
  assign n10585 = n10549 ^ n8898 ;
  assign n10586 = n10585 ^ n10549 ;
  assign n10587 = ~n10572 & n10586 ;
  assign n10588 = n10587 ^ n10549 ;
  assign n10589 = n8899 & ~n10588 ;
  assign n10841 = n10840 ^ n10589 ;
  assign n8935 = n8917 ^ n8859 ;
  assign n8936 = n8935 ^ n8847 ;
  assign n8937 = n8936 ^ n8856 ;
  assign n8938 = n8937 ^ n8916 ;
  assign n8939 = n8938 ^ n8906 ;
  assign n8940 = n8907 ^ n8580 ;
  assign n8941 = n8940 ^ n8861 ;
  assign n8944 = ~n8938 & ~n8941 ;
  assign n8945 = n8944 ^ n8861 ;
  assign n8946 = ~n8939 & ~n8945 ;
  assign n8947 = n8946 ^ n8906 ;
  assign n10842 = n10841 ^ n8947 ;
  assign n10843 = n10842 ^ n8078 ;
  assign n10827 = n8856 ^ n8845 ;
  assign n10828 = n10827 ^ n8920 ;
  assign n10829 = n10828 ^ n8912 ;
  assign n10830 = n8905 & n10829 ;
  assign n10844 = n10843 ^ n10830 ;
  assign n10849 = n10848 ^ n10844 ;
  assign n10826 = ~n8907 & ~n8937 ;
  assign n10850 = n10849 ^ n10826 ;
  assign n10821 = n8915 ^ n8580 ;
  assign n10822 = n10821 ^ n8915 ;
  assign n10823 = ~n10548 & n10822 ;
  assign n10824 = n10823 ^ n8915 ;
  assign n10825 = n8899 & ~n10824 ;
  assign n10851 = n10850 ^ n10825 ;
  assign n10852 = n10851 ^ x75 ;
  assign n8113 = n8112 ^ n8107 ;
  assign n8114 = n8113 ^ n8102 ;
  assign n8092 = n8087 ^ n8085 ;
  assign n8115 = n8114 ^ n8092 ;
  assign n8118 = n8115 ^ n8105 ;
  assign n8119 = n8118 ^ n8115 ;
  assign n8120 = ~n8110 & ~n8119 ;
  assign n8121 = n8120 ^ n8115 ;
  assign n8122 = ~n7958 & n8121 ;
  assign n8123 = n8122 ^ n8115 ;
  assign n8090 = n7958 & n8089 ;
  assign n8091 = n8090 ^ n8082 ;
  assign n8124 = n8123 ^ n8091 ;
  assign n8125 = ~n7957 & ~n8124 ;
  assign n8126 = n8125 ^ n8123 ;
  assign n8127 = n8126 ^ n7957 ;
  assign n8128 = n8127 ^ n8123 ;
  assign n8129 = n8128 ^ n8091 ;
  assign n8130 = n8129 ^ n4573 ;
  assign n8131 = n8130 ^ x85 ;
  assign n8322 = ~n8253 & n8284 ;
  assign n8323 = n8322 ^ n6192 ;
  assign n8305 = n8252 ^ n8234 ;
  assign n8307 = n8306 ^ n8305 ;
  assign n8308 = n8307 ^ n8252 ;
  assign n8309 = n8252 ^ n8159 ;
  assign n8310 = n8309 ^ n8252 ;
  assign n8311 = n8308 & ~n8310 ;
  assign n8312 = n8311 ^ n8252 ;
  assign n8313 = n8271 & ~n8312 ;
  assign n8314 = n8313 ^ n8252 ;
  assign n8299 = n8298 ^ n8278 ;
  assign n8300 = n8278 ^ n8271 ;
  assign n8301 = n8300 ^ n8278 ;
  assign n8302 = ~n8299 & ~n8301 ;
  assign n8303 = n8302 ^ n8278 ;
  assign n8304 = n8159 & n8303 ;
  assign n8315 = n8314 ^ n8304 ;
  assign n8289 = n8260 ^ n8253 ;
  assign n8290 = n8289 ^ n8285 ;
  assign n8291 = n8237 ^ n8234 ;
  assign n8287 = n8286 ^ n8271 ;
  assign n8292 = n8291 ^ n8287 ;
  assign n8293 = n8291 ^ n8289 ;
  assign n8294 = n8293 ^ n8291 ;
  assign n8295 = ~n8292 & ~n8294 ;
  assign n8296 = n8295 ^ n8291 ;
  assign n8297 = n8290 & ~n8296 ;
  assign n8316 = n8315 ^ n8297 ;
  assign n8288 = n8257 & n8287 ;
  assign n8317 = n8316 ^ n8288 ;
  assign n8320 = n8319 ^ n8317 ;
  assign n8321 = ~n8283 & n8320 ;
  assign n8324 = n8323 ^ n8321 ;
  assign n8325 = n8324 ^ x102 ;
  assign n5398 = n5397 ^ x88 ;
  assign n5966 = n5965 ^ x114 ;
  assign n5967 = n5398 & ~n5966 ;
  assign n6625 = n6624 ^ x120 ;
  assign n6817 = n6816 ^ x64 ;
  assign n6818 = n6625 & n6817 ;
  assign n6820 = n6818 ^ n6817 ;
  assign n6821 = n6820 ^ n6625 ;
  assign n6822 = n6821 ^ n6817 ;
  assign n6162 = n6112 ^ n5187 ;
  assign n6152 = n6102 & ~n6146 ;
  assign n6153 = n6152 ^ n6101 ;
  assign n6163 = n6162 ^ n6153 ;
  assign n6154 = n6153 ^ n6146 ;
  assign n6155 = n6154 ^ n6153 ;
  assign n6159 = n6155 & n6156 ;
  assign n6160 = n6159 ^ n6153 ;
  assign n6161 = ~n5968 & ~n6160 ;
  assign n6164 = n6163 ^ n6161 ;
  assign n6113 = n6112 ^ n6078 ;
  assign n6114 = n6113 ^ n6112 ;
  assign n6149 = n6114 & ~n6146 ;
  assign n6150 = n6149 ^ n6112 ;
  assign n6151 = ~n5968 & n6150 ;
  assign n6165 = n6164 ^ n6151 ;
  assign n6166 = n6165 ^ x82 ;
  assign n6358 = n6357 ^ n6333 ;
  assign n6359 = ~n6193 & n6358 ;
  assign n6360 = n6359 ^ n6355 ;
  assign n6367 = n6366 ^ n6360 ;
  assign n6364 = n6330 ^ n6303 ;
  assign n6368 = n6367 ^ n6364 ;
  assign n6369 = n6368 ^ n6360 ;
  assign n6370 = ~n6193 & n6369 ;
  assign n6371 = n6370 ^ n6367 ;
  assign n6372 = ~n6194 & n6371 ;
  assign n6362 = n6193 & n6350 ;
  assign n6352 = n6351 ^ n6350 ;
  assign n6353 = n6352 ^ n6303 ;
  assign n6354 = n6194 & n6353 ;
  assign n6361 = n6360 ^ n6354 ;
  assign n6363 = n6362 ^ n6361 ;
  assign n6373 = n6372 ^ n6363 ;
  assign n6375 = n6374 ^ n6373 ;
  assign n6376 = n6375 ^ n6349 ;
  assign n6377 = n6376 ^ n6341 ;
  assign n6378 = n6377 ^ n6319 ;
  assign n6393 = n6392 ^ n6378 ;
  assign n6394 = ~n6310 & ~n6393 ;
  assign n6395 = n6394 ^ n5166 ;
  assign n6396 = n6395 ^ x81 ;
  assign n6397 = n6166 & n6396 ;
  assign n6825 = n6397 ^ n6166 ;
  assign n6828 = n6825 ^ n6396 ;
  assign n6829 = n6828 ^ n6166 ;
  assign n6836 = n6822 & n6829 ;
  assign n6834 = n6822 & n6825 ;
  assign n6830 = ~n6821 & n6829 ;
  assign n6831 = n6830 ^ n6821 ;
  assign n6826 = ~n6821 & n6825 ;
  assign n6824 = n6397 & ~n6821 ;
  assign n6827 = n6826 ^ n6824 ;
  assign n6832 = n6831 ^ n6827 ;
  assign n6835 = n6834 ^ n6832 ;
  assign n6837 = n6836 ^ n6835 ;
  assign n6838 = n6837 ^ n6822 ;
  assign n6823 = n6397 & n6822 ;
  assign n6833 = n6832 ^ n6823 ;
  assign n6839 = n6838 ^ n6833 ;
  assign n6819 = n6397 & n6818 ;
  assign n6840 = n6839 ^ n6819 ;
  assign n6841 = n5967 & n6840 ;
  assign n6850 = n5967 ^ n5398 ;
  assign n6851 = n6819 & n6850 ;
  assign n6842 = n6397 & n6820 ;
  assign n6843 = n6842 ^ n6830 ;
  assign n6844 = n6843 ^ n6819 ;
  assign n6845 = n6843 ^ n5966 ;
  assign n6846 = n6845 ^ n6843 ;
  assign n6847 = n6844 & n6846 ;
  assign n6848 = n6847 ^ n6843 ;
  assign n6849 = ~n5398 & n6848 ;
  assign n6852 = n6851 ^ n6849 ;
  assign n6861 = n6818 & n6825 ;
  assign n6886 = n6850 ^ n5966 ;
  assign n6887 = n6861 & n6886 ;
  assign n6860 = n5966 ^ n5398 ;
  assign n6854 = n6818 & ~n6828 ;
  assign n6874 = n6854 ^ n6839 ;
  assign n6873 = n6832 ^ n6828 ;
  assign n6875 = n6874 ^ n6873 ;
  assign n6880 = n6875 ^ n6820 ;
  assign n6867 = n6820 & n6829 ;
  assign n6879 = n6867 ^ n6842 ;
  assign n6881 = n6880 ^ n6879 ;
  assign n6882 = n6860 & n6881 ;
  assign n6866 = n6832 ^ n6824 ;
  assign n6868 = n6867 ^ n6866 ;
  assign n6883 = n6882 ^ n6868 ;
  assign n6876 = n6875 ^ n6826 ;
  assign n6872 = n6843 ^ n6836 ;
  assign n6877 = n6876 ^ n6872 ;
  assign n6878 = n6850 & n6877 ;
  assign n6884 = n6883 ^ n6878 ;
  assign n6869 = n6868 ^ n6823 ;
  assign n6862 = n6861 ^ n6836 ;
  assign n6863 = n6862 ^ n6854 ;
  assign n6864 = n6863 ^ n6835 ;
  assign n6865 = ~n5398 & ~n6864 ;
  assign n6870 = n6869 ^ n6865 ;
  assign n6871 = ~n6860 & ~n6870 ;
  assign n6885 = n6884 ^ n6871 ;
  assign n6888 = n6887 ^ n6885 ;
  assign n6858 = n6818 & n6829 ;
  assign n6859 = n5967 & n6858 ;
  assign n6889 = n6888 ^ n6859 ;
  assign n6855 = n6854 ^ n6834 ;
  assign n6856 = n5966 & n6855 ;
  assign n6853 = n5398 & n6834 ;
  assign n6857 = n6856 ^ n6853 ;
  assign n6890 = n6889 ^ n6857 ;
  assign n6891 = ~n6852 & n6890 ;
  assign n6892 = ~n6841 & n6891 ;
  assign n6893 = n6892 ^ n6224 ;
  assign n6894 = n6893 ^ x124 ;
  assign n7358 = n7357 ^ n7211 ;
  assign n7359 = n7166 & n7358 ;
  assign n7363 = n7155 ^ n7150 ;
  assign n7361 = n6966 & n7149 ;
  assign n7362 = n7361 ^ n7150 ;
  assign n7364 = n7363 ^ n7362 ;
  assign n7365 = n7363 ^ n7356 ;
  assign n7366 = n7365 ^ n7363 ;
  assign n7367 = n7364 & ~n7366 ;
  assign n7368 = n7367 ^ n7363 ;
  assign n7369 = n7360 & n7368 ;
  assign n7370 = n7369 ^ n7150 ;
  assign n7415 = n7155 & ~n7360 ;
  assign n7404 = n7165 ^ n6968 ;
  assign n7405 = n7404 ^ n7158 ;
  assign n7406 = n7405 ^ n7162 ;
  assign n7408 = n7407 ^ n7406 ;
  assign n7409 = n7408 ^ n7361 ;
  assign n7410 = ~n7211 & ~n7409 ;
  assign n7403 = n7378 ^ n7162 ;
  assign n7411 = n7410 ^ n7403 ;
  assign n7412 = n7356 & n7411 ;
  assign n7386 = n7385 ^ n7374 ;
  assign n7388 = n7387 ^ n7386 ;
  assign n7373 = n7159 ^ n7150 ;
  assign n7389 = n7388 ^ n7373 ;
  assign n7390 = ~n7356 & n7389 ;
  assign n7391 = n7390 ^ n7388 ;
  assign n7401 = n7391 ^ n7378 ;
  assign n7392 = n7391 ^ n7384 ;
  assign n7394 = n7393 ^ n7392 ;
  assign n7395 = n7394 ^ n7391 ;
  assign n7398 = ~n7356 & n7395 ;
  assign n7399 = n7398 ^ n7391 ;
  assign n7400 = ~n7211 & n7399 ;
  assign n7402 = n7401 ^ n7400 ;
  assign n7413 = n7412 ^ n7402 ;
  assign n7372 = n7357 & n7371 ;
  assign n7414 = n7413 ^ n7372 ;
  assign n7416 = n7415 ^ n7414 ;
  assign n7425 = ~n7416 & ~n7424 ;
  assign n7426 = ~n7370 & n7425 ;
  assign n7434 = n7426 & ~n7433 ;
  assign n7435 = ~n7359 & n7434 ;
  assign n7436 = n7435 ^ n6294 ;
  assign n7437 = n7436 ^ x78 ;
  assign n7438 = n6894 & n7437 ;
  assign n7913 = n7438 ^ n7437 ;
  assign n7597 = n7596 ^ x85 ;
  assign n7439 = n6931 ^ x67 ;
  assign n7626 = n7597 ^ n7439 ;
  assign n7453 = n7452 ^ n7451 ;
  assign n7454 = n6537 & ~n6565 ;
  assign n7455 = n7453 & n7454 ;
  assign n7456 = n7455 ^ n6565 ;
  assign n7459 = ~n7456 & n7458 ;
  assign n7464 = n6539 & ~n6558 ;
  assign n7465 = n7459 & n7464 ;
  assign n7462 = n7461 ^ n7459 ;
  assign n7463 = n7462 ^ n7455 ;
  assign n7466 = n7465 ^ n7463 ;
  assign n7449 = n6582 ^ n6542 ;
  assign n7450 = n6563 & n7449 ;
  assign n7467 = n7466 ^ n7450 ;
  assign n7442 = n6588 ^ n6468 ;
  assign n7443 = n7442 ^ n6591 ;
  assign n7444 = n6591 ^ n6537 ;
  assign n7445 = n7444 ^ n6591 ;
  assign n7446 = n7443 & n7445 ;
  assign n7447 = n7446 ^ n6591 ;
  assign n7448 = ~n6536 & ~n7447 ;
  assign n7468 = n7467 ^ n7448 ;
  assign n7469 = ~n6607 & ~n7468 ;
  assign n7470 = ~n7441 & n7469 ;
  assign n7471 = ~n6610 & n7470 ;
  assign n7472 = ~n6621 & n7471 ;
  assign n7473 = n7472 ^ n5020 ;
  assign n7474 = n7473 ^ x116 ;
  assign n7475 = n7210 ^ x68 ;
  assign n7476 = n7474 & n7475 ;
  assign n7509 = n7508 ^ n7275 ;
  assign n7493 = n7492 ^ n7338 ;
  assign n7494 = n7493 ^ n7282 ;
  assign n7495 = n7212 & n7494 ;
  assign n7496 = n7495 ^ n7492 ;
  assign n7510 = n7509 ^ n7496 ;
  assign n7491 = n7332 ^ n7262 ;
  assign n7497 = n7496 ^ n7491 ;
  assign n7498 = n7497 ^ n7336 ;
  assign n7499 = n7498 ^ n7262 ;
  assign n7500 = n7499 ^ n7497 ;
  assign n7501 = n7497 ^ n7213 ;
  assign n7502 = n7501 ^ n7497 ;
  assign n7503 = n7500 & n7502 ;
  assign n7504 = n7503 ^ n7497 ;
  assign n7505 = n7323 & ~n7504 ;
  assign n7511 = n7510 ^ n7505 ;
  assign n7489 = n7266 ^ n7263 ;
  assign n7490 = ~n7215 & n7489 ;
  assign n7512 = n7511 ^ n7490 ;
  assign n7488 = n7216 & n7327 ;
  assign n7513 = n7512 ^ n7488 ;
  assign n7514 = n7262 ^ n7214 ;
  assign n7515 = n7514 ^ n7513 ;
  assign n7516 = n7307 ^ n7213 ;
  assign n7517 = ~n7214 & ~n7516 ;
  assign n7518 = n7517 ^ n7307 ;
  assign n7519 = ~n7515 & ~n7518 ;
  assign n7520 = n7519 ^ n7214 ;
  assign n7521 = n7513 & ~n7520 ;
  assign n7522 = ~n7487 & n7521 ;
  assign n7523 = ~n7485 & n7522 ;
  assign n7524 = ~n7296 & n7523 ;
  assign n7525 = n7524 ^ n4954 ;
  assign n7526 = n7525 ^ x102 ;
  assign n7552 = n7551 ^ x109 ;
  assign n7553 = n7526 & n7552 ;
  assign n7554 = n7553 ^ n7526 ;
  assign n7555 = n7554 ^ n7552 ;
  assign n7606 = n7476 & ~n7555 ;
  assign n7477 = n7476 ^ n7475 ;
  assign n7556 = n7555 ^ n7526 ;
  assign n7557 = n7477 & n7556 ;
  assign n7610 = n7606 ^ n7557 ;
  assign n7561 = n7477 ^ n7474 ;
  assign n7563 = n7561 ^ n7475 ;
  assign n7568 = ~n7555 & n7563 ;
  assign n7567 = n7553 & n7563 ;
  assign n7569 = n7568 ^ n7567 ;
  assign n7565 = n7556 & n7563 ;
  assign n7562 = ~n7555 & ~n7561 ;
  assign n7566 = n7565 ^ n7562 ;
  assign n7570 = n7569 ^ n7566 ;
  assign n7564 = n7563 ^ n7562 ;
  assign n7571 = n7570 ^ n7564 ;
  assign n7572 = n7571 ^ n7565 ;
  assign n7611 = n7610 ^ n7572 ;
  assign n7575 = n7554 & ~n7561 ;
  assign n7576 = n7575 ^ n7568 ;
  assign n7608 = n7576 ^ n7566 ;
  assign n7609 = n7608 ^ n7552 ;
  assign n7612 = n7611 ^ n7609 ;
  assign n7633 = n7612 ^ n7569 ;
  assign n7615 = n7476 & n7556 ;
  assign n7613 = n7612 ^ n7477 ;
  assign n7604 = n7477 & n7553 ;
  assign n7614 = n7613 ^ n7604 ;
  assign n7616 = n7615 ^ n7614 ;
  assign n7607 = n7606 ^ n7476 ;
  assign n7617 = n7616 ^ n7607 ;
  assign n7627 = n7617 ^ n7614 ;
  assign n7628 = n7627 ^ n7612 ;
  assign n7629 = n7627 ^ n7439 ;
  assign n7630 = n7626 & n7629 ;
  assign n7631 = n7630 ^ n7439 ;
  assign n7632 = ~n7628 & ~n7631 ;
  assign n7634 = n7633 ^ n7632 ;
  assign n7635 = n7634 ^ n7616 ;
  assign n7636 = n7635 ^ n7611 ;
  assign n7637 = n7636 ^ n7634 ;
  assign n7638 = n7634 ^ n7597 ;
  assign n7639 = n7638 ^ n7634 ;
  assign n7640 = ~n7637 & ~n7639 ;
  assign n7641 = n7640 ^ n7634 ;
  assign n7642 = n7626 & ~n7641 ;
  assign n7643 = n7642 ^ n7634 ;
  assign n7646 = n7606 ^ n7575 ;
  assign n7644 = n7615 ^ n7562 ;
  assign n7645 = n7644 ^ n7606 ;
  assign n7647 = n7646 ^ n7645 ;
  assign n7648 = n7647 ^ n7606 ;
  assign n7649 = n7606 ^ n7439 ;
  assign n7650 = n7649 ^ n7606 ;
  assign n7651 = n7648 & ~n7650 ;
  assign n7652 = n7651 ^ n7606 ;
  assign n7653 = n7597 & n7652 ;
  assign n7654 = n7643 & ~n7653 ;
  assign n7574 = n7553 & ~n7561 ;
  assign n7657 = n7439 & n7574 ;
  assign n7658 = n7654 & n7657 ;
  assign n7577 = n7576 ^ n7574 ;
  assign n7573 = n7569 ^ n7562 ;
  assign n7578 = n7577 ^ n7573 ;
  assign n7579 = n7578 ^ n7561 ;
  assign n7580 = n7579 ^ n7567 ;
  assign n7605 = n7604 ^ n7580 ;
  assign n7618 = n7617 ^ n7605 ;
  assign n7558 = n7477 & n7554 ;
  assign n7559 = n7558 ^ n7557 ;
  assign n7560 = n7559 ^ n7477 ;
  assign n7619 = n7618 ^ n7560 ;
  assign n7620 = n7597 & n7619 ;
  assign n7621 = n7620 ^ n7580 ;
  assign n7622 = ~n7439 & ~n7621 ;
  assign n7603 = n7575 & ~n7597 ;
  assign n7623 = n7622 ^ n7603 ;
  assign n7624 = n7623 ^ n5121 ;
  assign n7581 = n7580 ^ n7572 ;
  assign n7582 = n7581 ^ n7560 ;
  assign n7598 = n7597 ^ n7581 ;
  assign n7599 = n7598 ^ n7581 ;
  assign n7600 = ~n7582 & ~n7599 ;
  assign n7601 = n7600 ^ n7581 ;
  assign n7602 = ~n7439 & ~n7601 ;
  assign n7625 = n7624 ^ n7602 ;
  assign n7655 = n7654 ^ n7625 ;
  assign n7659 = n7658 ^ n7655 ;
  assign n7660 = n7659 ^ x68 ;
  assign n7907 = n7906 ^ n6254 ;
  assign n7899 = n7867 ^ n7843 ;
  assign n7900 = n7843 ^ n7699 ;
  assign n7901 = n7900 ^ n7843 ;
  assign n7902 = ~n7899 & ~n7901 ;
  assign n7903 = n7902 ^ n7843 ;
  assign n7904 = n7698 & ~n7903 ;
  assign n7908 = n7907 ^ n7904 ;
  assign n7887 = n7886 ^ n7831 ;
  assign n7883 = n7882 ^ n7852 ;
  assign n7884 = n7883 ^ n7846 ;
  assign n7874 = ~n7836 & ~n7873 ;
  assign n7875 = n7840 ^ n7837 ;
  assign n7876 = ~n7874 & n7875 ;
  assign n7877 = n7876 ^ n7839 ;
  assign n7871 = n7819 & n7862 ;
  assign n7878 = n7877 ^ n7871 ;
  assign n7885 = n7884 ^ n7878 ;
  assign n7888 = n7887 ^ n7885 ;
  assign n7889 = n7888 ^ n7878 ;
  assign n7890 = n7878 ^ n7699 ;
  assign n7891 = n7890 ^ n7878 ;
  assign n7892 = n7889 & n7891 ;
  assign n7893 = n7892 ^ n7878 ;
  assign n7894 = n7870 & n7893 ;
  assign n7895 = n7894 ^ n7878 ;
  assign n7864 = n7863 ^ n7828 ;
  assign n7868 = n7867 ^ n7864 ;
  assign n7869 = ~n7862 & n7868 ;
  assign n7896 = n7895 ^ n7869 ;
  assign n7848 = n7847 ^ n7843 ;
  assign n7849 = n7848 ^ n7835 ;
  assign n7853 = n7852 ^ n7849 ;
  assign n7856 = n7855 ^ n7853 ;
  assign n7857 = n7855 ^ n7699 ;
  assign n7858 = n7857 ^ n7855 ;
  assign n7859 = n7856 & ~n7858 ;
  assign n7860 = n7859 ^ n7855 ;
  assign n7861 = n7698 & ~n7860 ;
  assign n7897 = n7896 ^ n7861 ;
  assign n7898 = ~n7826 & ~n7897 ;
  assign n7909 = n7908 ^ n7898 ;
  assign n7910 = n7909 ^ x126 ;
  assign n7911 = n7660 & n7910 ;
  assign n7914 = n7911 ^ n7660 ;
  assign n8339 = n7914 ^ n7910 ;
  assign n8360 = n7913 & ~n8339 ;
  assign n8330 = n7913 ^ n6894 ;
  assign n8331 = n8330 ^ n7437 ;
  assign n8332 = n7914 & n8331 ;
  assign n7915 = n7913 & n7914 ;
  assign n7912 = n7438 & n7911 ;
  assign n7916 = n7915 ^ n7912 ;
  assign n8344 = n8332 ^ n7916 ;
  assign n8345 = n8344 ^ n7660 ;
  assign n8346 = n7438 & n8345 ;
  assign n10867 = n8360 ^ n8346 ;
  assign n10868 = ~n8325 & n10867 ;
  assign n8395 = n8325 ^ n8131 ;
  assign n8368 = n8346 ^ n7915 ;
  assign n8369 = n8368 ^ n8332 ;
  assign n8366 = n7911 & n7913 ;
  assign n8342 = n8339 ^ n7660 ;
  assign n8336 = n7910 ^ n7660 ;
  assign n8337 = n7660 ^ n7437 ;
  assign n8338 = n8336 & ~n8337 ;
  assign n8352 = n8342 ^ n8338 ;
  assign n8353 = n8352 ^ n7915 ;
  assign n8343 = n7438 & n8342 ;
  assign n8347 = n8346 ^ n8343 ;
  assign n8354 = n8353 ^ n8347 ;
  assign n8351 = ~n8330 & n8342 ;
  assign n8355 = n8354 ^ n8351 ;
  assign n8356 = n8355 ^ n8343 ;
  assign n8363 = n8356 ^ n8342 ;
  assign n8359 = n8331 & ~n8339 ;
  assign n8361 = n8360 ^ n8359 ;
  assign n8348 = n8347 ^ n7912 ;
  assign n8349 = n8348 ^ n7438 ;
  assign n8358 = n8349 ^ n8339 ;
  assign n8362 = n8361 ^ n8358 ;
  assign n8364 = n8363 ^ n8362 ;
  assign n8365 = n8364 ^ n8354 ;
  assign n8367 = n8366 ^ n8365 ;
  assign n8370 = n8369 ^ n8367 ;
  assign n8414 = n8361 ^ n8325 ;
  assign n8415 = n8414 ^ n8361 ;
  assign n10862 = ~n8370 & n8415 ;
  assign n10863 = n10862 ^ n8361 ;
  assign n10864 = n8395 & n10863 ;
  assign n10865 = n10864 ^ n8361 ;
  assign n10859 = n8346 ^ n7912 ;
  assign n10860 = n10859 ^ n8343 ;
  assign n10866 = n10865 ^ n10860 ;
  assign n10869 = n10868 ^ n10866 ;
  assign n10870 = n10869 ^ n10865 ;
  assign n8334 = n7660 ^ n6894 ;
  assign n8335 = n8334 ^ n7910 ;
  assign n8340 = n8339 ^ n8338 ;
  assign n8341 = n8335 & n8340 ;
  assign n10871 = n10870 ^ n8341 ;
  assign n10872 = n10871 ^ n10870 ;
  assign n10875 = ~n8325 & n10872 ;
  assign n10876 = n10875 ^ n10870 ;
  assign n10877 = ~n8131 & n10876 ;
  assign n10878 = n10877 ^ n10869 ;
  assign n10879 = n8364 ^ n8351 ;
  assign n10880 = n8351 ^ n8131 ;
  assign n10881 = n10880 ^ n8351 ;
  assign n10882 = ~n10879 & n10881 ;
  assign n10883 = n10882 ^ n8351 ;
  assign n10884 = n8325 & n10883 ;
  assign n10885 = ~n10878 & ~n10884 ;
  assign n8326 = n8131 & n8325 ;
  assign n8384 = n8326 ^ n8131 ;
  assign n8371 = n8370 ^ n8361 ;
  assign n8350 = n8349 ^ n8341 ;
  assign n8357 = n8356 ^ n8350 ;
  assign n8372 = n8371 ^ n8357 ;
  assign n10854 = n8372 ^ n8332 ;
  assign n10855 = n8384 & n10854 ;
  assign n8327 = n8326 ^ n8325 ;
  assign n8328 = n8327 ^ n8131 ;
  assign n10099 = ~n8328 & n8349 ;
  assign n10856 = n10855 ^ n10099 ;
  assign n10857 = n10856 ^ n8183 ;
  assign n8397 = n8369 ^ n7914 ;
  assign n8396 = n8372 ^ n8364 ;
  assign n8398 = n8397 ^ n8396 ;
  assign n8399 = n8398 ^ n8372 ;
  assign n8400 = n8372 ^ n8325 ;
  assign n8401 = n8400 ^ n8372 ;
  assign n8402 = ~n8399 & ~n8401 ;
  assign n8403 = n8402 ^ n8372 ;
  assign n8404 = n8395 & n8403 ;
  assign n8405 = n8404 ^ n8372 ;
  assign n10858 = n10857 ^ n8405 ;
  assign n10886 = n10885 ^ n10858 ;
  assign n10887 = n10886 ^ x76 ;
  assign n9068 = ~n7360 & n7385 ;
  assign n9066 = n8638 ^ n8636 ;
  assign n9062 = n7407 ^ n7378 ;
  assign n9063 = n9062 ^ n7151 ;
  assign n9064 = n7358 & n9063 ;
  assign n9065 = n9064 ^ n7406 ;
  assign n9067 = n9066 ^ n9065 ;
  assign n9069 = n9068 ^ n9067 ;
  assign n9057 = n7375 ^ n7356 ;
  assign n9058 = n9057 ^ n7375 ;
  assign n9059 = n7377 & ~n9058 ;
  assign n9060 = n9059 ^ n7375 ;
  assign n9061 = ~n7211 & n9060 ;
  assign n9070 = n9069 ^ n9061 ;
  assign n9048 = n7406 ^ n7381 ;
  assign n9049 = n9048 ^ n7406 ;
  assign n9050 = n7406 ^ n7211 ;
  assign n9051 = n9050 ^ n7406 ;
  assign n9052 = ~n9049 & n9051 ;
  assign n9053 = n9052 ^ n7406 ;
  assign n9054 = ~n7356 & ~n9053 ;
  assign n9071 = n9070 ^ n9054 ;
  assign n9072 = n9071 ^ n7359 ;
  assign n9073 = n9072 ^ n6535 ;
  assign n10336 = n9073 ^ x115 ;
  assign n10287 = n8554 ^ n8492 ;
  assign n10288 = n10287 ^ n8507 ;
  assign n9740 = n8525 ^ n8517 ;
  assign n10289 = n10288 ^ n9740 ;
  assign n9712 = n8552 ^ n8491 ;
  assign n10285 = n9712 ^ n8563 ;
  assign n10286 = n10285 ^ n9740 ;
  assign n10290 = n10289 ^ n10286 ;
  assign n10292 = n10285 ^ n8499 ;
  assign n10293 = n8505 & ~n10292 ;
  assign n10294 = n10293 ^ n8499 ;
  assign n10295 = ~n10290 & n10294 ;
  assign n10296 = n10295 ^ n10289 ;
  assign n10297 = ~n8521 & n10296 ;
  assign n10298 = n8515 & n10297 ;
  assign n10282 = n8525 ^ n8519 ;
  assign n10283 = n10282 ^ n8493 ;
  assign n10284 = ~n8499 & n10283 ;
  assign n10299 = n10298 ^ n10284 ;
  assign n10300 = n8505 & ~n10299 ;
  assign n10301 = n10300 ^ n10298 ;
  assign n10275 = n8553 ^ n8512 ;
  assign n10276 = n10275 ^ n8523 ;
  assign n10277 = n8523 ^ n8499 ;
  assign n10278 = n10277 ^ n8523 ;
  assign n10279 = ~n10276 & n10278 ;
  assign n10280 = n10279 ^ n8523 ;
  assign n10281 = ~n8498 & n10280 ;
  assign n10302 = n10301 ^ n10281 ;
  assign n10303 = n10302 ^ n8547 ;
  assign n10304 = n10303 ^ n8565 ;
  assign n9004 = n8545 ^ n8492 ;
  assign n9005 = n8558 & n9004 ;
  assign n9006 = n9005 ^ n8545 ;
  assign n9007 = n8505 & n9006 ;
  assign n10305 = n10304 ^ n9007 ;
  assign n10306 = n10305 ^ n6432 ;
  assign n10307 = n10306 ^ x74 ;
  assign n9271 = n8779 ^ n8765 ;
  assign n9272 = n9271 ^ n8684 ;
  assign n9273 = ~n8683 & ~n9272 ;
  assign n9263 = n8788 ^ n8726 ;
  assign n9241 = ~n8725 & n8754 ;
  assign n9264 = n9263 ^ n9241 ;
  assign n9267 = n9264 ^ n8765 ;
  assign n9262 = n8769 ^ n8764 ;
  assign n9265 = n9264 ^ n9262 ;
  assign n9266 = ~n8683 & n9265 ;
  assign n9268 = n9267 ^ n9266 ;
  assign n9269 = ~n8684 & ~n9268 ;
  assign n9110 = n8790 ^ n8683 ;
  assign n9111 = n8782 ^ n8768 ;
  assign n9112 = n9110 & n9111 ;
  assign n9261 = n9112 ^ n8805 ;
  assign n9270 = n9269 ^ n9261 ;
  assign n9274 = n9273 ^ n9270 ;
  assign n9242 = n9241 ^ n8687 ;
  assign n9243 = n8725 ^ n8723 ;
  assign n9244 = ~n8686 & ~n9243 ;
  assign n9245 = n9242 & n9244 ;
  assign n9246 = n9245 ^ n8686 ;
  assign n9251 = n8781 & n8790 ;
  assign n9252 = n9251 ^ n8776 ;
  assign n9253 = n9246 & ~n9252 ;
  assign n9254 = n9253 ^ n8686 ;
  assign n9255 = n8818 ^ n8790 ;
  assign n9258 = ~n9253 & n9255 ;
  assign n9259 = n9258 ^ n8790 ;
  assign n9260 = n9254 & ~n9259 ;
  assign n9275 = n9274 ^ n9260 ;
  assign n9240 = n8786 & n9110 ;
  assign n9276 = n9275 ^ n9240 ;
  assign n9277 = n8832 ^ n8759 ;
  assign n9278 = n8759 ^ n8684 ;
  assign n9279 = n9278 ^ n8759 ;
  assign n9280 = n9277 & ~n9279 ;
  assign n9281 = n9280 ^ n8759 ;
  assign n9282 = n8683 & n9281 ;
  assign n9283 = n9276 & ~n9282 ;
  assign n9284 = n9283 ^ n5876 ;
  assign n10308 = n9284 ^ x89 ;
  assign n10309 = n10307 & n10308 ;
  assign n10310 = n10309 ^ n10307 ;
  assign n10311 = n10310 ^ n10308 ;
  assign n10266 = n8885 ^ n8233 ;
  assign n10247 = n8298 ^ n8262 ;
  assign n10248 = n10247 ^ n8285 ;
  assign n10249 = n10248 ^ n8885 ;
  assign n10250 = ~n8252 & ~n10249 ;
  assign n10251 = n10250 ^ n8285 ;
  assign n10252 = n8287 ^ n8252 ;
  assign n10253 = ~n10251 & n10252 ;
  assign n10234 = n8874 ^ n8268 ;
  assign n10235 = n10234 ^ n8291 ;
  assign n10236 = ~n8159 & n10235 ;
  assign n10237 = n10236 ^ n8268 ;
  assign n10238 = n10237 ^ n8271 ;
  assign n10239 = n10238 ^ n10237 ;
  assign n10240 = n10237 ^ n8255 ;
  assign n10241 = n10240 ^ n8240 ;
  assign n10242 = n10241 ^ n10237 ;
  assign n10243 = ~n10239 & ~n10242 ;
  assign n10244 = n10243 ^ n10237 ;
  assign n10245 = ~n8281 & ~n10244 ;
  assign n10246 = n10245 ^ n10237 ;
  assign n10254 = n10253 ^ n10246 ;
  assign n10255 = ~n8322 & ~n10254 ;
  assign n10256 = n8281 ^ n8256 ;
  assign n10257 = n8256 ^ n8186 ;
  assign n10258 = n10257 ^ n8253 ;
  assign n10259 = ~n8159 & ~n10258 ;
  assign n10260 = n10259 ^ n8257 ;
  assign n10261 = n10256 & n10260 ;
  assign n10262 = n10261 ^ n8256 ;
  assign n10263 = n10255 & ~n10262 ;
  assign n10264 = ~n8891 & n10263 ;
  assign n10267 = ~n8285 & n10264 ;
  assign n10268 = n10266 & n10267 ;
  assign n10265 = n10264 ^ n6502 ;
  assign n10269 = n10268 ^ n10265 ;
  assign n10270 = n10269 ^ x64 ;
  assign n8961 = n8671 ^ n8658 ;
  assign n8962 = n7957 & n8961 ;
  assign n8963 = n8962 ^ n8658 ;
  assign n8964 = n8963 ^ n8102 ;
  assign n8965 = n8964 ^ n8114 ;
  assign n8966 = n8965 ^ n8964 ;
  assign n8969 = ~n7957 & ~n8966 ;
  assign n8970 = n8969 ^ n8964 ;
  assign n8971 = n7958 & n8970 ;
  assign n8972 = n8971 ^ n8963 ;
  assign n8973 = ~n8107 & ~n8972 ;
  assign n8974 = n8973 ^ n6467 ;
  assign n10271 = n8974 ^ x120 ;
  assign n10272 = ~n10270 & ~n10271 ;
  assign n10273 = n10272 ^ n10271 ;
  assign n10274 = n10273 ^ n10270 ;
  assign n10323 = n10274 ^ n10271 ;
  assign n10325 = ~n10311 & ~n10323 ;
  assign n10320 = ~n10274 & n10310 ;
  assign n9355 = ~n7439 & n7597 ;
  assign n9375 = n9355 ^ n7597 ;
  assign n9370 = n9355 ^ n7439 ;
  assign n9376 = n9375 ^ n9370 ;
  assign n9377 = n7617 ^ n7560 ;
  assign n9378 = ~n9376 & ~n9377 ;
  assign n9371 = n7581 ^ n7562 ;
  assign n9372 = ~n9370 & ~n9371 ;
  assign n9360 = n7580 ^ n7439 ;
  assign n9361 = n7577 ^ n7439 ;
  assign n9362 = n9361 ^ n7597 ;
  assign n9363 = n9362 ^ n9361 ;
  assign n9364 = n9361 ^ n7578 ;
  assign n9365 = n9364 ^ n9361 ;
  assign n9366 = n9363 & n9365 ;
  assign n9367 = n9366 ^ n9361 ;
  assign n9368 = ~n9360 & ~n9367 ;
  assign n9369 = n9368 ^ n7580 ;
  assign n9373 = n9372 ^ n9369 ;
  assign n9356 = n7615 ^ n7558 ;
  assign n9357 = n9356 ^ n7574 ;
  assign n9358 = n9357 ^ n7611 ;
  assign n9359 = n9355 & n9358 ;
  assign n9374 = n9373 ^ n9359 ;
  assign n9379 = n9378 ^ n9374 ;
  assign n9380 = ~n7597 & n7644 ;
  assign n9381 = n9380 ^ n7562 ;
  assign n9382 = n9381 ^ n7439 ;
  assign n9383 = n9382 ^ n9381 ;
  assign n9384 = ~n7597 & n7627 ;
  assign n9385 = n9384 ^ n9381 ;
  assign n9386 = n9383 & n9385 ;
  assign n9387 = n9386 ^ n9381 ;
  assign n9388 = n9379 & n9387 ;
  assign n9389 = n9388 ^ n9379 ;
  assign n9393 = ~n7597 & n7615 ;
  assign n9394 = n9393 ^ n7558 ;
  assign n9395 = n7439 & n9394 ;
  assign n9396 = n9389 & ~n9395 ;
  assign n9397 = n9396 ^ n5472 ;
  assign n10313 = n9397 ^ x122 ;
  assign n10691 = n10320 ^ n10313 ;
  assign n10692 = n10691 ^ n10320 ;
  assign n10693 = n10325 & n10692 ;
  assign n10694 = n10693 ^ n10320 ;
  assign n10695 = ~n10336 & n10694 ;
  assign n10342 = n10336 ^ n10313 ;
  assign n10345 = n10311 ^ n10307 ;
  assign n10346 = ~n10273 & n10345 ;
  assign n10315 = ~n10273 & n10309 ;
  assign n10889 = n10346 ^ n10315 ;
  assign n10326 = n10307 ^ n10270 ;
  assign n10327 = n10308 ^ n10307 ;
  assign n10328 = ~n10326 & n10327 ;
  assign n10365 = n10328 ^ n10310 ;
  assign n10330 = n10328 ^ n10320 ;
  assign n10329 = ~n10271 & n10328 ;
  assign n10331 = n10330 ^ n10329 ;
  assign n10332 = n10331 ^ n10325 ;
  assign n10317 = n10271 ^ n10270 ;
  assign n10318 = n10317 ^ n10308 ;
  assign n10319 = n10307 & ~n10318 ;
  assign n10321 = n10320 ^ n10319 ;
  assign n10314 = n10272 & n10310 ;
  assign n10316 = n10315 ^ n10314 ;
  assign n10322 = n10321 ^ n10316 ;
  assign n10324 = n10323 ^ n10322 ;
  assign n10333 = n10332 ^ n10324 ;
  assign n10334 = n10333 ^ n10331 ;
  assign n10366 = n10365 ^ n10334 ;
  assign n10367 = n10366 ^ n10272 ;
  assign n10343 = n10272 & ~n10311 ;
  assign n10368 = n10367 ^ n10343 ;
  assign n10388 = n10368 ^ n10329 ;
  assign n10389 = n10388 ^ n10343 ;
  assign n10372 = n10308 & n10326 ;
  assign n10373 = n10372 ^ n10368 ;
  assign n10347 = n10346 ^ n10322 ;
  assign n10374 = n10373 ^ n10347 ;
  assign n10375 = n10374 ^ n10325 ;
  assign n10378 = n10375 ^ n10331 ;
  assign n10379 = n10378 ^ n10320 ;
  assign n10390 = n10389 ^ n10379 ;
  assign n10391 = n10390 ^ n10321 ;
  assign n10380 = n10379 ^ n10274 ;
  assign n10312 = ~n10274 & ~n10311 ;
  assign n10377 = n10332 ^ n10312 ;
  assign n10381 = n10380 ^ n10377 ;
  assign n10385 = n10381 ^ n10346 ;
  assign n10386 = n10385 ^ n10333 ;
  assign n10387 = n10386 ^ n10312 ;
  assign n10392 = n10391 ^ n10387 ;
  assign n10890 = n10889 ^ n10392 ;
  assign n10369 = n10313 & ~n10336 ;
  assign n10370 = ~n10368 & n10369 ;
  assign n10891 = n10890 ^ n10370 ;
  assign n10395 = n10369 ^ n10313 ;
  assign n10888 = n10343 & n10395 ;
  assign n10892 = n10891 ^ n10888 ;
  assign n10893 = n10892 ^ n10325 ;
  assign n10684 = n10392 ^ n10329 ;
  assign n10685 = n10684 ^ n10315 ;
  assign n10894 = n10893 ^ n10685 ;
  assign n10895 = n10894 ^ n10892 ;
  assign n10896 = n10892 ^ n10336 ;
  assign n10897 = n10896 ^ n10892 ;
  assign n10898 = n10895 & ~n10897 ;
  assign n10899 = n10898 ^ n10892 ;
  assign n10900 = ~n10313 & n10899 ;
  assign n10901 = n10900 ^ n10892 ;
  assign n10909 = n10901 ^ n10322 ;
  assign n10902 = n10374 ^ n10313 ;
  assign n10903 = n10902 ^ n10374 ;
  assign n10376 = n10375 ^ n10366 ;
  assign n10904 = n10387 ^ n10376 ;
  assign n10905 = n10904 ^ n10374 ;
  assign n10906 = ~n10903 & n10905 ;
  assign n10907 = n10906 ^ n10374 ;
  assign n10908 = ~n10901 & n10907 ;
  assign n10910 = n10909 ^ n10908 ;
  assign n10911 = n10342 & ~n10910 ;
  assign n10912 = n10911 ^ n10909 ;
  assign n10913 = n10331 ^ n10313 ;
  assign n10914 = n10913 ^ n10331 ;
  assign n10915 = n10333 ^ n10312 ;
  assign n10916 = n10915 ^ n10331 ;
  assign n10917 = n10914 & ~n10916 ;
  assign n10918 = n10917 ^ n10331 ;
  assign n10919 = n10336 & n10918 ;
  assign n10920 = n10919 ^ n10331 ;
  assign n10921 = ~n10912 & ~n10920 ;
  assign n10922 = ~n10695 & n10921 ;
  assign n10923 = n10922 ^ n7956 ;
  assign n10924 = n10923 ^ x117 ;
  assign n10925 = ~n10887 & n10924 ;
  assign n10926 = n10925 ^ n10887 ;
  assign n10927 = n10926 ^ n10924 ;
  assign n9286 = n8616 ^ x82 ;
  assign n9285 = n9284 ^ x73 ;
  assign n9287 = n9286 ^ n9285 ;
  assign n9398 = n9397 ^ x97 ;
  assign n9313 = n7152 & n8634 ;
  assign n9310 = n8639 ^ n7370 ;
  assign n9305 = n7158 ^ n7155 ;
  assign n9306 = n9305 ^ n7387 ;
  assign n9307 = n7211 & n9306 ;
  assign n9311 = n9310 ^ n9307 ;
  assign n9301 = n7387 ^ n7378 ;
  assign n9302 = n9301 ^ n7361 ;
  assign n9303 = ~n7211 & n9302 ;
  assign n9300 = n7418 ^ n7374 ;
  assign n9304 = n9303 ^ n9300 ;
  assign n9308 = n9307 ^ n9304 ;
  assign n9309 = n7356 & n9308 ;
  assign n9312 = n9311 ^ n9309 ;
  assign n9314 = n9313 ^ n9312 ;
  assign n9299 = n7357 & n7407 ;
  assign n9315 = n9314 ^ n9299 ;
  assign n9291 = n7406 ^ n7156 ;
  assign n9292 = n9291 ^ n7380 ;
  assign n9293 = n9292 ^ n9291 ;
  assign n9294 = n9291 ^ n7356 ;
  assign n9295 = n9294 ^ n9291 ;
  assign n9296 = n9293 & ~n9295 ;
  assign n9297 = n9296 ^ n9291 ;
  assign n9298 = ~n7360 & ~n9297 ;
  assign n9316 = n9315 ^ n9298 ;
  assign n9317 = n9316 ^ n7359 ;
  assign n9318 = n9317 ^ n5644 ;
  assign n9319 = n9318 ^ x114 ;
  assign n9290 = n8897 ^ x88 ;
  assign n9333 = n6867 ^ n6862 ;
  assign n9334 = n9333 ^ n6876 ;
  assign n9344 = n9334 ^ n6841 ;
  assign n9338 = n6874 ^ n6842 ;
  assign n9339 = n6874 ^ n5398 ;
  assign n9340 = n9339 ^ n6874 ;
  assign n9341 = n9338 & n9340 ;
  assign n9342 = n9341 ^ n6874 ;
  assign n9343 = ~n6860 & n9342 ;
  assign n9345 = n9344 ^ n9343 ;
  assign n9346 = n9345 ^ n6849 ;
  assign n9123 = n6858 ^ n6834 ;
  assign n9332 = n9123 ^ n6824 ;
  assign n9335 = n9334 ^ n9332 ;
  assign n9328 = n6824 ^ n6396 ;
  assign n9329 = n9328 ^ n6874 ;
  assign n9330 = n9329 ^ n6881 ;
  assign n9331 = n5398 & ~n9330 ;
  assign n9336 = n9335 ^ n9331 ;
  assign n9337 = ~n6860 & n9336 ;
  assign n9347 = n9346 ^ n9337 ;
  assign n9132 = n6839 & n6850 ;
  assign n9348 = n9347 ^ n9132 ;
  assign n9349 = n9348 ^ n5506 ;
  assign n9350 = n9349 ^ n6881 ;
  assign n9320 = n6881 ^ n6823 ;
  assign n9321 = n9320 ^ n5398 ;
  assign n9322 = n9321 ^ n9320 ;
  assign n9323 = n9320 ^ n6832 ;
  assign n9324 = n9323 ^ n9320 ;
  assign n9325 = ~n9322 & ~n9324 ;
  assign n9326 = n9325 ^ n9320 ;
  assign n9327 = n5966 & n9326 ;
  assign n9351 = n9350 ^ n9327 ;
  assign n9352 = n9351 ^ x107 ;
  assign n9402 = ~n9290 & ~n9352 ;
  assign n9403 = n9402 ^ n9352 ;
  assign n9404 = ~n9319 & ~n9403 ;
  assign n9405 = n9404 ^ n9403 ;
  assign n9406 = n9398 & ~n9405 ;
  assign n9421 = n9406 ^ n9405 ;
  assign n9399 = ~n9290 & ~n9398 ;
  assign n9422 = n9421 ^ n9399 ;
  assign n9418 = n9403 ^ n9290 ;
  assign n9419 = ~n9398 & ~n9418 ;
  assign n9420 = n9419 ^ n9398 ;
  assign n9423 = n9422 ^ n9420 ;
  assign n9424 = n9423 ^ n9404 ;
  assign n9408 = n9319 & n9398 ;
  assign n9413 = n9408 ^ n9398 ;
  assign n9431 = n9424 ^ n9413 ;
  assign n9430 = ~n9290 & n9413 ;
  assign n9432 = n9431 ^ n9430 ;
  assign n9465 = n9432 ^ n9285 ;
  assign n9466 = n9465 ^ n9432 ;
  assign n9414 = n9402 & n9413 ;
  assign n9487 = n9430 ^ n9414 ;
  assign n9977 = n9487 ^ n9432 ;
  assign n9980 = ~n9466 & n9977 ;
  assign n9981 = n9980 ^ n9432 ;
  assign n9982 = ~n9287 & n9981 ;
  assign n9353 = n9319 & n9352 ;
  assign n9354 = ~n9290 & n9353 ;
  assign n9450 = n9354 ^ n9353 ;
  assign n9410 = n9352 & n9399 ;
  assign n9411 = n9410 ^ n9399 ;
  assign n9412 = n9411 ^ n9402 ;
  assign n9415 = n9414 ^ n9412 ;
  assign n9400 = n9353 & n9399 ;
  assign n9401 = n9400 ^ n9354 ;
  assign n9407 = n9406 ^ n9401 ;
  assign n9409 = n9408 ^ n9407 ;
  assign n9416 = n9415 ^ n9409 ;
  assign n9451 = n9450 ^ n9416 ;
  assign n9452 = n9451 ^ n9419 ;
  assign n9453 = n9452 ^ n9411 ;
  assign n10945 = n9453 ^ n9451 ;
  assign n10943 = n9414 ^ n9413 ;
  assign n10944 = n10943 ^ n9401 ;
  assign n10946 = n10945 ^ n10944 ;
  assign n10947 = ~n9285 & n10946 ;
  assign n10948 = n10947 ^ n10945 ;
  assign n10941 = n9453 ^ n9423 ;
  assign n10942 = n9285 & n10941 ;
  assign n10951 = n10948 ^ n10942 ;
  assign n10952 = ~n9286 & n10951 ;
  assign n9488 = n9487 ^ n9424 ;
  assign n9489 = n9424 ^ n9285 ;
  assign n9490 = n9489 ^ n9424 ;
  assign n9491 = n9488 & n9490 ;
  assign n9492 = n9491 ^ n9424 ;
  assign n9493 = ~n9287 & n9492 ;
  assign n10949 = n10948 ^ n9493 ;
  assign n10953 = n10952 ^ n10949 ;
  assign n10938 = ~n9286 & ~n9420 ;
  assign n10936 = n9421 ^ n9411 ;
  assign n10937 = n10936 ^ n9451 ;
  assign n10939 = n10938 ^ n10937 ;
  assign n10940 = ~n9285 & ~n10939 ;
  assign n10954 = n10953 ^ n10940 ;
  assign n9288 = ~n9285 & n9286 ;
  assign n9429 = n9288 ^ n9286 ;
  assign n9440 = n9429 ^ n9285 ;
  assign n10935 = n9408 & n9440 ;
  assign n10955 = n10954 ^ n10935 ;
  assign n9425 = n9424 ^ n9415 ;
  assign n9417 = n9416 ^ n9414 ;
  assign n9426 = n9425 ^ n9417 ;
  assign n10930 = n9425 ^ n9285 ;
  assign n10931 = n10930 ^ n9425 ;
  assign n10932 = n9426 & ~n10931 ;
  assign n10933 = n10932 ^ n9425 ;
  assign n10934 = ~n9287 & n10933 ;
  assign n10956 = n10955 ^ n10934 ;
  assign n10957 = ~n9982 & ~n10956 ;
  assign n10958 = n10957 ^ n8228 ;
  assign n10959 = n10958 ^ x124 ;
  assign n9524 = n8648 ^ x99 ;
  assign n9626 = n8579 ^ x106 ;
  assign n9546 = n6867 ^ n5398 ;
  assign n9547 = n9546 ^ n6867 ;
  assign n9548 = n6879 ^ n6867 ;
  assign n9549 = n9547 & n9548 ;
  assign n9550 = n9549 ^ n6867 ;
  assign n9551 = ~n5966 & n9550 ;
  assign n9552 = n9551 ^ n9343 ;
  assign n9535 = n6625 ^ n6166 ;
  assign n9536 = n6818 ^ n6396 ;
  assign n9537 = ~n5398 & n9536 ;
  assign n9538 = ~n9535 & n9537 ;
  assign n9545 = n9538 ^ n6867 ;
  assign n9553 = n9552 ^ n9545 ;
  assign n9540 = n9123 ^ n6823 ;
  assign n9122 = n6875 ^ n6830 ;
  assign n9541 = n9540 ^ n9122 ;
  assign n9539 = n9538 ^ n6819 ;
  assign n9542 = n9541 ^ n9539 ;
  assign n9532 = n9123 ^ n6837 ;
  assign n9533 = n9532 ^ n6823 ;
  assign n9534 = ~n5966 & ~n9533 ;
  assign n9543 = n9542 ^ n9534 ;
  assign n9544 = n6860 & n9543 ;
  assign n9554 = n9553 ^ n9544 ;
  assign n9555 = n9554 ^ n9132 ;
  assign n9527 = n6827 ^ n5966 ;
  assign n9528 = n9527 ^ n6827 ;
  assign n9529 = n6863 & n9528 ;
  assign n9530 = n9529 ^ n6827 ;
  assign n9531 = ~n6860 & n9530 ;
  assign n9556 = n9555 ^ n9531 ;
  assign n9557 = ~n6882 & ~n9556 ;
  assign n9558 = n9557 ^ n5285 ;
  assign n9559 = n9558 ^ x123 ;
  assign n9648 = n9626 ^ n9559 ;
  assign n9583 = n8289 ^ n8252 ;
  assign n9584 = n8286 & ~n9583 ;
  assign n9566 = ~n8271 & ~n8873 ;
  assign n9567 = n9566 ^ n8872 ;
  assign n9561 = n8277 ^ n8249 ;
  assign n9562 = n9561 ^ n8271 ;
  assign n9563 = n8238 & ~n9562 ;
  assign n9564 = ~n9561 & n9563 ;
  assign n9565 = n9564 ^ n9562 ;
  assign n9568 = n9567 ^ n9565 ;
  assign n9576 = n9567 ^ n8159 ;
  assign n9573 = n8261 & ~n8271 ;
  assign n9574 = n9573 ^ n8240 ;
  assign n9575 = n8159 & n9574 ;
  assign n9577 = n9576 ^ n9575 ;
  assign n9578 = n9577 ^ n8271 ;
  assign n9579 = n9578 ^ n9565 ;
  assign n9580 = n9579 ^ n9575 ;
  assign n9581 = n9568 & n9580 ;
  assign n9582 = n9581 ^ n9577 ;
  assign n9587 = n9584 ^ n9582 ;
  assign n9588 = ~n8288 & ~n9587 ;
  assign n9560 = n8322 ^ n6021 ;
  assign n9589 = n9588 ^ n9560 ;
  assign n9590 = n9589 ^ x105 ;
  assign n9640 = n9626 ^ n9590 ;
  assign n9595 = n7610 ^ n7560 ;
  assign n9606 = n9595 ^ n7555 ;
  assign n9607 = n9606 ^ n7613 ;
  assign n9605 = n7552 ^ n7474 ;
  assign n9608 = n9607 ^ n9605 ;
  assign n9609 = n9608 ^ n7627 ;
  assign n9610 = ~n7597 & n9609 ;
  assign n9611 = n9610 ^ n7627 ;
  assign n9612 = n7439 & n9611 ;
  assign n9592 = n7572 ^ n7567 ;
  assign n9593 = n9592 ^ n7646 ;
  assign n9594 = ~n7439 & n9593 ;
  assign n9597 = n9594 ^ n7608 ;
  assign n9596 = n9595 ^ n9594 ;
  assign n9598 = n9597 ^ n9596 ;
  assign n9601 = ~n7439 & n9598 ;
  assign n9602 = n9601 ^ n9597 ;
  assign n9603 = n7597 & n9602 ;
  assign n9604 = n9603 ^ n9594 ;
  assign n9613 = n9612 ^ n9604 ;
  assign n9616 = n7567 & n7597 ;
  assign n9617 = n9616 ^ n7557 ;
  assign n9618 = n7626 & n9617 ;
  assign n9619 = n9618 ^ n7557 ;
  assign n9620 = ~n9613 & n9619 ;
  assign n9621 = n9620 ^ n9613 ;
  assign n9622 = ~n9395 & ~n9621 ;
  assign n9623 = ~n7602 & n9622 ;
  assign n9624 = n9623 ^ n5987 ;
  assign n9625 = n9624 ^ x96 ;
  assign n9649 = n9640 ^ n9625 ;
  assign n9652 = ~n9559 & n9649 ;
  assign n9591 = n9590 ^ n9559 ;
  assign n9639 = n9591 ^ n9559 ;
  assign n9643 = n9626 ^ n9591 ;
  assign n9644 = n9639 & ~n9643 ;
  assign n9645 = n9644 ^ n9591 ;
  assign n9646 = n9625 & ~n9645 ;
  assign n9641 = n9640 ^ n9559 ;
  assign n9647 = n9646 ^ n9641 ;
  assign n9650 = n9649 ^ n9647 ;
  assign n9651 = n9650 ^ n9590 ;
  assign n9653 = n9652 ^ n9651 ;
  assign n9654 = n9653 ^ n9647 ;
  assign n9655 = ~n9648 & n9654 ;
  assign n9656 = n9655 ^ n9650 ;
  assign n9657 = n9524 & ~n9656 ;
  assign n9658 = n9657 ^ n9647 ;
  assign n9512 = n7883 ^ n7867 ;
  assign n9513 = n9512 ^ n7828 ;
  assign n9504 = n7854 ^ n7844 ;
  assign n9505 = n9504 ^ n8599 ;
  assign n9506 = n9505 ^ n7887 ;
  assign n9507 = ~n7698 & ~n9506 ;
  assign n9514 = n9513 ^ n9507 ;
  assign n9508 = n7839 ^ n7828 ;
  assign n9509 = n9508 ^ n7882 ;
  assign n9510 = n9509 ^ n7849 ;
  assign n9511 = ~n7698 & n9510 ;
  assign n9515 = n9514 ^ n9511 ;
  assign n9516 = n7699 & ~n9515 ;
  assign n9517 = n9516 ^ n9507 ;
  assign n9501 = n8590 ^ n7854 ;
  assign n9502 = n9501 ^ n7863 ;
  assign n9503 = n7872 & ~n9502 ;
  assign n9518 = n9517 ^ n9503 ;
  assign n9519 = n9518 ^ n7906 ;
  assign n9500 = n7837 & n7873 ;
  assign n9520 = n9519 ^ n9500 ;
  assign n9521 = ~n7904 & ~n9520 ;
  assign n9522 = n9521 ^ n4302 ;
  assign n9523 = n9522 ^ x81 ;
  assign n10960 = n9658 ^ n9523 ;
  assign n9636 = n9626 ^ n9625 ;
  assign n9632 = n9625 ^ n9590 ;
  assign n9633 = ~n9590 & n9626 ;
  assign n9634 = n9633 ^ n9559 ;
  assign n9635 = n9632 & ~n9634 ;
  assign n9637 = n9636 ^ n9635 ;
  assign n9627 = ~n9625 & n9626 ;
  assign n9628 = n9627 ^ n9590 ;
  assign n9629 = n9591 & n9628 ;
  assign n9630 = n9629 ^ n9590 ;
  assign n9631 = ~n9524 & ~n9630 ;
  assign n9638 = n9637 ^ n9631 ;
  assign n9659 = n9658 ^ n9638 ;
  assign n9660 = n9523 & n9659 ;
  assign n9661 = n9660 ^ n9658 ;
  assign n10961 = n10960 ^ n9661 ;
  assign n10962 = n10961 ^ n9638 ;
  assign n10963 = n10962 ^ n8189 ;
  assign n10964 = n10963 ^ x94 ;
  assign n10965 = n10959 & n10964 ;
  assign n10966 = n10965 ^ n10964 ;
  assign n10992 = n10927 & n10966 ;
  assign n10991 = n10927 & n10965 ;
  assign n10993 = n10992 ^ n10991 ;
  assign n10967 = n10966 ^ n10959 ;
  assign n10968 = n10927 & ~n10967 ;
  assign n10990 = n10968 ^ n10927 ;
  assign n10994 = n10993 ^ n10990 ;
  assign n10973 = n10967 ^ n10964 ;
  assign n10995 = n10994 ^ n10973 ;
  assign n10987 = n10927 ^ n10887 ;
  assign n10988 = n10973 & n10987 ;
  assign n10974 = n10925 & n10973 ;
  assign n10989 = n10988 ^ n10974 ;
  assign n10996 = n10995 ^ n10989 ;
  assign n10971 = n10925 & n10965 ;
  assign n11047 = n10996 ^ n10971 ;
  assign n9041 = n7839 ^ n7834 ;
  assign n9042 = n9041 ^ n7843 ;
  assign n9043 = ~n7699 & ~n9042 ;
  assign n9044 = n9043 ^ n7854 ;
  assign n9045 = n7870 & n9044 ;
  assign n9039 = n7873 & n7884 ;
  assign n9034 = n7864 & n7872 ;
  assign n9028 = n7874 ^ n7818 ;
  assign n9029 = ~n7870 & n9028 ;
  assign n9027 = ~n7874 & n7905 ;
  assign n9030 = n9029 ^ n9027 ;
  assign n9031 = n9030 ^ n7904 ;
  assign n9026 = n7843 & ~n7862 ;
  assign n9032 = n9031 ^ n9026 ;
  assign n9023 = n7841 ^ n7830 ;
  assign n9024 = n9023 ^ n7850 ;
  assign n9025 = n7700 & ~n9024 ;
  assign n9033 = n9032 ^ n9025 ;
  assign n9035 = n9034 ^ n9033 ;
  assign n9021 = n7867 ^ n7847 ;
  assign n9022 = ~n7862 & ~n9021 ;
  assign n9036 = n9035 ^ n9022 ;
  assign n9037 = n9036 ^ n7854 ;
  assign n9038 = n9037 ^ n6993 ;
  assign n9040 = n9039 ^ n9038 ;
  assign n9046 = n9045 ^ n9040 ;
  assign n9047 = n9046 ^ x100 ;
  assign n9074 = n9073 ^ x93 ;
  assign n9075 = n9047 & ~n9074 ;
  assign n9161 = n9075 ^ n9047 ;
  assign n9171 = n9161 ^ n9074 ;
  assign n9114 = n8811 ^ n8684 ;
  assign n9094 = n8786 & ~n8790 ;
  assign n9092 = n8776 ^ n8759 ;
  assign n9083 = n8684 ^ n8683 ;
  assign n9084 = n8788 ^ n8772 ;
  assign n9085 = n9084 ^ n8817 ;
  assign n9086 = n9085 ^ n8772 ;
  assign n9087 = n8772 ^ n8684 ;
  assign n9088 = n9087 ^ n8772 ;
  assign n9089 = n9086 & ~n9088 ;
  assign n9090 = n9089 ^ n8772 ;
  assign n9091 = n9083 & n9090 ;
  assign n9093 = n9092 ^ n9091 ;
  assign n9095 = n9094 ^ n9093 ;
  assign n9115 = n9114 ^ n9095 ;
  assign n9113 = n9112 ^ n8835 ;
  assign n9116 = n9115 ^ n9113 ;
  assign n9104 = n8819 ^ n8769 ;
  assign n9105 = n8769 ^ n8684 ;
  assign n9106 = n9105 ^ n8769 ;
  assign n9107 = n9104 & n9106 ;
  assign n9108 = n9107 ^ n8769 ;
  assign n9109 = n8683 & n9108 ;
  assign n9117 = n9116 ^ n9109 ;
  assign n9118 = n9117 ^ n6659 ;
  assign n9096 = n9095 ^ n9091 ;
  assign n9097 = n9096 ^ n8766 ;
  assign n9098 = n9097 ^ n9096 ;
  assign n9099 = n9096 ^ n8684 ;
  assign n9100 = n9099 ^ n9096 ;
  assign n9101 = ~n9098 & n9100 ;
  assign n9102 = n9101 ^ n9096 ;
  assign n9103 = n8683 & ~n9102 ;
  assign n9119 = n9118 ^ n9103 ;
  assign n9076 = n8790 ^ n8780 ;
  assign n9077 = n8765 ^ n8686 ;
  assign n9080 = n8790 & ~n9077 ;
  assign n9081 = n9080 ^ n8765 ;
  assign n9082 = n9076 & ~n9081 ;
  assign n9120 = n9119 ^ n9082 ;
  assign n9121 = n9120 ^ x83 ;
  assign n9154 = n5967 & ~n6833 ;
  assign n9136 = n6876 ^ n6842 ;
  assign n9137 = n9136 ^ n6867 ;
  assign n9138 = n9137 ^ n9136 ;
  assign n9139 = n9136 ^ n5966 ;
  assign n9140 = n9139 ^ n9136 ;
  assign n9141 = ~n9138 & n9140 ;
  assign n9142 = n9141 ^ n9136 ;
  assign n9145 = n6842 ^ n5398 ;
  assign n9146 = n9145 ^ n6852 ;
  assign n9143 = n6842 ^ n5966 ;
  assign n9144 = n9143 ^ n6852 ;
  assign n9147 = n9146 ^ n9144 ;
  assign n9148 = ~n9142 & ~n9147 ;
  assign n9149 = n9148 ^ n9146 ;
  assign n9133 = n6858 ^ n6839 ;
  assign n9134 = n9133 ^ n6862 ;
  assign n9135 = ~n5966 & n9134 ;
  assign n9150 = n9149 ^ n9135 ;
  assign n9151 = n9150 ^ n9132 ;
  assign n9152 = n9151 ^ n6882 ;
  assign n9124 = n9123 ^ n9122 ;
  assign n9125 = n9123 ^ n6886 ;
  assign n9126 = n9125 ^ n9123 ;
  assign n9127 = ~n9124 & n9126 ;
  assign n9128 = n9127 ^ n9123 ;
  assign n9129 = n6854 ^ n6832 ;
  assign n9130 = n9129 ^ n5966 ;
  assign n9131 = n9128 & ~n9130 ;
  assign n9153 = n9152 ^ n9131 ;
  assign n9155 = n9154 ^ n9153 ;
  assign n9156 = ~n6836 & n9155 ;
  assign n9157 = n9156 ^ n7027 ;
  assign n9158 = n9157 ^ x86 ;
  assign n9159 = n9121 & ~n9158 ;
  assign n9181 = n9159 ^ n9158 ;
  assign n9191 = n9171 & ~n9181 ;
  assign n9166 = n9075 ^ n9074 ;
  assign n9162 = n9159 ^ n9121 ;
  assign n9184 = n9162 ^ n9158 ;
  assign n9187 = ~n9166 & n9184 ;
  assign n9198 = n9191 ^ n9187 ;
  assign n8975 = n8974 ^ x69 ;
  assign n9008 = n9007 ^ n8504 ;
  assign n9009 = n9008 ^ n8508 ;
  assign n9001 = n8525 ^ n8523 ;
  assign n9000 = n8563 ^ n8491 ;
  assign n9002 = n9001 ^ n9000 ;
  assign n9003 = ~n8502 & n9002 ;
  assign n9010 = n9009 ^ n9003 ;
  assign n8992 = n8545 ^ n8508 ;
  assign n8993 = n8992 ^ n8554 ;
  assign n8994 = n8993 ^ n8508 ;
  assign n8995 = n8508 ^ n8498 ;
  assign n8996 = n8995 ^ n8508 ;
  assign n8997 = ~n8994 & ~n8996 ;
  assign n8998 = n8997 ^ n8508 ;
  assign n8999 = n8499 & n8998 ;
  assign n9011 = n9010 ^ n8999 ;
  assign n8985 = n8513 ^ n8497 ;
  assign n8986 = n8985 ^ n8524 ;
  assign n8987 = n8524 ^ n8499 ;
  assign n8988 = n8987 ^ n8524 ;
  assign n8989 = ~n8986 & n8988 ;
  assign n8990 = n8989 ^ n8524 ;
  assign n8991 = n8498 & n8990 ;
  assign n9012 = n9011 ^ n8991 ;
  assign n9013 = n9012 ^ n8552 ;
  assign n9014 = n9013 ^ n8544 ;
  assign n9015 = n9014 ^ n6718 ;
  assign n8984 = n8503 & n8529 ;
  assign n9016 = n9015 ^ n8984 ;
  assign n8983 = n8501 & ~n8554 ;
  assign n9017 = n9016 ^ n8983 ;
  assign n8976 = n8552 ^ n8502 ;
  assign n8977 = n8515 ^ n8500 ;
  assign n8980 = ~n8502 & n8977 ;
  assign n8981 = n8980 ^ n8500 ;
  assign n8982 = ~n8976 & ~n8981 ;
  assign n9018 = n9017 ^ n8982 ;
  assign n9019 = n9018 ^ x118 ;
  assign n10814 = n8975 & n9019 ;
  assign n10815 = n10814 ^ n8975 ;
  assign n10816 = n9198 & n10815 ;
  assign n9186 = n9161 & n9184 ;
  assign n9188 = n9187 ^ n9186 ;
  assign n9185 = n9075 & n9184 ;
  assign n9189 = n9188 ^ n9185 ;
  assign n9190 = n9189 ^ n9184 ;
  assign n9182 = n9075 & ~n9181 ;
  assign n9223 = n9190 ^ n9182 ;
  assign n9169 = n9075 & n9162 ;
  assign n9163 = n9161 & n9162 ;
  assign n9174 = n9169 ^ n9163 ;
  assign n9172 = n9162 & n9171 ;
  assign n9175 = n9174 ^ n9172 ;
  assign n9176 = n9175 ^ n9162 ;
  assign n9168 = n9159 & n9161 ;
  assign n9170 = n9169 ^ n9168 ;
  assign n9173 = n9172 ^ n9170 ;
  assign n9177 = n9176 ^ n9173 ;
  assign n9167 = n9159 & ~n9166 ;
  assign n9178 = n9177 ^ n9167 ;
  assign n9160 = n9075 & n9159 ;
  assign n9164 = n9163 ^ n9160 ;
  assign n9165 = n9164 ^ n9121 ;
  assign n9179 = n9178 ^ n9165 ;
  assign n9180 = n9179 ^ n9176 ;
  assign n9224 = n9223 ^ n9180 ;
  assign n9225 = n8975 & n9224 ;
  assign n9226 = n9225 ^ n9180 ;
  assign n9229 = n9226 ^ n9170 ;
  assign n9230 = n9229 ^ n9226 ;
  assign n9231 = ~n8975 & n9230 ;
  assign n9232 = n9231 ^ n9226 ;
  assign n9233 = ~n9019 & n9232 ;
  assign n9234 = n9233 ^ n9226 ;
  assign n10808 = n9234 ^ n9167 ;
  assign n10788 = n9188 ^ n9179 ;
  assign n10789 = n10788 ^ n9185 ;
  assign n10790 = n10789 ^ n9179 ;
  assign n10791 = n9019 & n10790 ;
  assign n10792 = n10791 ^ n10788 ;
  assign n10809 = n10808 ^ n10792 ;
  assign n9193 = n9161 & ~n9181 ;
  assign n9206 = n9193 ^ n9185 ;
  assign n9194 = n9193 ^ n9182 ;
  assign n9192 = n9191 ^ n9181 ;
  assign n9195 = n9194 ^ n9192 ;
  assign n9196 = n9195 ^ n9190 ;
  assign n10802 = n9206 ^ n9196 ;
  assign n10803 = n9196 ^ n9019 ;
  assign n10804 = n10803 ^ n9196 ;
  assign n10805 = ~n10802 & ~n10804 ;
  assign n10806 = n10805 ^ n9196 ;
  assign n10807 = ~n8975 & ~n10806 ;
  assign n10810 = n10809 ^ n10807 ;
  assign n10811 = n10810 ^ n8158 ;
  assign n9020 = n9019 ^ n8975 ;
  assign n10798 = n9223 ^ n9186 ;
  assign n10799 = ~n9019 & n10798 ;
  assign n10794 = n10792 ^ n9193 ;
  assign n10795 = n10794 ^ n9164 ;
  assign n10793 = n10792 ^ n9182 ;
  assign n10796 = n10795 ^ n10793 ;
  assign n10797 = n10796 ^ n10792 ;
  assign n10800 = n10799 ^ n10797 ;
  assign n10801 = n9020 & n10800 ;
  assign n10812 = n10811 ^ n10801 ;
  assign n10785 = n8975 & n9177 ;
  assign n10786 = n10785 ^ n9167 ;
  assign n10787 = n9019 & n10786 ;
  assign n10813 = n10812 ^ n10787 ;
  assign n10817 = n10816 ^ n10813 ;
  assign n10818 = n10817 ^ x93 ;
  assign n11048 = n10971 ^ n10818 ;
  assign n11049 = n11048 ^ n10971 ;
  assign n11050 = n11047 & ~n11049 ;
  assign n11051 = n11050 ^ n10971 ;
  assign n11052 = ~n10852 & n11051 ;
  assign n10983 = ~n10818 & ~n10852 ;
  assign n10984 = n10983 ^ n10852 ;
  assign n10985 = n10984 ^ n10818 ;
  assign n10998 = ~n10967 & n10987 ;
  assign n10999 = n10998 ^ n10992 ;
  assign n11013 = n10999 ^ n10971 ;
  assign n11007 = n10959 ^ n10925 ;
  assign n11010 = n10959 ^ n10887 ;
  assign n11008 = n10925 ^ n10924 ;
  assign n11009 = n11008 ^ n10964 ;
  assign n11011 = n11010 ^ n11009 ;
  assign n11012 = ~n11007 & ~n11011 ;
  assign n11014 = n11013 ^ n11012 ;
  assign n11015 = n11014 ^ n10991 ;
  assign n11004 = n10965 & n10987 ;
  assign n11005 = n11004 ^ n10998 ;
  assign n11003 = n10988 ^ n10987 ;
  assign n11006 = n11005 ^ n11003 ;
  assign n11016 = n11015 ^ n11006 ;
  assign n11017 = n11016 ^ n10959 ;
  assign n10975 = n10925 & n10966 ;
  assign n11000 = n10999 ^ n10975 ;
  assign n10976 = n10975 ^ n10974 ;
  assign n10972 = n10971 ^ n10925 ;
  assign n10977 = n10976 ^ n10972 ;
  assign n11001 = n11000 ^ n10977 ;
  assign n10997 = n10991 ^ n10968 ;
  assign n11002 = n11001 ^ n10997 ;
  assign n11018 = n11017 ^ n11002 ;
  assign n11019 = n11018 ^ n10996 ;
  assign n11063 = n11019 ^ n11015 ;
  assign n11064 = n11063 ^ n10993 ;
  assign n11062 = n10992 ^ n10926 ;
  assign n11065 = n11064 ^ n11062 ;
  assign n12745 = ~n10985 & n11065 ;
  assign n12738 = n11002 ^ n10974 ;
  assign n11035 = n11004 ^ n10977 ;
  assign n12739 = n12738 ^ n11035 ;
  assign n11770 = n11065 ^ n10968 ;
  assign n11771 = n11770 ^ n10992 ;
  assign n11772 = n11771 ^ n10994 ;
  assign n12740 = n12739 ^ n11772 ;
  assign n12741 = n10818 & n12740 ;
  assign n12732 = n11005 ^ n10976 ;
  assign n12733 = n12732 ^ n11018 ;
  assign n12734 = n12733 ^ n11014 ;
  assign n11021 = n10988 ^ n10975 ;
  assign n11022 = n11021 ^ n11006 ;
  assign n12726 = n11022 ^ n10974 ;
  assign n12727 = n12726 ^ n10818 ;
  assign n10853 = n10852 ^ n10818 ;
  assign n12728 = n10853 ^ n10818 ;
  assign n12729 = n12727 & ~n12728 ;
  assign n12730 = n12729 ^ n10818 ;
  assign n12731 = n10987 & ~n12730 ;
  assign n12735 = n12734 ^ n12731 ;
  assign n12737 = n12735 ^ n11002 ;
  assign n12742 = n12741 ^ n12737 ;
  assign n12743 = ~n10852 & ~n12742 ;
  assign n12736 = n12735 ^ n10994 ;
  assign n12744 = n12743 ^ n12736 ;
  assign n12746 = n12745 ^ n12744 ;
  assign n12719 = n11770 ^ n10994 ;
  assign n12720 = n12719 ^ n10994 ;
  assign n12721 = n10994 ^ n10818 ;
  assign n12722 = n12721 ^ n10994 ;
  assign n12723 = n12720 & ~n12722 ;
  assign n12724 = n12723 ^ n10994 ;
  assign n12725 = n10853 & n12724 ;
  assign n12747 = n12746 ^ n12725 ;
  assign n12748 = ~n11052 & n12747 ;
  assign n12749 = n12748 ^ n8324 ;
  assign n12750 = n12749 ^ x78 ;
  assign n10125 = n7606 ^ n7604 ;
  assign n10121 = ~n7559 & n9370 ;
  assign n10124 = ~n7616 & ~n10121 ;
  assign n10126 = n10125 ^ n10124 ;
  assign n10127 = n10126 ^ n7570 ;
  assign n10128 = n10127 ^ n7615 ;
  assign n10129 = n10128 ^ n9377 ;
  assign n10130 = n10129 ^ n10126 ;
  assign n10131 = n7439 & ~n10130 ;
  assign n10132 = n10131 ^ n10127 ;
  assign n10133 = n9376 & n10132 ;
  assign n10134 = n10133 ^ n10126 ;
  assign n10120 = n7567 ^ n7566 ;
  assign n10122 = n10121 ^ n10120 ;
  assign n10123 = n9375 & ~n10122 ;
  assign n10135 = n10134 ^ n10123 ;
  assign n10119 = n7571 & ~n9376 ;
  assign n10136 = n10135 ^ n10119 ;
  assign n10137 = n7574 ^ n7559 ;
  assign n10138 = n7597 & n10137 ;
  assign n10139 = n10138 ^ n7574 ;
  assign n10140 = n10139 ^ n7439 ;
  assign n10141 = n10140 ^ n10139 ;
  assign n10142 = ~n7581 & ~n7597 ;
  assign n10143 = n10142 ^ n10139 ;
  assign n10144 = n10141 & n10143 ;
  assign n10145 = n10144 ^ n10139 ;
  assign n10146 = ~n10136 & n10145 ;
  assign n10147 = n10146 ^ n10136 ;
  assign n10148 = ~n7623 & ~n10147 ;
  assign n10149 = n10148 ^ n6681 ;
  assign n10150 = n10149 ^ x101 ;
  assign n10116 = n8324 ^ x94 ;
  assign n10151 = n9018 ^ x116 ;
  assign n10117 = n8126 ^ n6724 ;
  assign n10118 = n10117 ^ x76 ;
  assign n10164 = n10151 ^ n10118 ;
  assign n10163 = ~n10118 & ~n10151 ;
  assign n10165 = n10164 ^ n10163 ;
  assign n10166 = n10165 ^ n10118 ;
  assign n10167 = n10116 & ~n10166 ;
  assign n10168 = ~n10150 & n10167 ;
  assign n10161 = n10116 & ~n10118 ;
  assign n10162 = ~n10150 & n10161 ;
  assign n10169 = n10168 ^ n10162 ;
  assign n10159 = ~n10116 & ~n10150 ;
  assign n10160 = n10159 ^ n10150 ;
  assign n10170 = n10169 ^ n10160 ;
  assign n10155 = n6893 ^ x67 ;
  assign n10156 = n9120 ^ x125 ;
  assign n10171 = n10155 & n10156 ;
  assign n10172 = n10171 ^ n10156 ;
  assign n10173 = ~n10170 & n10172 ;
  assign n10152 = n10150 & n10151 ;
  assign n10153 = ~n10118 & n10152 ;
  assign n10154 = ~n10116 & n10153 ;
  assign n10157 = n10156 ^ n10155 ;
  assign n10158 = n10154 & ~n10157 ;
  assign n10174 = n10173 ^ n10158 ;
  assign n10206 = n10154 ^ n10153 ;
  assign n10211 = n10206 ^ n10161 ;
  assign n10183 = ~n10151 & n10161 ;
  assign n10212 = n10211 ^ n10183 ;
  assign n10179 = n10159 & ~n10165 ;
  assign n10213 = n10212 ^ n10179 ;
  assign n10205 = n10168 ^ n10167 ;
  assign n10214 = n10213 ^ n10205 ;
  assign n10207 = n10206 ^ n10205 ;
  assign n10208 = n10207 ^ n10162 ;
  assign n10209 = n10208 ^ n10161 ;
  assign n10210 = n10209 ^ n10167 ;
  assign n10215 = n10214 ^ n10210 ;
  assign n10216 = n10156 & n10215 ;
  assign n10180 = n10159 & n10163 ;
  assign n10181 = n10180 ^ n10179 ;
  assign n10176 = n10159 & ~n10166 ;
  assign n10178 = n10176 ^ n10159 ;
  assign n10182 = n10181 ^ n10178 ;
  assign n10217 = n10216 ^ n10182 ;
  assign n10201 = n10159 ^ n10151 ;
  assign n10202 = n10201 ^ n10150 ;
  assign n10184 = n10183 ^ n10163 ;
  assign n10203 = n10202 ^ n10184 ;
  assign n10204 = ~n10156 & n10203 ;
  assign n10218 = n10217 ^ n10204 ;
  assign n10219 = ~n10157 & n10218 ;
  assign n10220 = n10219 ^ n10216 ;
  assign n10189 = n10153 ^ n10152 ;
  assign n10190 = ~n10116 & n10189 ;
  assign n10191 = n10190 ^ n10189 ;
  assign n10192 = n10191 ^ n10183 ;
  assign n10193 = n10192 ^ n10170 ;
  assign n10185 = n10184 ^ n10180 ;
  assign n10186 = n10185 ^ n10182 ;
  assign n10187 = n10186 ^ n10168 ;
  assign n10175 = n10167 ^ n10166 ;
  assign n10177 = n10176 ^ n10175 ;
  assign n10188 = n10187 ^ n10177 ;
  assign n10194 = n10193 ^ n10188 ;
  assign n10195 = n10194 ^ n10193 ;
  assign n10196 = n10193 ^ n10156 ;
  assign n10197 = n10196 ^ n10193 ;
  assign n10198 = n10195 & ~n10197 ;
  assign n10199 = n10198 ^ n10193 ;
  assign n10200 = n10155 & ~n10199 ;
  assign n10221 = n10220 ^ n10200 ;
  assign n10222 = ~n10174 & ~n10221 ;
  assign n10224 = n10190 ^ n10185 ;
  assign n10223 = n10179 ^ n10177 ;
  assign n10225 = n10224 ^ n10223 ;
  assign n10226 = n10224 ^ n10155 ;
  assign n10227 = n10226 ^ n10224 ;
  assign n10228 = ~n10225 & n10227 ;
  assign n10229 = n10228 ^ n10224 ;
  assign n10230 = n10156 & n10229 ;
  assign n10231 = n10222 & ~n10230 ;
  assign n10232 = n10231 ^ n6816 ;
  assign n12132 = n10232 ^ x112 ;
  assign n12131 = n10923 ^ x65 ;
  assign n12133 = n12132 ^ n12131 ;
  assign n9481 = n9451 ^ n9400 ;
  assign n9482 = n9286 & n9481 ;
  assign n9483 = n9482 ^ n9400 ;
  assign n9994 = n9285 & n9483 ;
  assign n9433 = n9432 ^ n9415 ;
  assign n9434 = ~n9429 & ~n9433 ;
  assign n9289 = n9288 ^ n9285 ;
  assign n9966 = n9289 & ~n9414 ;
  assign n9967 = ~n9434 & ~n9966 ;
  assign n9476 = n9423 ^ n9400 ;
  assign n9461 = ~n9319 & n9411 ;
  assign n9462 = n9461 ^ n9411 ;
  assign n9964 = n9476 ^ n9462 ;
  assign n9960 = n9424 & n9440 ;
  assign n9951 = n9487 ^ n9423 ;
  assign n9463 = n9462 ^ n9451 ;
  assign n9952 = n9951 ^ n9463 ;
  assign n9953 = n9952 ^ n9487 ;
  assign n9954 = n9487 ^ n9286 ;
  assign n9955 = n9954 ^ n9487 ;
  assign n9956 = n9953 & n9955 ;
  assign n9470 = n9407 ^ n9285 ;
  assign n9471 = n9470 ^ n9407 ;
  assign n9444 = n9410 ^ n9400 ;
  assign n9945 = n9444 ^ n9407 ;
  assign n9946 = ~n9471 & n9945 ;
  assign n9947 = n9946 ^ n9407 ;
  assign n9948 = n9287 & n9947 ;
  assign n9949 = n9948 ^ n9487 ;
  assign n9950 = n9949 ^ n9948 ;
  assign n9957 = n9956 ^ n9950 ;
  assign n9958 = ~n9285 & n9957 ;
  assign n9959 = n9958 ^ n9949 ;
  assign n9961 = n9960 ^ n9959 ;
  assign n9943 = n9424 ^ n9414 ;
  assign n9944 = n9288 & n9943 ;
  assign n9962 = n9961 ^ n9944 ;
  assign n9963 = n9962 ^ n9416 ;
  assign n9965 = n9964 ^ n9963 ;
  assign n9968 = n9967 ^ n9965 ;
  assign n9472 = n9452 ^ n9407 ;
  assign n9473 = n9471 & n9472 ;
  assign n9474 = n9473 ^ n9407 ;
  assign n9475 = n9287 & n9474 ;
  assign n9989 = n9968 ^ n9475 ;
  assign n9983 = n9452 ^ n9421 ;
  assign n9984 = n9421 ^ n9285 ;
  assign n9985 = n9984 ^ n9421 ;
  assign n9986 = ~n9983 & ~n9985 ;
  assign n9987 = n9986 ^ n9421 ;
  assign n9988 = ~n9286 & ~n9987 ;
  assign n9990 = n9989 ^ n9988 ;
  assign n9991 = n9990 ^ n9982 ;
  assign n9992 = n9991 ^ n5965 ;
  assign n9969 = n9968 ^ n9962 ;
  assign n9970 = n9969 ^ n9461 ;
  assign n9971 = n9970 ^ n9969 ;
  assign n9974 = n9285 & n9971 ;
  assign n9975 = n9974 ^ n9969 ;
  assign n9976 = n9287 & n9975 ;
  assign n9993 = n9992 ^ n9976 ;
  assign n9995 = n9994 ^ n9993 ;
  assign n12202 = n9995 ^ x90 ;
  assign n9681 = n8768 ^ n8764 ;
  assign n9680 = n8817 ^ n8808 ;
  assign n9682 = n9681 ^ n9680 ;
  assign n9683 = ~n8684 & n9682 ;
  assign n9684 = n9683 ^ n9681 ;
  assign n9688 = n9684 ^ n8833 ;
  assign n9666 = n8809 ^ n8787 ;
  assign n9665 = n8783 ^ n8776 ;
  assign n9667 = n9666 ^ n9665 ;
  assign n9668 = n9665 ^ n8684 ;
  assign n9669 = n9668 ^ n9665 ;
  assign n9670 = ~n9667 & n9669 ;
  assign n9671 = n9670 ^ n9665 ;
  assign n9672 = ~n8797 & ~n9671 ;
  assign n9689 = n9688 ^ n9672 ;
  assign n9678 = n8819 ^ n8785 ;
  assign n9679 = n9678 ^ n8788 ;
  assign n9685 = n9684 ^ n9679 ;
  assign n9674 = n8785 ^ n8764 ;
  assign n9675 = n9674 ^ n8807 ;
  assign n9676 = n9675 ^ n8819 ;
  assign n9677 = ~n8684 & n9676 ;
  assign n9686 = n9685 ^ n9677 ;
  assign n9687 = n8797 & n9686 ;
  assign n9690 = n9689 ^ n9687 ;
  assign n9673 = n8770 & n9110 ;
  assign n9691 = n9690 ^ n9673 ;
  assign n9692 = n9691 ^ n9672 ;
  assign n9695 = n9691 ^ n8683 ;
  assign n9696 = n9695 ^ n9691 ;
  assign n9697 = n9691 ^ n8772 ;
  assign n9698 = n9697 ^ n9691 ;
  assign n9699 = ~n9696 & n9698 ;
  assign n9700 = ~n9692 & n9699 ;
  assign n9701 = n9700 ^ n9692 ;
  assign n9702 = n9701 ^ n9672 ;
  assign n9703 = ~n9109 & ~n9702 ;
  assign n9704 = ~n9282 & n9703 ;
  assign n9705 = n9704 ^ n4890 ;
  assign n9706 = n9705 ^ x92 ;
  assign n9707 = n9522 ^ x70 ;
  assign n9708 = ~n9706 & n9707 ;
  assign n9709 = n9708 ^ n9707 ;
  assign n9710 = n9709 ^ n9706 ;
  assign n9711 = n8130 ^ x110 ;
  assign n9727 = ~n8502 & n8525 ;
  assign n9724 = n8519 ^ n8502 ;
  assign n9725 = ~n8546 & ~n9724 ;
  assign n9716 = n9001 ^ n8522 ;
  assign n9715 = n8552 ^ n8493 ;
  assign n9717 = n9716 ^ n9715 ;
  assign n9718 = n9716 ^ n8499 ;
  assign n9719 = n9718 ^ n9716 ;
  assign n9720 = n9717 & ~n9719 ;
  assign n9721 = n9720 ^ n9716 ;
  assign n9722 = ~n8505 & n9721 ;
  assign n9723 = n9722 ^ n8528 ;
  assign n9726 = n9725 ^ n9723 ;
  assign n9728 = n9727 ^ n9726 ;
  assign n9737 = n9728 ^ n9008 ;
  assign n9729 = n9728 ^ n9722 ;
  assign n9732 = n9729 ^ n9712 ;
  assign n9733 = n9732 ^ n9729 ;
  assign n9734 = ~n8498 & n9733 ;
  assign n9735 = n9734 ^ n9729 ;
  assign n9736 = n8499 & n9735 ;
  assign n9738 = n9737 ^ n9736 ;
  assign n9713 = n9712 ^ n8508 ;
  assign n9714 = n8500 & n9713 ;
  assign n9739 = n9738 ^ n9714 ;
  assign n9741 = n9740 ^ n8563 ;
  assign n9742 = n9741 ^ n8495 ;
  assign n9745 = n8499 & n9742 ;
  assign n9746 = n9745 ^ n8495 ;
  assign n9747 = n8505 & n9746 ;
  assign n9748 = ~n9739 & ~n9747 ;
  assign n9749 = ~n8561 & n9748 ;
  assign n9751 = ~n8499 & ~n8515 ;
  assign n9752 = n9749 & n9751 ;
  assign n9750 = n9749 ^ n3846 ;
  assign n9753 = n9752 ^ n9750 ;
  assign n9754 = n9753 ^ x77 ;
  assign n9755 = ~n9711 & ~n9754 ;
  assign n9763 = n9755 ^ n9754 ;
  assign n9767 = n9763 ^ n9711 ;
  assign n9768 = n9710 & ~n9767 ;
  assign n9758 = n9710 ^ n9707 ;
  assign n9764 = ~n9758 & ~n9763 ;
  assign n9761 = n9755 ^ n9711 ;
  assign n9762 = ~n9758 & ~n9761 ;
  assign n9765 = n9764 ^ n9762 ;
  assign n9759 = n9755 & ~n9758 ;
  assign n9760 = n9759 ^ n9758 ;
  assign n9766 = n9765 ^ n9760 ;
  assign n9769 = n9768 ^ n9766 ;
  assign n9798 = n9769 ^ n9767 ;
  assign n9775 = n9709 & n9755 ;
  assign n9776 = n9775 ^ n9709 ;
  assign n9777 = n9776 ^ n9707 ;
  assign n9778 = n9767 & n9777 ;
  assign n9790 = n9778 ^ n9777 ;
  assign n9799 = n9798 ^ n9790 ;
  assign n10009 = n9799 ^ n9775 ;
  assign n10010 = n10009 ^ n9790 ;
  assign n9756 = n9710 & n9755 ;
  assign n9815 = n9756 ^ n9710 ;
  assign n9788 = n9710 & ~n9761 ;
  assign n9789 = n9788 ^ n9768 ;
  assign n9816 = n9815 ^ n9789 ;
  assign n10001 = n9816 ^ n9766 ;
  assign n12176 = n10010 ^ n10001 ;
  assign n9795 = n9708 & ~n9761 ;
  assign n10006 = n9795 ^ n9708 ;
  assign n9774 = n9708 & n9755 ;
  assign n9792 = n9790 ^ n9774 ;
  assign n10007 = n10006 ^ n9792 ;
  assign n12194 = n12176 ^ n10007 ;
  assign n9770 = n7659 ^ x109 ;
  assign n9664 = n9558 ^ x91 ;
  assign n9773 = n9770 ^ n9664 ;
  assign n9794 = n9788 ^ n9764 ;
  assign n9796 = n9795 ^ n9794 ;
  assign n9793 = n9765 ^ n9761 ;
  assign n9797 = n9796 ^ n9793 ;
  assign n11406 = n9797 ^ n9759 ;
  assign n11407 = n9759 ^ n9664 ;
  assign n11408 = n11407 ^ n9759 ;
  assign n11409 = ~n11406 & n11408 ;
  assign n11410 = n11409 ^ n9759 ;
  assign n11411 = ~n9773 & n11410 ;
  assign n12195 = n12194 ^ n11411 ;
  assign n9771 = n9664 & n9770 ;
  assign n9824 = n9759 & n9771 ;
  assign n12193 = n9824 ^ n7980 ;
  assign n12196 = n12195 ^ n12193 ;
  assign n12185 = n10007 ^ n9768 ;
  assign n9800 = n9799 ^ n9797 ;
  assign n9801 = n9800 ^ n9776 ;
  assign n9802 = n9801 ^ n9792 ;
  assign n12186 = n12185 ^ n9802 ;
  assign n12187 = n12186 ^ n10007 ;
  assign n12188 = n10007 ^ n9664 ;
  assign n12189 = n12188 ^ n10007 ;
  assign n12190 = ~n12187 & n12189 ;
  assign n12191 = n12190 ^ n10007 ;
  assign n12192 = ~n9770 & n12191 ;
  assign n12197 = n12196 ^ n12192 ;
  assign n11398 = n9801 ^ n9797 ;
  assign n12179 = n11398 ^ n9794 ;
  assign n12180 = n9794 ^ n9770 ;
  assign n12181 = n12180 ^ n9794 ;
  assign n12182 = n12179 & n12181 ;
  assign n12183 = n12182 ^ n9794 ;
  assign n12184 = ~n9664 & n12183 ;
  assign n12198 = n12197 ^ n12184 ;
  assign n12170 = n9768 ^ n9765 ;
  assign n12173 = n12170 ^ n9756 ;
  assign n12169 = n9788 ^ n9759 ;
  assign n12171 = n12170 ^ n12169 ;
  assign n12172 = n9664 & n12171 ;
  assign n12174 = n12173 ^ n12172 ;
  assign n12175 = n12174 ^ n9795 ;
  assign n12177 = n12176 ^ n12175 ;
  assign n12178 = n9773 & ~n12177 ;
  assign n12199 = n12198 ^ n12178 ;
  assign n12200 = n12199 ^ x89 ;
  assign n12205 = n10851 ^ x107 ;
  assign n12164 = n9194 & n10815 ;
  assign n12148 = n9176 ^ n9172 ;
  assign n9205 = n9168 ^ n9167 ;
  assign n12149 = n12148 ^ n9205 ;
  assign n12150 = ~n9019 & n12149 ;
  assign n12160 = n12150 ^ n8026 ;
  assign n9217 = n9198 ^ n9185 ;
  assign n9218 = n9198 ^ n8975 ;
  assign n9219 = n9218 ^ n9198 ;
  assign n9220 = n9217 & ~n9219 ;
  assign n9221 = n9220 ^ n9198 ;
  assign n9222 = ~n9019 & n9221 ;
  assign n12161 = n12160 ^ n9222 ;
  assign n12147 = n9179 ^ n9175 ;
  assign n12151 = n12150 ^ n12147 ;
  assign n12134 = n9170 ^ n9160 ;
  assign n12152 = n12151 ^ n12134 ;
  assign n12153 = n12152 ^ n9175 ;
  assign n12154 = n12153 ^ n12151 ;
  assign n12157 = n9019 & n12154 ;
  assign n12158 = n12157 ^ n12151 ;
  assign n12159 = n9020 & n12158 ;
  assign n12162 = n12161 ^ n12159 ;
  assign n12143 = n9196 ^ n9188 ;
  assign n12146 = n10814 & ~n12143 ;
  assign n12163 = n12162 ^ n12146 ;
  assign n12165 = n12164 ^ n12163 ;
  assign n12144 = n10814 ^ n9019 ;
  assign n12145 = ~n12143 & n12144 ;
  assign n12166 = n12165 ^ n12145 ;
  assign n9203 = n9195 ^ n9186 ;
  assign n12136 = n9203 ^ n9191 ;
  assign n12135 = n12134 ^ n9176 ;
  assign n12137 = n12136 ^ n12135 ;
  assign n12138 = n12135 ^ n9019 ;
  assign n12139 = n12138 ^ n12135 ;
  assign n12140 = ~n12137 & ~n12139 ;
  assign n12141 = n12140 ^ n12135 ;
  assign n12142 = ~n9020 & n12141 ;
  assign n12167 = n12166 ^ n12142 ;
  assign n12168 = n12167 ^ x80 ;
  assign n12219 = n12205 ^ n12168 ;
  assign n12208 = n12168 & ~n12205 ;
  assign n12220 = n12219 ^ n12208 ;
  assign n12228 = n12220 ^ n12168 ;
  assign n12229 = n12200 & n12228 ;
  assign n12230 = n12229 ^ n12168 ;
  assign n12231 = ~n12202 & n12230 ;
  assign n12223 = n12200 & n12202 ;
  assign n12224 = n12223 ^ n12202 ;
  assign n12225 = n12224 ^ n12200 ;
  assign n12226 = ~n12208 & n12225 ;
  assign n12227 = n12226 ^ n12200 ;
  assign n12232 = n12231 ^ n12227 ;
  assign n12233 = n12232 ^ n12225 ;
  assign n12221 = n12220 ^ n12202 ;
  assign n12210 = n12168 & n12202 ;
  assign n12222 = n12221 ^ n12210 ;
  assign n12234 = n12233 ^ n12222 ;
  assign n12235 = n12234 ^ n12210 ;
  assign n12236 = n12235 ^ n12234 ;
  assign n12237 = n12234 ^ n12205 ;
  assign n12238 = n12237 ^ n12234 ;
  assign n12239 = n12236 & n12238 ;
  assign n12240 = n12239 ^ n12234 ;
  assign n12241 = n12132 & n12240 ;
  assign n12242 = n12241 ^ n12232 ;
  assign n12211 = n12210 ^ n12205 ;
  assign n12209 = n12208 ^ n12202 ;
  assign n12212 = n12211 ^ n12209 ;
  assign n12213 = ~n12200 & n12212 ;
  assign n12214 = n12213 ^ n12211 ;
  assign n12203 = n12202 ^ n12200 ;
  assign n12215 = n12214 ^ n12203 ;
  assign n12201 = n12200 ^ n12168 ;
  assign n12204 = ~n12168 & n12203 ;
  assign n12206 = n12205 ^ n12204 ;
  assign n12207 = ~n12201 & n12206 ;
  assign n12216 = n12215 ^ n12207 ;
  assign n12217 = ~n12132 & n12216 ;
  assign n12218 = n12217 ^ n12214 ;
  assign n12243 = n12242 ^ n12218 ;
  assign n12244 = ~n12133 & ~n12243 ;
  assign n12245 = n12244 ^ n12218 ;
  assign n12246 = n12245 ^ n8130 ;
  assign n12751 = n12246 ^ x124 ;
  assign n12752 = n12750 & ~n12751 ;
  assign n12753 = n12752 ^ n12751 ;
  assign n12754 = n12753 ^ n12750 ;
  assign n12755 = n12754 ^ n12751 ;
  assign n12756 = n12755 ^ n12753 ;
  assign n10601 = n8905 & ~n8935 ;
  assign n10597 = n8913 ^ n8849 ;
  assign n10598 = n10597 ^ n8924 ;
  assign n10599 = n8906 & ~n10598 ;
  assign n10590 = n8848 & n8905 ;
  assign n8950 = n8949 ^ n8925 ;
  assign n8951 = ~n8907 & n8950 ;
  assign n10591 = n10590 ^ n8951 ;
  assign n10592 = n10591 ^ n7525 ;
  assign n10593 = n10592 ^ n10589 ;
  assign n10554 = n8916 ^ n8854 ;
  assign n10555 = n10554 ^ n8936 ;
  assign n10556 = n8907 & n10555 ;
  assign n10551 = n8917 ^ n8848 ;
  assign n10552 = n10551 ^ n8938 ;
  assign n10553 = n10552 ^ n8898 ;
  assign n10557 = n10556 ^ n10553 ;
  assign n10558 = n10557 ^ n8898 ;
  assign n10559 = n10558 ^ n10557 ;
  assign n10560 = n10557 ^ n8949 ;
  assign n10561 = n10560 ^ n10557 ;
  assign n10562 = n10559 & n10561 ;
  assign n10563 = n10562 ^ n10557 ;
  assign n10564 = n8580 & ~n10563 ;
  assign n10565 = n10564 ^ n10557 ;
  assign n10594 = n10593 ^ n10565 ;
  assign n10574 = n10573 ^ n8861 ;
  assign n10568 = n8935 ^ n8848 ;
  assign n10575 = n10574 ^ n10568 ;
  assign n10576 = n10575 ^ n10574 ;
  assign n10577 = n10576 ^ n10574 ;
  assign n10578 = n10574 ^ n8580 ;
  assign n10579 = n10578 ^ n10574 ;
  assign n10580 = n10577 & n10579 ;
  assign n10581 = n10580 ^ n10574 ;
  assign n10582 = ~n8898 & ~n10581 ;
  assign n10595 = n10594 ^ n10582 ;
  assign n10550 = n10549 ^ n8925 ;
  assign n10566 = n8940 & n10565 ;
  assign n10567 = ~n10550 & n10566 ;
  assign n10596 = n10595 ^ n10567 ;
  assign n10600 = n10599 ^ n10596 ;
  assign n10602 = n10601 ^ n10600 ;
  assign n10603 = n10602 ^ x70 ;
  assign n8329 = n7916 & ~n8328 ;
  assign n8379 = n7911 & n8331 ;
  assign n8380 = n8326 & n8379 ;
  assign n8333 = n8332 ^ n8327 ;
  assign n8373 = n8372 ^ n8131 ;
  assign n8375 = n8327 & n8373 ;
  assign n8376 = n8375 ^ n8131 ;
  assign n8377 = n8333 & n8376 ;
  assign n8378 = n8377 ^ n8332 ;
  assign n8381 = n8380 ^ n8378 ;
  assign n8409 = n8366 ^ n8351 ;
  assign n8410 = n8409 ^ n8379 ;
  assign n8411 = n8327 & n8410 ;
  assign n8388 = n8361 ^ n8339 ;
  assign n8389 = n8328 & n8388 ;
  assign n8390 = n8389 ^ n8343 ;
  assign n8391 = n8365 ^ n8360 ;
  assign n8392 = ~n8328 & n8391 ;
  assign n8393 = n8392 ^ n8131 ;
  assign n8394 = ~n8390 & ~n8393 ;
  assign n8406 = n8405 ^ n8394 ;
  assign n8385 = n8351 ^ n8347 ;
  assign n8386 = n8385 ^ n8359 ;
  assign n8387 = n8384 & n8386 ;
  assign n8407 = n8406 ^ n8387 ;
  assign n8382 = n8354 ^ n8344 ;
  assign n8383 = n8326 & n8382 ;
  assign n8408 = n8407 ^ n8383 ;
  assign n8412 = n8411 ^ n8408 ;
  assign n8413 = ~n8381 & ~n8412 ;
  assign n8416 = n8366 ^ n8361 ;
  assign n8417 = ~n8415 & n8416 ;
  assign n8418 = n8417 ^ n8361 ;
  assign n8419 = n8131 & n8418 ;
  assign n8420 = n8413 & ~n8419 ;
  assign n8421 = ~n8329 & n8420 ;
  assign n8422 = n8421 ^ n7210 ;
  assign n10604 = n8422 ^ x67 ;
  assign n10605 = n10603 & ~n10604 ;
  assign n10606 = n10605 ^ n10604 ;
  assign n10637 = n10230 ^ n10173 ;
  assign n10620 = n10206 ^ n10170 ;
  assign n10621 = n10620 ^ n10152 ;
  assign n10622 = n10621 ^ n10224 ;
  assign n10623 = n10622 ^ n10150 ;
  assign n10608 = n10207 ^ n10191 ;
  assign n10609 = n10608 ^ n10187 ;
  assign n10626 = n10623 ^ n10609 ;
  assign n10627 = n10156 & ~n10626 ;
  assign n10610 = n10182 ^ n10176 ;
  assign n10611 = n10610 ^ n10172 ;
  assign n10612 = n10171 ^ n10155 ;
  assign n10613 = n10612 ^ n10192 ;
  assign n10616 = n10610 & ~n10613 ;
  assign n10617 = n10616 ^ n10192 ;
  assign n10618 = n10611 & ~n10617 ;
  assign n10619 = n10618 ^ n10172 ;
  assign n10624 = n10623 ^ n10619 ;
  assign n10628 = n10627 ^ n10624 ;
  assign n10638 = n10637 ^ n10628 ;
  assign n10639 = n10638 ^ n7551 ;
  assign n10629 = n10628 ^ n10619 ;
  assign n10630 = n10629 ^ n10194 ;
  assign n10631 = n10630 ^ n10629 ;
  assign n10634 = ~n10156 & ~n10631 ;
  assign n10635 = n10634 ^ n10629 ;
  assign n10636 = ~n10155 & ~n10635 ;
  assign n10640 = n10639 ^ n10636 ;
  assign n10641 = n10640 ^ x77 ;
  assign n10642 = n10343 & n10369 ;
  assign n10643 = n10642 ^ n10370 ;
  assign n10356 = n10346 ^ n10331 ;
  assign n10359 = ~n10336 & n10356 ;
  assign n10360 = n10359 ^ n10331 ;
  assign n10361 = ~n10313 & n10360 ;
  assign n10686 = n10395 & n10685 ;
  assign n10671 = n10372 ^ n10270 ;
  assign n10672 = n10317 ^ n10307 ;
  assign n10673 = n10672 ^ n10308 ;
  assign n10674 = n10671 & ~n10673 ;
  assign n10666 = n10374 ^ n10333 ;
  assign n10670 = n10666 ^ n10325 ;
  assign n10675 = n10674 ^ n10670 ;
  assign n10676 = n10675 ^ n10666 ;
  assign n10677 = n10666 ^ n10336 ;
  assign n10678 = n10677 ^ n10666 ;
  assign n10679 = n10676 & n10678 ;
  assign n10344 = n10343 ^ n10315 ;
  assign n10348 = n10347 ^ n10344 ;
  assign n10349 = n10348 ^ n10329 ;
  assign n10350 = n10349 ^ n10344 ;
  assign n10351 = n10344 ^ n10313 ;
  assign n10352 = n10351 ^ n10344 ;
  assign n10353 = n10350 & ~n10352 ;
  assign n10354 = n10353 ^ n10344 ;
  assign n10355 = n10342 & n10354 ;
  assign n10662 = n10346 & n10355 ;
  assign n10663 = n10662 ^ n10313 ;
  assign n10664 = ~n10392 & ~n10663 ;
  assign n10665 = n10664 ^ n10313 ;
  assign n10667 = n10666 ^ n10665 ;
  assign n10655 = ~n10336 & n10377 ;
  assign n10656 = n10655 ^ n10332 ;
  assign n10657 = n10313 & n10656 ;
  assign n10668 = n10667 ^ n10657 ;
  assign n10669 = n10668 ^ n10665 ;
  assign n10680 = n10679 ^ n10669 ;
  assign n10681 = n10680 ^ n10657 ;
  assign n10682 = n10342 & n10681 ;
  assign n10683 = n10682 ^ n10668 ;
  assign n10687 = n10686 ^ n10683 ;
  assign n10644 = n10366 ^ n10322 ;
  assign n10645 = n10644 ^ n10386 ;
  assign n10646 = n10386 ^ n10313 ;
  assign n10647 = n10646 ^ n10386 ;
  assign n10648 = n10645 & ~n10647 ;
  assign n10649 = n10648 ^ n10386 ;
  assign n10650 = ~n10336 & ~n10649 ;
  assign n10688 = n10687 ^ n10650 ;
  assign n10696 = n10688 & ~n10695 ;
  assign n10697 = ~n10361 & n10696 ;
  assign n10698 = ~n10643 & n10697 ;
  assign n10699 = n10698 ^ n7473 ;
  assign n10700 = n10699 ^ x84 ;
  assign n10701 = n10641 & ~n10700 ;
  assign n10702 = n10701 ^ n10700 ;
  assign n10741 = ~n10606 & ~n10702 ;
  assign n10742 = n10741 ^ n10606 ;
  assign n10704 = n10701 ^ n10641 ;
  assign n10607 = n10606 ^ n10603 ;
  assign n10708 = n10607 ^ n10604 ;
  assign n10713 = n10704 & n10708 ;
  assign n10703 = n10607 & ~n10702 ;
  assign n10726 = n10713 ^ n10703 ;
  assign n10727 = n10726 ^ n10704 ;
  assign n10724 = n10605 & n10704 ;
  assign n10705 = n10607 & n10704 ;
  assign n10706 = n10705 ^ n10703 ;
  assign n10725 = n10724 ^ n10706 ;
  assign n10728 = n10727 ^ n10725 ;
  assign n10778 = n10742 ^ n10728 ;
  assign n10744 = n10605 & ~n10702 ;
  assign n12255 = n10778 ^ n10744 ;
  assign n10047 = ~n9559 & ~n9590 ;
  assign n10052 = n9636 & n10047 ;
  assign n10528 = n9524 ^ n9523 ;
  assign n10058 = n9647 ^ n9635 ;
  assign n10055 = n9652 ^ n9590 ;
  assign n10056 = n9648 & ~n10055 ;
  assign n10057 = n10056 ^ n9649 ;
  assign n10059 = n10058 ^ n10057 ;
  assign n10054 = n9625 ^ n9559 ;
  assign n10060 = n10059 ^ n10054 ;
  assign n10074 = n10060 ^ n10057 ;
  assign n10529 = ~n9523 & n10074 ;
  assign n10530 = n10529 ^ n10057 ;
  assign n10046 = n9633 ^ n9590 ;
  assign n10048 = n10047 ^ n10046 ;
  assign n10049 = n10048 ^ n9559 ;
  assign n10050 = ~n9625 & ~n10049 ;
  assign n10051 = n10050 ^ n9641 ;
  assign n10532 = n10530 ^ n10051 ;
  assign n10068 = n9632 ^ n9625 ;
  assign n10069 = ~n9649 & ~n10068 ;
  assign n10070 = n10069 ^ n9625 ;
  assign n10071 = n9641 & n10070 ;
  assign n10072 = n10071 ^ n9559 ;
  assign n10531 = n10530 ^ n10072 ;
  assign n10533 = n10532 ^ n10531 ;
  assign n10536 = ~n9523 & ~n10533 ;
  assign n10537 = n10536 ^ n10532 ;
  assign n10538 = ~n10528 & ~n10537 ;
  assign n10539 = n10538 ^ n10530 ;
  assign n10540 = ~n10052 & ~n10539 ;
  assign n10541 = n10540 ^ n7596 ;
  assign n10542 = n10541 ^ x116 ;
  assign n9484 = n9483 ^ n9476 ;
  assign n9485 = n9285 & n9484 ;
  assign n9445 = n9444 ^ n9421 ;
  assign n9435 = n9434 ^ n9401 ;
  assign n9446 = n9445 ^ n9435 ;
  assign n9441 = n9408 ^ n9399 ;
  assign n9442 = n9441 ^ n9290 ;
  assign n9443 = n9440 & ~n9442 ;
  assign n9447 = n9446 ^ n9443 ;
  assign n9437 = ~n9426 & ~n9434 ;
  assign n9438 = n9437 ^ n9401 ;
  assign n9439 = n9289 & n9438 ;
  assign n9448 = n9447 ^ n9439 ;
  assign n9477 = n9476 ^ n9448 ;
  assign n9478 = n9477 ^ n9475 ;
  assign n9464 = n9463 ^ n9432 ;
  assign n9467 = n9464 & n9466 ;
  assign n9468 = n9467 ^ n9432 ;
  assign n9469 = n9287 & n9468 ;
  assign n9479 = n9478 ^ n9469 ;
  assign n9449 = n9448 ^ n9443 ;
  assign n9456 = n9449 ^ n9285 ;
  assign n9457 = n9456 ^ n9449 ;
  assign n9458 = n9453 & ~n9457 ;
  assign n9459 = n9458 ^ n9449 ;
  assign n9460 = n9287 & n9459 ;
  assign n9480 = n9479 ^ n9460 ;
  assign n9486 = n9485 ^ n9480 ;
  assign n9494 = ~n9486 & ~n9493 ;
  assign n9495 = n9494 ^ n6931 ;
  assign n10543 = n9495 ^ x102 ;
  assign n10544 = ~n10542 & ~n10543 ;
  assign n11718 = n10544 ^ n10543 ;
  assign n11719 = n10728 & ~n11718 ;
  assign n10709 = ~n10702 & n10708 ;
  assign n10714 = n10709 ^ n10607 ;
  assign n10707 = n10607 & n10701 ;
  assign n10710 = n10709 ^ n10707 ;
  assign n10711 = n10710 ^ n10706 ;
  assign n10715 = n10714 ^ n10711 ;
  assign n10716 = n10715 ^ n10713 ;
  assign n10752 = n10544 & n10716 ;
  assign n11720 = n11719 ^ n10752 ;
  assign n10545 = n10544 ^ n10542 ;
  assign n12275 = ~n10545 & n10711 ;
  assign n12266 = n10724 ^ n10543 ;
  assign n10740 = ~n10606 & n10700 ;
  assign n10743 = n10742 ^ n10740 ;
  assign n10776 = n10743 ^ n10701 ;
  assign n10717 = ~n10641 & n10708 ;
  assign n10718 = n10717 ^ n10709 ;
  assign n10719 = n10718 ^ n10716 ;
  assign n10712 = n10711 ^ n10604 ;
  assign n10720 = n10719 ^ n10712 ;
  assign n10721 = n10720 ^ n10707 ;
  assign n10777 = n10776 ^ n10721 ;
  assign n12258 = n10777 ^ n10741 ;
  assign n12269 = n12258 ^ n10703 ;
  assign n10745 = n10744 ^ n10743 ;
  assign n10722 = n10702 ^ n10641 ;
  assign n10723 = n10605 & n10722 ;
  assign n12267 = n10745 ^ n10723 ;
  assign n12270 = n12269 ^ n12267 ;
  assign n12271 = n10542 & n12270 ;
  assign n12268 = n12267 ^ n10724 ;
  assign n12272 = n12271 ^ n12268 ;
  assign n12273 = n12266 & n12272 ;
  assign n12274 = n12273 ^ n10543 ;
  assign n12276 = n12275 ^ n12274 ;
  assign n10729 = n10728 ^ n10723 ;
  assign n12259 = n12258 ^ n10729 ;
  assign n12256 = n10721 ^ n10715 ;
  assign n12257 = n12256 ^ n10723 ;
  assign n12260 = n12259 ^ n12257 ;
  assign n12261 = n12257 ^ n10542 ;
  assign n12262 = n12261 ^ n12257 ;
  assign n12263 = ~n12260 & ~n12262 ;
  assign n12264 = n12263 ^ n12257 ;
  assign n12265 = ~n10543 & n12264 ;
  assign n12277 = n12276 ^ n12265 ;
  assign n12278 = n10709 ^ n10544 ;
  assign n12279 = n12278 ^ n12277 ;
  assign n12280 = n11718 ^ n10542 ;
  assign n12281 = n12280 ^ n10720 ;
  assign n12282 = ~n10544 & n12281 ;
  assign n12283 = n12282 ^ n10720 ;
  assign n12284 = n12279 & ~n12283 ;
  assign n12285 = n12284 ^ n10544 ;
  assign n12286 = ~n12277 & ~n12285 ;
  assign n12287 = ~n11720 & n12286 ;
  assign n12288 = ~n11718 & n12287 ;
  assign n12289 = ~n12255 & n12288 ;
  assign n12290 = n12289 ^ n12287 ;
  assign n12294 = n12290 ^ n7659 ;
  assign n11690 = n10718 ^ n10705 ;
  assign n12291 = n11690 ^ n10715 ;
  assign n12292 = ~n12280 & n12291 ;
  assign n12293 = n12290 & n12292 ;
  assign n12295 = n12294 ^ n12293 ;
  assign n12757 = n12295 ^ x75 ;
  assign n9998 = n9816 ^ n9790 ;
  assign n9826 = n9771 ^ n9770 ;
  assign n9827 = n9826 ^ n9664 ;
  assign n9828 = n9827 ^ n9770 ;
  assign n9999 = ~n9766 & n9828 ;
  assign n10000 = n9999 ^ n9824 ;
  assign n9829 = n9828 ^ n9762 ;
  assign n9830 = n9826 ^ n9768 ;
  assign n9833 = ~n9828 & ~n9830 ;
  assign n9834 = n9833 ^ n9768 ;
  assign n9835 = n9829 & n9834 ;
  assign n9836 = n9835 ^ n9762 ;
  assign n10014 = n10010 ^ n9795 ;
  assign n10008 = n10007 ^ n9797 ;
  assign n10011 = n10010 ^ n10008 ;
  assign n10012 = n10011 ^ n9756 ;
  assign n10013 = ~n9770 & ~n10012 ;
  assign n10015 = n10014 ^ n10013 ;
  assign n10016 = n9664 & ~n9795 ;
  assign n10017 = ~n10015 & n10016 ;
  assign n10018 = n10017 ^ n9664 ;
  assign n10004 = n9799 ^ n9709 ;
  assign n10005 = n9826 & n10004 ;
  assign n10019 = n10018 ^ n10005 ;
  assign n10002 = n10001 ^ n9788 ;
  assign n10003 = ~n9827 & ~n10002 ;
  assign n10020 = n10019 ^ n10003 ;
  assign n10021 = n10007 ^ n9762 ;
  assign n10024 = n9770 & n10021 ;
  assign n10025 = n10024 ^ n9762 ;
  assign n10026 = ~n9664 & n10025 ;
  assign n10027 = ~n10020 & ~n10026 ;
  assign n9804 = n9794 ^ n9756 ;
  assign n10030 = n9770 & n9804 ;
  assign n10031 = n10030 ^ n9759 ;
  assign n10032 = ~n9773 & n10031 ;
  assign n10033 = n10032 ^ n9759 ;
  assign n10034 = n10027 & n10033 ;
  assign n10035 = n10034 ^ n10027 ;
  assign n10036 = ~n9836 & n10035 ;
  assign n10037 = ~n10000 & n10036 ;
  assign n10038 = n9826 & n10037 ;
  assign n10039 = n9998 & n10038 ;
  assign n10040 = n10039 ^ n10037 ;
  assign n10043 = n10040 ^ n5397 ;
  assign n9997 = n9776 ^ n9774 ;
  assign n10041 = ~n9827 & n10040 ;
  assign n10042 = n9997 & n10041 ;
  assign n10044 = n10043 ^ n10042 ;
  assign n10045 = n10044 ^ x121 ;
  assign n10233 = n10232 ^ x97 ;
  assign n10400 = n10320 & ~n10342 ;
  assign n10396 = n10375 ^ n10368 ;
  assign n10397 = n10396 ^ n10333 ;
  assign n10398 = n10395 & ~n10397 ;
  assign n10393 = ~n10336 & n10392 ;
  assign n10382 = n10381 ^ n10376 ;
  assign n10383 = n10369 & n10382 ;
  assign n10362 = n10361 ^ n10344 ;
  assign n10363 = n10362 ^ n10355 ;
  assign n10335 = n10334 ^ n10316 ;
  assign n10339 = ~n10335 & ~n10336 ;
  assign n10340 = n10339 ^ n10316 ;
  assign n10341 = ~n10313 & n10340 ;
  assign n10364 = n10363 ^ n10341 ;
  assign n10371 = n10370 ^ n10364 ;
  assign n10384 = n10383 ^ n10371 ;
  assign n10394 = n10393 ^ n10384 ;
  assign n10399 = n10398 ^ n10394 ;
  assign n10401 = n10400 ^ n10399 ;
  assign n10402 = ~n10312 & ~n10401 ;
  assign n10403 = n10402 ^ n6624 ;
  assign n10404 = n10403 ^ x88 ;
  assign n10405 = ~n10233 & n10404 ;
  assign n10410 = n10405 ^ n10233 ;
  assign n10081 = n10052 ^ n6165 ;
  assign n10082 = n10081 ^ n10060 ;
  assign n10073 = n10072 ^ n10060 ;
  assign n10075 = n10074 ^ n10073 ;
  assign n10076 = n10074 ^ n9523 ;
  assign n10077 = n10076 ^ n10074 ;
  assign n10078 = ~n10075 & n10077 ;
  assign n10079 = n10078 ^ n10074 ;
  assign n10080 = ~n9524 & ~n10079 ;
  assign n10083 = n10082 ^ n10080 ;
  assign n10053 = n10052 ^ n10051 ;
  assign n10061 = n10060 ^ n10053 ;
  assign n10062 = n10061 ^ n10052 ;
  assign n10063 = n10052 ^ n9524 ;
  assign n10064 = n10063 ^ n10052 ;
  assign n10065 = n10062 & n10064 ;
  assign n10066 = n10065 ^ n10052 ;
  assign n10067 = ~n9523 & n10066 ;
  assign n10084 = n10083 ^ n10067 ;
  assign n10085 = n10084 ^ x115 ;
  assign n10093 = n8389 ^ n8359 ;
  assign n10094 = ~n8327 & ~n8356 ;
  assign n10095 = ~n8354 & ~n10094 ;
  assign n10096 = n10093 & n10095 ;
  assign n10097 = n10096 ^ n10094 ;
  assign n10106 = n10097 ^ n8338 ;
  assign n10102 = n8369 ^ n7437 ;
  assign n10103 = n10102 ^ n8335 ;
  assign n10104 = n10103 ^ n8338 ;
  assign n10105 = ~n8325 & ~n10104 ;
  assign n10107 = n10106 ^ n10105 ;
  assign n10108 = n8131 & ~n10107 ;
  assign n10098 = n10097 ^ n8397 ;
  assign n10100 = n10099 ^ n10098 ;
  assign n10101 = n10100 ^ n8381 ;
  assign n10109 = n10108 ^ n10101 ;
  assign n10086 = n8397 ^ n7916 ;
  assign n10087 = n10086 ^ n8397 ;
  assign n10088 = n8397 ^ n8325 ;
  assign n10089 = n10088 ^ n8397 ;
  assign n10090 = n10087 & n10089 ;
  assign n10091 = n10090 ^ n8397 ;
  assign n10092 = n8395 & n10091 ;
  assign n10110 = n10109 ^ n10092 ;
  assign n10111 = ~n8419 & n10110 ;
  assign n10112 = ~n8329 & n10111 ;
  assign n10113 = n10112 ^ n6395 ;
  assign n10114 = n10113 ^ x114 ;
  assign n10115 = n10085 & n10114 ;
  assign n10417 = n10115 ^ n10085 ;
  assign n10418 = ~n10410 & n10417 ;
  assign n10406 = n10405 ^ n10404 ;
  assign n10407 = n10406 ^ n10233 ;
  assign n10408 = n10115 & n10407 ;
  assign n10435 = n10418 ^ n10408 ;
  assign n10414 = n10115 ^ n10114 ;
  assign n10415 = n10414 ^ n10085 ;
  assign n10416 = n10407 & ~n10415 ;
  assign n10436 = n10435 ^ n10416 ;
  assign n10432 = n10114 ^ n10085 ;
  assign n10433 = ~n10404 & ~n10432 ;
  assign n10434 = n10433 ^ n10410 ;
  assign n10437 = n10436 ^ n10434 ;
  assign n10515 = n10437 ^ n10416 ;
  assign n10411 = ~n10114 & n10407 ;
  assign n10412 = n10411 ^ n10410 ;
  assign n10420 = ~n10085 & ~n10412 ;
  assign n10516 = n10515 ^ n10420 ;
  assign n10431 = n10416 ^ n10411 ;
  assign n10517 = n10516 ^ n10431 ;
  assign n10442 = n10405 & n10414 ;
  assign n10428 = n10405 & ~n10415 ;
  assign n10438 = n10437 ^ n10428 ;
  assign n10439 = n10438 ^ n10415 ;
  assign n10440 = n10439 ^ n10420 ;
  assign n10443 = n10442 ^ n10440 ;
  assign n10444 = n10443 ^ n10428 ;
  assign n10424 = n10115 & n10405 ;
  assign n10445 = n10444 ^ n10424 ;
  assign n10441 = n10440 ^ n10405 ;
  assign n10446 = n10445 ^ n10441 ;
  assign n10447 = n10446 ^ n10431 ;
  assign n10430 = n10418 ^ n10417 ;
  assign n10448 = n10447 ^ n10430 ;
  assign n10518 = n10517 ^ n10448 ;
  assign n9996 = n9995 ^ x82 ;
  assign n10519 = n10448 ^ n9996 ;
  assign n10520 = n10519 ^ n10448 ;
  assign n10521 = ~n10518 & n10520 ;
  assign n10522 = n10521 ^ n10448 ;
  assign n10523 = n10045 & n10522 ;
  assign n10492 = n10448 ^ n10446 ;
  assign n10493 = n10446 ^ n9996 ;
  assign n10494 = n10493 ^ n10446 ;
  assign n10495 = n10492 & n10494 ;
  assign n10496 = n10495 ^ n10446 ;
  assign n10497 = ~n10045 & n10496 ;
  assign n10468 = n10045 ^ n9996 ;
  assign n12779 = n10424 & n10468 ;
  assign n10498 = ~n9996 & n10045 ;
  assign n11724 = n10498 ^ n10045 ;
  assign n12434 = n10446 ^ n10437 ;
  assign n12776 = n11724 & ~n12434 ;
  assign n10421 = n10420 ^ n10410 ;
  assign n10419 = n10418 ^ n10416 ;
  assign n10422 = n10421 ^ n10419 ;
  assign n10409 = n10408 ^ n10404 ;
  assign n10413 = n10412 ^ n10409 ;
  assign n10423 = n10422 ^ n10413 ;
  assign n10425 = n10424 ^ n10423 ;
  assign n10509 = n10424 ^ n10045 ;
  assign n10510 = n10509 ^ n10424 ;
  assign n10511 = ~n10425 & ~n10510 ;
  assign n10512 = n10511 ^ n10424 ;
  assign n10513 = ~n10468 & n10512 ;
  assign n10476 = n10423 ^ n10115 ;
  assign n10449 = n10423 ^ n10416 ;
  assign n10450 = n10449 ^ n10448 ;
  assign n10429 = n10428 ^ n10416 ;
  assign n10451 = n10450 ^ n10429 ;
  assign n10452 = n10451 ^ n10404 ;
  assign n10453 = n10452 ^ n10434 ;
  assign n10426 = n10233 ^ n10085 ;
  assign n10427 = n10426 ^ n10114 ;
  assign n10454 = n10453 ^ n10427 ;
  assign n10455 = n10454 ^ n10425 ;
  assign n10456 = n10455 ^ n10408 ;
  assign n10477 = n10476 ^ n10456 ;
  assign n10478 = n10477 ^ n10454 ;
  assign n10479 = n10478 ^ n10422 ;
  assign n10499 = ~n10479 & n10498 ;
  assign n12774 = n10513 ^ n10499 ;
  assign n12759 = n10456 ^ n10045 ;
  assign n12760 = n12759 ^ n10456 ;
  assign n10489 = n10479 ^ n10428 ;
  assign n12761 = n10455 & ~n10489 ;
  assign n12762 = n12761 ^ n10456 ;
  assign n12763 = n12760 & ~n12762 ;
  assign n12764 = n12763 ^ n10456 ;
  assign n12765 = n9996 & ~n12764 ;
  assign n12766 = n12765 ^ n10455 ;
  assign n12769 = ~n9996 & ~n10453 ;
  assign n12770 = n12769 ^ n10434 ;
  assign n12771 = ~n10468 & ~n12770 ;
  assign n12772 = n12771 ^ n10434 ;
  assign n12773 = n12766 & n12772 ;
  assign n12775 = n12774 ^ n12773 ;
  assign n12777 = n12776 ^ n12775 ;
  assign n11725 = n11724 ^ n9996 ;
  assign n12758 = n10443 & n11725 ;
  assign n12778 = n12777 ^ n12758 ;
  assign n12780 = n12779 ^ n12778 ;
  assign n12781 = ~n10497 & n12780 ;
  assign n12782 = ~n10523 & n12781 ;
  assign n12783 = n12782 ^ n6893 ;
  assign n12784 = n12783 ^ x100 ;
  assign n12785 = n12757 & ~n12784 ;
  assign n11295 = n10640 ^ x99 ;
  assign n11284 = n9182 ^ n9019 ;
  assign n11285 = n9191 ^ n8975 ;
  assign n11288 = ~n9182 & n11285 ;
  assign n11289 = n11288 ^ n8975 ;
  assign n11290 = ~n11284 & ~n11289 ;
  assign n11275 = n9196 ^ n9185 ;
  assign n11276 = n9185 ^ n8975 ;
  assign n11277 = n11276 ^ n9185 ;
  assign n11278 = ~n11275 & n11277 ;
  assign n11279 = n11278 ^ n9185 ;
  assign n11270 = n10785 ^ n9177 ;
  assign n9200 = n9172 ^ n9164 ;
  assign n11266 = n9200 ^ n9176 ;
  assign n11263 = n9172 ^ n9160 ;
  assign n11264 = n11263 ^ n9179 ;
  assign n11265 = ~n8975 & n11264 ;
  assign n11267 = n11266 ^ n11265 ;
  assign n11271 = n11270 ^ n11267 ;
  assign n11272 = n9019 & ~n11271 ;
  assign n11260 = n9191 ^ n9189 ;
  assign n11261 = n11260 ^ n9173 ;
  assign n11262 = n10814 & n11261 ;
  assign n11268 = n11267 ^ n11262 ;
  assign n11269 = n11268 ^ n9167 ;
  assign n11273 = n11272 ^ n11269 ;
  assign n11274 = n11273 ^ n11268 ;
  assign n11280 = n11279 ^ n11274 ;
  assign n11281 = n11280 ^ n11272 ;
  assign n11282 = n9020 & n11281 ;
  assign n11283 = n11282 ^ n11273 ;
  assign n11291 = n11290 ^ n11283 ;
  assign n11292 = ~n10807 & n11291 ;
  assign n11293 = n11292 ^ n7697 ;
  assign n11294 = n11293 ^ x106 ;
  assign n11466 = n11295 ^ n11294 ;
  assign n11387 = n9768 & n9771 ;
  assign n11382 = n9816 ^ n9788 ;
  assign n11383 = n11382 ^ n9816 ;
  assign n11384 = n9796 & n9826 ;
  assign n11385 = ~n11383 & n11384 ;
  assign n11386 = n11385 ^ n11382 ;
  assign n11388 = n11387 ^ n11386 ;
  assign n11412 = n11388 ^ n9775 ;
  assign n9817 = n9816 ^ n9795 ;
  assign n9818 = n9795 ^ n9664 ;
  assign n9819 = n9818 ^ n9795 ;
  assign n9820 = n9817 & ~n9819 ;
  assign n9821 = n9820 ^ n9795 ;
  assign n9822 = ~n9773 & n9821 ;
  assign n11413 = n11412 ^ n9822 ;
  assign n11414 = n11413 ^ n11411 ;
  assign n11415 = n11414 ^ n10026 ;
  assign n11397 = n9828 ^ n9775 ;
  assign n9805 = n9804 ^ n9795 ;
  assign n11399 = n11398 ^ n9805 ;
  assign n11400 = n11399 ^ n9826 ;
  assign n11403 = n9828 & ~n11400 ;
  assign n11404 = n11403 ^ n9826 ;
  assign n11405 = n11397 & ~n11404 ;
  assign n11416 = n11415 ^ n11405 ;
  assign n11389 = n11388 ^ n10006 ;
  assign n11390 = n11389 ^ n9799 ;
  assign n11391 = n11390 ^ n11388 ;
  assign n11392 = n11388 ^ n9664 ;
  assign n11393 = n11392 ^ n11388 ;
  assign n11394 = n11391 & ~n11393 ;
  assign n11395 = n11394 ^ n11388 ;
  assign n11396 = ~n9770 & n11395 ;
  assign n11417 = n11416 ^ n11396 ;
  assign n11381 = ~n9800 & n9826 ;
  assign n11418 = n11417 ^ n11381 ;
  assign n11375 = n9792 ^ n9756 ;
  assign n11376 = n9792 ^ n9770 ;
  assign n11377 = n11376 ^ n9792 ;
  assign n11378 = n11375 & ~n11377 ;
  assign n11379 = n11378 ^ n9792 ;
  assign n11380 = ~n9773 & n11379 ;
  assign n11419 = n11418 ^ n11380 ;
  assign n11420 = ~n10000 & ~n11419 ;
  assign n11421 = n11420 ^ n7773 ;
  assign n11422 = n11421 ^ x113 ;
  assign n11333 = n9406 ^ n9403 ;
  assign n11334 = n11333 ^ n9415 ;
  assign n11335 = n9286 & ~n11334 ;
  assign n11336 = n11335 ^ n9423 ;
  assign n11337 = n9287 & n11336 ;
  assign n11317 = n9461 ^ n9400 ;
  assign n11318 = n11317 ^ n9451 ;
  assign n11305 = n9424 ^ n9421 ;
  assign n11306 = ~n9966 & ~n11305 ;
  assign n11304 = n9429 ^ n9415 ;
  assign n11307 = n11306 ^ n11304 ;
  assign n11308 = n9414 ^ n9406 ;
  assign n11309 = n11308 ^ n9966 ;
  assign n11310 = n11309 ^ n11308 ;
  assign n11311 = n11308 ^ n9415 ;
  assign n11312 = n11311 ^ n11308 ;
  assign n11313 = n11310 & n11312 ;
  assign n11314 = n11313 ^ n11308 ;
  assign n11315 = n11307 & ~n11314 ;
  assign n11302 = n9982 ^ n9429 ;
  assign n11303 = n11302 ^ n9948 ;
  assign n11316 = n11315 ^ n11303 ;
  assign n11319 = n11318 ^ n11316 ;
  assign n11330 = n11319 ^ n9988 ;
  assign n11320 = n11319 ^ n9977 ;
  assign n11321 = n11320 ^ n11316 ;
  assign n11322 = n11321 ^ n9964 ;
  assign n11323 = n11322 ^ n9977 ;
  assign n11324 = n11323 ^ n11321 ;
  assign n11325 = n11321 ^ n9286 ;
  assign n11326 = n11325 ^ n11321 ;
  assign n11327 = n11324 & n11326 ;
  assign n11328 = n11327 ^ n11321 ;
  assign n11329 = n9287 & n11328 ;
  assign n11331 = n11330 ^ n11329 ;
  assign n11301 = n9429 & n9444 ;
  assign n11332 = n11331 ^ n11301 ;
  assign n11338 = n11337 ^ n11332 ;
  assign n11339 = ~n9469 & ~n11338 ;
  assign n11340 = n11339 ^ n7815 ;
  assign n11341 = n11340 ^ x123 ;
  assign n11350 = n10094 ^ n8362 ;
  assign n11351 = n8354 ^ n8346 ;
  assign n11352 = n11351 ^ n10854 ;
  assign n11353 = n8327 & n11352 ;
  assign n11354 = n11353 ^ n8384 ;
  assign n11355 = n11350 & n11354 ;
  assign n11358 = n8361 ^ n8343 ;
  assign n11359 = n8327 & n11358 ;
  assign n11360 = ~n11355 & n11359 ;
  assign n11343 = n8410 ^ n8363 ;
  assign n11344 = n11343 ^ n8350 ;
  assign n11345 = n8350 ^ n8325 ;
  assign n11346 = n11345 ^ n8350 ;
  assign n11347 = n11344 & ~n11346 ;
  assign n11348 = n11347 ^ n8350 ;
  assign n11349 = ~n8395 & n11348 ;
  assign n11356 = n11355 ^ n11349 ;
  assign n11361 = n11360 ^ n11356 ;
  assign n11364 = ~n8325 & n8368 ;
  assign n11365 = n11364 ^ n8360 ;
  assign n11366 = n8395 & n11365 ;
  assign n11367 = n11366 ^ n8360 ;
  assign n11368 = ~n11361 & n11367 ;
  assign n11369 = n11368 ^ n11361 ;
  assign n11370 = ~n10884 & ~n11369 ;
  assign n11371 = ~n10856 & n11370 ;
  assign n11372 = ~n8329 & n11371 ;
  assign n11373 = n11372 ^ n7735 ;
  assign n11374 = n11373 ^ x73 ;
  assign n11300 = n10541 ^ x104 ;
  assign n11428 = n11374 ^ n11300 ;
  assign n11427 = n11300 & ~n11374 ;
  assign n11429 = n11428 ^ n11427 ;
  assign n11430 = n11341 & n11429 ;
  assign n11431 = n11430 ^ n11341 ;
  assign n11342 = n11300 & n11341 ;
  assign n11432 = n11431 ^ n11342 ;
  assign n11447 = n11422 & n11432 ;
  assign n11437 = ~n11341 & n11422 ;
  assign n11445 = n11429 & n11437 ;
  assign n11423 = n11374 & ~n11422 ;
  assign n11425 = n11300 & n11423 ;
  assign n11443 = n11425 ^ n11423 ;
  assign n11444 = n11443 ^ n11429 ;
  assign n11446 = n11445 ^ n11444 ;
  assign n11448 = n11447 ^ n11446 ;
  assign n11439 = ~n11341 & n11427 ;
  assign n11440 = n11439 ^ n11427 ;
  assign n11441 = n11440 ^ n11342 ;
  assign n11424 = n11342 & n11423 ;
  assign n11442 = n11441 ^ n11424 ;
  assign n11449 = n11448 ^ n11442 ;
  assign n11438 = n11437 ^ n11422 ;
  assign n11450 = n11449 ^ n11438 ;
  assign n11469 = n11450 ^ n11440 ;
  assign n11467 = n11446 ^ n11430 ;
  assign n11468 = n11467 ^ n11443 ;
  assign n11470 = n11469 ^ n11468 ;
  assign n11471 = n11469 ^ n11294 ;
  assign n11472 = n11471 ^ n11469 ;
  assign n11473 = n11470 & ~n11472 ;
  assign n11474 = n11473 ^ n11469 ;
  assign n11475 = n11466 & n11474 ;
  assign n12470 = n11448 ^ n11294 ;
  assign n12471 = n12470 ^ n11448 ;
  assign n12472 = n11449 & ~n12471 ;
  assign n12473 = n12472 ^ n11448 ;
  assign n12474 = n11466 & n12473 ;
  assign n11296 = ~n11294 & n11295 ;
  assign n11433 = n11429 ^ n11300 ;
  assign n11434 = n11433 ^ n11432 ;
  assign n11606 = n11296 & ~n11434 ;
  assign n11435 = ~n11422 & ~n11434 ;
  assign n12807 = ~n11294 & n11435 ;
  assign n11297 = n11296 ^ n11295 ;
  assign n11298 = n11297 ^ n11294 ;
  assign n11299 = n11298 ^ n11295 ;
  assign n11454 = n11435 ^ n11434 ;
  assign n11455 = n11454 ^ n11445 ;
  assign n12803 = n11455 ^ n11447 ;
  assign n12804 = ~n11299 & ~n12803 ;
  assign n12789 = n11446 ^ n11440 ;
  assign n11426 = n11425 ^ n11424 ;
  assign n12790 = n12789 ^ n11426 ;
  assign n11452 = n11427 & n11437 ;
  assign n11502 = n11452 ^ n11424 ;
  assign n12488 = n11502 ^ n11469 ;
  assign n12489 = n12488 ^ n11442 ;
  assign n12791 = n12790 ^ n12489 ;
  assign n12792 = n11294 & n12791 ;
  assign n12793 = n12792 ^ n12489 ;
  assign n11499 = n11452 ^ n11439 ;
  assign n11453 = n11452 ^ n11437 ;
  assign n11456 = n11455 ^ n11453 ;
  assign n12491 = n11499 ^ n11456 ;
  assign n12799 = n12793 ^ n12491 ;
  assign n12796 = n12491 ^ n11454 ;
  assign n11451 = n11450 ^ n11424 ;
  assign n11457 = n11456 ^ n11451 ;
  assign n12797 = n12796 ^ n11457 ;
  assign n12798 = n11294 & ~n12797 ;
  assign n12800 = n12799 ^ n12798 ;
  assign n12801 = n11466 & ~n12800 ;
  assign n11501 = n11447 ^ n11432 ;
  assign n11618 = n11501 ^ n11445 ;
  assign n11619 = n11297 & n11618 ;
  assign n12794 = n12793 ^ n11619 ;
  assign n11481 = n11468 ^ n11450 ;
  assign n11482 = n11450 ^ n11294 ;
  assign n11483 = n11482 ^ n11450 ;
  assign n11484 = n11481 & n11483 ;
  assign n11485 = n11484 ^ n11450 ;
  assign n11486 = n11466 & n11485 ;
  assign n12795 = n12794 ^ n11486 ;
  assign n12802 = n12801 ^ n12795 ;
  assign n12805 = n12804 ^ n12802 ;
  assign n12787 = n11467 ^ n11435 ;
  assign n12788 = n11295 & n12787 ;
  assign n12806 = n12805 ^ n12788 ;
  assign n12808 = n12807 ^ n12806 ;
  assign n12809 = ~n11606 & ~n12808 ;
  assign n12810 = ~n12474 & n12809 ;
  assign n12811 = ~n11475 & n12810 ;
  assign n12812 = n12811 ^ n7909 ;
  assign n12813 = n12812 ^ x102 ;
  assign n8423 = n8422 ^ x109 ;
  assign n8948 = n8947 ^ n8911 ;
  assign n8952 = n8951 ^ n8948 ;
  assign n8927 = n8926 ^ n8854 ;
  assign n8928 = n8927 ^ n8617 ;
  assign n8929 = n8928 ^ n8926 ;
  assign n8930 = n8926 ^ n8898 ;
  assign n8931 = n8930 ^ n8926 ;
  assign n8932 = ~n8929 & n8931 ;
  assign n8933 = n8932 ^ n8926 ;
  assign n8934 = ~n8899 & n8933 ;
  assign n8953 = n8952 ^ n8934 ;
  assign n8918 = n8917 ^ n8913 ;
  assign n8919 = ~n8907 & ~n8918 ;
  assign n8954 = n8953 ^ n8919 ;
  assign n8900 = n8859 ^ n8580 ;
  assign n8901 = n8900 ^ n8859 ;
  assign n8902 = ~n8860 & n8901 ;
  assign n8903 = n8902 ^ n8859 ;
  assign n8904 = n8899 & ~n8903 ;
  assign n8955 = n8954 ^ n8904 ;
  assign n8956 = n8955 ^ n7355 ;
  assign n8862 = n8861 ^ n8856 ;
  assign n8863 = ~n8580 & n8862 ;
  assign n8957 = n8956 ^ n8863 ;
  assign n8958 = n8957 ^ x118 ;
  assign n8959 = n8423 & ~n8958 ;
  assign n9235 = n9234 ^ n9222 ;
  assign n9207 = n9206 ^ n9205 ;
  assign n9202 = n9173 ^ n9160 ;
  assign n9208 = n9207 ^ n9202 ;
  assign n9209 = n9019 & n9208 ;
  assign n9204 = n9203 ^ n9202 ;
  assign n9210 = n9209 ^ n9204 ;
  assign n9236 = n9235 ^ n9210 ;
  assign n9237 = n9236 ^ n7129 ;
  assign n9199 = n9198 ^ n9169 ;
  assign n9201 = n9200 ^ n9199 ;
  assign n9211 = n9210 ^ n9201 ;
  assign n9212 = n9211 ^ n9210 ;
  assign n9183 = n9182 ^ n9180 ;
  assign n9197 = n9196 ^ n9183 ;
  assign n9213 = n9212 ^ n9197 ;
  assign n9214 = ~n9019 & ~n9213 ;
  assign n9215 = n9214 ^ n9211 ;
  assign n9216 = ~n9020 & ~n9215 ;
  assign n9238 = n9237 ^ n9216 ;
  assign n9239 = n9238 ^ x85 ;
  assign n9496 = n9495 ^ x100 ;
  assign n9497 = ~n9239 & n9496 ;
  assign n9498 = n9497 ^ n9496 ;
  assign n9499 = n9498 ^ n9239 ;
  assign n9662 = n9661 ^ n7146 ;
  assign n9663 = n9662 ^ x91 ;
  assign n9825 = n9824 ^ n6963 ;
  assign n9837 = n9836 ^ n9825 ;
  assign n9803 = n9802 ^ n9764 ;
  assign n9806 = n9805 ^ n9803 ;
  assign n9809 = n9806 ^ n9776 ;
  assign n9791 = n9790 ^ n9789 ;
  assign n9807 = n9806 ^ n9791 ;
  assign n9808 = n9770 & ~n9807 ;
  assign n9810 = n9809 ^ n9808 ;
  assign n9811 = ~n9664 & ~n9810 ;
  assign n9786 = n9764 & ~n9770 ;
  assign n9779 = n9778 ^ n9774 ;
  assign n9780 = n9778 ^ n9770 ;
  assign n9781 = n9780 ^ n9778 ;
  assign n9782 = n9779 & ~n9781 ;
  assign n9783 = n9782 ^ n9778 ;
  assign n9784 = n9773 & n9783 ;
  assign n9785 = n9784 ^ n9776 ;
  assign n9787 = n9786 ^ n9785 ;
  assign n9812 = n9811 ^ n9787 ;
  assign n9772 = ~n9769 & n9771 ;
  assign n9813 = n9812 ^ n9772 ;
  assign n9757 = n9664 & n9756 ;
  assign n9814 = n9813 ^ n9757 ;
  assign n9823 = ~n9814 & ~n9822 ;
  assign n9838 = n9837 ^ n9823 ;
  assign n9839 = n9838 ^ x78 ;
  assign n9840 = ~n9663 & ~n9839 ;
  assign n9861 = n9499 & n9840 ;
  assign n9860 = n9497 & n9840 ;
  assign n9862 = n9861 ^ n9860 ;
  assign n9846 = n9840 ^ n9839 ;
  assign n9856 = n9498 & ~n9846 ;
  assign n9859 = n9856 ^ n9846 ;
  assign n9863 = n9862 ^ n9859 ;
  assign n9845 = n9497 ^ n9239 ;
  assign n9855 = n9840 & ~n9845 ;
  assign n9857 = n9856 ^ n9855 ;
  assign n9858 = n9857 ^ n9839 ;
  assign n9864 = n9863 ^ n9858 ;
  assign n9865 = n9864 ^ n9855 ;
  assign n12422 = n8959 & n9865 ;
  assign n12836 = n12422 ^ n7436 ;
  assign n9877 = n9499 & ~n9846 ;
  assign n9870 = n9497 & ~n9846 ;
  assign n9878 = n9877 ^ n9870 ;
  assign n9879 = n9878 ^ n9859 ;
  assign n9880 = n9879 ^ n9857 ;
  assign n9841 = n9840 ^ n9663 ;
  assign n9843 = n9497 & ~n9841 ;
  assign n9866 = n9865 ^ n9843 ;
  assign n9851 = ~n9239 & ~n9839 ;
  assign n9852 = n9851 ^ n9496 ;
  assign n9853 = n9663 & n9852 ;
  assign n9854 = n9853 ^ n9852 ;
  assign n9867 = n9866 ^ n9854 ;
  assign n9847 = n9846 ^ n9663 ;
  assign n9848 = ~n9845 & ~n9847 ;
  assign n9868 = n9867 ^ n9848 ;
  assign n9871 = n9870 ^ n9868 ;
  assign n9872 = n9871 ^ n9861 ;
  assign n9869 = n9868 ^ n9866 ;
  assign n9873 = n9872 ^ n9869 ;
  assign n9850 = n9840 ^ n9497 ;
  assign n9874 = n9873 ^ n9850 ;
  assign n9881 = n9880 ^ n9874 ;
  assign n9876 = n9855 ^ n9853 ;
  assign n9882 = n9881 ^ n9876 ;
  assign n9888 = n8959 & ~n9882 ;
  assign n8960 = n8959 ^ n8423 ;
  assign n9842 = n9499 & ~n9841 ;
  assign n9844 = n9843 ^ n9842 ;
  assign n9883 = n9882 ^ n9844 ;
  assign n9884 = n9883 ^ n9847 ;
  assign n9849 = n9848 ^ n9844 ;
  assign n9875 = n9874 ^ n9849 ;
  assign n9885 = n9884 ^ n9875 ;
  assign n9886 = n9885 ^ n9856 ;
  assign n9887 = n8960 & n9886 ;
  assign n9889 = n9888 ^ n9887 ;
  assign n9899 = n8959 ^ n8958 ;
  assign n11675 = n9899 ^ n8960 ;
  assign n12830 = n9885 ^ n9879 ;
  assign n12831 = n12830 ^ n9860 ;
  assign n9891 = n9867 ^ n9841 ;
  assign n9892 = n9891 ^ n9844 ;
  assign n9907 = n9892 ^ n9867 ;
  assign n12819 = n9907 ^ n9874 ;
  assign n12832 = n12831 ^ n12819 ;
  assign n12833 = n11675 & n12832 ;
  assign n12815 = n9870 ^ n9861 ;
  assign n12814 = n9883 ^ n9867 ;
  assign n12816 = n12815 ^ n12814 ;
  assign n12817 = ~n8423 & ~n12816 ;
  assign n12818 = n12817 ^ n12815 ;
  assign n11658 = n9860 ^ n9842 ;
  assign n12826 = n12818 ^ n11658 ;
  assign n12823 = n9848 ^ n9843 ;
  assign n12824 = n12823 ^ n11658 ;
  assign n12825 = n8423 & n12824 ;
  assign n12827 = n12826 ^ n12825 ;
  assign n12828 = ~n8958 & n12827 ;
  assign n12820 = n12819 ^ n12818 ;
  assign n12416 = n9870 ^ n8958 ;
  assign n12417 = n12416 ^ n9870 ;
  assign n12418 = n9878 & ~n12417 ;
  assign n12419 = n12418 ^ n9870 ;
  assign n12420 = ~n8423 & n12419 ;
  assign n12821 = n12820 ^ n12420 ;
  assign n11676 = n9857 ^ n8423 ;
  assign n11677 = n11676 ^ n9857 ;
  assign n11680 = ~n9880 & n11677 ;
  assign n11681 = n11680 ^ n9857 ;
  assign n11682 = ~n11675 & n11681 ;
  assign n12822 = n12821 ^ n11682 ;
  assign n12829 = n12828 ^ n12822 ;
  assign n12834 = n12833 ^ n12829 ;
  assign n12835 = ~n9889 & n12834 ;
  assign n12837 = n12836 ^ n12835 ;
  assign n12838 = n12837 ^ x117 ;
  assign n12839 = n12813 & n12838 ;
  assign n12846 = n12839 ^ n12813 ;
  assign n12852 = n12846 ^ n12838 ;
  assign n12876 = n12785 & ~n12852 ;
  assign n12786 = n12785 ^ n12757 ;
  assign n12842 = n12786 & n12839 ;
  assign n12877 = n12876 ^ n12842 ;
  assign n12848 = n12785 ^ n12784 ;
  assign n12859 = n12846 & ~n12848 ;
  assign n12849 = n12839 & ~n12848 ;
  assign n12869 = n12859 ^ n12849 ;
  assign n12840 = n12839 ^ n12838 ;
  assign n12867 = n12840 & ~n12848 ;
  assign n12868 = n12867 ^ n12848 ;
  assign n12870 = n12869 ^ n12868 ;
  assign n12844 = n12786 ^ n12784 ;
  assign n12847 = n12844 & n12846 ;
  assign n12871 = n12870 ^ n12847 ;
  assign n12865 = n12785 & n12840 ;
  assign n12872 = n12871 ^ n12865 ;
  assign n12873 = n12872 ^ n12846 ;
  assign n12861 = ~n12785 & n12846 ;
  assign n12874 = n12873 ^ n12861 ;
  assign n12875 = n12874 ^ n12872 ;
  assign n12878 = n12877 ^ n12875 ;
  assign n12879 = n12878 ^ n12757 ;
  assign n12860 = n12859 ^ n12847 ;
  assign n12862 = n12861 ^ n12860 ;
  assign n12853 = n12844 & ~n12852 ;
  assign n12854 = n12853 ^ n12849 ;
  assign n12855 = n12854 ^ n12844 ;
  assign n12850 = n12849 ^ n12847 ;
  assign n12845 = n12840 & n12844 ;
  assign n12851 = n12850 ^ n12845 ;
  assign n12856 = n12855 ^ n12851 ;
  assign n12857 = n12856 ^ n12849 ;
  assign n12843 = n12842 ^ n12839 ;
  assign n12858 = n12857 ^ n12843 ;
  assign n12863 = n12862 ^ n12858 ;
  assign n12841 = n12786 & n12840 ;
  assign n12864 = n12863 ^ n12841 ;
  assign n12866 = n12865 ^ n12864 ;
  assign n12880 = n12879 ^ n12866 ;
  assign n12881 = n12880 ^ n12850 ;
  assign n12882 = n12850 ^ n12750 ;
  assign n12883 = n12882 ^ n12850 ;
  assign n12884 = n12881 & ~n12883 ;
  assign n12885 = n12884 ^ n12850 ;
  assign n12886 = n12756 & n12885 ;
  assign n13615 = ~n12753 & n12854 ;
  assign n13632 = n12867 ^ n12850 ;
  assign n13633 = n12754 & n13632 ;
  assign n13628 = n12867 ^ n12853 ;
  assign n13629 = n12755 & n13628 ;
  assign n13621 = n12871 ^ n12859 ;
  assign n13622 = n13621 ^ n12874 ;
  assign n13623 = n13622 ^ n12876 ;
  assign n13624 = n12750 & n13623 ;
  assign n13619 = n12878 ^ n12862 ;
  assign n13620 = n13619 ^ n12856 ;
  assign n13625 = n13624 ^ n13620 ;
  assign n13626 = n13625 ^ n12870 ;
  assign n13630 = n13629 ^ n13626 ;
  assign n13616 = n12880 ^ n12859 ;
  assign n13617 = n13616 ^ n12858 ;
  assign n13618 = n13617 ^ n12841 ;
  assign n13627 = n13626 ^ n13618 ;
  assign n13631 = n13630 ^ n13627 ;
  assign n13634 = n13633 ^ n13631 ;
  assign n12920 = n12870 ^ n12845 ;
  assign n12905 = n12876 ^ n12841 ;
  assign n13635 = n12920 ^ n12905 ;
  assign n13636 = n12920 ^ n12750 ;
  assign n13637 = n13636 ^ n12920 ;
  assign n13638 = ~n13635 & ~n13637 ;
  assign n13639 = n13638 ^ n12920 ;
  assign n13640 = ~n13634 & n13639 ;
  assign n13641 = n13640 ^ n13630 ;
  assign n13642 = n12756 & n13641 ;
  assign n13643 = n13642 ^ n13630 ;
  assign n13644 = ~n13615 & n13643 ;
  assign n13645 = ~n12886 & n13644 ;
  assign n13646 = n13645 ^ n11373 ;
  assign n13647 = n13646 ^ x98 ;
  assign n11053 = n11018 ^ n10994 ;
  assign n11054 = ~n10984 & ~n11053 ;
  assign n13369 = n11054 ^ n10269 ;
  assign n10986 = n10985 ^ n10983 ;
  assign n13340 = n11014 ^ n10968 ;
  assign n13341 = n13340 ^ n10994 ;
  assign n13339 = n10989 ^ n10971 ;
  assign n13342 = n13341 ^ n13339 ;
  assign n13343 = n13341 ^ n10818 ;
  assign n13344 = n13343 ^ n13341 ;
  assign n13345 = n13342 & n13344 ;
  assign n13346 = n13345 ^ n13341 ;
  assign n13347 = n10986 & n13346 ;
  assign n11040 = n10998 ^ n10818 ;
  assign n11041 = n11040 ^ n10998 ;
  assign n11044 = n10999 & ~n11041 ;
  assign n11045 = n11044 ^ n10998 ;
  assign n11046 = n10986 & n11045 ;
  assign n13348 = n13347 ^ n11046 ;
  assign n13336 = n10971 ^ n10968 ;
  assign n10978 = n10977 ^ n10968 ;
  assign n13334 = n11021 ^ n10978 ;
  assign n13335 = n10852 & n13334 ;
  assign n13337 = n13336 ^ n13335 ;
  assign n13338 = ~n10818 & n13337 ;
  assign n13349 = n13348 ^ n13338 ;
  assign n13350 = ~n10852 & ~n13349 ;
  assign n13351 = n10993 ^ n10818 ;
  assign n13352 = n13351 ^ n10993 ;
  assign n13355 = ~n11064 & ~n13352 ;
  assign n13356 = n13355 ^ n10993 ;
  assign n13357 = n13350 & n13356 ;
  assign n13358 = n13357 ^ n13349 ;
  assign n13359 = n11035 ^ n10985 ;
  assign n13360 = n11012 ^ n11010 ;
  assign n13361 = n13360 ^ n10983 ;
  assign n13364 = ~n11035 & ~n13361 ;
  assign n13365 = n13364 ^ n10983 ;
  assign n13366 = ~n13359 & n13365 ;
  assign n13367 = n13366 ^ n10985 ;
  assign n13368 = ~n13358 & n13367 ;
  assign n13370 = n13369 ^ n13368 ;
  assign n13371 = n13370 ^ x105 ;
  assign n11799 = n11373 ^ x122 ;
  assign n11850 = n11293 ^ x81 ;
  assign n11851 = n10044 ^ x72 ;
  assign n11852 = n11850 & n11851 ;
  assign n11853 = n11852 ^ n11850 ;
  assign n11854 = n11853 ^ n11851 ;
  assign n11139 = n10210 ^ n10180 ;
  assign n11140 = n10180 ^ n10156 ;
  assign n11141 = n11140 ^ n10180 ;
  assign n11142 = n11139 & n11141 ;
  assign n11143 = n11142 ^ n10180 ;
  assign n11144 = ~n10157 & n11143 ;
  assign n11809 = n10185 ^ n10170 ;
  assign n11810 = n11809 ^ n10223 ;
  assign n11811 = ~n10172 & ~n11810 ;
  assign n11814 = n11811 ^ n10208 ;
  assign n11114 = n10177 & ~n10612 ;
  assign n11812 = ~n10186 & ~n11811 ;
  assign n11813 = n11114 & n11812 ;
  assign n11815 = n11814 ^ n11813 ;
  assign n11819 = n11815 ^ n10174 ;
  assign n11806 = n10210 ^ n10191 ;
  assign n11804 = n10184 ^ n10179 ;
  assign n11805 = n10171 & n11804 ;
  assign n11807 = n11806 ^ n11805 ;
  assign n11808 = n11807 ^ n10212 ;
  assign n11816 = n11815 ^ n11808 ;
  assign n11801 = n10212 ^ n10190 ;
  assign n11802 = n11801 ^ n10610 ;
  assign n11803 = ~n10156 & n11802 ;
  assign n11817 = n11816 ^ n11803 ;
  assign n11818 = ~n10157 & ~n11817 ;
  assign n11820 = n11819 ^ n11818 ;
  assign n11821 = ~n11144 & n11820 ;
  assign n11822 = n11821 ^ n8486 ;
  assign n11823 = n11822 ^ x98 ;
  assign n11828 = n8935 ^ n8858 ;
  assign n11829 = n8898 & n11828 ;
  assign n11830 = n11829 ^ n8912 ;
  assign n11831 = n11830 ^ n8849 ;
  assign n11839 = n11831 ^ n10839 ;
  assign n11833 = n10571 ^ n8861 ;
  assign n11834 = n11833 ^ n8936 ;
  assign n11825 = n10597 ^ n10546 ;
  assign n11826 = n11825 ^ n10575 ;
  assign n11824 = n8842 ^ n8617 ;
  assign n11827 = n11826 ^ n11824 ;
  assign n11835 = n11834 ^ n11827 ;
  assign n11836 = ~n8898 & ~n11835 ;
  assign n11832 = n11831 ^ n11827 ;
  assign n11837 = n11836 ^ n11832 ;
  assign n11838 = n8580 & n11837 ;
  assign n11840 = n11839 ^ n11838 ;
  assign n11841 = ~n10591 & ~n11840 ;
  assign n11842 = ~n10589 & n11841 ;
  assign n11844 = n8899 & ~n10846 ;
  assign n11845 = n11842 & n11844 ;
  assign n11843 = n11842 ^ n8447 ;
  assign n11846 = n11845 ^ n11843 ;
  assign n11847 = n11846 ^ x120 ;
  assign n11848 = n11823 & n11847 ;
  assign n11858 = n11848 ^ n11823 ;
  assign n11859 = n11858 ^ n11847 ;
  assign n11895 = ~n11854 & ~n11859 ;
  assign n11849 = n11848 ^ n11847 ;
  assign n11875 = n11849 & n11852 ;
  assign n11865 = n11851 ^ n11850 ;
  assign n11866 = n11858 ^ n11851 ;
  assign n11867 = n11865 & ~n11866 ;
  assign n11868 = n11867 ^ n11853 ;
  assign n11863 = n11854 ^ n11850 ;
  assign n11864 = n11858 & n11863 ;
  assign n11869 = n11868 ^ n11864 ;
  assign n11862 = n11848 & n11853 ;
  assign n11870 = n11869 ^ n11862 ;
  assign n11876 = n11875 ^ n11870 ;
  assign n11856 = n11848 & n11852 ;
  assign n11877 = n11876 ^ n11856 ;
  assign n11873 = n11852 & n11858 ;
  assign n11860 = n11853 & ~n11859 ;
  assign n11871 = n11860 ^ n11853 ;
  assign n11872 = n11871 ^ n11870 ;
  assign n11874 = n11873 ^ n11872 ;
  assign n11878 = n11877 ^ n11874 ;
  assign n11861 = n11860 ^ n11850 ;
  assign n11879 = n11878 ^ n11861 ;
  assign n11896 = n11895 ^ n11879 ;
  assign n11894 = n11860 ^ n11859 ;
  assign n11897 = n11896 ^ n11894 ;
  assign n11890 = n11873 ^ n11858 ;
  assign n11891 = n11890 ^ n11868 ;
  assign n11887 = n11849 & n11863 ;
  assign n11888 = n11887 ^ n11869 ;
  assign n11855 = n11849 & ~n11854 ;
  assign n11889 = n11888 ^ n11855 ;
  assign n11892 = n11891 ^ n11889 ;
  assign n11893 = n11892 ^ n11875 ;
  assign n11898 = n11897 ^ n11893 ;
  assign n11899 = n11898 ^ n11866 ;
  assign n11857 = n11856 ^ n11855 ;
  assign n11880 = n11879 ^ n11857 ;
  assign n11900 = n11899 ^ n11880 ;
  assign n11886 = n11869 ^ n11856 ;
  assign n11901 = n11900 ^ n11886 ;
  assign n11885 = n11870 ^ n11848 ;
  assign n11902 = n11901 ^ n11885 ;
  assign n11921 = n11902 ^ n11864 ;
  assign n11922 = n11921 ^ n11887 ;
  assign n11798 = n10403 ^ x66 ;
  assign n11923 = n11887 ^ n11798 ;
  assign n11924 = n11923 ^ n11887 ;
  assign n11925 = ~n11922 & n11924 ;
  assign n11926 = n11925 ^ n11887 ;
  assign n11927 = ~n11799 & n11926 ;
  assign n13403 = n11891 ^ n11856 ;
  assign n13389 = n11873 ^ n11871 ;
  assign n12120 = n11897 ^ n11891 ;
  assign n13390 = n13389 ^ n12120 ;
  assign n13391 = n13390 ^ n11855 ;
  assign n13392 = n11798 & ~n13391 ;
  assign n13393 = n13392 ^ n11871 ;
  assign n13404 = n13403 ^ n13393 ;
  assign n11944 = ~n11798 & ~n11799 ;
  assign n11945 = n11944 ^ n11799 ;
  assign n12085 = n11945 ^ n11798 ;
  assign n12086 = n12085 ^ n11799 ;
  assign n12087 = n11897 ^ n11873 ;
  assign n12088 = ~n12086 & ~n12087 ;
  assign n11939 = n11879 ^ n11799 ;
  assign n11940 = n11939 ^ n11879 ;
  assign n11941 = n11896 & ~n11940 ;
  assign n11942 = n11941 ^ n11879 ;
  assign n11943 = ~n11798 & n11942 ;
  assign n13402 = n12088 ^ n11943 ;
  assign n13405 = n13404 ^ n13402 ;
  assign n11800 = n11799 ^ n11798 ;
  assign n12096 = n11887 ^ n11879 ;
  assign n12097 = ~n11798 & n12096 ;
  assign n12098 = n12097 ^ n11879 ;
  assign n12101 = n12098 ^ n11862 ;
  assign n12102 = n12101 ^ n11856 ;
  assign n12103 = n12102 ^ n12098 ;
  assign n12104 = n11798 & n12103 ;
  assign n12105 = n12104 ^ n12098 ;
  assign n12106 = ~n11800 & n12105 ;
  assign n12107 = n12106 ^ n12098 ;
  assign n13406 = n13405 ^ n12107 ;
  assign n13394 = n13393 ^ n11873 ;
  assign n13395 = n13394 ^ n11889 ;
  assign n13396 = n13395 ^ n13393 ;
  assign n13399 = n11798 & n13396 ;
  assign n13400 = n13399 ^ n13393 ;
  assign n13401 = ~n11799 & n13400 ;
  assign n13407 = n13406 ^ n13401 ;
  assign n13382 = n11944 ^ n11891 ;
  assign n13383 = n12086 ^ n11867 ;
  assign n13386 = n11891 & n13383 ;
  assign n13387 = n13386 ^ n11867 ;
  assign n13388 = n13382 & n13387 ;
  assign n13408 = n13407 ^ n13388 ;
  assign n11951 = n11875 ^ n11860 ;
  assign n13375 = n11856 ^ n11798 ;
  assign n13376 = n13375 ^ n11856 ;
  assign n13379 = n11951 & n13376 ;
  assign n13380 = n13379 ^ n11856 ;
  assign n13381 = n11799 & n13380 ;
  assign n13409 = n13408 ^ n13381 ;
  assign n13410 = ~n11927 & ~n13409 ;
  assign n13411 = n13410 ^ n10306 ;
  assign n13412 = n13411 ^ x115 ;
  assign n13422 = ~n13371 & ~n13412 ;
  assign n11145 = n11144 ^ n8753 ;
  assign n11119 = n10190 ^ n10180 ;
  assign n11118 = n10212 ^ n10192 ;
  assign n11120 = n11119 ^ n11118 ;
  assign n11121 = ~n10156 & n11120 ;
  assign n11122 = n11121 ^ n11119 ;
  assign n11127 = n11122 ^ n10230 ;
  assign n11123 = n11122 ^ n10176 ;
  assign n11115 = n10186 ^ n10154 ;
  assign n11116 = n11115 ^ n10172 ;
  assign n11117 = ~n11114 & n11116 ;
  assign n11124 = n11123 ^ n11117 ;
  assign n11111 = n10170 ^ n10167 ;
  assign n11112 = n11111 ^ n10212 ;
  assign n11113 = n10155 & ~n11112 ;
  assign n11125 = n11124 ^ n11113 ;
  assign n11126 = n10157 & n11125 ;
  assign n11128 = n11127 ^ n11126 ;
  assign n11110 = n10171 & ~n10620 ;
  assign n11129 = n11128 ^ n11110 ;
  assign n11131 = n10169 ^ n10154 ;
  assign n11130 = n10223 ^ n10154 ;
  assign n11132 = n11131 ^ n11130 ;
  assign n11133 = n11131 ^ n10156 ;
  assign n11134 = n11133 ^ n11131 ;
  assign n11135 = ~n11132 & ~n11134 ;
  assign n11136 = n11135 ^ n11131 ;
  assign n11137 = ~n10155 & n11136 ;
  assign n11138 = ~n11129 & ~n11137 ;
  assign n11146 = n11145 ^ n11138 ;
  assign n11147 = n11146 ^ x125 ;
  assign n11160 = n10665 ^ n10379 ;
  assign n11161 = n11160 ^ n10657 ;
  assign n11162 = n11161 ^ n10643 ;
  assign n11163 = n11162 ^ n10341 ;
  assign n11164 = n11163 ^ n8722 ;
  assign n11159 = ~n10336 & n10390 ;
  assign n11165 = n11164 ^ n11159 ;
  assign n11153 = n10889 ^ n10390 ;
  assign n11154 = n11153 ^ n10674 ;
  assign n11155 = n10336 & n11154 ;
  assign n11157 = n11155 ^ n10389 ;
  assign n11158 = n10313 & ~n11157 ;
  assign n11166 = n11165 ^ n11158 ;
  assign n11148 = n10374 ^ n10319 ;
  assign n11149 = n11148 ^ n10374 ;
  assign n11150 = n10903 & n11149 ;
  assign n11151 = n11150 ^ n10374 ;
  assign n11152 = ~n10336 & ~n11151 ;
  assign n11167 = n11166 ^ n11152 ;
  assign n11168 = n11167 ^ x110 ;
  assign n11169 = ~n11147 & ~n11168 ;
  assign n11170 = n11169 ^ n11147 ;
  assign n11106 = n8957 ^ x108 ;
  assign n11107 = n10817 ^ x83 ;
  assign n11108 = ~n11106 & n11107 ;
  assign n11173 = n11108 ^ n11107 ;
  assign n11174 = n11173 ^ n11106 ;
  assign n11175 = ~n11170 & n11174 ;
  assign n11109 = n11108 ^ n11106 ;
  assign n11171 = n11170 ^ n11168 ;
  assign n11172 = ~n11109 & ~n11171 ;
  assign n11176 = n11175 ^ n11172 ;
  assign n11103 = n10963 ^ x69 ;
  assign n11104 = n9838 ^ x86 ;
  assign n11226 = ~n11103 & n11104 ;
  assign n11256 = n11176 & n11226 ;
  assign n11227 = n11226 ^ n11103 ;
  assign n11252 = n11227 ^ n11104 ;
  assign n11200 = n11169 & n11174 ;
  assign n11211 = n11200 ^ n11172 ;
  assign n11203 = ~n11109 & n11169 ;
  assign n11212 = n11211 ^ n11203 ;
  assign n11213 = n11212 ^ n11109 ;
  assign n11179 = n11169 ^ n11168 ;
  assign n11189 = n11173 & ~n11179 ;
  assign n11180 = n11108 & ~n11179 ;
  assign n11197 = n11189 ^ n11180 ;
  assign n11195 = n11174 & ~n11179 ;
  assign n11196 = n11195 ^ n11179 ;
  assign n11198 = n11197 ^ n11196 ;
  assign n11201 = n11200 ^ n11198 ;
  assign n11214 = n11213 ^ n11201 ;
  assign n11253 = n11214 ^ n11195 ;
  assign n11254 = n11252 & n11253 ;
  assign n11184 = n11108 & n11169 ;
  assign n11229 = n11184 ^ n11108 ;
  assign n11230 = ~n11104 & n11229 ;
  assign n11185 = n11184 ^ n11176 ;
  assign n11182 = n11108 & ~n11170 ;
  assign n11178 = ~n11171 & n11173 ;
  assign n11183 = n11182 ^ n11178 ;
  assign n11186 = n11185 ^ n11183 ;
  assign n11181 = n11180 ^ n11178 ;
  assign n11187 = n11186 ^ n11181 ;
  assign n11177 = n11176 ^ n11108 ;
  assign n11188 = n11187 ^ n11177 ;
  assign n11193 = n11188 ^ n11178 ;
  assign n11192 = n11172 ^ n11171 ;
  assign n11194 = n11193 ^ n11192 ;
  assign n11202 = n11201 ^ n11194 ;
  assign n11204 = n11203 ^ n11202 ;
  assign n11205 = n11204 ^ n11184 ;
  assign n11206 = n11205 ^ n11169 ;
  assign n11199 = n11198 ^ n11194 ;
  assign n11207 = n11206 ^ n11199 ;
  assign n11208 = n11207 ^ n11193 ;
  assign n11231 = n11230 ^ n11208 ;
  assign n11215 = n11214 ^ n11200 ;
  assign n11216 = n11215 ^ n11172 ;
  assign n11190 = n11189 ^ n11188 ;
  assign n11191 = n11190 ^ n11173 ;
  assign n11209 = n11208 ^ n11191 ;
  assign n11217 = n11216 ^ n11209 ;
  assign n11218 = ~n11104 & n11217 ;
  assign n11219 = n11218 ^ n11215 ;
  assign n11247 = n11231 ^ n11219 ;
  assign n11105 = n11104 ^ n11103 ;
  assign n11240 = n11207 ^ n11190 ;
  assign n11241 = n11240 ^ n11184 ;
  assign n11242 = n11184 ^ n11104 ;
  assign n11243 = n11242 ^ n11184 ;
  assign n11244 = n11241 & ~n11243 ;
  assign n11245 = n11244 ^ n11184 ;
  assign n11246 = n11105 & n11245 ;
  assign n11248 = n11247 ^ n11246 ;
  assign n11232 = n11231 ^ n11184 ;
  assign n11233 = n11232 ^ n11205 ;
  assign n11234 = n11233 ^ n11232 ;
  assign n11237 = n11104 & n11234 ;
  assign n11238 = n11237 ^ n11232 ;
  assign n11239 = n11103 & n11238 ;
  assign n11249 = n11248 ^ n11239 ;
  assign n11228 = n11199 & ~n11227 ;
  assign n11250 = n11249 ^ n11228 ;
  assign n11251 = n11250 ^ n9284 ;
  assign n11255 = n11254 ^ n11251 ;
  assign n11257 = n11256 ^ n11255 ;
  assign n11221 = n11203 ^ n11189 ;
  assign n11222 = n11221 ^ n11183 ;
  assign n11223 = n11104 & n11222 ;
  assign n11210 = n11209 ^ n11203 ;
  assign n11220 = n11219 ^ n11210 ;
  assign n11224 = n11223 ^ n11220 ;
  assign n11225 = ~n11105 & n11224 ;
  assign n11258 = n11257 ^ n11225 ;
  assign n13333 = n11258 ^ x65 ;
  assign n12548 = n12205 ^ n12202 ;
  assign n12549 = n12548 ^ n12214 ;
  assign n12550 = n12549 ^ n12227 ;
  assign n12545 = n12222 ^ n12205 ;
  assign n12546 = n12545 ^ n12207 ;
  assign n12542 = n12202 & n12220 ;
  assign n12547 = n12546 ^ n12542 ;
  assign n12551 = n12550 ^ n12547 ;
  assign n12552 = n12551 ^ n12200 ;
  assign n12543 = n12542 ^ n12208 ;
  assign n12544 = n12543 ^ n12225 ;
  assign n12553 = n12552 ^ n12544 ;
  assign n12561 = n12552 ^ n12550 ;
  assign n12562 = ~n12132 & n12561 ;
  assign n12563 = n12562 ^ n12550 ;
  assign n12556 = n12546 ^ n12223 ;
  assign n12555 = n12229 ^ n12204 ;
  assign n12557 = n12556 ^ n12555 ;
  assign n12554 = n12233 ^ n12211 ;
  assign n12558 = n12557 ^ n12554 ;
  assign n12559 = n12132 & n12558 ;
  assign n12560 = n12559 ^ n12557 ;
  assign n12564 = n12563 ^ n12560 ;
  assign n12565 = n12563 ^ n12131 ;
  assign n12566 = n12565 ^ n12563 ;
  assign n12567 = n12564 & ~n12566 ;
  assign n12568 = n12567 ^ n12563 ;
  assign n12569 = ~n12553 & n12568 ;
  assign n12570 = n12569 ^ n8974 ;
  assign n13373 = n12570 ^ x96 ;
  assign n13421 = n13333 & ~n13373 ;
  assign n13428 = n13421 ^ n13373 ;
  assign n13442 = n13428 ^ n13333 ;
  assign n13443 = n13422 & n13442 ;
  assign n13453 = n13443 ^ n13422 ;
  assign n13423 = n13422 ^ n13412 ;
  assign n13424 = n13423 ^ n13371 ;
  assign n13437 = ~n13424 & ~n13428 ;
  assign n13433 = n13421 & n13422 ;
  assign n13429 = n13422 ^ n13371 ;
  assign n13430 = ~n13428 & ~n13429 ;
  assign n13425 = n13421 & ~n13424 ;
  assign n13432 = n13430 ^ n13425 ;
  assign n13434 = n13433 ^ n13432 ;
  assign n13435 = n13434 ^ n13421 ;
  assign n13427 = n13421 & ~n13423 ;
  assign n13431 = n13430 ^ n13427 ;
  assign n13436 = n13435 ^ n13431 ;
  assign n13438 = n13437 ^ n13436 ;
  assign n13372 = n13371 ^ n13333 ;
  assign n13417 = n13373 ^ n13371 ;
  assign n13418 = ~n13372 & ~n13417 ;
  assign n13419 = n13418 ^ n13373 ;
  assign n13420 = n13412 & ~n13419 ;
  assign n13426 = n13425 ^ n13420 ;
  assign n13439 = n13438 ^ n13426 ;
  assign n13447 = n13443 ^ n13439 ;
  assign n13413 = n13412 ^ n13373 ;
  assign n13414 = ~n13372 & n13413 ;
  assign n13444 = n13443 ^ n13414 ;
  assign n13445 = n13444 ^ n13432 ;
  assign n13446 = n13445 ^ n13443 ;
  assign n13448 = n13447 ^ n13446 ;
  assign n13441 = n13430 ^ n13418 ;
  assign n13449 = n13448 ^ n13441 ;
  assign n13452 = n13449 ^ n13433 ;
  assign n13454 = n13453 ^ n13452 ;
  assign n10779 = n10778 ^ n10777 ;
  assign n10780 = n10543 & n10779 ;
  assign n10781 = n10780 ^ n10778 ;
  assign n10782 = n10542 & ~n10781 ;
  assign n10732 = n10543 ^ n10542 ;
  assign n10771 = n10741 ^ n10717 ;
  assign n10759 = n10740 ^ n10712 ;
  assign n10754 = n10721 ^ n10712 ;
  assign n10755 = n10721 ^ n10543 ;
  assign n10756 = n10732 & n10755 ;
  assign n10757 = n10756 ^ n10543 ;
  assign n10758 = n10754 & ~n10757 ;
  assign n10760 = n10759 ^ n10758 ;
  assign n10772 = n10771 ^ n10760 ;
  assign n10767 = n10744 ^ n10707 ;
  assign n10768 = n10767 ^ n10718 ;
  assign n10765 = n10724 ^ n10717 ;
  assign n10766 = n10765 ^ n10741 ;
  assign n10769 = n10768 ^ n10766 ;
  assign n10770 = ~n10543 & n10769 ;
  assign n10773 = n10772 ^ n10770 ;
  assign n10774 = n10732 & n10773 ;
  assign n10746 = n10745 ^ n10741 ;
  assign n10747 = n10741 ^ n10543 ;
  assign n10748 = n10747 ^ n10741 ;
  assign n10749 = ~n10746 & ~n10748 ;
  assign n10750 = n10749 ^ n10741 ;
  assign n10751 = ~n10732 & n10750 ;
  assign n10753 = n10752 ^ n10751 ;
  assign n10761 = n10760 ^ n10753 ;
  assign n10733 = n10706 ^ n10543 ;
  assign n10734 = n10733 ^ n10706 ;
  assign n10737 = n10725 & n10734 ;
  assign n10738 = n10737 ^ n10706 ;
  assign n10739 = n10732 & n10738 ;
  assign n10762 = n10761 ^ n10739 ;
  assign n10730 = n10729 ^ n10721 ;
  assign n10731 = ~n10545 & n10730 ;
  assign n10763 = n10762 ^ n10731 ;
  assign n10764 = n10763 ^ n9397 ;
  assign n10775 = n10774 ^ n10764 ;
  assign n10783 = n10782 ^ n10775 ;
  assign n13329 = n10783 ^ x98 ;
  assign n13668 = ~n13329 & n13437 ;
  assign n13512 = n13424 ^ n13420 ;
  assign n13513 = n13512 ^ n13436 ;
  assign n13653 = n13513 ^ n13432 ;
  assign n13487 = ~n13423 & ~n13428 ;
  assign n13488 = n13487 ^ n13436 ;
  assign n13654 = n13653 ^ n13488 ;
  assign n13655 = n13329 & ~n13654 ;
  assign n13475 = n13421 ^ n13333 ;
  assign n13476 = n13475 ^ n13454 ;
  assign n13477 = n13476 ^ n13448 ;
  assign n13478 = n13477 ^ n13449 ;
  assign n12423 = n12422 ^ n9073 ;
  assign n9893 = n9892 ^ n9882 ;
  assign n9894 = n9882 ^ n8958 ;
  assign n9895 = n9894 ^ n9882 ;
  assign n9896 = n9893 & ~n9895 ;
  assign n9897 = n9896 ^ n9882 ;
  assign n9898 = ~n8423 & ~n9897 ;
  assign n12424 = n12423 ^ n9898 ;
  assign n12411 = n9844 & n11675 ;
  assign n12407 = n9868 ^ n9856 ;
  assign n12408 = n12407 ^ n9877 ;
  assign n12409 = n8959 & n12408 ;
  assign n12394 = n9861 ^ n9857 ;
  assign n12395 = n12394 ^ n9848 ;
  assign n12396 = n12395 ^ n9864 ;
  assign n11660 = n9882 ^ n9862 ;
  assign n11661 = n11660 ^ n9868 ;
  assign n12397 = n12396 ^ n11661 ;
  assign n12398 = ~n8958 & ~n12397 ;
  assign n12399 = n12398 ^ n12395 ;
  assign n12410 = n12409 ^ n12399 ;
  assign n12412 = n12411 ^ n12410 ;
  assign n11664 = n11661 ^ n9870 ;
  assign n11665 = n11664 ^ n9857 ;
  assign n12400 = n12399 ^ n11665 ;
  assign n12401 = n12400 ^ n12399 ;
  assign n12402 = n12399 ^ n8958 ;
  assign n12403 = n12402 ^ n12399 ;
  assign n12404 = n12401 & n12403 ;
  assign n12405 = n12404 ^ n12399 ;
  assign n12406 = n8423 & n12405 ;
  assign n12413 = n12412 ^ n12406 ;
  assign n12421 = ~n12413 & ~n12420 ;
  assign n12425 = n12424 ^ n12421 ;
  assign n13330 = n12425 ^ x120 ;
  assign n13507 = n13449 ^ n13330 ;
  assign n13508 = n13507 ^ n13449 ;
  assign n13509 = n13478 & ~n13508 ;
  assign n13510 = n13509 ^ n13449 ;
  assign n13511 = n13329 & n13510 ;
  assign n13665 = n13655 ^ n13511 ;
  assign n13374 = n13373 ^ n13372 ;
  assign n13658 = n13420 ^ n13374 ;
  assign n13415 = n13414 ^ n13374 ;
  assign n13472 = n13412 ^ n13333 ;
  assign n13473 = ~n13415 & ~n13472 ;
  assign n13474 = n13473 ^ n13443 ;
  assign n13479 = n13478 ^ n13474 ;
  assign n13521 = n13479 ^ n13439 ;
  assign n13656 = n13521 ^ n13452 ;
  assign n13657 = n13656 ^ n13655 ;
  assign n13659 = n13658 ^ n13657 ;
  assign n13660 = n13657 ^ n13329 ;
  assign n13661 = n13660 ^ n13657 ;
  assign n13662 = n13659 & ~n13661 ;
  assign n13663 = n13662 ^ n13657 ;
  assign n13664 = ~n13330 & n13663 ;
  assign n13666 = n13665 ^ n13664 ;
  assign n13331 = ~n13329 & n13330 ;
  assign n13650 = n13446 ^ n13439 ;
  assign n13651 = n13650 ^ n13477 ;
  assign n13652 = n13331 & n13651 ;
  assign n13667 = n13666 ^ n13652 ;
  assign n13669 = n13668 ^ n13667 ;
  assign n13458 = n13330 ^ n13329 ;
  assign n13470 = n13430 ^ n13329 ;
  assign n13471 = n13470 ^ n13430 ;
  assign n13672 = n13431 & ~n13471 ;
  assign n13673 = n13672 ^ n13430 ;
  assign n13674 = n13458 & n13673 ;
  assign n13675 = ~n13669 & ~n13674 ;
  assign n13466 = n13331 ^ n13330 ;
  assign n13514 = n13466 ^ n13329 ;
  assign n13648 = n13427 & n13514 ;
  assign n13480 = n13479 ^ n13430 ;
  assign n13481 = n13471 & n13480 ;
  assign n13482 = n13481 ^ n13430 ;
  assign n13483 = n13330 & n13482 ;
  assign n13649 = n13648 ^ n13483 ;
  assign n13676 = n13675 ^ n13649 ;
  assign n13677 = ~n13454 & n13676 ;
  assign n13678 = n13677 ^ n10403 ;
  assign n13679 = n13678 ^ x107 ;
  assign n13680 = n13647 & n13679 ;
  assign n13681 = n13680 ^ n13679 ;
  assign n11881 = ~n11798 & n11880 ;
  assign n11882 = n11881 ^ n11879 ;
  assign n11903 = n11902 ^ n11882 ;
  assign n11904 = n11903 ^ n11882 ;
  assign n11905 = ~n11798 & ~n11904 ;
  assign n11906 = n11905 ^ n11882 ;
  assign n11907 = n11800 & n11906 ;
  assign n11908 = n11907 ^ n11882 ;
  assign n11956 = n11879 ^ n11870 ;
  assign n11934 = ~n11798 & ~n11901 ;
  assign n11935 = n11934 ^ n11900 ;
  assign n11957 = n11956 ^ n11935 ;
  assign n11952 = n11951 ^ n11873 ;
  assign n11953 = n11952 ^ n11869 ;
  assign n11954 = n11953 ^ n11879 ;
  assign n11955 = n11798 & n11954 ;
  assign n11958 = n11957 ^ n11955 ;
  assign n11959 = ~n11799 & ~n11958 ;
  assign n11946 = n11855 & ~n11945 ;
  assign n11947 = n11946 ^ n11943 ;
  assign n11909 = n11799 & ~n11898 ;
  assign n11910 = n11909 ^ n11897 ;
  assign n11936 = n11935 ^ n11910 ;
  assign n11948 = n11947 ^ n11936 ;
  assign n11928 = n11864 ^ n11862 ;
  assign n11929 = n11864 ^ n11798 ;
  assign n11930 = n11929 ^ n11864 ;
  assign n11931 = n11928 & n11930 ;
  assign n11932 = n11931 ^ n11864 ;
  assign n11933 = n11799 & n11932 ;
  assign n11949 = n11948 ^ n11933 ;
  assign n11950 = n11949 ^ n11927 ;
  assign n11960 = n11959 ^ n11950 ;
  assign n11914 = n11910 ^ n11900 ;
  assign n11911 = n11895 ^ n11872 ;
  assign n11912 = n11911 ^ n11897 ;
  assign n11913 = n11912 ^ n11910 ;
  assign n11915 = n11914 ^ n11913 ;
  assign n11916 = n11914 ^ n11799 ;
  assign n11917 = n11916 ^ n11914 ;
  assign n11918 = n11915 & n11917 ;
  assign n11919 = n11918 ^ n11914 ;
  assign n11920 = ~n11798 & n11919 ;
  assign n11961 = n11960 ^ n11920 ;
  assign n11962 = ~n11908 & ~n11961 ;
  assign n11963 = n11962 ^ n8579 ;
  assign n12925 = n11963 ^ x74 ;
  assign n11055 = n11054 ^ n10968 ;
  assign n11024 = n11013 ^ n10988 ;
  assign n11030 = n11024 ^ n11015 ;
  assign n11023 = n11022 ^ n10998 ;
  assign n11025 = n11024 ^ n11023 ;
  assign n11026 = n11024 ^ n10818 ;
  assign n11027 = n10853 & n11026 ;
  assign n11028 = n11027 ^ n10818 ;
  assign n11029 = n11025 & n11028 ;
  assign n11031 = n11030 ^ n11029 ;
  assign n11056 = n11055 ^ n11031 ;
  assign n11057 = n11056 ^ n11052 ;
  assign n11058 = n11057 ^ n11046 ;
  assign n11033 = n10989 ^ n10926 ;
  assign n11034 = n11033 ^ n11019 ;
  assign n11036 = n11035 ^ n11034 ;
  assign n11037 = ~n10818 & n11036 ;
  assign n11020 = n11019 ^ n10926 ;
  assign n11032 = n11031 ^ n11020 ;
  assign n11038 = n11037 ^ n11032 ;
  assign n11039 = n10986 & n11038 ;
  assign n11059 = n11058 ^ n11039 ;
  assign n10969 = n10968 ^ n10818 ;
  assign n10970 = n10969 ^ n10968 ;
  assign n10980 = n10970 & n10977 ;
  assign n10981 = n10980 ^ n10968 ;
  assign n10982 = ~n10852 & n10981 ;
  assign n11060 = n11059 ^ n10982 ;
  assign n11061 = n11060 ^ n10974 ;
  assign n11066 = n11065 ^ n11061 ;
  assign n11067 = n11066 ^ n11060 ;
  assign n11068 = ~n10852 & n11067 ;
  assign n11069 = n11068 ^ n11061 ;
  assign n11080 = n11069 ^ n8897 ;
  assign n11070 = n11069 ^ n11060 ;
  assign n11071 = n11070 ^ n11069 ;
  assign n11072 = n11019 ^ n11006 ;
  assign n11073 = ~n10818 & ~n11072 ;
  assign n11074 = n11073 ^ n11006 ;
  assign n11077 = ~n11071 & ~n11074 ;
  assign n11078 = n11077 ^ n11069 ;
  assign n11079 = n10853 & ~n11078 ;
  assign n11081 = n11080 ^ n11079 ;
  assign n12926 = n11081 ^ x113 ;
  assign n12927 = ~n12925 & ~n12926 ;
  assign n13007 = n12927 ^ n12925 ;
  assign n13008 = n13007 ^ n12926 ;
  assign n9904 = n8960 ^ n8958 ;
  assign n9905 = n9879 ^ n9864 ;
  assign n9906 = n9904 & ~n9905 ;
  assign n11683 = n9906 ^ n9887 ;
  assign n11657 = n9892 ^ n9870 ;
  assign n11659 = n11658 ^ n11657 ;
  assign n11662 = n11661 ^ n11659 ;
  assign n11663 = ~n8423 & ~n11662 ;
  assign n11666 = n11665 ^ n11663 ;
  assign n11684 = n11683 ^ n11666 ;
  assign n11685 = n11684 ^ n11682 ;
  assign n9900 = n9885 & ~n9899 ;
  assign n9901 = ~n9898 & n9900 ;
  assign n9902 = n9901 ^ n9898 ;
  assign n11686 = n11685 ^ n9902 ;
  assign n11687 = n11686 ^ n8648 ;
  assign n9910 = n8958 ^ n8423 ;
  assign n11667 = n11666 ^ n9872 ;
  assign n11668 = n11667 ^ n8958 ;
  assign n11669 = n11668 ^ n11667 ;
  assign n11670 = n11667 ^ n9873 ;
  assign n11671 = n11670 ^ n11667 ;
  assign n11672 = n11669 & n11671 ;
  assign n11673 = n11672 ^ n11667 ;
  assign n11674 = ~n9910 & n11673 ;
  assign n11688 = n11687 ^ n11674 ;
  assign n12936 = n11688 ^ x89 ;
  assign n12043 = n11180 ^ n11103 ;
  assign n12044 = n12043 ^ n11180 ;
  assign n12045 = n11197 & ~n12044 ;
  assign n12046 = n12045 ^ n11180 ;
  assign n12047 = ~n11104 & n12046 ;
  assign n12952 = n11226 ^ n11193 ;
  assign n12957 = n11212 ^ n11195 ;
  assign n12953 = n11212 ^ n11104 ;
  assign n12954 = ~n11105 & n12953 ;
  assign n12955 = n12954 ^ n11104 ;
  assign n12956 = ~n11109 & n12955 ;
  assign n12958 = n12957 ^ n12956 ;
  assign n12961 = ~n12952 & ~n12958 ;
  assign n12962 = n12961 ^ n11226 ;
  assign n12939 = n11209 ^ n11184 ;
  assign n12965 = n12939 ^ n11104 ;
  assign n12963 = n12939 ^ n11227 ;
  assign n12964 = n12963 ^ n12958 ;
  assign n12966 = n12965 ^ n12964 ;
  assign n12967 = n12962 & n12966 ;
  assign n12968 = n12967 ^ n12965 ;
  assign n12524 = n11203 ^ n11175 ;
  assign n12525 = n12524 ^ n11207 ;
  assign n12526 = n11207 ^ n11104 ;
  assign n12527 = n12526 ^ n11207 ;
  assign n12528 = n12525 & n12527 ;
  assign n12529 = n12528 ^ n11207 ;
  assign n12530 = n11103 & n12529 ;
  assign n12969 = n12968 ^ n12530 ;
  assign n12940 = n11183 ^ n11180 ;
  assign n12941 = n12940 ^ n11215 ;
  assign n12942 = ~n11104 & ~n12941 ;
  assign n12943 = n12942 ^ n11183 ;
  assign n12970 = n12969 ^ n12943 ;
  assign n12036 = n11214 ^ n11194 ;
  assign n12945 = n12943 ^ n12036 ;
  assign n12944 = n12943 ^ n12939 ;
  assign n12946 = n12945 ^ n12944 ;
  assign n12949 = ~n11104 & ~n12946 ;
  assign n12950 = n12949 ^ n12945 ;
  assign n12951 = n11103 & ~n12950 ;
  assign n12971 = n12970 ^ n12951 ;
  assign n12972 = ~n12047 & n12971 ;
  assign n12937 = n11228 ^ n8841 ;
  assign n12034 = n11252 ^ n11103 ;
  assign n12035 = n11190 & n12034 ;
  assign n12938 = n12937 ^ n12035 ;
  assign n12973 = n12972 ^ n12938 ;
  assign n12974 = n12973 ^ x106 ;
  assign n12975 = n12936 & n12974 ;
  assign n13009 = n12975 ^ n12936 ;
  assign n12931 = n12560 ^ n8681 ;
  assign n12928 = n12563 ^ n12553 ;
  assign n12929 = n12928 ^ n12560 ;
  assign n12930 = ~n12131 & ~n12929 ;
  assign n12932 = n12931 ^ n12930 ;
  assign n12933 = n12932 ^ x107 ;
  assign n11505 = n11501 ^ n11455 ;
  assign n11508 = n11505 ^ n11499 ;
  assign n11493 = n11467 ^ n11454 ;
  assign n11476 = n11469 ^ n11426 ;
  assign n11477 = n11476 ^ n11442 ;
  assign n11478 = n11477 ^ n11456 ;
  assign n11494 = n11493 ^ n11478 ;
  assign n11479 = n11466 ^ n11442 ;
  assign n11480 = ~n11478 & ~n11479 ;
  assign n11492 = n11294 & n11480 ;
  assign n11495 = n11494 ^ n11492 ;
  assign n11509 = n11508 ^ n11495 ;
  assign n11503 = n11502 ^ n11501 ;
  assign n11500 = n11499 ^ n11435 ;
  assign n11504 = n11503 ^ n11500 ;
  assign n11506 = n11505 ^ n11504 ;
  assign n11507 = ~n11294 & ~n11506 ;
  assign n11510 = n11509 ^ n11507 ;
  assign n11511 = n11466 & ~n11510 ;
  assign n11487 = n11298 & n11447 ;
  assign n11488 = n11487 ^ n11486 ;
  assign n11489 = n11488 ^ n11480 ;
  assign n11490 = n11489 ^ n11475 ;
  assign n11491 = n11490 ^ n8616 ;
  assign n11496 = n11495 ^ n11491 ;
  assign n11460 = n11446 ^ n11294 ;
  assign n11461 = n11460 ^ n11446 ;
  assign n11463 = n11447 & n11461 ;
  assign n11464 = n11463 ^ n11446 ;
  assign n11465 = n11295 & n11464 ;
  assign n11497 = n11496 ^ n11465 ;
  assign n11436 = n11435 ^ n11426 ;
  assign n11458 = n11457 ^ n11436 ;
  assign n11459 = ~n11299 & ~n11458 ;
  assign n11498 = n11497 ^ n11459 ;
  assign n11512 = n11511 ^ n11498 ;
  assign n12934 = n11512 ^ x80 ;
  assign n12935 = n12933 & n12934 ;
  assign n12981 = n12935 ^ n12934 ;
  assign n12984 = n12975 ^ n12974 ;
  assign n12985 = n12984 ^ n12936 ;
  assign n12988 = n12981 & ~n12985 ;
  assign n12976 = n12935 & n12975 ;
  assign n12995 = n12988 ^ n12976 ;
  assign n12982 = n12981 ^ n12933 ;
  assign n12986 = ~n12982 & ~n12985 ;
  assign n12983 = n12975 & ~n12982 ;
  assign n12987 = n12986 ^ n12983 ;
  assign n12989 = n12988 ^ n12987 ;
  assign n12978 = n12974 ^ n12936 ;
  assign n12979 = ~n12933 & n12978 ;
  assign n12980 = n12979 ^ n12933 ;
  assign n12990 = n12989 ^ n12980 ;
  assign n12996 = n12995 ^ n12990 ;
  assign n12994 = n12981 & n12984 ;
  assign n12997 = n12996 ^ n12994 ;
  assign n12993 = n12981 ^ n12976 ;
  assign n12998 = n12997 ^ n12993 ;
  assign n13020 = n13009 ^ n12998 ;
  assign n13015 = n12935 & n12984 ;
  assign n13016 = n13015 ^ n12935 ;
  assign n13003 = n12935 & ~n12985 ;
  assign n13004 = n13003 ^ n12976 ;
  assign n13017 = n13016 ^ n13004 ;
  assign n13011 = n12935 ^ n12933 ;
  assign n13012 = n12984 & n13011 ;
  assign n13013 = n13012 ^ n12983 ;
  assign n13010 = ~n12982 & n13009 ;
  assign n13014 = n13013 ^ n13010 ;
  assign n13018 = n13017 ^ n13014 ;
  assign n13019 = n13018 ^ n13013 ;
  assign n13021 = n13020 ^ n13019 ;
  assign n13022 = n13021 ^ n12986 ;
  assign n13023 = ~n13008 & ~n13022 ;
  assign n13002 = n12926 ^ n12925 ;
  assign n13029 = n12979 ^ n12936 ;
  assign n13030 = ~n12934 & ~n13029 ;
  assign n13031 = n13030 ^ n13014 ;
  assign n13032 = n13031 ^ n12987 ;
  assign n13689 = n13032 ^ n13015 ;
  assign n13687 = n13004 ^ n12983 ;
  assign n13690 = n13689 ^ n13687 ;
  assign n13691 = n12925 & n13690 ;
  assign n12999 = n12998 ^ n12994 ;
  assign n13686 = n13014 ^ n12999 ;
  assign n13688 = n13687 ^ n13686 ;
  assign n13692 = n13691 ^ n13688 ;
  assign n13693 = ~n13002 & ~n13692 ;
  assign n13694 = n13693 ^ n13014 ;
  assign n13039 = n13010 ^ n12982 ;
  assign n13040 = n13039 ^ n12987 ;
  assign n13685 = ~n12925 & ~n13040 ;
  assign n13695 = n13694 ^ n13685 ;
  assign n13000 = n12927 ^ n12926 ;
  assign n13683 = n13017 ^ n12994 ;
  assign n13684 = ~n13000 & n13683 ;
  assign n13696 = n13695 ^ n13684 ;
  assign n13682 = n12995 & n13002 ;
  assign n13697 = n13696 ^ n13682 ;
  assign n13033 = n13032 ^ n13011 ;
  assign n13025 = n13021 ^ n13012 ;
  assign n13034 = n13033 ^ n13025 ;
  assign n13698 = n13034 ^ n12925 ;
  assign n13699 = n13698 ^ n13034 ;
  assign n13052 = n13017 ^ n13003 ;
  assign n13700 = n12926 & n13052 ;
  assign n13701 = n13700 ^ n13034 ;
  assign n13702 = ~n13699 & ~n13701 ;
  assign n13703 = n13702 ^ n13034 ;
  assign n13704 = ~n13697 & ~n13703 ;
  assign n13705 = n13704 ^ n13697 ;
  assign n13706 = ~n13023 & ~n13705 ;
  assign n13709 = n13706 ^ n11846 ;
  assign n13026 = n13025 ^ n12990 ;
  assign n13027 = ~n12925 & n13026 ;
  assign n13028 = n13027 ^ n12990 ;
  assign n13707 = ~n13002 & n13706 ;
  assign n13708 = ~n13028 & n13707 ;
  assign n13710 = n13709 ^ n13708 ;
  assign n13711 = n13710 ^ x96 ;
  assign n12598 = n11933 ^ n11874 ;
  assign n12599 = n12598 ^ n11908 ;
  assign n12600 = n12599 ^ n11900 ;
  assign n12601 = n12600 ^ n12120 ;
  assign n12591 = n11888 ^ n11874 ;
  assign n12592 = n12591 ^ n11878 ;
  assign n12593 = n11878 ^ n11799 ;
  assign n12594 = n12593 ^ n11878 ;
  assign n12595 = n12592 & n12594 ;
  assign n12596 = n12595 ^ n11878 ;
  assign n12597 = n11800 & n12596 ;
  assign n12602 = n12601 ^ n12597 ;
  assign n12589 = n11895 ^ n11864 ;
  assign n12590 = ~n11945 & n12589 ;
  assign n12603 = n12602 ^ n12590 ;
  assign n12581 = n11900 ^ n11887 ;
  assign n12582 = n12581 ^ n11902 ;
  assign n12583 = n12582 ^ n11900 ;
  assign n12584 = n11900 ^ n11798 ;
  assign n12585 = n12584 ^ n11900 ;
  assign n12586 = ~n12583 & n12585 ;
  assign n12587 = n12586 ^ n11900 ;
  assign n12588 = n11799 & ~n12587 ;
  assign n12604 = n12603 ^ n12588 ;
  assign n12573 = n12120 ^ n11951 ;
  assign n12574 = n12573 ^ n11862 ;
  assign n12575 = n12574 ^ n12120 ;
  assign n12576 = n12120 ^ n11799 ;
  assign n12577 = n12576 ^ n12120 ;
  assign n12578 = n12575 & n12577 ;
  assign n12579 = n12578 ^ n12120 ;
  assign n12580 = n11800 & ~n12579 ;
  assign n12605 = n12604 ^ n12580 ;
  assign n12606 = ~n11947 & ~n12605 ;
  assign n12607 = n12606 ^ n9018 ;
  assign n12608 = n12607 ^ x94 ;
  assign n12571 = n12570 ^ x108 ;
  assign n12426 = n12425 ^ x69 ;
  assign n12430 = n10489 ^ n10443 ;
  assign n12440 = n12430 ^ n10423 ;
  assign n12441 = ~n10045 & n12440 ;
  assign n12442 = n12441 ^ n10423 ;
  assign n11729 = n10516 ^ n10413 ;
  assign n12431 = n11729 ^ n10450 ;
  assign n12432 = n10045 & n12431 ;
  assign n12433 = n12432 ^ n10450 ;
  assign n12449 = n12442 ^ n12433 ;
  assign n12450 = n12449 ^ n10523 ;
  assign n12451 = n12450 ^ n9157 ;
  assign n12435 = n12434 ^ n12433 ;
  assign n12436 = n12435 ^ n12430 ;
  assign n12437 = n12436 ^ n12433 ;
  assign n12438 = n10045 & n12437 ;
  assign n12439 = n12438 ^ n12435 ;
  assign n12452 = n12451 ^ n12439 ;
  assign n12447 = n10431 ^ n10408 ;
  assign n12448 = n10468 & n12447 ;
  assign n12453 = n12452 ^ n12448 ;
  assign n12443 = n12442 ^ n10445 ;
  assign n12444 = n12443 ^ n12439 ;
  assign n12427 = n10445 ^ n10438 ;
  assign n12428 = n12427 ^ n10455 ;
  assign n12429 = n10045 & n12428 ;
  assign n12445 = n12444 ^ n12429 ;
  assign n12446 = ~n9996 & ~n12445 ;
  assign n12454 = n12453 ^ n12446 ;
  assign n12455 = n12454 ^ x125 ;
  assign n12456 = n12426 & ~n12455 ;
  assign n12610 = n12456 ^ n12455 ;
  assign n12611 = n12610 ^ n12426 ;
  assign n12477 = n11467 ^ n11447 ;
  assign n12478 = n12477 ^ n11436 ;
  assign n12475 = n11468 ^ n11448 ;
  assign n12476 = n12475 ^ n11501 ;
  assign n12479 = n12478 ^ n12476 ;
  assign n12480 = ~n11294 & n12479 ;
  assign n12481 = n12480 ^ n12476 ;
  assign n12490 = n12489 ^ n12481 ;
  assign n11624 = n11505 ^ n11446 ;
  assign n12495 = n12490 ^ n11624 ;
  assign n12496 = n12495 ^ n12481 ;
  assign n12497 = n12496 ^ n11499 ;
  assign n12498 = ~n11294 & ~n12497 ;
  assign n12492 = n12491 ^ n12490 ;
  assign n12499 = n12498 ^ n12492 ;
  assign n12500 = ~n11295 & ~n12499 ;
  assign n12486 = n11294 & n11499 ;
  assign n12458 = n11450 ^ n11426 ;
  assign n12482 = n12481 ^ n12458 ;
  assign n12483 = n12482 ^ n12474 ;
  assign n12484 = n12483 ^ n9046 ;
  assign n12485 = n12484 ^ n11456 ;
  assign n12487 = n12486 ^ n12485 ;
  assign n12501 = n12500 ^ n12487 ;
  assign n12466 = n11445 ^ n11435 ;
  assign n12467 = n11298 & n12466 ;
  assign n12502 = n12501 ^ n12467 ;
  assign n12459 = n12458 ^ n11295 ;
  assign n12460 = n12459 ^ n12458 ;
  assign n12461 = n12458 ^ n11502 ;
  assign n12462 = n12461 ^ n12458 ;
  assign n12463 = n12460 & n12462 ;
  assign n12464 = n12463 ^ n12458 ;
  assign n12465 = n11466 & n12464 ;
  assign n12503 = n12502 ^ n12465 ;
  assign n11615 = n11469 ^ n11424 ;
  assign n12457 = ~n11299 & n11615 ;
  assign n12504 = n12503 ^ n12457 ;
  assign n12505 = n12504 ^ x76 ;
  assign n12531 = n12530 ^ n11219 ;
  assign n12048 = n11209 & n11226 ;
  assign n12049 = n12048 ^ n12047 ;
  assign n12037 = n11252 & ~n12036 ;
  assign n12038 = n12037 ^ n12035 ;
  assign n12523 = n12049 ^ n12038 ;
  assign n12532 = n12531 ^ n12523 ;
  assign n12533 = n12532 ^ n11228 ;
  assign n12534 = n12533 ^ n9120 ;
  assign n12516 = n11195 ^ n11182 ;
  assign n12517 = n12516 ^ n11201 ;
  assign n12518 = n11201 ^ n11104 ;
  assign n12519 = n12518 ^ n11201 ;
  assign n12520 = ~n12517 & n12519 ;
  assign n12521 = n12520 ^ n11201 ;
  assign n12522 = n11103 & ~n12521 ;
  assign n12535 = n12534 ^ n12522 ;
  assign n12514 = n11240 ^ n11199 ;
  assign n12515 = n11226 & n12514 ;
  assign n12536 = n12535 ^ n12515 ;
  assign n12506 = n11219 ^ n11181 ;
  assign n12507 = n12506 ^ n11103 ;
  assign n12508 = n12507 ^ n12506 ;
  assign n12509 = n12506 ^ n11187 ;
  assign n12510 = n12509 ^ n12506 ;
  assign n12511 = ~n12508 & n12510 ;
  assign n12512 = n12511 ^ n12506 ;
  assign n12513 = ~n11105 & n12512 ;
  assign n12537 = n12536 ^ n12513 ;
  assign n12538 = n12537 ^ x126 ;
  assign n12539 = ~n12505 & ~n12538 ;
  assign n12636 = n12539 ^ n12538 ;
  assign n12639 = n12611 & ~n12636 ;
  assign n12676 = n12639 ^ n12636 ;
  assign n12612 = n12611 ^ n12455 ;
  assign n12540 = n12539 ^ n12505 ;
  assign n12617 = n12540 ^ n12538 ;
  assign n12648 = n12612 & ~n12617 ;
  assign n12613 = ~n12540 & n12612 ;
  assign n12643 = n12613 ^ n12540 ;
  assign n12625 = ~n12540 & ~n12610 ;
  assign n12541 = n12456 & ~n12540 ;
  assign n12642 = n12625 ^ n12541 ;
  assign n12644 = n12643 ^ n12642 ;
  assign n12638 = n12456 & ~n12617 ;
  assign n12645 = n12644 ^ n12638 ;
  assign n12618 = n12611 & ~n12617 ;
  assign n12646 = n12645 ^ n12618 ;
  assign n12652 = n12648 ^ n12646 ;
  assign n12651 = n12644 ^ n12617 ;
  assign n12653 = n12652 ^ n12651 ;
  assign n12660 = n12653 ^ n12638 ;
  assign n12661 = n12660 ^ n12541 ;
  assign n12662 = n12661 ^ n12618 ;
  assign n12655 = ~n12610 & ~n12636 ;
  assign n12654 = n12653 ^ n12648 ;
  assign n12656 = n12655 ^ n12654 ;
  assign n12649 = n12648 ^ n12625 ;
  assign n12650 = n12649 ^ n12610 ;
  assign n12657 = n12656 ^ n12650 ;
  assign n12628 = n12539 & n12612 ;
  assign n12658 = n12657 ^ n12628 ;
  assign n12640 = n12639 ^ n12638 ;
  assign n12641 = n12640 ^ n12611 ;
  assign n12647 = n12646 ^ n12641 ;
  assign n12659 = n12658 ^ n12647 ;
  assign n12663 = n12662 ^ n12659 ;
  assign n12633 = n12538 ^ n12426 ;
  assign n12634 = ~n12505 & n12633 ;
  assign n12635 = n12634 ^ n12612 ;
  assign n12637 = n12636 ^ n12635 ;
  assign n12664 = n12663 ^ n12637 ;
  assign n12665 = n12664 ^ n12655 ;
  assign n12677 = n12676 ^ n12665 ;
  assign n12678 = n12677 ^ n12658 ;
  assign n13719 = n12678 ^ n12646 ;
  assign n13720 = n12571 & n13719 ;
  assign n13721 = n13720 ^ n12646 ;
  assign n13715 = n12652 ^ n12635 ;
  assign n13716 = ~n12571 & ~n13715 ;
  assign n13717 = n13716 ^ n12652 ;
  assign n13718 = n13717 ^ n12639 ;
  assign n13722 = n13721 ^ n13718 ;
  assign n13723 = n13722 ^ n12625 ;
  assign n13724 = n13723 ^ n12639 ;
  assign n13725 = n13724 ^ n13722 ;
  assign n13728 = ~n12571 & n13725 ;
  assign n13729 = n13728 ^ n13722 ;
  assign n13730 = n12608 & n13729 ;
  assign n13731 = n13730 ^ n13717 ;
  assign n12670 = n12608 ^ n12571 ;
  assign n12697 = n12655 ^ n12608 ;
  assign n12698 = n12697 ^ n12655 ;
  assign n12701 = ~n12656 & n12698 ;
  assign n12702 = n12701 ^ n12655 ;
  assign n12703 = ~n12670 & n12702 ;
  assign n13742 = n13731 ^ n12703 ;
  assign n13739 = ~n12678 & n12698 ;
  assign n13740 = n13739 ^ n12655 ;
  assign n13741 = n12670 & n13740 ;
  assign n13743 = n13742 ^ n13741 ;
  assign n12688 = n12659 ^ n12539 ;
  assign n12689 = n12688 ^ n12647 ;
  assign n12690 = n12689 ^ n12677 ;
  assign n13713 = n12690 ^ n12608 ;
  assign n13714 = n13713 ^ n12690 ;
  assign n13732 = n12642 & n13731 ;
  assign n13733 = n13732 ^ n12690 ;
  assign n13734 = n13714 & ~n13733 ;
  assign n13735 = n13734 ^ n12690 ;
  assign n13736 = n12571 & ~n13735 ;
  assign n13744 = n13743 ^ n13736 ;
  assign n12629 = ~n12571 & n12608 ;
  assign n12630 = n12629 ^ n12608 ;
  assign n12631 = n12630 ^ n12571 ;
  assign n12667 = n12631 ^ n12608 ;
  assign n13712 = n12639 & ~n12667 ;
  assign n13745 = n13744 ^ n13712 ;
  assign n13746 = n13745 ^ n11293 ;
  assign n13747 = n13746 ^ x122 ;
  assign n13748 = n13711 & ~n13747 ;
  assign n12296 = n12295 ^ x85 ;
  assign n10457 = n10045 & ~n10456 ;
  assign n10458 = n10457 ^ n10408 ;
  assign n10460 = n10458 ^ n10446 ;
  assign n10459 = n10458 ^ n10431 ;
  assign n10461 = n10460 ^ n10459 ;
  assign n10464 = ~n10045 & n10461 ;
  assign n10465 = n10464 ^ n10460 ;
  assign n10466 = ~n9996 & n10465 ;
  assign n10467 = n10466 ^ n10458 ;
  assign n11738 = ~n10045 & ~n10421 ;
  assign n11730 = n10477 ^ n10431 ;
  assign n11731 = n11730 ^ n10233 ;
  assign n11732 = n11731 ^ n10431 ;
  assign n11733 = n10431 ^ n10045 ;
  assign n11734 = n11733 ^ n10431 ;
  assign n11735 = n11732 & n11734 ;
  assign n11736 = n11735 ^ n10431 ;
  assign n11737 = n11729 & ~n11736 ;
  assign n11739 = n11738 ^ n11737 ;
  assign n11740 = n10468 & ~n11739 ;
  assign n11741 = n11740 ^ n11738 ;
  assign n11726 = n10448 ^ n10438 ;
  assign n11727 = n11726 ^ n10424 ;
  assign n11728 = n11725 & ~n11727 ;
  assign n11742 = n11741 ^ n11728 ;
  assign n11743 = n10468 ^ n10442 ;
  assign n11746 = n10516 ^ n10479 ;
  assign n11745 = n10446 ^ n10421 ;
  assign n11747 = n11746 ^ n11745 ;
  assign n11750 = n11747 ^ n10442 ;
  assign n11744 = n10489 ^ n10455 ;
  assign n11748 = n11747 ^ n11744 ;
  assign n11749 = ~n9996 & ~n11748 ;
  assign n11751 = n11750 ^ n11749 ;
  assign n11752 = ~n11743 & n11751 ;
  assign n11753 = n11752 ^ n10468 ;
  assign n11754 = ~n11742 & n11753 ;
  assign n11755 = ~n10467 & n11754 ;
  assign n11756 = n11755 ^ n9558 ;
  assign n12297 = n11756 ^ x67 ;
  assign n12298 = n12296 & ~n12297 ;
  assign n12247 = n12246 ^ x86 ;
  assign n12052 = n12036 ^ n11195 ;
  assign n12050 = n11209 ^ n11193 ;
  assign n12051 = n12050 ^ n11198 ;
  assign n12053 = n12052 ^ n12051 ;
  assign n12054 = n11104 & n12053 ;
  assign n12055 = n12054 ^ n12050 ;
  assign n12060 = n12055 ^ n11207 ;
  assign n12061 = n12060 ^ n11180 ;
  assign n12062 = n12061 ^ n12055 ;
  assign n12065 = n11104 & n12062 ;
  assign n12066 = n12065 ^ n12055 ;
  assign n12067 = n11105 & n12066 ;
  assign n12056 = n12055 ^ n12049 ;
  assign n12057 = n12056 ^ n11246 ;
  assign n12068 = n12067 ^ n12057 ;
  assign n12069 = n11203 ^ n11201 ;
  assign n12070 = n12069 ^ n11175 ;
  assign n12071 = n12070 ^ n11203 ;
  assign n12072 = n11203 ^ n11103 ;
  assign n12073 = n12072 ^ n11203 ;
  assign n12074 = ~n12071 & ~n12073 ;
  assign n12075 = n12074 ^ n11203 ;
  assign n12076 = ~n11104 & n12075 ;
  assign n12077 = ~n12068 & ~n12076 ;
  assign n12080 = n12052 ^ n11172 ;
  assign n12081 = n11226 & ~n12080 ;
  assign n12082 = n12077 & n12081 ;
  assign n12039 = n12038 ^ n9705 ;
  assign n12029 = n11182 ^ n11104 ;
  assign n12030 = n12029 ^ n11182 ;
  assign n12031 = n11207 & n12030 ;
  assign n12032 = n12031 ^ n11182 ;
  assign n12033 = n11103 & n12032 ;
  assign n12040 = n12039 ^ n12033 ;
  assign n12078 = n12077 ^ n12040 ;
  assign n12083 = n12082 ^ n12078 ;
  assign n12084 = n12083 ^ x68 ;
  assign n12128 = n11799 & ~n11935 ;
  assign n12121 = n12120 ^ n11912 ;
  assign n12122 = n12120 ^ n11798 ;
  assign n12123 = n12122 ^ n12120 ;
  assign n12124 = n12121 & n12123 ;
  assign n12125 = n12124 ^ n12120 ;
  assign n12126 = ~n11800 & ~n12125 ;
  assign n12112 = n12085 ^ n11860 ;
  assign n12113 = n12085 ^ n11855 ;
  assign n12114 = n12113 ^ n12085 ;
  assign n12115 = n12112 & ~n12114 ;
  assign n12116 = n12115 ^ n12085 ;
  assign n12117 = n12086 ^ n11855 ;
  assign n12118 = ~n12116 & ~n12117 ;
  assign n12092 = n11900 ^ n11891 ;
  assign n12093 = ~n11945 & ~n12092 ;
  assign n12090 = n11951 ^ n11869 ;
  assign n12091 = ~n11799 & n12090 ;
  assign n12094 = n12093 ^ n12091 ;
  assign n12089 = n12088 ^ n12086 ;
  assign n12095 = n12094 ^ n12089 ;
  assign n12108 = n12107 ^ n12095 ;
  assign n12109 = n12108 ^ n11927 ;
  assign n12110 = n12109 ^ n11908 ;
  assign n12111 = n12110 ^ n9753 ;
  assign n12119 = n12118 ^ n12111 ;
  assign n12127 = n12126 ^ n12119 ;
  assign n12129 = n12128 ^ n12127 ;
  assign n12130 = n12129 ^ x116 ;
  assign n12314 = n12084 & n12130 ;
  assign n12317 = n12314 ^ n12084 ;
  assign n12318 = n12247 & n12317 ;
  assign n12303 = ~n12084 & n12247 ;
  assign n12316 = n12303 ^ n12247 ;
  assign n12319 = n12318 ^ n12316 ;
  assign n12323 = n12319 ^ n12314 ;
  assign n11616 = n11615 ^ n11456 ;
  assign n11617 = n11616 ^ n11294 ;
  assign n11620 = n11619 ^ n11493 ;
  assign n11621 = n11620 ^ n11448 ;
  assign n11622 = n11505 ^ n11448 ;
  assign n11623 = n11622 ^ n11294 ;
  assign n11625 = n11624 ^ n11295 ;
  assign n11628 = ~n11622 & ~n11625 ;
  assign n11629 = n11628 ^ n11295 ;
  assign n11630 = n11623 & n11629 ;
  assign n11631 = n11630 ^ n11294 ;
  assign n11632 = ~n11621 & ~n11631 ;
  assign n11635 = ~n11617 & ~n11632 ;
  assign n11636 = n11635 ^ n11294 ;
  assign n11607 = n11477 ^ n11440 ;
  assign n11608 = n11607 ^ n11503 ;
  assign n11609 = n11608 ^ n11477 ;
  assign n11610 = n11477 ^ n11294 ;
  assign n11611 = n11610 ^ n11477 ;
  assign n11612 = n11609 & n11611 ;
  assign n11613 = n11612 ^ n11477 ;
  assign n11614 = ~n11295 & n11613 ;
  assign n11638 = n11614 ^ n11295 ;
  assign n11637 = n11632 ^ n11614 ;
  assign n11639 = n11638 ^ n11637 ;
  assign n11640 = ~n11636 & n11639 ;
  assign n11641 = n11640 ^ n11638 ;
  assign n11642 = n11641 ^ n11614 ;
  assign n11645 = n11641 ^ n11466 ;
  assign n11646 = n11645 ^ n11641 ;
  assign n11647 = n11641 ^ n11499 ;
  assign n11648 = n11647 ^ n11641 ;
  assign n11649 = ~n11646 & n11648 ;
  assign n11650 = ~n11642 & n11649 ;
  assign n11651 = n11650 ^ n11642 ;
  assign n11652 = n11651 ^ n11614 ;
  assign n11653 = ~n11606 & ~n11652 ;
  assign n11654 = ~n11488 & n11653 ;
  assign n11655 = n11654 ^ n9522 ;
  assign n12248 = n11655 ^ x109 ;
  assign n12249 = n12247 & ~n12248 ;
  assign n12250 = n12249 ^ n12248 ;
  assign n12251 = n12250 ^ n12247 ;
  assign n12252 = n12130 & n12251 ;
  assign n12253 = ~n12084 & n12252 ;
  assign n12254 = n12253 ^ n12252 ;
  assign n12324 = n12323 ^ n12254 ;
  assign n12308 = ~n12084 & ~n12250 ;
  assign n12322 = n12308 ^ n12250 ;
  assign n12325 = n12324 ^ n12322 ;
  assign n13752 = n12298 & ~n12325 ;
  assign n12299 = n12298 ^ n12297 ;
  assign n12309 = n12130 & n12308 ;
  assign n12310 = n12309 ^ n12308 ;
  assign n12311 = ~n12299 & n12310 ;
  assign n13753 = n13752 ^ n12311 ;
  assign n12300 = n12299 ^ n12296 ;
  assign n12363 = n12324 ^ n12309 ;
  assign n12315 = n12249 & n12314 ;
  assign n13779 = n12363 ^ n12315 ;
  assign n12342 = n12252 ^ n12251 ;
  assign n12321 = n12318 ^ n12317 ;
  assign n12326 = n12325 ^ n12321 ;
  assign n12343 = n12342 ^ n12326 ;
  assign n12304 = n12248 & n12303 ;
  assign n12338 = ~n12130 & n12304 ;
  assign n12344 = n12343 ^ n12338 ;
  assign n12320 = n12319 ^ n12315 ;
  assign n12327 = n12326 ^ n12320 ;
  assign n12345 = n12344 ^ n12327 ;
  assign n12339 = n12338 ^ n12304 ;
  assign n12340 = n12339 ^ n12252 ;
  assign n12341 = n12340 ^ n12248 ;
  assign n12346 = n12345 ^ n12341 ;
  assign n12357 = n12346 ^ n12318 ;
  assign n13776 = n12357 ^ n12324 ;
  assign n13777 = n13776 ^ n12130 ;
  assign n12347 = n12346 ^ n12339 ;
  assign n12348 = n12347 ^ n12343 ;
  assign n12349 = n12348 ^ n12253 ;
  assign n12305 = n12304 ^ n12303 ;
  assign n12306 = n12130 & n12305 ;
  assign n12334 = n12306 ^ n12305 ;
  assign n12335 = n12334 ^ n12325 ;
  assign n12336 = n12335 ^ n12324 ;
  assign n12337 = n12336 ^ n12310 ;
  assign n12350 = n12349 ^ n12337 ;
  assign n13778 = n13777 ^ n12350 ;
  assign n13780 = n13779 ^ n13778 ;
  assign n13781 = n12300 & ~n13780 ;
  assign n13758 = n12299 ^ n12252 ;
  assign n13759 = n13758 ^ n12346 ;
  assign n13760 = n12324 ^ n12299 ;
  assign n12383 = n12325 ^ n12315 ;
  assign n12384 = n12383 ^ n12306 ;
  assign n13761 = n13760 ^ n12384 ;
  assign n13762 = ~n13759 & n13761 ;
  assign n13763 = n13762 ^ n12299 ;
  assign n13765 = n12343 ^ n12320 ;
  assign n13766 = n13765 ^ n12339 ;
  assign n12358 = n12357 ^ n12309 ;
  assign n12359 = n12358 ^ n12254 ;
  assign n12360 = n12359 ^ n12310 ;
  assign n13767 = n13766 ^ n12360 ;
  assign n13764 = n12336 ^ n12320 ;
  assign n13768 = n13767 ^ n13764 ;
  assign n13769 = n13764 ^ n12297 ;
  assign n13770 = n13769 ^ n13764 ;
  assign n13771 = n13768 & ~n13770 ;
  assign n13772 = n13771 ^ n13764 ;
  assign n13773 = n12296 & ~n13772 ;
  assign n13774 = n13763 & ~n13773 ;
  assign n12301 = n12300 ^ n12297 ;
  assign n13754 = n12346 ^ n12338 ;
  assign n13755 = n13754 ^ n12253 ;
  assign n13756 = n12301 & n13755 ;
  assign n12374 = n12343 ^ n12334 ;
  assign n12375 = n12343 ^ n12296 ;
  assign n12376 = n12375 ^ n12343 ;
  assign n12377 = ~n12374 & ~n12376 ;
  assign n12378 = n12377 ^ n12343 ;
  assign n12379 = n12297 & ~n12378 ;
  assign n13757 = n13756 ^ n12379 ;
  assign n13775 = n13774 ^ n13757 ;
  assign n13782 = n13781 ^ n13775 ;
  assign n13783 = ~n13753 & n13782 ;
  assign n13784 = n13783 ^ n10044 ;
  assign n13785 = n13784 ^ x113 ;
  assign n13175 = n12537 ^ x101 ;
  assign n13176 = n12783 ^ x110 ;
  assign n13177 = n13175 & n13176 ;
  assign n13178 = n13177 ^ n13176 ;
  assign n13179 = n13178 ^ n13175 ;
  assign n13200 = n12291 ^ n10741 ;
  assign n13201 = n13200 ^ n10720 ;
  assign n13202 = ~n10543 & n13201 ;
  assign n13187 = n10744 ^ n10726 ;
  assign n13203 = n13202 ^ n13187 ;
  assign n13204 = n10732 & n13203 ;
  assign n11709 = n10745 ^ n10716 ;
  assign n13196 = n11709 ^ n10781 ;
  assign n13192 = n10724 ^ n10710 ;
  assign n13193 = n13192 ^ n10729 ;
  assign n13194 = n13193 ^ n11709 ;
  assign n13195 = ~n10543 & ~n13194 ;
  assign n13197 = n13196 ^ n13195 ;
  assign n13198 = ~n10542 & n13197 ;
  assign n11691 = n11690 ^ n10778 ;
  assign n11692 = n11691 ^ n10777 ;
  assign n11693 = n10777 ^ n10543 ;
  assign n11694 = n11693 ^ n10777 ;
  assign n11695 = n11692 & n11694 ;
  assign n11696 = n11695 ^ n10777 ;
  assign n11697 = n10542 & ~n11696 ;
  assign n13188 = n13187 ^ n11697 ;
  assign n13189 = n13188 ^ n10781 ;
  assign n13190 = n13189 ^ n10731 ;
  assign n13191 = n13190 ^ n10149 ;
  assign n13199 = n13198 ^ n13191 ;
  assign n13205 = n13204 ^ n13199 ;
  assign n13206 = n13205 ^ x77 ;
  assign n13207 = n12607 ^ x92 ;
  assign n13208 = ~n13206 & n13207 ;
  assign n13180 = n12749 ^ x70 ;
  assign n13181 = n12242 ^ n12131 ;
  assign n13182 = n13181 ^ n12244 ;
  assign n13183 = n13182 ^ n10117 ;
  assign n13184 = n13183 ^ x83 ;
  assign n13185 = n13180 & ~n13184 ;
  assign n13186 = n13185 ^ n13180 ;
  assign n13216 = n13186 ^ n13184 ;
  assign n13245 = n13208 & n13216 ;
  assign n13237 = n13207 ^ n13206 ;
  assign n13240 = n13237 ^ n13180 ;
  assign n13213 = n13207 ^ n13180 ;
  assign n13214 = n13184 & n13213 ;
  assign n13215 = n13214 ^ n13207 ;
  assign n13232 = n13206 ^ n13184 ;
  assign n13239 = n13215 & ~n13232 ;
  assign n13241 = n13240 ^ n13239 ;
  assign n13233 = ~n13180 & ~n13232 ;
  assign n13238 = n13237 ^ n13233 ;
  assign n13242 = n13241 ^ n13238 ;
  assign n13235 = n13232 ^ n13180 ;
  assign n13211 = n13208 ^ n13206 ;
  assign n13222 = n13185 & ~n13211 ;
  assign n13236 = n13235 ^ n13222 ;
  assign n13243 = n13242 ^ n13236 ;
  assign n13226 = n13185 ^ n13184 ;
  assign n13209 = n13208 ^ n13207 ;
  assign n13227 = n13209 ^ n13206 ;
  assign n13228 = ~n13226 & n13227 ;
  assign n13244 = n13243 ^ n13228 ;
  assign n13246 = n13245 ^ n13244 ;
  assign n13247 = n13246 ^ n13216 ;
  assign n13230 = ~n13211 & ~n13226 ;
  assign n13231 = n13230 ^ n13228 ;
  assign n13234 = n13233 ^ n13231 ;
  assign n13248 = n13247 ^ n13234 ;
  assign n13249 = n13248 ^ n13244 ;
  assign n13217 = n13209 & n13216 ;
  assign n13250 = n13249 ^ n13217 ;
  assign n13251 = n13250 ^ n13247 ;
  assign n13252 = n13251 ^ n13245 ;
  assign n13221 = n13185 & n13209 ;
  assign n13223 = n13222 ^ n13221 ;
  assign n13219 = n13185 & n13208 ;
  assign n13220 = n13219 ^ n13185 ;
  assign n13224 = n13223 ^ n13220 ;
  assign n13210 = n13186 & n13209 ;
  assign n13225 = n13224 ^ n13210 ;
  assign n13229 = n13228 ^ n13225 ;
  assign n13253 = n13252 ^ n13229 ;
  assign n13218 = n13217 ^ n13215 ;
  assign n13254 = n13253 ^ n13218 ;
  assign n13212 = n13211 ^ n13210 ;
  assign n13255 = n13254 ^ n13212 ;
  assign n13256 = ~n13179 & ~n13255 ;
  assign n13278 = n13210 ^ n13186 ;
  assign n13275 = n13241 ^ n13180 ;
  assign n13276 = n13275 ^ n13253 ;
  assign n13277 = n13276 ^ n13255 ;
  assign n13279 = n13278 ^ n13277 ;
  assign n13792 = n13279 ^ n13221 ;
  assign n13793 = n13792 ^ n13222 ;
  assign n13811 = n13793 ^ n13276 ;
  assign n13812 = n13178 & ~n13811 ;
  assign n13806 = n13244 ^ n13225 ;
  assign n13807 = n13806 ^ n13277 ;
  assign n13808 = n13177 & ~n13807 ;
  assign n13805 = n13176 & ~n13251 ;
  assign n13809 = n13808 ^ n13805 ;
  assign n13798 = n13248 ^ n13243 ;
  assign n13799 = n13798 ^ n13253 ;
  assign n13800 = n13253 ^ n13176 ;
  assign n13801 = n13800 ^ n13253 ;
  assign n13802 = ~n13799 & n13801 ;
  assign n13803 = n13802 ^ n13253 ;
  assign n13804 = ~n13175 & ~n13803 ;
  assign n13810 = n13809 ^ n13804 ;
  assign n13813 = n13812 ^ n13810 ;
  assign n13791 = n13177 ^ n13175 ;
  assign n13260 = n13245 ^ n13230 ;
  assign n13288 = n13260 ^ n13180 ;
  assign n13289 = n13288 ^ n13247 ;
  assign n13795 = n13289 ^ n13248 ;
  assign n13794 = n13793 ^ n13260 ;
  assign n13796 = n13795 ^ n13794 ;
  assign n13797 = n13791 & ~n13796 ;
  assign n13814 = n13813 ^ n13797 ;
  assign n13786 = n13219 ^ n13217 ;
  assign n13789 = n13176 & n13786 ;
  assign n13790 = n13789 ^ n13217 ;
  assign n13815 = n13814 ^ n13790 ;
  assign n13788 = ~n13179 & ~n13276 ;
  assign n13816 = n13815 ^ n13788 ;
  assign n13787 = ~n13175 & n13786 ;
  assign n13817 = n13816 ^ n13787 ;
  assign n13818 = ~n13256 & ~n13817 ;
  assign n13819 = n13818 ^ n11822 ;
  assign n13820 = n13819 ^ x74 ;
  assign n13821 = ~n13785 & ~n13820 ;
  assign n13822 = n13821 ^ n13820 ;
  assign n13847 = n13748 & ~n13822 ;
  assign n13830 = n13821 ^ n13785 ;
  assign n13832 = n13830 ^ n13820 ;
  assign n13846 = n13748 & ~n13832 ;
  assign n13848 = n13847 ^ n13846 ;
  assign n15121 = n13848 ^ n13822 ;
  assign n13749 = n13748 ^ n13711 ;
  assign n13750 = n13749 ^ n13747 ;
  assign n13833 = n13750 & ~n13832 ;
  assign n13831 = n13750 & ~n13830 ;
  assign n13834 = n13833 ^ n13831 ;
  assign n13828 = n13750 & ~n13822 ;
  assign n13829 = n13828 ^ n13750 ;
  assign n13835 = n13834 ^ n13829 ;
  assign n13751 = n13750 ^ n13711 ;
  assign n13823 = ~n13751 & ~n13822 ;
  assign n13918 = n13835 ^ n13823 ;
  assign n15122 = n15121 ^ n13918 ;
  assign n15123 = n13681 & ~n15122 ;
  assign n13827 = n13749 & n13821 ;
  assign n13836 = n13835 ^ n13827 ;
  assign n14805 = n13836 ^ n13821 ;
  assign n14806 = n13681 & n14805 ;
  assign n15124 = n15123 ^ n14806 ;
  assign n13838 = ~n13751 & ~n13830 ;
  assign n13868 = n13847 ^ n13838 ;
  assign n13869 = n13868 ^ n13823 ;
  assign n15111 = n13680 & n13869 ;
  assign n13842 = n13679 ^ n13647 ;
  assign n13825 = n13748 & n13821 ;
  assign n13826 = n13825 ^ n13821 ;
  assign n13837 = n13836 ^ n13826 ;
  assign n14807 = n13846 ^ n13837 ;
  assign n15104 = n14807 ^ n13847 ;
  assign n15105 = n13847 ^ n13679 ;
  assign n15106 = n15105 ^ n13847 ;
  assign n15107 = n15104 & ~n15106 ;
  assign n15108 = n15107 ^ n13847 ;
  assign n15109 = ~n13842 & n15108 ;
  assign n13885 = n13825 ^ n13748 ;
  assign n13886 = n13885 ^ n13848 ;
  assign n15102 = n13886 ^ n13827 ;
  assign n15101 = n13847 ^ n13833 ;
  assign n15103 = n15102 ^ n15101 ;
  assign n15110 = n15109 ^ n15103 ;
  assign n15112 = n15111 ^ n15110 ;
  assign n15125 = n15124 ^ n15112 ;
  assign n13861 = n13681 ^ n13647 ;
  assign n13862 = n13861 ^ n13679 ;
  assign n13870 = n13838 ^ n13828 ;
  assign n13871 = n13870 ^ n13822 ;
  assign n13872 = n13871 ^ n13869 ;
  assign n14803 = n13862 & ~n13872 ;
  assign n13839 = n13838 ^ n13837 ;
  assign n13824 = n13823 ^ n13751 ;
  assign n13840 = n13839 ^ n13824 ;
  assign n13884 = ~n13840 & ~n13861 ;
  assign n14804 = n14803 ^ n13884 ;
  assign n15126 = n15125 ^ n14804 ;
  assign n13919 = n13647 & n13918 ;
  assign n13920 = n13919 ^ n13835 ;
  assign n13865 = n13846 ^ n13827 ;
  assign n13866 = n13865 ^ n13847 ;
  assign n13863 = n13785 ^ n13747 ;
  assign n13864 = n13711 & n13863 ;
  assign n13867 = n13866 ^ n13864 ;
  assign n13917 = n13867 ^ n13828 ;
  assign n13921 = n13920 ^ n13917 ;
  assign n13922 = n13921 ^ n13920 ;
  assign n13923 = n13920 ^ n13647 ;
  assign n13924 = n13923 ^ n13920 ;
  assign n13925 = n13922 & n13924 ;
  assign n13926 = n13925 ^ n13920 ;
  assign n13927 = n13679 & n13926 ;
  assign n13928 = n13927 ^ n13920 ;
  assign n13916 = n13825 & n13862 ;
  assign n13929 = n13928 ^ n13916 ;
  assign n15127 = n15126 ^ n13929 ;
  assign n13873 = n13872 ^ n13867 ;
  assign n13887 = n13873 ^ n13827 ;
  assign n13888 = n13887 ^ n13749 ;
  assign n14817 = n13888 ^ n13838 ;
  assign n14818 = n13862 & ~n14817 ;
  assign n13895 = n13681 & n13831 ;
  assign n14819 = n14818 ^ n13895 ;
  assign n15128 = n15127 ^ n14819 ;
  assign n13841 = n13681 & ~n13840 ;
  assign n15129 = n15128 ^ n13841 ;
  assign n15130 = n15129 ^ n12607 ;
  assign n15113 = n15112 ^ n13917 ;
  assign n15114 = n15113 ^ n13831 ;
  assign n15115 = n15114 ^ n15112 ;
  assign n15118 = n13647 & n15115 ;
  assign n15119 = n15118 ^ n15112 ;
  assign n15120 = n13842 & n15119 ;
  assign n15131 = n15130 ^ n15120 ;
  assign n15132 = n15131 ^ x125 ;
  assign n12683 = n12631 & ~n12654 ;
  assign n12682 = ~n12571 & n12618 ;
  assign n12684 = n12683 ^ n12682 ;
  assign n12632 = ~n12628 & ~n12631 ;
  assign n14735 = n12688 ^ n12664 ;
  assign n14736 = n14735 ^ n12667 ;
  assign n14737 = n14736 ^ n12657 ;
  assign n14738 = ~n12632 & n14737 ;
  assign n14739 = n14738 ^ n12677 ;
  assign n13986 = n12655 ^ n12613 ;
  assign n13987 = n12613 ^ n12608 ;
  assign n13988 = n13987 ^ n12613 ;
  assign n13989 = n13986 & n13988 ;
  assign n13990 = n13989 ^ n12613 ;
  assign n13991 = n12571 & n13990 ;
  assign n14747 = n14739 ^ n13991 ;
  assign n14740 = n14739 ^ n12663 ;
  assign n14741 = n14740 ^ n12647 ;
  assign n12668 = n12664 ^ n12658 ;
  assign n14742 = n14741 ^ n12668 ;
  assign n14743 = n14742 ^ n14739 ;
  assign n14744 = ~n12571 & ~n14743 ;
  assign n14745 = n14744 ^ n14740 ;
  assign n14746 = n12608 & ~n14745 ;
  assign n14748 = n14747 ^ n14746 ;
  assign n14727 = n12649 ^ n12541 ;
  assign n14728 = n14727 ^ n12655 ;
  assign n14729 = n14728 ^ n12541 ;
  assign n14732 = ~n12608 & n14729 ;
  assign n14733 = n14732 ^ n12541 ;
  assign n14734 = ~n12571 & n14733 ;
  assign n14749 = n14748 ^ n14734 ;
  assign n14721 = n12660 ^ n12644 ;
  assign n14722 = n12644 ^ n12608 ;
  assign n14723 = n14722 ^ n12644 ;
  assign n14724 = n14721 & n14723 ;
  assign n14725 = n14724 ^ n12644 ;
  assign n14726 = n12670 & ~n14725 ;
  assign n14750 = n14749 ^ n14726 ;
  assign n14751 = ~n12684 & n14750 ;
  assign n14752 = ~n13712 & n14751 ;
  assign n14753 = n14752 ^ n12167 ;
  assign n14754 = n14753 ^ x121 ;
  assign n13965 = n12997 ^ n12934 ;
  assign n13966 = ~n13007 & ~n13965 ;
  assign n13963 = ~n13008 & n13030 ;
  assign n13296 = n13017 ^ n12988 ;
  assign n13297 = n13296 ^ n13040 ;
  assign n13298 = ~n12927 & n13297 ;
  assign n13301 = n13298 ^ n13015 ;
  assign n13960 = n12927 & n12997 ;
  assign n13961 = n13960 ^ n12926 ;
  assign n13962 = ~n13301 & ~n13961 ;
  assign n13964 = n13963 ^ n13962 ;
  assign n13967 = n13966 ^ n13964 ;
  assign n13955 = n13004 ^ n12994 ;
  assign n13956 = ~n13008 & n13955 ;
  assign n13968 = n13967 ^ n13956 ;
  assign n13969 = n13968 ^ n13010 ;
  assign n13950 = n13010 ^ n12926 ;
  assign n13951 = n13950 ^ n13010 ;
  assign n13952 = ~n13021 & ~n13951 ;
  assign n13953 = n13952 ^ n13010 ;
  assign n13954 = n12925 & n13953 ;
  assign n13970 = n13969 ^ n13954 ;
  assign n13971 = n13970 ^ n12987 ;
  assign n13035 = n13034 ^ n13028 ;
  assign n13036 = ~n13002 & n13035 ;
  assign n13037 = n13036 ^ n13034 ;
  assign n13972 = n13971 ^ n13037 ;
  assign n13973 = n13972 ^ n10851 ;
  assign n13943 = n12987 ^ n12926 ;
  assign n13944 = n13943 ^ n12987 ;
  assign n13945 = n13032 & ~n13944 ;
  assign n13946 = n13945 ^ n12987 ;
  assign n13947 = ~n13002 & n13946 ;
  assign n13974 = n13973 ^ n13947 ;
  assign n14716 = n13974 ^ x112 ;
  assign n12381 = n12306 ^ n12296 ;
  assign n12382 = n12381 ^ n12306 ;
  assign n12387 = n12382 & ~n12384 ;
  assign n12388 = n12387 ^ n12306 ;
  assign n12389 = ~n12297 & n12388 ;
  assign n12307 = n12301 & n12306 ;
  assign n12312 = n12311 ^ n12307 ;
  assign n14706 = n12325 ^ n12309 ;
  assign n14707 = ~n12299 & ~n14706 ;
  assign n14692 = n12315 ^ n12250 ;
  assign n14693 = ~n12296 & ~n14692 ;
  assign n14691 = n13776 ^ n12310 ;
  assign n14694 = n14693 ^ n14691 ;
  assign n14697 = n14694 ^ n12349 ;
  assign n14700 = n14697 ^ n12248 ;
  assign n14701 = n14700 ^ n14697 ;
  assign n14702 = ~n12296 & n14701 ;
  assign n14703 = n14702 ^ n14697 ;
  assign n14704 = ~n12297 & ~n14703 ;
  assign n12302 = n12254 & n12301 ;
  assign n14695 = n14694 ^ n12302 ;
  assign n14696 = n14695 ^ n13756 ;
  assign n14705 = n14704 ^ n14696 ;
  assign n14708 = n14707 ^ n14705 ;
  assign n14709 = n14708 ^ n12334 ;
  assign n14690 = n12298 & n12320 ;
  assign n14710 = n14709 ^ n14690 ;
  assign n14683 = n12334 ^ n12300 ;
  assign n14684 = n13766 ^ n12298 ;
  assign n14685 = n12334 ^ n12298 ;
  assign n14686 = n14685 ^ n12298 ;
  assign n14687 = n14684 & ~n14686 ;
  assign n14688 = n14687 ^ n12298 ;
  assign n14689 = n14683 & ~n14688 ;
  assign n14711 = n14710 ^ n14689 ;
  assign n14712 = ~n12312 & ~n14711 ;
  assign n14713 = ~n12389 & n14712 ;
  assign n14714 = n14713 ^ n12199 ;
  assign n14715 = n14714 ^ x65 ;
  assign n14759 = n14716 ^ n14715 ;
  assign n10784 = n10783 ^ x73 ;
  assign n11082 = n11081 ^ x64 ;
  assign n11083 = n10784 & ~n11082 ;
  assign n9918 = n9855 ^ n8958 ;
  assign n9919 = n9918 ^ n9855 ;
  assign n9920 = n9876 ^ n9855 ;
  assign n9921 = ~n9919 & n9920 ;
  assign n9922 = n9921 ^ n9855 ;
  assign n9923 = ~n9910 & n9922 ;
  assign n9924 = n9923 ^ n9855 ;
  assign n9925 = n9924 ^ n9859 ;
  assign n9911 = n9863 ^ n8958 ;
  assign n9912 = n9911 ^ n9863 ;
  assign n9915 = n9875 & n9912 ;
  assign n9916 = n9915 ^ n9863 ;
  assign n9917 = ~n9910 & ~n9916 ;
  assign n9926 = n9925 ^ n9917 ;
  assign n9908 = n9907 ^ n9864 ;
  assign n9909 = n8959 & ~n9908 ;
  assign n9927 = n9926 ^ n9909 ;
  assign n9930 = n9927 ^ n9871 ;
  assign n9931 = n9930 ^ n9927 ;
  assign n9928 = n9927 ^ n9924 ;
  assign n9934 = n9927 ^ n9904 ;
  assign n9935 = n9934 ^ n9927 ;
  assign n9936 = n9928 & n9935 ;
  assign n9937 = n9931 & n9936 ;
  assign n9938 = n9937 ^ n9931 ;
  assign n9939 = n9938 ^ n9930 ;
  assign n9940 = ~n9906 & n9939 ;
  assign n9890 = n9889 ^ n9318 ;
  assign n9903 = n9902 ^ n9890 ;
  assign n9941 = n9940 ^ n9903 ;
  assign n9942 = n9941 ^ x90 ;
  assign n10500 = n10499 ^ n10479 ;
  assign n10501 = n10500 ^ n10497 ;
  assign n10488 = n10449 ^ n10437 ;
  assign n10490 = n10489 ^ n10488 ;
  assign n10491 = n10468 & ~n10490 ;
  assign n10502 = n10501 ^ n10491 ;
  assign n10487 = ~n10045 & ~n10437 ;
  assign n10503 = n10502 ^ n10487 ;
  assign n10480 = n10479 ^ n10045 ;
  assign n10481 = n10480 ^ n10479 ;
  assign n10482 = n10479 ^ n10442 ;
  assign n10483 = n10482 ^ n10479 ;
  assign n10484 = ~n10481 & n10483 ;
  assign n10485 = n10484 ^ n10479 ;
  assign n10486 = n9996 & ~n10485 ;
  assign n10504 = n10503 ^ n10486 ;
  assign n10469 = n10443 ^ n10435 ;
  assign n10470 = n10469 ^ n10443 ;
  assign n10471 = n10443 ^ n9996 ;
  assign n10472 = n10471 ^ n10443 ;
  assign n10473 = n10470 & n10472 ;
  assign n10474 = n10473 ^ n10443 ;
  assign n10475 = ~n10468 & n10474 ;
  assign n10505 = n10504 ^ n10475 ;
  assign n10506 = ~n10467 & n10505 ;
  assign n10514 = n10506 & ~n10513 ;
  assign n10524 = n10514 & ~n10523 ;
  assign n10525 = n10524 ^ n9351 ;
  assign n10526 = n10525 ^ x112 ;
  assign n10527 = ~n9942 & n10526 ;
  assign n11092 = n10527 ^ n10526 ;
  assign n11093 = n11092 ^ n9942 ;
  assign n11094 = n11093 ^ n10526 ;
  assign n11095 = n11083 & ~n11094 ;
  assign n11259 = n11258 ^ x114 ;
  assign n11513 = n11512 ^ x123 ;
  assign n11514 = n11259 & ~n11513 ;
  assign n11515 = n11514 ^ n11259 ;
  assign n11584 = n11095 & n11515 ;
  assign n11087 = n11083 ^ n11082 ;
  assign n11088 = n11087 ^ n10784 ;
  assign n11526 = n11088 & n11092 ;
  assign n14223 = n11514 & n11526 ;
  assign n11084 = n11083 ^ n10784 ;
  assign n11531 = n11084 & ~n11094 ;
  assign n11549 = n11515 ^ n11513 ;
  assign n11550 = n11549 ^ n11259 ;
  assign n11586 = n11531 & ~n11550 ;
  assign n14224 = n14223 ^ n11586 ;
  assign n11090 = n9942 & n11083 ;
  assign n11091 = n11090 ^ n11083 ;
  assign n11096 = n11095 ^ n11091 ;
  assign n11532 = n11531 ^ n11096 ;
  assign n14047 = n11514 & n11532 ;
  assign n11517 = ~n11087 & n11093 ;
  assign n11572 = n11517 & ~n11550 ;
  assign n14048 = n14047 ^ n11572 ;
  assign n11089 = n10527 & n11088 ;
  assign n11551 = n11089 ^ n11088 ;
  assign n11099 = n11088 & n11093 ;
  assign n11527 = n11526 ^ n11099 ;
  assign n11552 = n11551 ^ n11527 ;
  assign n11553 = ~n11550 & n11552 ;
  assign n11516 = n11513 ^ n11259 ;
  assign n11534 = n11526 ^ n11517 ;
  assign n11097 = n11096 ^ n11089 ;
  assign n11085 = n10527 & n11084 ;
  assign n11086 = n11085 ^ n10527 ;
  assign n11098 = n11097 ^ n11086 ;
  assign n11535 = n11534 ^ n11098 ;
  assign n11536 = n11535 ^ n11085 ;
  assign n11518 = n11084 & n11092 ;
  assign n11530 = n11518 ^ n11099 ;
  assign n11533 = n11532 ^ n11530 ;
  assign n11537 = n11536 ^ n11533 ;
  assign n11529 = n11093 ^ n11084 ;
  assign n11538 = n11537 ^ n11529 ;
  assign n11528 = n11527 ^ n11095 ;
  assign n11539 = n11538 ^ n11528 ;
  assign n11100 = n11099 ^ n11098 ;
  assign n11525 = n11100 ^ n11083 ;
  assign n11540 = n11539 ^ n11525 ;
  assign n11541 = n11540 ^ n11534 ;
  assign n11519 = n11518 ^ n11517 ;
  assign n11524 = n11519 ^ n11092 ;
  assign n11542 = n11541 ^ n11524 ;
  assign n11545 = ~n11513 & n11542 ;
  assign n11520 = n11513 & n11519 ;
  assign n11521 = n11520 ^ n11518 ;
  assign n11546 = n11545 ^ n11521 ;
  assign n11547 = ~n11516 & n11546 ;
  assign n11548 = n11547 ^ n11521 ;
  assign n11554 = n11553 ^ n11548 ;
  assign n11589 = n11084 & n11093 ;
  assign n14242 = n11515 & n11589 ;
  assign n11567 = n11540 ^ n11090 ;
  assign n14231 = n11567 ^ n11542 ;
  assign n14232 = n14231 ^ n11089 ;
  assign n14236 = n14232 ^ n11096 ;
  assign n14233 = n14232 ^ n11526 ;
  assign n11590 = n11589 ^ n11540 ;
  assign n11591 = n11590 ^ n11095 ;
  assign n14234 = n14233 ^ n11591 ;
  assign n14235 = n11513 & n14234 ;
  assign n14237 = n14236 ^ n14235 ;
  assign n14238 = n11516 & n14237 ;
  assign n11101 = ~n11087 & ~n11094 ;
  assign n14055 = n11101 ^ n11089 ;
  assign n14056 = n11549 & n14055 ;
  assign n14229 = n14056 ^ n11096 ;
  assign n11573 = n11518 ^ n11101 ;
  assign n11576 = n11513 & n11573 ;
  assign n11577 = n11576 ^ n11101 ;
  assign n11578 = n11259 & n11577 ;
  assign n14230 = n14229 ^ n11578 ;
  assign n14239 = n14238 ^ n14230 ;
  assign n14226 = n11552 ^ n11517 ;
  assign n14227 = n14226 ^ n11100 ;
  assign n14228 = n11515 & n14227 ;
  assign n14240 = n14239 ^ n14228 ;
  assign n14225 = n11530 & ~n11550 ;
  assign n14241 = n14240 ^ n14225 ;
  assign n14243 = n14242 ^ n14241 ;
  assign n14244 = n11095 ^ n11085 ;
  assign n14247 = n11513 & n14244 ;
  assign n14248 = n14247 ^ n11095 ;
  assign n14249 = ~n11259 & n14248 ;
  assign n14250 = ~n14243 & ~n14249 ;
  assign n14251 = ~n11554 & n14250 ;
  assign n14252 = ~n14048 & n14251 ;
  assign n14253 = ~n14224 & n14252 ;
  assign n14254 = ~n11584 & n14253 ;
  assign n14255 = n14254 ^ n9995 ;
  assign n14717 = n14255 ^ x66 ;
  assign n14762 = n14759 ^ n14717 ;
  assign n14718 = n14717 ^ n14716 ;
  assign n14719 = n14715 & n14718 ;
  assign n14720 = n14719 ^ n14717 ;
  assign n14763 = n14762 ^ n14720 ;
  assign n14764 = ~n14754 & ~n14763 ;
  assign n14755 = n14754 ^ n14715 ;
  assign n14765 = n14755 ^ n14716 ;
  assign n14766 = n14718 & n14765 ;
  assign n14767 = n14717 & ~n14766 ;
  assign n14768 = n14766 ^ n14715 ;
  assign n14769 = n14768 ^ n14716 ;
  assign n14770 = n14767 & n14769 ;
  assign n14771 = n14770 ^ n14768 ;
  assign n14772 = ~n14764 & n14771 ;
  assign n15133 = n14772 ^ n14771 ;
  assign n13290 = n13289 ^ n13251 ;
  assign n13291 = ~n13179 & ~n13290 ;
  assign n13280 = n13279 ^ n13246 ;
  assign n13281 = n13246 ^ n13176 ;
  assign n13282 = n13281 ^ n13246 ;
  assign n13283 = ~n13280 & ~n13282 ;
  assign n13284 = n13283 ^ n13246 ;
  assign n13285 = ~n13175 & ~n13284 ;
  assign n14312 = n13789 ^ n13219 ;
  assign n14311 = n13255 ^ n13221 ;
  assign n14315 = n14312 ^ n14311 ;
  assign n14308 = ~n13176 & ~n13242 ;
  assign n14309 = n14308 ^ n13241 ;
  assign n14304 = n13222 ^ n13219 ;
  assign n14305 = n14304 ^ n13279 ;
  assign n14306 = n13176 & n14305 ;
  assign n14307 = n14306 ^ n13222 ;
  assign n14310 = n14309 ^ n14307 ;
  assign n14316 = n14315 ^ n14310 ;
  assign n14300 = n13243 ^ n13221 ;
  assign n14301 = n14300 ^ n13224 ;
  assign n14302 = n14301 ^ n13255 ;
  assign n14303 = ~n13176 & n14302 ;
  assign n14317 = n14316 ^ n14303 ;
  assign n14318 = ~n13175 & n14317 ;
  assign n14319 = n14318 ^ n14309 ;
  assign n14320 = ~n13285 & n14319 ;
  assign n14321 = ~n13788 & n14320 ;
  assign n14322 = ~n13291 & n14321 ;
  assign n14323 = n14322 ^ n10232 ;
  assign n14682 = n14323 ^ x88 ;
  assign n14038 = n13445 ^ n13433 ;
  assign n14039 = n14038 ^ n13479 ;
  assign n14040 = ~n13330 & n14039 ;
  assign n14029 = n13452 ^ n13430 ;
  assign n14041 = n14040 ^ n14029 ;
  assign n14042 = n13329 & n14041 ;
  assign n14023 = n13488 ^ n13443 ;
  assign n14024 = n13443 ^ n13330 ;
  assign n14025 = n14024 ^ n13443 ;
  assign n14026 = n14023 & ~n14025 ;
  assign n14027 = n14026 ^ n13443 ;
  assign n14028 = n13329 & n14027 ;
  assign n14030 = n14029 ^ n14028 ;
  assign n13522 = n13521 ^ n13477 ;
  assign n13523 = n13477 ^ n13330 ;
  assign n13524 = n13523 ^ n13477 ;
  assign n13525 = n13522 & n13524 ;
  assign n13526 = n13525 ^ n13477 ;
  assign n13527 = ~n13329 & n13526 ;
  assign n14031 = n14030 ^ n13527 ;
  assign n14032 = n14031 ^ n13674 ;
  assign n13515 = ~n13513 & n13514 ;
  assign n13516 = n13515 ^ n13511 ;
  assign n14033 = n14032 ^ n13516 ;
  assign n13440 = n13439 ^ n13427 ;
  assign n13450 = n13449 ^ n13440 ;
  assign n13416 = n13415 ^ n13373 ;
  assign n13451 = n13450 ^ n13416 ;
  assign n13455 = n13454 ^ n13451 ;
  assign n13496 = ~n13455 & n13466 ;
  assign n13490 = n13445 ^ n13437 ;
  assign n13491 = n13445 ^ n13329 ;
  assign n13492 = n13491 ^ n13445 ;
  assign n13493 = n13490 & ~n13492 ;
  assign n13494 = n13493 ^ n13445 ;
  assign n13495 = ~n13458 & n13494 ;
  assign n13497 = n13496 ^ n13495 ;
  assign n14034 = n14033 ^ n13497 ;
  assign n14035 = n14034 ^ n10923 ;
  assign n14016 = n13479 ^ n13446 ;
  assign n14015 = n13513 ^ n13454 ;
  assign n14017 = n14016 ^ n14015 ;
  assign n14018 = n14016 ^ n13330 ;
  assign n14019 = n14018 ^ n14016 ;
  assign n14020 = ~n14017 & n14019 ;
  assign n14021 = n14020 ^ n14016 ;
  assign n14022 = ~n13329 & n14021 ;
  assign n14036 = n14035 ^ n14022 ;
  assign n14012 = n13487 ^ n13420 ;
  assign n14013 = n14012 ^ n13438 ;
  assign n14014 = n13466 & n14013 ;
  assign n14037 = n14036 ^ n14014 ;
  assign n14043 = n14042 ^ n14037 ;
  assign n14681 = n14043 ^ x106 ;
  assign n15134 = n14682 ^ n14681 ;
  assign n15141 = n14764 ^ n14762 ;
  assign n14760 = n14759 ^ n14754 ;
  assign n15135 = ~n14717 & n14760 ;
  assign n14778 = n14754 ^ n14716 ;
  assign n14790 = ~n14717 & ~n14754 ;
  assign n14791 = n14778 & ~n14790 ;
  assign n15136 = n15135 ^ n14791 ;
  assign n14756 = ~n14717 & n14755 ;
  assign n14757 = n14756 ^ n14754 ;
  assign n14758 = ~n14718 & ~n14757 ;
  assign n14761 = n14760 ^ n14758 ;
  assign n15137 = n15136 ^ n14761 ;
  assign n15138 = n14681 & n15137 ;
  assign n15139 = n15138 ^ n15136 ;
  assign n15142 = n15141 ^ n15139 ;
  assign n15140 = n15139 ^ n14771 ;
  assign n15143 = n15142 ^ n15140 ;
  assign n15144 = n15142 ^ n14682 ;
  assign n15145 = n15144 ^ n15142 ;
  assign n15146 = n15143 & n15145 ;
  assign n15147 = n15146 ^ n15142 ;
  assign n15148 = n15134 & ~n15147 ;
  assign n15149 = n15148 ^ n15139 ;
  assign n15150 = ~n15133 & ~n15149 ;
  assign n15151 = n15150 ^ n12570 ;
  assign n15152 = n15151 ^ x76 ;
  assign n15153 = n15132 & n15152 ;
  assign n13053 = n13052 ^ n12989 ;
  assign n13054 = n12927 & n13053 ;
  assign n13046 = n13014 ^ n12982 ;
  assign n13047 = n13046 ^ n13030 ;
  assign n13041 = n13040 ^ n13003 ;
  assign n13038 = n13015 ^ n12995 ;
  assign n13042 = n13041 ^ n13038 ;
  assign n13043 = n12925 & ~n13042 ;
  assign n13049 = n13047 ^ n13043 ;
  assign n13050 = n13002 & ~n13049 ;
  assign n13044 = n13043 ^ n13037 ;
  assign n13024 = n13023 ^ n8957 ;
  assign n13045 = n13044 ^ n13024 ;
  assign n13051 = n13050 ^ n13045 ;
  assign n13055 = n13054 ^ n13051 ;
  assign n13005 = n13004 ^ n12935 ;
  assign n13006 = n13002 & n13005 ;
  assign n13056 = n13055 ^ n13006 ;
  assign n13001 = ~n12999 & ~n13000 ;
  assign n13057 = n13056 ^ n13001 ;
  assign n12991 = n12990 ^ n12976 ;
  assign n12992 = ~n12925 & ~n12991 ;
  assign n13058 = n13057 ^ n12992 ;
  assign n12977 = n12927 & n12976 ;
  assign n13059 = n13058 ^ n12977 ;
  assign n13060 = n13059 ^ x94 ;
  assign n12695 = ~n12645 & ~n12670 ;
  assign n12691 = n12690 ^ n12657 ;
  assign n12692 = n12630 & ~n12691 ;
  assign n12572 = n12571 ^ n12541 ;
  assign n12609 = n12608 ^ n12572 ;
  assign n12614 = n12613 ^ n12541 ;
  assign n12615 = n12614 ^ n12608 ;
  assign n12616 = n12615 ^ n12614 ;
  assign n12619 = n12618 ^ n12541 ;
  assign n12620 = n12619 ^ n12614 ;
  assign n12621 = ~n12616 & n12620 ;
  assign n12622 = n12621 ^ n12614 ;
  assign n12623 = n12609 & n12622 ;
  assign n12624 = n12623 ^ n12541 ;
  assign n12685 = n12684 ^ n12624 ;
  assign n12666 = n12665 ^ n12632 ;
  assign n12669 = ~n12667 & n12668 ;
  assign n12671 = n12670 ^ n12669 ;
  assign n12672 = n12671 ^ n12669 ;
  assign n12673 = ~n12639 & n12672 ;
  assign n12674 = n12666 & n12673 ;
  assign n12675 = n12674 ^ n12671 ;
  assign n12686 = n12685 ^ n12675 ;
  assign n12679 = n12678 ^ n12647 ;
  assign n12680 = n12571 & ~n12679 ;
  assign n12681 = n12675 & n12680 ;
  assign n12687 = n12686 ^ n12681 ;
  assign n12693 = n12692 ^ n12687 ;
  assign n12626 = ~n12571 & n12625 ;
  assign n12627 = ~n12624 & n12626 ;
  assign n12694 = n12693 ^ n12627 ;
  assign n12696 = n12695 ^ n12694 ;
  assign n12704 = ~n12696 & ~n12703 ;
  assign n12705 = n12704 ^ n9238 ;
  assign n12706 = n12705 ^ x124 ;
  assign n11557 = n11526 ^ n11513 ;
  assign n11558 = n11557 ^ n11526 ;
  assign n11559 = n11552 & n11558 ;
  assign n11560 = n11559 ^ n11526 ;
  assign n11561 = n11516 & n11560 ;
  assign n11562 = n11561 ^ n11526 ;
  assign n11579 = n11099 & n11514 ;
  assign n11580 = n11579 ^ n11578 ;
  assign n11581 = n11580 ^ n11572 ;
  assign n11568 = n11567 ^ n11085 ;
  assign n11582 = n11581 ^ n11568 ;
  assign n11569 = n11568 ^ n11097 ;
  assign n11563 = n10784 ^ n10526 ;
  assign n11564 = n11563 ^ n11097 ;
  assign n11565 = n11564 ^ n11538 ;
  assign n11566 = ~n11259 & n11565 ;
  assign n11570 = n11569 ^ n11566 ;
  assign n11571 = n11516 & n11570 ;
  assign n11583 = n11582 ^ n11571 ;
  assign n11585 = n11584 ^ n11583 ;
  assign n11587 = n11586 ^ n11585 ;
  assign n11588 = ~n11513 & ~n11587 ;
  assign n11592 = n11591 ^ n11098 ;
  assign n11595 = n11259 & n11592 ;
  assign n11596 = n11595 ^ n11098 ;
  assign n11597 = n11588 & n11596 ;
  assign n11598 = n11597 ^ n11587 ;
  assign n11599 = ~n11562 & ~n11598 ;
  assign n11600 = ~n11554 & n11599 ;
  assign n11603 = n11600 ^ n9495 ;
  assign n11102 = n11101 ^ n11100 ;
  assign n11601 = n11515 & n11600 ;
  assign n11602 = n11102 & n11601 ;
  assign n11604 = n11603 ^ n11602 ;
  assign n11605 = n11604 ^ x76 ;
  assign n13096 = n12706 ^ n11605 ;
  assign n11656 = n11655 ^ x122 ;
  assign n11689 = n11688 ^ x104 ;
  assign n11964 = n11963 ^ x82 ;
  assign n11780 = ~n10984 & n11035 ;
  assign n11769 = n10992 ^ n10971 ;
  assign n11773 = n11772 ^ n11769 ;
  assign n11767 = n11014 ^ n10990 ;
  assign n11768 = ~n10852 & n11767 ;
  assign n11774 = n11773 ^ n11768 ;
  assign n11776 = n11769 ^ n10818 ;
  assign n11775 = n11769 ^ n10852 ;
  assign n11777 = n11776 ^ n11775 ;
  assign n11778 = n11774 & ~n11777 ;
  assign n11779 = n11778 ^ n11775 ;
  assign n11781 = n11780 ^ n11779 ;
  assign n11761 = n10988 ^ n10852 ;
  assign n11762 = n10988 ^ n10818 ;
  assign n11763 = n11016 ^ n10818 ;
  assign n11764 = ~n11762 & ~n11763 ;
  assign n11765 = n11764 ^ n10818 ;
  assign n11766 = n11761 & n11765 ;
  assign n11782 = n11781 ^ n11766 ;
  assign n11783 = n11782 ^ n10976 ;
  assign n11759 = n11074 ^ n10976 ;
  assign n11760 = n10986 & n11759 ;
  assign n11784 = n11783 ^ n11760 ;
  assign n11785 = n11019 ^ n10977 ;
  assign n11786 = ~n10852 & ~n11785 ;
  assign n11787 = n11786 ^ n10977 ;
  assign n11788 = n11787 ^ n10818 ;
  assign n11789 = n11788 ^ n11787 ;
  assign n11790 = ~n10852 & n11005 ;
  assign n11791 = n11790 ^ n11787 ;
  assign n11792 = ~n11789 & n11791 ;
  assign n11793 = n11792 ^ n11787 ;
  assign n11794 = ~n11784 & ~n11793 ;
  assign n11795 = n11794 ^ n9589 ;
  assign n11796 = n11795 ^ x81 ;
  assign n11721 = n11720 ^ n9624 ;
  assign n11703 = n10740 ^ n10726 ;
  assign n11704 = n11703 ^ n10768 ;
  assign n11705 = n10543 & n11704 ;
  assign n11713 = n11705 ^ n10723 ;
  assign n11710 = ~n10543 & ~n11709 ;
  assign n11699 = n10777 ^ n10706 ;
  assign n11698 = n10720 ^ n10709 ;
  assign n11700 = n11699 ^ n11698 ;
  assign n11701 = ~n10543 & ~n11700 ;
  assign n11702 = n11701 ^ n11698 ;
  assign n11711 = n11710 ^ n11702 ;
  assign n11714 = n11713 ^ n11711 ;
  assign n11715 = ~n10732 & n11714 ;
  assign n11706 = n11705 ^ n11702 ;
  assign n11707 = n11706 ^ n11697 ;
  assign n11708 = n11707 ^ n10751 ;
  assign n11712 = n11711 ^ n11708 ;
  assign n11716 = n11715 ^ n11712 ;
  assign n11717 = ~n10739 & ~n11716 ;
  assign n11722 = n11721 ^ n11717 ;
  assign n11723 = n11722 ^ x72 ;
  assign n11966 = n11796 ^ n11723 ;
  assign n11967 = ~n11964 & ~n11966 ;
  assign n12016 = n11967 ^ n11964 ;
  assign n11757 = n11756 ^ x99 ;
  assign n11971 = ~n11723 & ~n11757 ;
  assign n11972 = n11971 ^ n11796 ;
  assign n11973 = n11972 ^ n11723 ;
  assign n11969 = n11757 & ~n11796 ;
  assign n11970 = n11969 ^ n11757 ;
  assign n11974 = n11973 ^ n11970 ;
  assign n11975 = ~n11964 & n11974 ;
  assign n12013 = n11975 ^ n11969 ;
  assign n11965 = n11964 ^ n11796 ;
  assign n11979 = n11965 ^ n11757 ;
  assign n11996 = n11969 & ~n11979 ;
  assign n12014 = n12013 ^ n11996 ;
  assign n11758 = n11757 ^ n11723 ;
  assign n12015 = n12014 ^ n11758 ;
  assign n12017 = n12016 ^ n12015 ;
  assign n11994 = n11965 ^ n11723 ;
  assign n11995 = n11979 ^ n11796 ;
  assign n11997 = n11996 ^ n11995 ;
  assign n11998 = ~n11994 & ~n11997 ;
  assign n11993 = n11970 ^ n11796 ;
  assign n11999 = n11998 ^ n11993 ;
  assign n12000 = n11999 ^ n11995 ;
  assign n12001 = n12000 ^ n11965 ;
  assign n11990 = n11723 & n11964 ;
  assign n11991 = ~n11969 & n11990 ;
  assign n11982 = ~n11796 & ~n11979 ;
  assign n11989 = n11982 ^ n11979 ;
  assign n11992 = n11991 ^ n11989 ;
  assign n12002 = n12001 ^ n11992 ;
  assign n12003 = n12002 ^ n11723 ;
  assign n12008 = n11966 & n12003 ;
  assign n12009 = n12008 ^ n11964 ;
  assign n12010 = n11758 & n12009 ;
  assign n12011 = n12010 ^ n12003 ;
  assign n12012 = n12011 ^ n11991 ;
  assign n12018 = n12017 ^ n12012 ;
  assign n12019 = ~n11689 & n12018 ;
  assign n12020 = n12019 ^ n12015 ;
  assign n11976 = n11975 ^ n11972 ;
  assign n11968 = n11967 ^ n11965 ;
  assign n11977 = n11976 ^ n11968 ;
  assign n11797 = n11796 ^ n11758 ;
  assign n11978 = n11977 ^ n11797 ;
  assign n11980 = n11979 ^ n11978 ;
  assign n11981 = n11980 ^ n11964 ;
  assign n11983 = n11982 ^ n11981 ;
  assign n11984 = n11983 ^ n11978 ;
  assign n11985 = ~n11723 & ~n11984 ;
  assign n11986 = n11985 ^ n11980 ;
  assign n11987 = n11689 & n11986 ;
  assign n11988 = n11987 ^ n11978 ;
  assign n12021 = n12020 ^ n11988 ;
  assign n12022 = ~n11656 & n12021 ;
  assign n12023 = n12022 ^ n12020 ;
  assign n12024 = n12023 ^ n9662 ;
  assign n12025 = n12024 ^ x67 ;
  assign n13073 = ~n12025 & ~n12706 ;
  assign n12313 = n12297 ^ n12296 ;
  assign n12371 = n12313 & n12338 ;
  assign n12364 = n12363 ^ n12327 ;
  assign n12365 = n12364 ^ n12346 ;
  assign n12366 = n12365 ^ n12360 ;
  assign n12367 = n12296 & ~n12366 ;
  assign n12352 = n12340 ^ n12310 ;
  assign n12351 = n12350 ^ n12130 ;
  assign n12353 = n12352 ^ n12351 ;
  assign n12354 = ~n12296 & ~n12353 ;
  assign n12355 = n12354 ^ n12352 ;
  assign n12361 = n12360 ^ n12355 ;
  assign n12368 = n12367 ^ n12361 ;
  assign n12369 = n12297 & n12368 ;
  assign n12328 = n12327 ^ n12306 ;
  assign n12329 = n12327 ^ n12296 ;
  assign n12330 = n12329 ^ n12327 ;
  assign n12331 = ~n12328 & n12330 ;
  assign n12332 = n12331 ^ n12327 ;
  assign n12333 = n12313 & ~n12332 ;
  assign n12356 = n12355 ^ n12333 ;
  assign n12370 = n12369 ^ n12356 ;
  assign n12372 = n12371 ^ n12370 ;
  assign n12373 = ~n12312 & ~n12372 ;
  assign n12380 = n12373 & ~n12379 ;
  assign n12390 = n12380 & ~n12389 ;
  assign n12391 = ~n12302 & n12390 ;
  assign n12392 = n12391 ^ n9838 ;
  assign n12393 = n12392 ^ x117 ;
  assign n13097 = n13073 ^ n12393 ;
  assign n13098 = ~n13096 & n13097 ;
  assign n12707 = n12393 & ~n12706 ;
  assign n12708 = n12707 ^ n12706 ;
  assign n12709 = n12708 ^ n12393 ;
  assign n12026 = ~n11605 & ~n12025 ;
  assign n12712 = n12026 ^ n12025 ;
  assign n12716 = n12709 & ~n12712 ;
  assign n12713 = n12712 ^ n11605 ;
  assign n12714 = n12713 ^ n12025 ;
  assign n12715 = n12709 & ~n12714 ;
  assign n12717 = n12716 ^ n12715 ;
  assign n12710 = n12026 & n12709 ;
  assign n12711 = n12710 ^ n12709 ;
  assign n12718 = n12717 ^ n12711 ;
  assign n13106 = n13098 ^ n12718 ;
  assign n13068 = ~n12708 & ~n12713 ;
  assign n13069 = n13068 ^ n12710 ;
  assign n13065 = ~n12708 & ~n12712 ;
  assign n13105 = n13069 ^ n13065 ;
  assign n13107 = n13106 ^ n13105 ;
  assign n12921 = n12755 & ~n12920 ;
  assign n12897 = n12838 ^ n12757 ;
  assign n12898 = n12897 ^ n12859 ;
  assign n12899 = n12898 ^ n12874 ;
  assign n12900 = n12750 & n12899 ;
  assign n12901 = n12900 ^ n12859 ;
  assign n12902 = n12756 & n12901 ;
  assign n12903 = n12902 ^ n12859 ;
  assign n12913 = n12877 ^ n12864 ;
  assign n12906 = n12905 ^ n12863 ;
  assign n12887 = n12867 ^ n12856 ;
  assign n12904 = n12887 ^ n12870 ;
  assign n12907 = n12906 ^ n12904 ;
  assign n12908 = ~n12750 & ~n12907 ;
  assign n12914 = n12913 ^ n12908 ;
  assign n12909 = n12877 ^ n12865 ;
  assign n12910 = n12909 ^ n12851 ;
  assign n12911 = n12910 ^ n12864 ;
  assign n12912 = ~n12750 & n12911 ;
  assign n12915 = n12914 ^ n12912 ;
  assign n12916 = n12751 & n12915 ;
  assign n12917 = n12916 ^ n12908 ;
  assign n12918 = ~n12903 & ~n12917 ;
  assign n12890 = n12875 ^ n12867 ;
  assign n12891 = n12867 ^ n12750 ;
  assign n12892 = n12891 ^ n12867 ;
  assign n12893 = n12890 & ~n12892 ;
  assign n12894 = n12893 ^ n12867 ;
  assign n12895 = n12756 & n12894 ;
  assign n12888 = n12754 & n12887 ;
  assign n12889 = n12888 ^ n12886 ;
  assign n12896 = n12895 ^ n12889 ;
  assign n12919 = n12918 ^ n12896 ;
  assign n12922 = n12921 ^ n12919 ;
  assign n12923 = n12922 ^ n8422 ;
  assign n12924 = n12923 ^ x85 ;
  assign n15263 = n13107 ^ n12924 ;
  assign n15264 = n15263 ^ n13107 ;
  assign n15266 = n13107 ^ n13069 ;
  assign n15267 = ~n15264 & ~n15266 ;
  assign n15268 = n15267 ^ n13107 ;
  assign n15269 = n13060 & ~n15268 ;
  assign n13064 = n13060 ^ n12924 ;
  assign n13087 = ~n11605 & ~n12706 ;
  assign n13070 = n12026 & ~n12708 ;
  assign n13077 = n13070 ^ n12716 ;
  assign n13075 = n12709 ^ n12706 ;
  assign n13076 = ~n12712 & n13075 ;
  assign n13078 = n13077 ^ n13076 ;
  assign n13074 = n13073 ^ n12712 ;
  assign n13079 = n13078 ^ n13074 ;
  assign n13080 = n13079 ^ n13076 ;
  assign n13100 = n13087 ^ n13080 ;
  assign n13071 = n13070 ^ n13069 ;
  assign n13066 = n13065 ^ n12710 ;
  assign n13067 = n13066 ^ n12708 ;
  assign n13072 = n13071 ^ n13067 ;
  assign n13099 = n13098 ^ n13072 ;
  assign n13101 = n13100 ^ n13099 ;
  assign n15253 = n13101 ^ n13080 ;
  assign n13112 = n12707 & ~n12712 ;
  assign n13092 = n12707 & ~n12713 ;
  assign n13093 = n13092 ^ n13080 ;
  assign n13088 = n13087 ^ n12025 ;
  assign n13089 = n12393 & n13088 ;
  assign n13090 = n13089 ^ n12393 ;
  assign n13091 = n13090 ^ n12707 ;
  assign n13094 = n13093 ^ n13091 ;
  assign n13095 = n13094 ^ n13076 ;
  assign n13113 = n13112 ^ n13095 ;
  assign n13114 = n13113 ^ n13090 ;
  assign n13130 = n13114 ^ n13112 ;
  assign n15251 = n13130 ^ n13070 ;
  assign n15252 = n15251 ^ n12718 ;
  assign n15254 = n15253 ^ n15252 ;
  assign n15255 = n15254 ^ n13066 ;
  assign n15256 = n15255 ^ n15252 ;
  assign n15257 = n15252 ^ n13060 ;
  assign n15258 = n15257 ^ n15252 ;
  assign n15259 = ~n15256 & ~n15258 ;
  assign n15260 = n15259 ^ n15252 ;
  assign n15261 = ~n13064 & ~n15260 ;
  assign n15262 = n15261 ^ n15252 ;
  assign n15270 = n15269 ^ n15262 ;
  assign n15279 = n15270 ^ n12425 ;
  assign n13115 = n13101 ^ n13094 ;
  assign n13116 = n13115 ^ n13114 ;
  assign n13117 = n13114 ^ n13060 ;
  assign n13118 = n13117 ^ n13114 ;
  assign n13119 = n13116 & n13118 ;
  assign n13120 = n13119 ^ n13114 ;
  assign n13121 = ~n12924 & ~n13120 ;
  assign n15280 = n15279 ^ n13121 ;
  assign n15271 = ~n13060 & n15270 ;
  assign n15276 = n12924 & ~n13095 ;
  assign n15277 = n15276 ^ n12717 ;
  assign n15278 = n15271 & n15277 ;
  assign n15281 = n15280 ^ n15278 ;
  assign n15282 = n15281 ^ x100 ;
  assign n14121 = n11988 ^ n11656 ;
  assign n14122 = n14121 ^ n12022 ;
  assign n14123 = n14122 ^ n10963 ;
  assign n14854 = n14123 ^ x108 ;
  assign n14876 = n13437 & n13514 ;
  assign n14871 = n14028 ^ n13495 ;
  assign n14866 = n13521 ^ n13432 ;
  assign n14867 = n14866 ^ n13443 ;
  assign n14868 = n13514 & ~n14867 ;
  assign n14869 = n14868 ^ n13434 ;
  assign n14870 = n13329 & ~n14869 ;
  assign n14872 = n14871 ^ n14870 ;
  assign n14865 = n13466 & ~n13478 ;
  assign n14873 = n14872 ^ n14865 ;
  assign n14861 = n13449 ^ n13438 ;
  assign n14862 = n14861 ^ n13479 ;
  assign n13456 = n13455 ^ n13445 ;
  assign n14863 = n14862 ^ n13456 ;
  assign n14864 = n13331 & ~n14863 ;
  assign n14874 = n14873 ^ n14864 ;
  assign n13332 = n13331 ^ n13329 ;
  assign n14858 = n13473 ^ n13374 ;
  assign n14859 = n14858 ^ n13477 ;
  assign n14860 = ~n13332 & ~n14859 ;
  assign n14875 = n14874 ^ n14860 ;
  assign n14877 = n14876 ^ n14875 ;
  assign n14878 = ~n13649 & ~n14877 ;
  assign n14879 = n14878 ^ n11167 ;
  assign n14880 = n14879 ^ x86 ;
  assign n13999 = n12629 & n12665 ;
  assign n13995 = n12689 ^ n12613 ;
  assign n13996 = ~n12571 & n13995 ;
  assign n13992 = n13991 ^ n12669 ;
  assign n13981 = n12668 ^ n12645 ;
  assign n13979 = n12653 ^ n12541 ;
  assign n13982 = n13981 ^ n13979 ;
  assign n13983 = n12608 & n13982 ;
  assign n13980 = n13979 ^ n12625 ;
  assign n13984 = n13983 ^ n13980 ;
  assign n13985 = ~n12670 & ~n13984 ;
  assign n13993 = n13992 ^ n13985 ;
  assign n13977 = n12640 ^ n12541 ;
  assign n13978 = n12631 & n13977 ;
  assign n13994 = n13993 ^ n13978 ;
  assign n13997 = n13996 ^ n13994 ;
  assign n13976 = ~n12608 & n12689 ;
  assign n13998 = n13997 ^ n13976 ;
  assign n14000 = n13999 ^ n13998 ;
  assign n14001 = ~n12683 & ~n14000 ;
  assign n14002 = n13712 ^ n12608 ;
  assign n14003 = n14002 ^ n13712 ;
  assign n14006 = ~n13721 & n14003 ;
  assign n14007 = n14006 ^ n13712 ;
  assign n14008 = n14001 & ~n14007 ;
  assign n14009 = n14008 ^ n10817 ;
  assign n14881 = n14009 ^ x126 ;
  assign n14882 = ~n14880 & ~n14881 ;
  assign n14883 = n14882 ^ n14881 ;
  assign n14884 = n14883 ^ n14880 ;
  assign n14885 = n13059 ^ x84 ;
  assign n14909 = n13276 ^ n13224 ;
  assign n14910 = n13175 & ~n14909 ;
  assign n14888 = n13175 & n13250 ;
  assign n14889 = n14888 ^ n13217 ;
  assign n14908 = n14889 ^ n13222 ;
  assign n14911 = n14910 ^ n14908 ;
  assign n14912 = n13176 & n14911 ;
  assign n14906 = n13178 & n13210 ;
  assign n14893 = n13792 ^ n13277 ;
  assign n14891 = n13245 ^ n13233 ;
  assign n14892 = n14891 ^ n13243 ;
  assign n14894 = n14893 ^ n14892 ;
  assign n14895 = n13176 & ~n14894 ;
  assign n14896 = n14895 ^ n14893 ;
  assign n14898 = n14896 ^ n13231 ;
  assign n14899 = n14898 ^ n13244 ;
  assign n14900 = n14899 ^ n13795 ;
  assign n14901 = n14900 ^ n14896 ;
  assign n14902 = n13176 & n14901 ;
  assign n14903 = n14902 ^ n14898 ;
  assign n14904 = ~n13175 & n14903 ;
  assign n14890 = n14889 ^ n13291 ;
  assign n14897 = n14896 ^ n14890 ;
  assign n14905 = n14904 ^ n14897 ;
  assign n14907 = n14906 ^ n14905 ;
  assign n14913 = n14912 ^ n14907 ;
  assign n14914 = n14913 ^ n13790 ;
  assign n14886 = n14307 ^ n13790 ;
  assign n14887 = ~n13175 & n14886 ;
  assign n14915 = n14914 ^ n14887 ;
  assign n14916 = ~n13788 & ~n14915 ;
  assign n14917 = ~n13256 & n14916 ;
  assign n14918 = n14917 ^ n11146 ;
  assign n14919 = n14918 ^ x101 ;
  assign n14920 = ~n14885 & n14919 ;
  assign n14921 = n14920 ^ n14919 ;
  assign n14929 = n14921 ^ n14885 ;
  assign n14942 = ~n14884 & n14929 ;
  assign n14941 = ~n14884 & n14920 ;
  assign n14943 = n14942 ^ n14941 ;
  assign n14922 = ~n14884 & n14921 ;
  assign n14940 = n14922 ^ n14884 ;
  assign n14944 = n14943 ^ n14940 ;
  assign n14925 = n14920 ^ n14885 ;
  assign n14948 = n14944 ^ n14925 ;
  assign n14935 = n14882 & ~n14925 ;
  assign n14926 = ~n14883 & ~n14925 ;
  assign n14947 = n14935 ^ n14926 ;
  assign n14949 = n14948 ^ n14947 ;
  assign n14950 = n14949 ^ n14943 ;
  assign n14951 = n14950 ^ n14881 ;
  assign n14930 = ~n14883 & n14929 ;
  assign n14928 = ~n14883 & n14920 ;
  assign n14931 = n14930 ^ n14928 ;
  assign n14927 = n14926 ^ n14883 ;
  assign n14932 = n14931 ^ n14927 ;
  assign n14924 = n14882 & n14921 ;
  assign n14933 = n14932 ^ n14924 ;
  assign n14923 = n14922 ^ n14921 ;
  assign n14934 = n14933 ^ n14923 ;
  assign n14945 = n14944 ^ n14934 ;
  assign n14937 = n14884 ^ n14881 ;
  assign n14938 = n14920 & ~n14937 ;
  assign n14939 = n14938 ^ n14922 ;
  assign n14946 = n14945 ^ n14939 ;
  assign n14952 = n14951 ^ n14946 ;
  assign n14963 = n14952 ^ n14944 ;
  assign n14971 = n14963 ^ n14949 ;
  assign n14853 = n12392 ^ x125 ;
  assign n14972 = n14949 ^ n14853 ;
  assign n14973 = n14972 ^ n14949 ;
  assign n14974 = ~n14971 & n14973 ;
  assign n14975 = n14974 ^ n14949 ;
  assign n14976 = n14854 & n14975 ;
  assign n14855 = n14853 & ~n14854 ;
  assign n14856 = n14855 ^ n14854 ;
  assign n15326 = n14935 ^ n14930 ;
  assign n15327 = ~n14856 & n15326 ;
  assign n14857 = n14856 ^ n14853 ;
  assign n15323 = n14857 ^ n14854 ;
  assign n14959 = n14882 & n14920 ;
  assign n15324 = n14959 ^ n14932 ;
  assign n15325 = n15323 & ~n15324 ;
  assign n15328 = n15327 ^ n15325 ;
  assign n14977 = n14854 ^ n14853 ;
  assign n15314 = n14924 ^ n14854 ;
  assign n15315 = n15314 ^ n14924 ;
  assign n15318 = n14952 & ~n15315 ;
  assign n15319 = n15318 ^ n14924 ;
  assign n15320 = ~n14977 & n15319 ;
  assign n15308 = n14935 ^ n14854 ;
  assign n15309 = n15308 ^ n14935 ;
  assign n15310 = n14947 & n15309 ;
  assign n15311 = n15310 ^ n14935 ;
  assign n15312 = n14977 & n15311 ;
  assign n15313 = n15312 ^ n14924 ;
  assign n15321 = n15320 ^ n15313 ;
  assign n15296 = n14933 ^ n14921 ;
  assign n15297 = n15296 ^ n14938 ;
  assign n15298 = n15297 ^ n14926 ;
  assign n15299 = n15298 ^ n15296 ;
  assign n15300 = n15296 ^ n14854 ;
  assign n15301 = n15300 ^ n15296 ;
  assign n15302 = n15299 & ~n15301 ;
  assign n15303 = n15302 ^ n15296 ;
  assign n15304 = ~n14977 & ~n15303 ;
  assign n15305 = n15304 ^ n15296 ;
  assign n15290 = n14949 ^ n14935 ;
  assign n15291 = n14935 ^ n14853 ;
  assign n15292 = n15291 ^ n14935 ;
  assign n15293 = n15290 & n15292 ;
  assign n15294 = n15293 ^ n14935 ;
  assign n15295 = n14854 & n15294 ;
  assign n15306 = n15305 ^ n15295 ;
  assign n15307 = n15306 ^ n14943 ;
  assign n15322 = n15321 ^ n15307 ;
  assign n15329 = n15328 ^ n15322 ;
  assign n14978 = n14932 ^ n14931 ;
  assign n14979 = n14978 ^ n14854 ;
  assign n14980 = n14979 ^ n14978 ;
  assign n14960 = n14959 ^ n14924 ;
  assign n14961 = n14960 ^ n14935 ;
  assign n14981 = n14961 ^ n14882 ;
  assign n14982 = n14981 ^ n14931 ;
  assign n14983 = n14982 ^ n14978 ;
  assign n14984 = n14980 & ~n14983 ;
  assign n14985 = n14984 ^ n14978 ;
  assign n14986 = ~n14977 & ~n14985 ;
  assign n14987 = n14986 ^ n14931 ;
  assign n15330 = n15329 ^ n14987 ;
  assign n15283 = n14943 ^ n14854 ;
  assign n15284 = n15283 ^ n14943 ;
  assign n15287 = ~n14963 & ~n15284 ;
  assign n15288 = n15287 ^ n14943 ;
  assign n15289 = n14977 & n15288 ;
  assign n15331 = n15330 ^ n15289 ;
  assign n15332 = ~n14976 & n15331 ;
  assign n15333 = n15332 ^ n12537 ;
  assign n15334 = n15333 ^ x94 ;
  assign n15335 = ~n15282 & ~n15334 ;
  assign n15336 = n15335 ^ n15334 ;
  assign n15337 = n15336 ^ n15282 ;
  assign n13292 = n13291 ^ n10640 ;
  assign n13258 = n13176 ^ n13175 ;
  assign n13261 = n13260 ^ n13221 ;
  assign n13262 = n13261 ^ n13219 ;
  assign n13259 = n13254 ^ n13235 ;
  assign n13263 = n13262 ^ n13259 ;
  assign n13264 = n13176 & n13263 ;
  assign n13265 = n13264 ^ n13262 ;
  assign n13266 = n13265 ^ n13241 ;
  assign n13267 = n13266 ^ n13251 ;
  assign n13268 = n13267 ^ n13223 ;
  assign n13269 = n13268 ^ n13265 ;
  assign n13270 = n13176 & n13269 ;
  assign n13271 = n13270 ^ n13266 ;
  assign n13272 = n13258 & ~n13271 ;
  assign n13273 = n13272 ^ n13265 ;
  assign n13257 = n13176 & n13225 ;
  assign n13274 = n13273 ^ n13257 ;
  assign n13286 = ~n13274 & ~n13285 ;
  assign n13287 = ~n13256 & n13286 ;
  assign n13293 = n13292 ^ n13287 ;
  assign n14442 = n13293 ^ x104 ;
  assign n14045 = n11515 & n11531 ;
  assign n14046 = n14045 ^ n11584 ;
  assign n14501 = n11259 & n11537 ;
  assign n14502 = n14501 ^ n11533 ;
  assign n14049 = n11100 ^ n11085 ;
  assign n14050 = n11259 ^ n11085 ;
  assign n14051 = n14050 ^ n11085 ;
  assign n14052 = n14049 & ~n14051 ;
  assign n14053 = n14052 ^ n11085 ;
  assign n14054 = ~n11513 & n14053 ;
  assign n14057 = n14056 ^ n14054 ;
  assign n14511 = n14502 ^ n14057 ;
  assign n14512 = n14511 ^ n14249 ;
  assign n14503 = n14502 ^ n11089 ;
  assign n14504 = n14503 ^ n11090 ;
  assign n14505 = n14504 ^ n14502 ;
  assign n14508 = ~n11259 & n14505 ;
  assign n14509 = n14508 ^ n14502 ;
  assign n14510 = ~n11513 & n14509 ;
  assign n14513 = n14512 ^ n14510 ;
  assign n14495 = n11590 ^ n11539 ;
  assign n14496 = n11539 ^ n11513 ;
  assign n14497 = n14496 ^ n11539 ;
  assign n14498 = n14495 & n14497 ;
  assign n14499 = n14498 ^ n11539 ;
  assign n14500 = n11259 & n14499 ;
  assign n14514 = n14513 ^ n14500 ;
  assign n14515 = ~n11548 & ~n14514 ;
  assign n14516 = ~n14224 & n14515 ;
  assign n14517 = ~n14046 & n14516 ;
  assign n14518 = n14517 ^ n11340 ;
  assign n14519 = n14518 ^ x99 ;
  assign n14520 = n13646 ^ x114 ;
  assign n14521 = n14519 & ~n14520 ;
  assign n14538 = n14521 ^ n14520 ;
  assign n14444 = n12358 ^ n12297 ;
  assign n14445 = n14444 ^ n12296 ;
  assign n14464 = n12300 & n12347 ;
  assign n14458 = n12349 ^ n12296 ;
  assign n14459 = n14458 ^ n12349 ;
  assign n14460 = n12350 & ~n14459 ;
  assign n14461 = n14460 ^ n12349 ;
  assign n14462 = n12297 & ~n14461 ;
  assign n14446 = n12297 ^ n12252 ;
  assign n14447 = n12327 ^ n12252 ;
  assign n14448 = n14447 ^ n12345 ;
  assign n14449 = n14448 ^ n14447 ;
  assign n14450 = n14447 ^ n12296 ;
  assign n14451 = n14450 ^ n14447 ;
  assign n14452 = n14449 & ~n14451 ;
  assign n14453 = n14452 ^ n14447 ;
  assign n14454 = ~n14446 & n14453 ;
  assign n14455 = n14454 ^ n12297 ;
  assign n14463 = n14462 ^ n14455 ;
  assign n14465 = n14464 ^ n14463 ;
  assign n14466 = ~n14445 & n14465 ;
  assign n14467 = n14466 ^ n14465 ;
  assign n14469 = n14467 ^ n12315 ;
  assign n14470 = n14469 ^ n14467 ;
  assign n14471 = n14467 ^ n12297 ;
  assign n14472 = n14471 ^ n14467 ;
  assign n14473 = n14470 & ~n14472 ;
  assign n14474 = n14466 & n14473 ;
  assign n14475 = n14474 ^ n14466 ;
  assign n14476 = n14475 ^ n14465 ;
  assign n14477 = ~n12313 & n14476 ;
  assign n14478 = n14477 ^ n14465 ;
  assign n14479 = n12296 & n14478 ;
  assign n14480 = n12334 ^ n12297 ;
  assign n14481 = n14480 ^ n12334 ;
  assign n14482 = n12334 ^ n12309 ;
  assign n14483 = n14482 ^ n12334 ;
  assign n14484 = ~n14481 & n14483 ;
  assign n14485 = n14484 ^ n12334 ;
  assign n14486 = n14479 & n14485 ;
  assign n14487 = n14486 ^ n14478 ;
  assign n14488 = ~n12333 & n14487 ;
  assign n14489 = ~n13753 & n14488 ;
  assign n14490 = ~n12302 & n14489 ;
  assign n14491 = n14490 ^ n11421 ;
  assign n14492 = n14491 ^ x89 ;
  assign n13149 = ~n11757 & n11990 ;
  assign n13150 = n13149 ^ n11991 ;
  assign n13159 = n11982 ^ n11964 ;
  assign n13160 = n11723 & n13159 ;
  assign n13161 = n13160 ^ n11979 ;
  assign n13152 = n13149 ^ n12011 ;
  assign n13153 = n13152 ^ n11976 ;
  assign n13154 = ~n11656 & ~n13153 ;
  assign n13155 = n13154 ^ n11976 ;
  assign n13162 = n13161 ^ n13155 ;
  assign n13151 = n12001 ^ n11723 ;
  assign n13156 = n13155 ^ n13151 ;
  assign n13163 = n13162 ^ n13156 ;
  assign n13164 = n11656 & n13163 ;
  assign n13165 = n13164 ^ n13156 ;
  assign n13166 = ~n11689 & ~n13165 ;
  assign n13167 = n13166 ^ n13155 ;
  assign n13168 = ~n13150 & ~n13167 ;
  assign n13169 = n13168 ^ n10541 ;
  assign n14493 = n13169 ^ x80 ;
  assign n14494 = n14492 & n14493 ;
  assign n14553 = n14494 ^ n14492 ;
  assign n14554 = n14553 ^ n14493 ;
  assign n14556 = ~n14538 & ~n14554 ;
  assign n14524 = n14494 & n14521 ;
  assign n15173 = n14556 ^ n14524 ;
  assign n14441 = n13746 ^ x82 ;
  assign n15174 = n14524 ^ n14441 ;
  assign n15175 = n15174 ^ n14524 ;
  assign n15176 = n15173 & ~n15175 ;
  assign n15177 = n15176 ^ n14524 ;
  assign n15178 = ~n14442 & n15177 ;
  assign n14539 = n14538 ^ n14519 ;
  assign n14564 = n14494 & n14539 ;
  assign n15160 = n14564 ^ n14553 ;
  assign n14571 = n14539 & n14553 ;
  assign n14561 = n14521 & n14553 ;
  assign n14572 = n14571 ^ n14561 ;
  assign n14555 = n14521 & ~n14554 ;
  assign n14584 = n14572 ^ n14555 ;
  assign n14558 = n14539 & ~n14554 ;
  assign n14559 = n14558 ^ n14554 ;
  assign n14557 = n14556 ^ n14555 ;
  assign n14560 = n14559 ^ n14557 ;
  assign n15159 = n14584 ^ n14560 ;
  assign n15161 = n15160 ^ n15159 ;
  assign n15162 = n15161 ^ n14584 ;
  assign n15163 = ~n14441 & ~n15162 ;
  assign n15164 = n15163 ^ n15159 ;
  assign n15179 = n15178 ^ n15164 ;
  assign n14522 = n14521 ^ n14519 ;
  assign n14527 = n14494 ^ n14493 ;
  assign n14528 = n14522 & n14527 ;
  assign n14523 = n14494 & n14522 ;
  assign n14526 = n14523 ^ n14494 ;
  assign n14529 = n14528 ^ n14526 ;
  assign n14575 = n14529 ^ n14493 ;
  assign n14540 = n14527 & n14539 ;
  assign n14537 = n14521 & n14527 ;
  assign n14541 = n14540 ^ n14537 ;
  assign n14542 = n14541 ^ n14523 ;
  assign n14576 = n14575 ^ n14542 ;
  assign n14603 = n14576 ^ n14523 ;
  assign n15155 = n14603 ^ n14528 ;
  assign n15166 = n15164 ^ n15155 ;
  assign n14562 = n14561 ^ n14560 ;
  assign n14563 = n14562 ^ n14558 ;
  assign n15165 = n15164 ^ n14563 ;
  assign n15167 = n15166 ^ n15165 ;
  assign n15170 = ~n14441 & ~n15167 ;
  assign n15171 = n15170 ^ n15166 ;
  assign n15172 = ~n14442 & ~n15171 ;
  assign n15180 = n15179 ^ n15172 ;
  assign n14443 = n14442 ^ n14441 ;
  assign n15157 = n14564 ^ n14537 ;
  assign n15158 = ~n14443 & n15157 ;
  assign n15181 = n15180 ^ n15158 ;
  assign n14551 = n14441 & ~n14442 ;
  assign n14552 = n14551 ^ n14441 ;
  assign n14599 = n14552 ^ n14442 ;
  assign n15156 = n14599 & n15155 ;
  assign n15182 = n15181 ^ n15156 ;
  assign n14565 = n14564 ^ n14524 ;
  assign n14566 = n14565 ^ n14526 ;
  assign n15190 = n14566 ^ n14558 ;
  assign n15191 = n15190 ^ n14555 ;
  assign n14577 = n14576 ^ n14538 ;
  assign n14574 = n14566 ^ n14556 ;
  assign n14578 = n14577 ^ n14574 ;
  assign n14585 = n14578 ^ n14560 ;
  assign n15192 = n15191 ^ n14585 ;
  assign n15193 = ~n14442 & n15192 ;
  assign n15194 = n15193 ^ n14566 ;
  assign n15195 = n14441 & n15194 ;
  assign n15196 = n15195 ^ n14540 ;
  assign n14525 = n14524 ^ n14523 ;
  assign n15183 = n14540 ^ n14525 ;
  assign n15184 = n15183 ^ n14540 ;
  assign n15185 = n14540 ^ n14441 ;
  assign n15186 = n15185 ^ n14540 ;
  assign n15187 = n15184 & ~n15186 ;
  assign n15188 = n15187 ^ n14540 ;
  assign n15189 = ~n14442 & n15188 ;
  assign n15197 = n15196 ^ n15189 ;
  assign n15198 = n15182 & ~n15197 ;
  assign n15199 = n15198 ^ n12504 ;
  assign n15200 = n15199 ^ x75 ;
  assign n14222 = n13784 ^ x97 ;
  assign n14290 = n12909 ^ n12880 ;
  assign n14291 = n12755 & n14290 ;
  assign n14278 = n12905 ^ n12861 ;
  assign n14287 = n14278 ^ n12845 ;
  assign n14288 = ~n12752 & n14287 ;
  assign n14279 = n14278 ^ n12857 ;
  assign n14280 = n14279 ^ n12863 ;
  assign n14281 = n14280 ^ n12880 ;
  assign n14282 = n14281 ^ n14278 ;
  assign n14283 = ~n12750 & n14282 ;
  assign n14284 = n14283 ^ n14279 ;
  assign n14285 = n12751 & n14284 ;
  assign n14286 = n14285 ^ n12845 ;
  assign n14289 = n14288 ^ n14286 ;
  assign n14292 = n14291 ^ n14289 ;
  assign n14091 = n12751 ^ n12750 ;
  assign n14080 = n12859 ^ n12853 ;
  assign n14271 = n14080 ^ n12906 ;
  assign n14272 = n14271 ^ n14080 ;
  assign n14273 = n14080 ^ n12751 ;
  assign n14274 = n14273 ^ n14080 ;
  assign n14275 = n14272 & ~n14274 ;
  assign n14276 = n14275 ^ n14080 ;
  assign n14277 = n14091 & n14276 ;
  assign n14293 = n14292 ^ n14277 ;
  assign n14294 = n14293 ^ n13615 ;
  assign n14295 = n14294 ^ n12895 ;
  assign n14089 = ~n12753 & n12865 ;
  assign n14090 = n14089 ^ n12888 ;
  assign n14296 = n14295 ^ n14090 ;
  assign n14297 = n14296 ^ n12921 ;
  assign n14298 = n14297 ^ n10113 ;
  assign n14299 = n14298 ^ x90 ;
  assign n14324 = n14323 ^ x73 ;
  assign n14325 = ~n14299 & ~n14324 ;
  assign n14326 = n14325 ^ n14324 ;
  assign n14327 = n14326 ^ n14299 ;
  assign n14258 = n13678 ^ x64 ;
  assign n14261 = n13161 ^ n11976 ;
  assign n14262 = ~n11689 & ~n14261 ;
  assign n14263 = n14262 ^ n11976 ;
  assign n14267 = n14263 ^ n10084 ;
  assign n14264 = n14263 ^ n12012 ;
  assign n14259 = n13152 ^ n13151 ;
  assign n14260 = ~n11689 & n14259 ;
  assign n14265 = n14264 ^ n14260 ;
  assign n14266 = n11656 & n14265 ;
  assign n14268 = n14267 ^ n14266 ;
  assign n14269 = n14268 ^ x120 ;
  assign n14270 = ~n14258 & n14269 ;
  assign n14329 = n14270 ^ n14269 ;
  assign n14330 = n14329 ^ n14258 ;
  assign n14348 = ~n14327 & n14330 ;
  assign n14331 = n14330 ^ n14269 ;
  assign n14336 = n14325 ^ n14299 ;
  assign n14344 = ~n14331 & ~n14336 ;
  assign n14339 = n14270 & n14325 ;
  assign n14345 = n14344 ^ n14339 ;
  assign n14328 = n14270 & ~n14327 ;
  assign n14340 = n14339 ^ n14328 ;
  assign n14337 = n14270 & ~n14336 ;
  assign n14338 = n14337 ^ n14270 ;
  assign n14341 = n14340 ^ n14338 ;
  assign n14335 = n14325 & ~n14331 ;
  assign n14342 = n14341 ^ n14335 ;
  assign n14343 = n14342 ^ n14337 ;
  assign n14346 = n14345 ^ n14343 ;
  assign n14332 = ~n14326 & ~n14331 ;
  assign n14333 = n14332 ^ n14328 ;
  assign n14334 = n14333 ^ n14258 ;
  assign n14347 = n14346 ^ n14334 ;
  assign n14349 = n14348 ^ n14347 ;
  assign n14256 = n14255 ^ x123 ;
  assign n14403 = n14348 ^ n14256 ;
  assign n14404 = n14403 ^ n14348 ;
  assign n14405 = ~n14349 & ~n14404 ;
  assign n14406 = n14405 ^ n14348 ;
  assign n14407 = ~n14222 & n14406 ;
  assign n14257 = n14256 ^ n14222 ;
  assign n15241 = n14222 & n14345 ;
  assign n14363 = ~n14326 & n14329 ;
  assign n14368 = n14363 ^ n14341 ;
  assign n14369 = n14368 ^ n14326 ;
  assign n14370 = n14369 ^ n14332 ;
  assign n14371 = n14370 ^ n14348 ;
  assign n14366 = n14330 & ~n14336 ;
  assign n14367 = n14366 ^ n14330 ;
  assign n14372 = n14371 ^ n14367 ;
  assign n14373 = n14372 ^ n14339 ;
  assign n14365 = n14335 ^ n14325 ;
  assign n14374 = n14373 ^ n14365 ;
  assign n15239 = n14374 ^ n14345 ;
  assign n15201 = n14363 ^ n14345 ;
  assign n15202 = ~n14222 & n15201 ;
  assign n15203 = n15202 ^ n14363 ;
  assign n15240 = n15239 ^ n15203 ;
  assign n15242 = n15241 ^ n15240 ;
  assign n15243 = n14257 & ~n15242 ;
  assign n15244 = n15243 ^ n14374 ;
  assign n14358 = n14222 & n14256 ;
  assign n14359 = n14347 ^ n14344 ;
  assign n14360 = n14358 & ~n14359 ;
  assign n15245 = n15244 ^ n14360 ;
  assign n15204 = n14256 & n15203 ;
  assign n14350 = n14328 ^ n14327 ;
  assign n14351 = n14350 ^ n14349 ;
  assign n15231 = n14366 ^ n14351 ;
  assign n15230 = n14345 ^ n14328 ;
  assign n15232 = n15231 ^ n15230 ;
  assign n14380 = n14374 ^ n14370 ;
  assign n15233 = n15232 ^ n14380 ;
  assign n15234 = ~n14222 & n15233 ;
  assign n15235 = n15234 ^ n14380 ;
  assign n15236 = ~n14256 & n15235 ;
  assign n14375 = n14374 ^ n14351 ;
  assign n14364 = n14363 ^ n14329 ;
  assign n14376 = n14375 ^ n14364 ;
  assign n15228 = n14257 & ~n14376 ;
  assign n15223 = n14374 ^ n14333 ;
  assign n15224 = n14256 & ~n15223 ;
  assign n15217 = n14337 ^ n14333 ;
  assign n15212 = n14376 ^ n14348 ;
  assign n15213 = n15212 ^ n14341 ;
  assign n15214 = n15213 ^ n14372 ;
  assign n15207 = n14363 ^ n14256 ;
  assign n15208 = n15207 ^ n14363 ;
  assign n15209 = n14368 & ~n15208 ;
  assign n15210 = n15209 ^ n14363 ;
  assign n15211 = ~n14222 & n15210 ;
  assign n15215 = n15214 ^ n15211 ;
  assign n15216 = n15215 ^ n14366 ;
  assign n15218 = n15217 ^ n15216 ;
  assign n15219 = n15218 ^ n15211 ;
  assign n15220 = ~n14256 & n15219 ;
  assign n15221 = n15220 ^ n15215 ;
  assign n15222 = n15221 ^ n15211 ;
  assign n15225 = n15224 ^ n15222 ;
  assign n15226 = ~n14222 & n15225 ;
  assign n15227 = n15226 ^ n15221 ;
  assign n15229 = n15228 ^ n15227 ;
  assign n15237 = n15236 ^ n15229 ;
  assign n15238 = ~n15204 & ~n15237 ;
  assign n15246 = n15245 ^ n15238 ;
  assign n15247 = ~n14407 & ~n15246 ;
  assign n15248 = n15247 ^ n12454 ;
  assign n15249 = n15248 ^ x93 ;
  assign n15250 = n15200 & ~n15249 ;
  assign n15341 = n15250 ^ n15249 ;
  assign n15356 = ~n15337 & ~n15341 ;
  assign n16636 = n15153 & n15356 ;
  assign n15349 = n15250 & ~n15337 ;
  assign n15408 = n15349 ^ n15337 ;
  assign n15346 = n15250 ^ n15200 ;
  assign n15379 = ~n15337 & n15346 ;
  assign n15393 = n15379 ^ n15356 ;
  assign n15409 = n15408 ^ n15393 ;
  assign n15338 = n15337 ^ n15334 ;
  assign n15390 = ~n15338 & ~n15341 ;
  assign n15410 = n15409 ^ n15390 ;
  assign n16627 = n15410 ^ n15349 ;
  assign n15375 = n15250 & ~n15336 ;
  assign n15347 = n15346 ^ n15249 ;
  assign n15348 = ~n15336 & n15347 ;
  assign n15383 = n15375 ^ n15348 ;
  assign n15365 = ~n15336 & n15346 ;
  assign n15382 = n15365 ^ n15336 ;
  assign n15384 = n15383 ^ n15382 ;
  assign n15366 = n15250 & n15335 ;
  assign n15367 = n15366 ^ n15365 ;
  assign n15385 = n15384 ^ n15367 ;
  assign n15342 = n15335 & ~n15341 ;
  assign n15381 = n15367 ^ n15342 ;
  assign n15386 = n15385 ^ n15381 ;
  assign n16629 = n16627 ^ n15386 ;
  assign n15374 = n15335 & n15346 ;
  assign n15376 = n15375 ^ n15374 ;
  assign n16630 = n16629 ^ n15376 ;
  assign n16631 = n15132 & n16630 ;
  assign n16618 = n15366 ^ n15336 ;
  assign n16619 = n16618 ^ n15342 ;
  assign n15364 = n15335 & n15347 ;
  assign n16620 = n16619 ^ n15364 ;
  assign n16621 = n15132 & ~n16620 ;
  assign n16622 = n16621 ^ n15385 ;
  assign n16628 = n16627 ^ n16622 ;
  assign n16632 = n16631 ^ n16628 ;
  assign n16633 = n15152 & n16632 ;
  assign n15355 = ~n15338 & n15346 ;
  assign n16607 = n15409 ^ n15355 ;
  assign n15406 = ~n15338 & n15347 ;
  assign n16616 = n16607 ^ n15406 ;
  assign n15154 = n15153 ^ n15152 ;
  assign n15343 = n15154 ^ n15132 ;
  assign n15344 = n15342 & ~n15343 ;
  assign n15339 = n15250 & ~n15338 ;
  assign n15340 = n15154 & n15339 ;
  assign n15345 = n15344 ^ n15340 ;
  assign n16617 = n16616 ^ n15345 ;
  assign n16623 = n16622 ^ n16617 ;
  assign n16624 = n16623 ^ n13746 ;
  assign n16608 = n16607 ^ n15339 ;
  assign n15357 = n15356 ^ n15355 ;
  assign n16609 = n16608 ^ n15357 ;
  assign n16610 = n16609 ^ n16607 ;
  assign n16611 = n16607 ^ n15152 ;
  assign n16612 = n16611 ^ n16607 ;
  assign n16613 = n16610 & ~n16612 ;
  assign n16614 = n16613 ^ n16607 ;
  assign n16615 = ~n15132 & ~n16614 ;
  assign n16625 = n16624 ^ n16615 ;
  assign n16599 = n15152 ^ n15132 ;
  assign n16600 = n15406 ^ n15152 ;
  assign n16601 = n16600 ^ n15406 ;
  assign n15392 = n15379 ^ n15339 ;
  assign n16602 = n15406 ^ n15392 ;
  assign n16603 = n16602 ^ n15406 ;
  assign n16604 = ~n16601 & n16603 ;
  assign n16605 = n16604 ^ n15406 ;
  assign n16606 = n16599 & n16605 ;
  assign n16626 = n16625 ^ n16606 ;
  assign n16634 = n16633 ^ n16626 ;
  assign n16596 = n15384 ^ n15366 ;
  assign n16595 = n15365 ^ n15364 ;
  assign n16597 = n16596 ^ n16595 ;
  assign n16598 = n15154 & ~n16597 ;
  assign n16635 = n16634 ^ n16598 ;
  assign n16637 = n16636 ^ n16635 ;
  assign n16638 = n16637 ^ x115 ;
  assign n15420 = n15333 ^ x69 ;
  assign n15456 = n15241 ^ n14343 ;
  assign n15457 = ~n14257 & n15456 ;
  assign n15451 = n14371 ^ n14345 ;
  assign n15440 = n14347 ^ n14333 ;
  assign n15441 = n14256 & ~n15440 ;
  assign n15442 = n15441 ^ n14333 ;
  assign n15452 = n15451 ^ n15442 ;
  assign n14392 = n14380 ^ n14351 ;
  assign n14393 = n14392 ^ n14371 ;
  assign n15450 = n14256 & ~n14393 ;
  assign n15453 = n15452 ^ n15450 ;
  assign n15454 = ~n14222 & ~n15453 ;
  assign n15446 = ~n14257 & n14366 ;
  assign n15447 = n15446 ^ n15204 ;
  assign n15448 = n15447 ^ n12783 ;
  assign n15443 = n15442 ^ n14345 ;
  assign n15444 = n15443 ^ n14407 ;
  assign n15432 = n14351 ^ n14222 ;
  assign n15445 = n15444 ^ n15432 ;
  assign n15449 = n15448 ^ n15445 ;
  assign n15455 = n15454 ^ n15449 ;
  assign n15458 = n15457 ^ n15455 ;
  assign n15437 = n14358 ^ n14222 ;
  assign n15438 = n14374 ^ n14366 ;
  assign n15439 = n15437 & ~n15438 ;
  assign n15459 = n15458 ^ n15439 ;
  assign n14377 = n14376 ^ n14370 ;
  assign n15433 = n15432 ^ n14351 ;
  assign n15434 = n14377 & n15433 ;
  assign n15435 = n15434 ^ n14351 ;
  assign n15436 = n14256 & ~n15435 ;
  assign n15460 = n15459 ^ n15436 ;
  assign n15421 = n14358 ^ n14257 ;
  assign n15422 = n15421 ^ n14256 ;
  assign n15423 = n15422 ^ n14257 ;
  assign n15424 = n14341 ^ n14256 ;
  assign n15427 = n15423 & ~n15424 ;
  assign n15428 = n15427 ^ n14257 ;
  assign n15429 = n14372 & n15428 ;
  assign n15461 = n15460 ^ n15429 ;
  assign n15462 = n15461 ^ x78 ;
  assign n15463 = ~n15420 & ~n15462 ;
  assign n15464 = n15463 ^ n15420 ;
  assign n14115 = n12880 ^ n12847 ;
  assign n14103 = ~n12751 & n12842 ;
  assign n14116 = n14115 ^ n14103 ;
  assign n14112 = n12875 ^ n12847 ;
  assign n14113 = n14112 ^ n12905 ;
  assign n14114 = ~n12751 & n14113 ;
  assign n14117 = n14116 ^ n14114 ;
  assign n14118 = n12750 & n14117 ;
  assign n14108 = n12871 ^ n12866 ;
  assign n14109 = n12754 & n14108 ;
  assign n14092 = n12921 ^ n12863 ;
  assign n14093 = n14092 ^ n12921 ;
  assign n14094 = n14093 ^ n12751 ;
  assign n14095 = n14094 ^ n14093 ;
  assign n14096 = n14093 ^ n12854 ;
  assign n14097 = n14096 ^ n14093 ;
  assign n14098 = ~n14095 & n14097 ;
  assign n14099 = n14098 ^ n14093 ;
  assign n14100 = n14091 & n14099 ;
  assign n14101 = n14100 ^ n14092 ;
  assign n14102 = n14101 ^ n12887 ;
  assign n14104 = n14103 ^ n14102 ;
  assign n14105 = n14104 ^ n14090 ;
  assign n14106 = n14105 ^ n10886 ;
  assign n14082 = n12887 ^ n12751 ;
  assign n14083 = n14082 ^ n12887 ;
  assign n14086 = n12920 & ~n14083 ;
  assign n14087 = n14086 ^ n12887 ;
  assign n14088 = ~n12750 & ~n14087 ;
  assign n14107 = n14106 ^ n14088 ;
  assign n14110 = n14109 ^ n14107 ;
  assign n14081 = ~n12751 & n14080 ;
  assign n14111 = n14110 ^ n14081 ;
  assign n14119 = n14118 ^ n14111 ;
  assign n14120 = n14119 ^ x83 ;
  assign n14124 = n14123 ^ x70 ;
  assign n14125 = ~n14120 & n14124 ;
  assign n14126 = n14125 ^ n14124 ;
  assign n14127 = n14126 ^ n14120 ;
  assign n14044 = n14043 ^ x93 ;
  assign n14071 = n11098 & n11549 ;
  assign n14064 = n11518 ^ n11092 ;
  assign n14065 = n14064 ^ n11552 ;
  assign n14066 = n14065 ^ n11567 ;
  assign n14067 = n11513 & n14066 ;
  assign n14059 = n11586 ^ n11096 ;
  assign n14060 = n14059 ^ n11590 ;
  assign n14058 = n11518 & n11549 ;
  assign n14061 = n14060 ^ n14058 ;
  assign n14063 = n14061 ^ n11541 ;
  assign n14068 = n14067 ^ n14063 ;
  assign n14069 = n11259 & n14068 ;
  assign n14062 = n14061 ^ n14057 ;
  assign n14070 = n14069 ^ n14062 ;
  assign n14072 = n14071 ^ n14070 ;
  assign n14073 = ~n11562 & ~n14072 ;
  assign n14074 = ~n14048 & n14073 ;
  assign n14075 = ~n11580 & n14074 ;
  assign n14076 = ~n14046 & n14075 ;
  assign n14077 = n14076 ^ n10958 ;
  assign n14078 = n14077 ^ x100 ;
  assign n14079 = n14044 & n14078 ;
  assign n14132 = n14079 ^ n14044 ;
  assign n14133 = n14132 ^ n14078 ;
  assign n14139 = n14133 ^ n14044 ;
  assign n14140 = n14127 & n14139 ;
  assign n13975 = n13974 ^ x118 ;
  assign n14010 = n14009 ^ x69 ;
  assign n14190 = ~n13975 & n14010 ;
  assign n14191 = n14190 ^ n14010 ;
  assign n14192 = n14191 ^ n13975 ;
  assign n14193 = n14192 ^ n14010 ;
  assign n15497 = n14140 & ~n14193 ;
  assign n14160 = n14044 & n14120 ;
  assign n14147 = n14079 & n14127 ;
  assign n14138 = n14126 & n14132 ;
  assign n14157 = n14147 ^ n14138 ;
  assign n14148 = n14147 ^ n14127 ;
  assign n14143 = n14125 & ~n14133 ;
  assign n14128 = n14127 ^ n14124 ;
  assign n14134 = ~n14128 & ~n14133 ;
  assign n14144 = n14143 ^ n14134 ;
  assign n14130 = ~n14044 & n14126 ;
  assign n14131 = n14078 & n14130 ;
  assign n14141 = n14131 ^ n14130 ;
  assign n14142 = n14141 ^ n14133 ;
  assign n14145 = n14144 ^ n14142 ;
  assign n14146 = n14145 ^ n14140 ;
  assign n14149 = n14148 ^ n14146 ;
  assign n14158 = n14157 ^ n14149 ;
  assign n14161 = n14160 ^ n14158 ;
  assign n14129 = n14079 & ~n14128 ;
  assign n14162 = n14161 ^ n14129 ;
  assign n14150 = n14125 & n14132 ;
  assign n14135 = n14134 ^ n14131 ;
  assign n14136 = n14135 ^ n14129 ;
  assign n14151 = n14150 ^ n14136 ;
  assign n14152 = n14151 ^ n14149 ;
  assign n14153 = n14152 ^ n14138 ;
  assign n14137 = n14136 ^ n14132 ;
  assign n14154 = n14153 ^ n14137 ;
  assign n14155 = n14154 ^ n14150 ;
  assign n14163 = n14162 ^ n14155 ;
  assign n14159 = n14158 ^ n14044 ;
  assign n14164 = n14163 ^ n14159 ;
  assign n14165 = n14164 ^ n14154 ;
  assign n14167 = n14165 ^ n14150 ;
  assign n14168 = n14167 ^ n14143 ;
  assign n14169 = n14168 ^ n14125 ;
  assign n14170 = n14169 ^ n14154 ;
  assign n14171 = n14170 ^ n14144 ;
  assign n14172 = n14171 ^ n14154 ;
  assign n14166 = n14165 ^ n14129 ;
  assign n14173 = n14172 ^ n14166 ;
  assign n14156 = n14155 ^ n14120 ;
  assign n14174 = n14173 ^ n14156 ;
  assign n15495 = ~n13975 & n14174 ;
  assign n15467 = n14167 ^ n14147 ;
  assign n15466 = n14140 ^ n14127 ;
  assign n15468 = n15467 ^ n15466 ;
  assign n14195 = n14143 ^ n14131 ;
  assign n15469 = n15468 ^ n14195 ;
  assign n15470 = n14010 & n15469 ;
  assign n15465 = n14146 ^ n14127 ;
  assign n15471 = n15470 ^ n15465 ;
  assign n14011 = n14010 ^ n13975 ;
  assign n14175 = n14174 ^ n14149 ;
  assign n14176 = n14010 & ~n14175 ;
  assign n14177 = n14176 ^ n14149 ;
  assign n14178 = ~n14011 & ~n14177 ;
  assign n15493 = n15471 ^ n14178 ;
  assign n14210 = n14144 ^ n14141 ;
  assign n14211 = n14210 ^ n14133 ;
  assign n14212 = n14211 ^ n14141 ;
  assign n14213 = n14141 ^ n13975 ;
  assign n14214 = n14213 ^ n14141 ;
  assign n14215 = ~n14212 & n14214 ;
  assign n14216 = n14215 ^ n14141 ;
  assign n14217 = ~n14010 & n14216 ;
  assign n15494 = n15493 ^ n14217 ;
  assign n15496 = n15495 ^ n15494 ;
  assign n15498 = n15497 ^ n15496 ;
  assign n15487 = n14170 ^ n14162 ;
  assign n15488 = n14162 ^ n14010 ;
  assign n15489 = n15488 ^ n14162 ;
  assign n15490 = n15487 & n15489 ;
  assign n15491 = n15490 ^ n14162 ;
  assign n15492 = n13975 & ~n15491 ;
  assign n15499 = n15498 ^ n15492 ;
  assign n15500 = n15499 ^ n12749 ;
  assign n14198 = n14164 ^ n14158 ;
  assign n15480 = n14198 ^ n14135 ;
  assign n15479 = n14144 ^ n14138 ;
  assign n15481 = n15480 ^ n15479 ;
  assign n15482 = n15479 ^ n14010 ;
  assign n15483 = n15482 ^ n15479 ;
  assign n15484 = n15481 & n15483 ;
  assign n15485 = n15484 ^ n15479 ;
  assign n15486 = n13975 & n15485 ;
  assign n15501 = n15500 ^ n15486 ;
  assign n15472 = n15471 ^ n14168 ;
  assign n15473 = n15472 ^ n15471 ;
  assign n15474 = n15471 ^ n13975 ;
  assign n15475 = n15474 ^ n15471 ;
  assign n15476 = n15473 & ~n15475 ;
  assign n15477 = n15476 ^ n15471 ;
  assign n15478 = ~n14011 & ~n15477 ;
  assign n15502 = n15501 ^ n15478 ;
  assign n15503 = n15502 ^ x101 ;
  assign n15504 = n15131 ^ x91 ;
  assign n13148 = n11604 ^ x78 ;
  assign n13170 = n13169 ^ x92 ;
  assign n13171 = n13148 & n13170 ;
  assign n13172 = n13171 ^ n13170 ;
  assign n13294 = n13293 ^ x116 ;
  assign n13320 = n13023 ^ n10602 ;
  assign n13310 = ~n12925 & n13019 ;
  assign n13311 = n13310 ^ n13013 ;
  assign n13321 = n13320 ^ n13311 ;
  assign n13305 = n13034 ^ n13021 ;
  assign n13306 = n13002 & n13305 ;
  assign n13299 = n13298 ^ n12990 ;
  assign n13300 = n13007 & n13299 ;
  assign n13302 = n13301 ^ n12981 ;
  assign n13303 = n13300 & ~n13302 ;
  assign n13304 = n13303 ^ n13299 ;
  assign n13307 = n13306 ^ n13304 ;
  assign n13322 = n13321 ^ n13307 ;
  assign n13313 = n13311 ^ n12987 ;
  assign n13312 = n13311 ^ n13041 ;
  assign n13314 = n13313 ^ n13312 ;
  assign n13317 = n12925 & ~n13314 ;
  assign n13318 = n13317 ^ n13313 ;
  assign n13319 = n13002 & n13318 ;
  assign n13323 = n13322 ^ n13319 ;
  assign n13295 = n12999 ^ n12995 ;
  assign n13308 = n12925 & ~n13307 ;
  assign n13309 = ~n13295 & n13308 ;
  assign n13324 = n13323 ^ n13309 ;
  assign n13325 = n13324 ^ x109 ;
  assign n13326 = n13294 & n13325 ;
  assign n13328 = n12923 ^ x110 ;
  assign n13489 = n13488 ^ n13433 ;
  assign n13498 = n13497 ^ n13489 ;
  assign n13499 = n13498 ^ n13483 ;
  assign n13484 = n13449 ^ n13436 ;
  assign n13485 = n13484 ^ n13425 ;
  assign n13486 = n13329 & n13485 ;
  assign n13500 = n13499 ^ n13486 ;
  assign n13517 = n13516 ^ n13500 ;
  assign n13501 = n13500 ^ n13497 ;
  assign n13502 = n13501 ^ n13483 ;
  assign n13469 = ~n13329 & n13450 ;
  assign n13503 = n13502 ^ n13469 ;
  assign n13504 = ~n13458 & n13503 ;
  assign n13518 = n13517 ^ n13504 ;
  assign n13467 = n13438 ^ n13433 ;
  assign n13468 = n13466 & n13467 ;
  assign n13519 = n13518 ^ n13468 ;
  assign n13461 = n13446 ^ n13330 ;
  assign n13462 = n13461 ^ n13446 ;
  assign n13463 = n13448 & ~n13462 ;
  assign n13464 = n13463 ^ n13446 ;
  assign n13465 = n13458 & n13464 ;
  assign n13520 = n13519 ^ n13465 ;
  assign n13528 = n13527 ^ n13520 ;
  assign n13529 = n13528 ^ n10699 ;
  assign n13457 = ~n13332 & ~n13456 ;
  assign n13530 = n13529 ^ n13457 ;
  assign n13531 = n13530 ^ x91 ;
  assign n13532 = n13328 & ~n13531 ;
  assign n13537 = n13532 ^ n13328 ;
  assign n13539 = n13326 & n13537 ;
  assign n13538 = n13325 & n13537 ;
  assign n13540 = n13539 ^ n13538 ;
  assign n13327 = n13326 ^ n13294 ;
  assign n13536 = n13327 & n13532 ;
  assign n13541 = n13540 ^ n13536 ;
  assign n14660 = n13172 & n13541 ;
  assign n13173 = n13172 ^ n13148 ;
  assign n13174 = n13173 ^ n13170 ;
  assign n13533 = n13532 ^ n13531 ;
  assign n13562 = n13326 ^ n13325 ;
  assign n13563 = ~n13533 & n13562 ;
  assign n13534 = n13327 & ~n13533 ;
  assign n13564 = n13563 ^ n13534 ;
  assign n13542 = n13327 ^ n13325 ;
  assign n13543 = n13537 & ~n13542 ;
  assign n13555 = n13543 ^ n13539 ;
  assign n13554 = n13326 & ~n13533 ;
  assign n13556 = n13555 ^ n13554 ;
  assign n13551 = n13326 & n13532 ;
  assign n13552 = n13551 ^ n13543 ;
  assign n13553 = n13552 ^ n13326 ;
  assign n13557 = n13556 ^ n13553 ;
  assign n13549 = n13537 ^ n13531 ;
  assign n13550 = ~n13542 & n13549 ;
  assign n13558 = n13557 ^ n13550 ;
  assign n13544 = n13543 ^ n13537 ;
  assign n13545 = n13544 ^ n13538 ;
  assign n13546 = n13545 ^ n13541 ;
  assign n13547 = n13546 ^ n13540 ;
  assign n13535 = n13534 ^ n13327 ;
  assign n13548 = n13547 ^ n13535 ;
  assign n13559 = n13558 ^ n13548 ;
  assign n13561 = n13559 ^ n13549 ;
  assign n13565 = n13564 ^ n13561 ;
  assign n13566 = n13565 ^ n13554 ;
  assign n13560 = n13559 ^ n13328 ;
  assign n13567 = n13566 ^ n13560 ;
  assign n13568 = n13174 & ~n13567 ;
  assign n14661 = n14660 ^ n13568 ;
  assign n13595 = n13170 ^ n13148 ;
  assign n14636 = n13567 ^ n13561 ;
  assign n14637 = n14636 ^ n13554 ;
  assign n15524 = n14637 ^ n13534 ;
  assign n15525 = n13171 & ~n15524 ;
  assign n14666 = n13536 ^ n13532 ;
  assign n13569 = n13325 ^ n13294 ;
  assign n13570 = ~n13328 & n13569 ;
  assign n13571 = n13570 ^ n13294 ;
  assign n13582 = n13571 ^ n13325 ;
  assign n13583 = n13582 ^ n13546 ;
  assign n14630 = n13583 ^ n13551 ;
  assign n14667 = n14666 ^ n14630 ;
  assign n15514 = n13174 & n14667 ;
  assign n15513 = n14667 ^ n13174 ;
  assign n15515 = n15514 ^ n15513 ;
  assign n15516 = n13546 ^ n13173 ;
  assign n15517 = n15516 ^ n13555 ;
  assign n15518 = n15515 & ~n15517 ;
  assign n15519 = n15518 ^ n13555 ;
  assign n15520 = n15519 ^ n13551 ;
  assign n13584 = n13583 ^ n13545 ;
  assign n15511 = n13584 ^ n13551 ;
  assign n15512 = n13170 & n15511 ;
  assign n15521 = n15520 ^ n15512 ;
  assign n15509 = n13584 ^ n13555 ;
  assign n15510 = ~n13148 & n15509 ;
  assign n15522 = n15521 ^ n15510 ;
  assign n15508 = n13172 & n13566 ;
  assign n15523 = n15522 ^ n15508 ;
  assign n15526 = n15525 ^ n15523 ;
  assign n15527 = n13566 ^ n13328 ;
  assign n15528 = n15527 ^ n13558 ;
  assign n15529 = n13558 ^ n13148 ;
  assign n15530 = n15529 ^ n13558 ;
  assign n15531 = ~n15528 & ~n15530 ;
  assign n15532 = n15531 ^ n13558 ;
  assign n15533 = ~n13170 & n15532 ;
  assign n15534 = ~n15526 & ~n15533 ;
  assign n15535 = n13595 & n15534 ;
  assign n15536 = n13554 ^ n13148 ;
  assign n15537 = n15536 ^ n13554 ;
  assign n15538 = n13556 & ~n15537 ;
  assign n15539 = n15538 ^ n13554 ;
  assign n15540 = n15535 & n15539 ;
  assign n15541 = n15540 ^ n15534 ;
  assign n15542 = ~n14661 & n15541 ;
  assign n15543 = n15542 ^ n13205 ;
  assign n15544 = n15543 ^ x108 ;
  assign n15563 = n15544 ^ n15504 ;
  assign n15564 = ~n15504 & ~n15563 ;
  assign n14792 = n14791 ^ n14790 ;
  assign n14793 = n14792 ^ n14717 ;
  assign n14794 = n14793 ^ n14772 ;
  assign n14795 = n14682 & ~n14794 ;
  assign n14776 = n14717 ^ n14715 ;
  assign n14774 = n14756 ^ n14715 ;
  assign n14775 = n14774 ^ n14772 ;
  assign n14777 = n14776 ^ n14775 ;
  assign n14796 = n14795 ^ n14777 ;
  assign n14779 = n14778 ^ n14777 ;
  assign n14773 = n14772 ^ n14761 ;
  assign n14780 = n14779 ^ n14773 ;
  assign n14781 = n14780 ^ n14762 ;
  assign n14782 = n14781 ^ n14720 ;
  assign n14783 = n14782 ^ n14781 ;
  assign n14784 = n14781 ^ n14754 ;
  assign n14785 = n14784 ^ n14781 ;
  assign n14786 = n14783 & n14785 ;
  assign n14787 = n14786 ^ n14781 ;
  assign n14788 = n14682 & ~n14787 ;
  assign n14789 = n14788 ^ n14780 ;
  assign n14797 = n14796 ^ n14789 ;
  assign n14798 = n14681 & ~n14797 ;
  assign n15545 = n14798 ^ n14789 ;
  assign n15546 = n15545 ^ n13183 ;
  assign n15547 = n15546 ^ x118 ;
  assign n15583 = n15564 ^ n15547 ;
  assign n15584 = n15503 & ~n15583 ;
  assign n15505 = n15503 & ~n15504 ;
  assign n15548 = ~n15544 & ~n15547 ;
  assign n15568 = n15505 & n15548 ;
  assign n15549 = n15548 ^ n15547 ;
  assign n15550 = n15549 ^ n15544 ;
  assign n15553 = n15505 & ~n15550 ;
  assign n15569 = n15568 ^ n15553 ;
  assign n15566 = n15505 & ~n15549 ;
  assign n15567 = n15566 ^ n15505 ;
  assign n15570 = n15569 ^ n15567 ;
  assign n15561 = n15503 & ~n15549 ;
  assign n15582 = n15570 ^ n15561 ;
  assign n15585 = n15584 ^ n15582 ;
  assign n15621 = ~n15464 & n15585 ;
  assign n15579 = n15563 ^ n15547 ;
  assign n15580 = n15579 ^ n15504 ;
  assign n15599 = n15582 ^ n15580 ;
  assign n15506 = n15505 ^ n15504 ;
  assign n15507 = n15506 ^ n15503 ;
  assign n15587 = n15507 & n15548 ;
  assign n15557 = n15507 & ~n15550 ;
  assign n15555 = n15505 ^ n15503 ;
  assign n15556 = ~n15550 & n15555 ;
  assign n15558 = n15557 ^ n15556 ;
  assign n15554 = n15553 ^ n15550 ;
  assign n15559 = n15558 ^ n15554 ;
  assign n15588 = n15587 ^ n15559 ;
  assign n15586 = n15585 ^ n15569 ;
  assign n15589 = n15588 ^ n15586 ;
  assign n15581 = n15580 ^ n15558 ;
  assign n15590 = n15589 ^ n15581 ;
  assign n15571 = n15570 ^ n15568 ;
  assign n15565 = n15564 ^ n15506 ;
  assign n15572 = n15571 ^ n15565 ;
  assign n15573 = n15572 ^ n15559 ;
  assign n15562 = n15561 ^ n15549 ;
  assign n15574 = n15573 ^ n15562 ;
  assign n15591 = n15590 ^ n15574 ;
  assign n15551 = n15550 ^ n15547 ;
  assign n15552 = n15507 & ~n15551 ;
  assign n15578 = n15573 ^ n15552 ;
  assign n15592 = n15591 ^ n15578 ;
  assign n15593 = n15592 ^ n15506 ;
  assign n15560 = n15559 ^ n15552 ;
  assign n15575 = n15574 ^ n15560 ;
  assign n15594 = n15593 ^ n15575 ;
  assign n15600 = n15599 ^ n15594 ;
  assign n15598 = n15562 ^ n15552 ;
  assign n15601 = n15600 ^ n15598 ;
  assign n16639 = n15601 ^ n15553 ;
  assign n16640 = n15463 & ~n16639 ;
  assign n15595 = n15594 ^ n15557 ;
  assign n16672 = n15463 & n15595 ;
  assign n15637 = n15566 ^ n15561 ;
  assign n16668 = n15637 ^ n15570 ;
  assign n16669 = ~n15464 & n16668 ;
  assign n16651 = n15582 ^ n15558 ;
  assign n16652 = n16651 ^ n15560 ;
  assign n16648 = n15566 ^ n15556 ;
  assign n16649 = n16648 ^ n15591 ;
  assign n15624 = n15462 ^ n15420 ;
  assign n16641 = n15590 ^ n15462 ;
  assign n16642 = n16641 ^ n15590 ;
  assign n16643 = n15590 ^ n15553 ;
  assign n16644 = n16643 ^ n15590 ;
  assign n16645 = n16642 & n16644 ;
  assign n16646 = n16645 ^ n15590 ;
  assign n16647 = n15624 & n16646 ;
  assign n16650 = n16649 ^ n16647 ;
  assign n16653 = n16652 ^ n16650 ;
  assign n16654 = n16653 ^ n16647 ;
  assign n16655 = n15420 & n16654 ;
  assign n16656 = n16655 ^ n16650 ;
  assign n16670 = n16669 ^ n16656 ;
  assign n16660 = n15547 ^ n15503 ;
  assign n16661 = n16660 ^ n15504 ;
  assign n16662 = n16661 ^ n15600 ;
  assign n16665 = n15420 & n16662 ;
  assign n16657 = n16656 ^ n16647 ;
  assign n16666 = n16665 ^ n16657 ;
  assign n16667 = n15462 & ~n16666 ;
  assign n16671 = n16670 ^ n16667 ;
  assign n16673 = n16672 ^ n16671 ;
  assign n16674 = ~n16640 & n16673 ;
  assign n15576 = ~n15464 & n15575 ;
  assign n16675 = n16674 ^ n15576 ;
  assign n16676 = ~n15621 & n16675 ;
  assign n16677 = n16676 ^ n13293 ;
  assign n16678 = n16677 ^ x72 ;
  assign n16703 = n16638 & ~n16678 ;
  assign n16704 = n16703 ^ n16638 ;
  assign n14181 = ~n14011 & n14140 ;
  assign n14202 = n14170 ^ n14138 ;
  assign n14197 = n14144 ^ n14140 ;
  assign n14199 = n14198 ^ n14197 ;
  assign n14203 = n14202 ^ n14199 ;
  assign n14196 = n14195 ^ n14174 ;
  assign n14200 = n14199 ^ n14196 ;
  assign n14201 = ~n14010 & n14200 ;
  assign n14204 = n14203 ^ n14201 ;
  assign n14205 = n14011 & ~n14204 ;
  assign n14206 = n14205 ^ n14202 ;
  assign n14194 = n14163 & ~n14193 ;
  assign n14207 = n14206 ^ n14194 ;
  assign n14183 = n14165 ^ n14161 ;
  assign n14182 = n14151 ^ n14141 ;
  assign n14184 = n14183 ^ n14182 ;
  assign n14185 = n14183 ^ n14010 ;
  assign n14186 = n14185 ^ n14183 ;
  assign n14187 = ~n14184 & n14186 ;
  assign n14188 = n14187 ^ n14183 ;
  assign n14189 = n13975 & ~n14188 ;
  assign n14208 = n14207 ^ n14189 ;
  assign n14209 = ~n14181 & n14208 ;
  assign n14218 = n14209 & ~n14217 ;
  assign n14179 = n14178 ^ n14177 ;
  assign n14180 = n14179 ^ n11795 ;
  assign n14219 = n14218 ^ n14180 ;
  assign n14220 = n14219 ^ x114 ;
  assign n13905 = n13865 ^ n13828 ;
  assign n13906 = n13905 ^ n13873 ;
  assign n13907 = n13906 ^ n13905 ;
  assign n13908 = n13905 ^ n13679 ;
  assign n13909 = n13908 ^ n13905 ;
  assign n13910 = ~n13907 & ~n13909 ;
  assign n13911 = n13910 ^ n13905 ;
  assign n13912 = ~n13647 & n13911 ;
  assign n13913 = n13912 ^ n13846 ;
  assign n13897 = n13872 ^ n13831 ;
  assign n13898 = n13897 ^ n13846 ;
  assign n13899 = n13898 ^ n13827 ;
  assign n13900 = n13827 ^ n13647 ;
  assign n13901 = n13900 ^ n13827 ;
  assign n13902 = ~n13899 & n13901 ;
  assign n13903 = n13902 ^ n13827 ;
  assign n13904 = ~n13842 & n13903 ;
  assign n13914 = n13913 ^ n13904 ;
  assign n13915 = n13914 ^ n13895 ;
  assign n13930 = n13929 ^ n13915 ;
  assign n13889 = n13888 ^ n13886 ;
  assign n13890 = n13888 ^ n13647 ;
  assign n13891 = n13890 ^ n13888 ;
  assign n13892 = ~n13889 & n13891 ;
  assign n13893 = n13892 ^ n13888 ;
  assign n13894 = n13842 & ~n13893 ;
  assign n13931 = n13930 ^ n13894 ;
  assign n13932 = n13931 ^ n13839 ;
  assign n13933 = n13932 ^ n13884 ;
  assign n13877 = n13847 ^ n13647 ;
  assign n13878 = n13877 ^ n13847 ;
  assign n13879 = n13848 ^ n13847 ;
  assign n13880 = n13879 ^ n13847 ;
  assign n13881 = ~n13878 & n13880 ;
  assign n13882 = n13881 ^ n13847 ;
  assign n13883 = ~n13842 & n13882 ;
  assign n13934 = n13933 ^ n13883 ;
  assign n13874 = n13873 ^ n13833 ;
  assign n13875 = n13862 & ~n13874 ;
  assign n13853 = n13839 ^ n13823 ;
  assign n13854 = n13853 ^ n13751 ;
  assign n13855 = n13854 ^ n13823 ;
  assign n13856 = n13823 ^ n13647 ;
  assign n13857 = n13856 ^ n13823 ;
  assign n13858 = ~n13855 & n13857 ;
  assign n13859 = n13858 ^ n13823 ;
  assign n13860 = n13679 & n13859 ;
  assign n13876 = n13875 ^ n13860 ;
  assign n13935 = n13934 ^ n13876 ;
  assign n13843 = n13839 ^ n13835 ;
  assign n13844 = n13843 ^ n13748 ;
  assign n13845 = n13844 ^ n13839 ;
  assign n13849 = n13848 ^ n13845 ;
  assign n13850 = ~n13647 & n13849 ;
  assign n13851 = n13850 ^ n13843 ;
  assign n13852 = n13842 & n13851 ;
  assign n13936 = n13935 ^ n13852 ;
  assign n13937 = ~n13841 & ~n13936 ;
  assign n13938 = n13937 ^ n11963 ;
  assign n13939 = n13938 ^ x115 ;
  assign n14395 = n14373 ^ n14337 ;
  assign n14396 = n14395 ^ n14393 ;
  assign n14397 = ~n14222 & n14396 ;
  assign n14389 = n14340 ^ n14332 ;
  assign n14390 = n14389 ^ n14363 ;
  assign n14391 = n14390 ^ n14335 ;
  assign n14394 = n14393 ^ n14391 ;
  assign n14398 = n14397 ^ n14394 ;
  assign n14399 = n14257 & ~n14398 ;
  assign n14387 = ~n14256 & n14337 ;
  assign n14381 = n14380 ^ n14341 ;
  assign n14378 = n14377 ^ n14372 ;
  assign n14382 = n14381 ^ n14378 ;
  assign n14383 = n14222 & ~n14382 ;
  assign n14379 = n14378 ^ n14366 ;
  assign n14384 = n14383 ^ n14379 ;
  assign n14385 = ~n14257 & ~n14384 ;
  assign n14361 = n14360 ^ n14340 ;
  assign n14352 = n14351 ^ n14344 ;
  assign n14353 = n14344 ^ n14222 ;
  assign n14354 = n14353 ^ n14344 ;
  assign n14355 = n14352 & ~n14354 ;
  assign n14356 = n14355 ^ n14344 ;
  assign n14357 = n14257 & n14356 ;
  assign n14362 = n14361 ^ n14357 ;
  assign n14386 = n14385 ^ n14362 ;
  assign n14388 = n14387 ^ n14386 ;
  assign n14400 = n14399 ^ n14388 ;
  assign n14408 = ~n14400 & ~n14407 ;
  assign n14409 = n14408 ^ n11756 ;
  assign n14410 = n14409 ^ x96 ;
  assign n14427 = ~n13939 & ~n14410 ;
  assign n13596 = n13550 & ~n13595 ;
  assign n13585 = n13584 ^ n13170 ;
  assign n13587 = n13584 ^ n13538 ;
  assign n13586 = n13584 ^ n13552 ;
  assign n13588 = n13587 ^ n13586 ;
  assign n13589 = n13587 ^ n13148 ;
  assign n13590 = n13589 ^ n13587 ;
  assign n13591 = n13588 & n13590 ;
  assign n13592 = n13591 ^ n13587 ;
  assign n13593 = ~n13585 & ~n13592 ;
  assign n13594 = n13593 ^ n13170 ;
  assign n13597 = n13596 ^ n13594 ;
  assign n13574 = n13567 ^ n13554 ;
  assign n13575 = n13574 ^ n13534 ;
  assign n13576 = n13575 ^ n13557 ;
  assign n13573 = n13328 ^ n13325 ;
  assign n13577 = n13576 ^ n13573 ;
  assign n13572 = n13531 & n13571 ;
  assign n13578 = n13577 ^ n13572 ;
  assign n13579 = n13148 & ~n13578 ;
  assign n13580 = n13579 ^ n13576 ;
  assign n13581 = n13170 & ~n13580 ;
  assign n13598 = n13597 ^ n13581 ;
  assign n13599 = n13557 ^ n13548 ;
  assign n13600 = ~n13170 & n13599 ;
  assign n13601 = n13600 ^ n13561 ;
  assign n13603 = n13601 ^ n13587 ;
  assign n13602 = n13601 ^ n13575 ;
  assign n13604 = n13603 ^ n13602 ;
  assign n13607 = ~n13170 & ~n13604 ;
  assign n13608 = n13607 ^ n13603 ;
  assign n13609 = ~n13148 & n13608 ;
  assign n13610 = n13609 ^ n13601 ;
  assign n13611 = n13598 & ~n13610 ;
  assign n13612 = ~n13568 & n13611 ;
  assign n13613 = n13612 ^ n11722 ;
  assign n13614 = n13613 ^ x105 ;
  assign n14412 = ~n13614 & ~n14410 ;
  assign n14428 = n14427 ^ n14412 ;
  assign n14433 = n14220 & n14428 ;
  assign n13102 = n13101 ^ n13075 ;
  assign n13103 = n13102 ^ n13095 ;
  assign n13139 = n13103 ^ n12718 ;
  assign n13140 = n13103 ^ n12924 ;
  assign n13141 = n13140 ^ n13103 ;
  assign n13142 = ~n13139 & ~n13141 ;
  assign n13143 = n13142 ^ n13103 ;
  assign n13144 = ~n13064 & ~n13143 ;
  assign n13145 = n13144 ^ n11688 ;
  assign n13061 = ~n12924 & n13060 ;
  assign n13062 = n13061 ^ n13060 ;
  assign n13063 = n12718 & n13062 ;
  assign n13104 = n13103 ^ n13071 ;
  assign n13108 = n13107 ^ n13104 ;
  assign n13109 = ~n12924 & n13108 ;
  assign n13110 = n13109 ^ n13107 ;
  assign n13126 = n13110 ^ n13078 ;
  assign n13123 = n13080 ^ n13065 ;
  assign n13124 = n13123 ^ n12718 ;
  assign n13125 = ~n12924 & ~n13124 ;
  assign n13127 = n13126 ^ n13125 ;
  assign n13128 = n13060 & ~n13127 ;
  assign n13081 = n13080 ^ n13072 ;
  assign n13082 = n13080 ^ n12924 ;
  assign n13083 = n13082 ^ n13080 ;
  assign n13084 = n13081 & n13083 ;
  assign n13085 = n13084 ^ n13080 ;
  assign n13086 = ~n13064 & ~n13085 ;
  assign n13111 = n13110 ^ n13086 ;
  assign n13122 = n13121 ^ n13111 ;
  assign n13129 = n13128 ^ n13122 ;
  assign n13131 = n13130 ^ n13072 ;
  assign n13132 = n13072 ^ n12924 ;
  assign n13133 = n13132 ^ n13072 ;
  assign n13134 = n13131 & n13133 ;
  assign n13135 = n13134 ^ n13072 ;
  assign n13136 = n13060 & ~n13135 ;
  assign n13137 = n13129 & ~n13136 ;
  assign n13138 = ~n13063 & n13137 ;
  assign n13146 = n13145 ^ n13138 ;
  assign n13147 = n13146 ^ x72 ;
  assign n14604 = n14603 ^ n14537 ;
  assign n14602 = n14564 ^ n14528 ;
  assign n14605 = n14604 ^ n14602 ;
  assign n14606 = n14441 & n14605 ;
  assign n14607 = n14606 ^ n14556 ;
  assign n14608 = ~n14442 & n14607 ;
  assign n14600 = n14555 & n14599 ;
  assign n14586 = n14585 ^ n14540 ;
  assign n14587 = ~n14441 & n14586 ;
  assign n14588 = n14587 ^ n14540 ;
  assign n14589 = n14588 ^ n14584 ;
  assign n14590 = n14589 ^ n14588 ;
  assign n14593 = n14441 & n14590 ;
  assign n14594 = n14593 ^ n14588 ;
  assign n14595 = ~n14442 & n14594 ;
  assign n14596 = n14595 ^ n14588 ;
  assign n14570 = n14551 ^ n14442 ;
  assign n14573 = n14572 ^ n14553 ;
  assign n14579 = n14578 ^ n14573 ;
  assign n14580 = n14579 ^ n14559 ;
  assign n14581 = ~n14570 & n14580 ;
  assign n14567 = n14566 ^ n14563 ;
  assign n14568 = n14552 & ~n14567 ;
  assign n14530 = n14529 ^ n14525 ;
  assign n14531 = n14441 & n14530 ;
  assign n14532 = n14531 ^ n14529 ;
  assign n14533 = n14532 ^ n14441 ;
  assign n14535 = n14533 ^ n14524 ;
  assign n14536 = n14535 ^ n14533 ;
  assign n14545 = ~n14536 & ~n14542 ;
  assign n14546 = ~n14441 & n14545 ;
  assign n14547 = n14546 ^ n14441 ;
  assign n14548 = n14547 ^ n14532 ;
  assign n14549 = n14443 & ~n14548 ;
  assign n14550 = n14549 ^ n14532 ;
  assign n14569 = n14568 ^ n14550 ;
  assign n14582 = n14581 ^ n14569 ;
  assign n14583 = n14582 ^ n14556 ;
  assign n14597 = n14596 ^ n14583 ;
  assign n14598 = n14597 ^ n11655 ;
  assign n14601 = n14600 ^ n14598 ;
  assign n14609 = n14608 ^ n14601 ;
  assign n14610 = n14609 ^ x90 ;
  assign n14221 = n14220 ^ n13939 ;
  assign n14417 = n14410 ^ n13614 ;
  assign n14424 = n14417 ^ n14220 ;
  assign n14425 = ~n14221 & n14424 ;
  assign n14426 = n14425 ^ n13939 ;
  assign n14431 = n14220 ^ n13614 ;
  assign n14432 = ~n14426 & n14431 ;
  assign n16176 = n14432 ^ n14417 ;
  assign n14411 = n14410 ^ n14221 ;
  assign n14413 = n14412 ^ n13939 ;
  assign n14414 = n14411 & n14413 ;
  assign n13940 = n13939 ^ n13614 ;
  assign n14415 = n14414 ^ n13940 ;
  assign n14416 = n14410 ^ n13939 ;
  assign n14420 = ~n14416 & n14417 ;
  assign n14421 = n14420 ^ n14410 ;
  assign n14422 = ~n14411 & n14421 ;
  assign n14423 = n14415 & ~n14422 ;
  assign n16177 = n16176 ^ n14423 ;
  assign n16178 = ~n14610 & n16177 ;
  assign n16179 = n16178 ^ n14423 ;
  assign n16175 = n14610 ^ n14423 ;
  assign n16180 = n16179 ^ n16175 ;
  assign n16181 = n16180 ^ n16176 ;
  assign n16183 = n16181 ^ n14415 ;
  assign n14613 = n14422 ^ n14410 ;
  assign n16182 = n16181 ^ n14613 ;
  assign n16184 = n16183 ^ n16182 ;
  assign n16187 = n14610 & ~n16184 ;
  assign n16188 = n16187 ^ n16183 ;
  assign n16189 = n13147 & ~n16188 ;
  assign n16190 = n16189 ^ n16181 ;
  assign n16191 = ~n14433 & ~n16190 ;
  assign n16192 = n16191 ^ n13169 ;
  assign n16193 = n16192 ^ x113 ;
  assign n16334 = n15502 ^ x109 ;
  assign n14799 = n14796 ^ n14681 ;
  assign n14800 = n14799 ^ n14798 ;
  assign n14801 = n14800 ^ n12246 ;
  assign n16335 = n14801 ^ x92 ;
  assign n16336 = ~n16334 & ~n16335 ;
  assign n16337 = n16336 ^ n16335 ;
  assign n16245 = n15461 ^ x68 ;
  assign n16247 = n13061 ^ n12924 ;
  assign n16248 = n16247 ^ n13060 ;
  assign n16249 = n13130 ^ n13103 ;
  assign n16257 = n13065 ^ n12924 ;
  assign n16262 = n13070 ^ n13065 ;
  assign n16263 = n16262 ^ n12715 ;
  assign n16258 = n13065 ^ n12708 ;
  assign n16259 = n16258 ^ n13103 ;
  assign n16260 = n16259 ^ n12715 ;
  assign n16261 = n13060 & n16260 ;
  assign n16264 = n16263 ^ n16261 ;
  assign n16265 = ~n16257 & ~n16264 ;
  assign n16266 = n16265 ^ n12924 ;
  assign n16256 = n13061 & ~n13113 ;
  assign n16267 = n16266 ^ n16256 ;
  assign n16250 = n12716 ^ n12708 ;
  assign n16251 = n16250 ^ n13068 ;
  assign n16252 = n16251 ^ n13093 ;
  assign n16253 = ~n13060 & n16252 ;
  assign n16254 = n16253 ^ n13093 ;
  assign n16255 = n12924 & ~n16254 ;
  assign n16268 = n16267 ^ n16255 ;
  assign n16269 = ~n13144 & n16268 ;
  assign n16270 = n16249 & n16269 ;
  assign n16271 = n16248 & n16270 ;
  assign n16272 = n16271 ^ n16269 ;
  assign n16273 = n13101 ^ n13064 ;
  assign n16274 = n16273 ^ n13101 ;
  assign n16275 = n13060 & n13069 ;
  assign n16276 = n16275 ^ n13101 ;
  assign n16277 = ~n16274 & n16276 ;
  assign n16278 = n16277 ^ n13101 ;
  assign n16279 = n16272 & n16278 ;
  assign n16280 = n16279 ^ n16272 ;
  assign n16281 = ~n13086 & n16280 ;
  assign n16282 = ~n13063 & n16281 ;
  assign n16285 = n16282 ^ n12837 ;
  assign n16246 = n13094 ^ n13092 ;
  assign n16283 = ~n16247 & n16282 ;
  assign n16284 = ~n16246 & n16283 ;
  assign n16286 = n16285 ^ n16284 ;
  assign n16287 = n16286 ^ x85 ;
  assign n16288 = ~n16245 & ~n16287 ;
  assign n16224 = n14579 ^ n14521 ;
  assign n16225 = n16224 ^ n14561 ;
  assign n16222 = n14493 ^ n14492 ;
  assign n16223 = n16222 ^ n14520 ;
  assign n16226 = n16225 ^ n16223 ;
  assign n16227 = n16226 ^ n14443 ;
  assign n16228 = n14578 & n16227 ;
  assign n16229 = n16228 ^ n14443 ;
  assign n16205 = n15155 ^ n14524 ;
  assign n16211 = n16205 ^ n14558 ;
  assign n16203 = n14565 ^ n14560 ;
  assign n16204 = n16203 ^ n14537 ;
  assign n16206 = n16205 ^ n16204 ;
  assign n16207 = n16204 ^ n14441 ;
  assign n16208 = n14443 & n16207 ;
  assign n16209 = n16208 ^ n14441 ;
  assign n16210 = ~n16206 & n16209 ;
  assign n16212 = n16211 ^ n16210 ;
  assign n16230 = n16212 ^ n14578 ;
  assign n16231 = n16230 ^ n14599 ;
  assign n16232 = n16231 ^ n16212 ;
  assign n16233 = n16229 & ~n16232 ;
  assign n16234 = n16233 ^ n16230 ;
  assign n16235 = n16234 ^ n14579 ;
  assign n16221 = n15178 ^ n12812 ;
  assign n16236 = n16235 ^ n16221 ;
  assign n16213 = n16212 ^ n14571 ;
  assign n16214 = n16213 ^ n14559 ;
  assign n16215 = n16214 ^ n16212 ;
  assign n16216 = n16212 ^ n14441 ;
  assign n16217 = n16216 ^ n16212 ;
  assign n16218 = ~n16215 & n16217 ;
  assign n16219 = n16218 ^ n16212 ;
  assign n16220 = n14443 & n16219 ;
  assign n16237 = n16236 ^ n16220 ;
  assign n16202 = n14552 & n14561 ;
  assign n16238 = n16237 ^ n16202 ;
  assign n16201 = n14542 & n14551 ;
  assign n16239 = n16238 ^ n16201 ;
  assign n16194 = n14579 ^ n14555 ;
  assign n16195 = n16194 ^ n14579 ;
  assign n16196 = n14579 ^ n14441 ;
  assign n16197 = n16196 ^ n14579 ;
  assign n16198 = n16195 & ~n16197 ;
  assign n16199 = n16198 ^ n14579 ;
  assign n16200 = ~n14442 & ~n16199 ;
  assign n16240 = n16239 ^ n16200 ;
  assign n16241 = n16240 ^ x70 ;
  assign n14673 = n14667 ^ n13564 ;
  assign n14671 = n13558 ^ n13551 ;
  assign n14648 = n13583 ^ n13548 ;
  assign n14672 = n14671 ^ n14648 ;
  assign n14674 = n14673 ^ n14672 ;
  assign n14675 = n13172 & n14674 ;
  assign n14662 = n14648 ^ n13564 ;
  assign n14663 = n14662 ^ n14661 ;
  assign n14657 = n13554 ^ n13548 ;
  assign n14658 = n14657 ^ n13564 ;
  assign n14659 = n13174 & n14658 ;
  assign n14664 = n14663 ^ n14659 ;
  assign n14649 = n14648 ^ n13550 ;
  assign n14650 = n14649 ^ n13148 ;
  assign n14651 = n14650 ^ n14649 ;
  assign n14652 = n14649 ^ n13557 ;
  assign n14653 = n14652 ^ n14649 ;
  assign n14654 = ~n14651 & n14653 ;
  assign n14655 = n14654 ^ n14649 ;
  assign n14656 = ~n13170 & n14655 ;
  assign n14665 = n14664 ^ n14656 ;
  assign n14668 = n14667 ^ n14665 ;
  assign n14638 = ~n13148 & n13547 ;
  assign n14639 = n14638 ^ n13540 ;
  assign n14640 = n14639 ^ n14637 ;
  assign n14641 = n14640 ^ n14639 ;
  assign n14642 = n14639 ^ n13170 ;
  assign n14643 = n14642 ^ n14639 ;
  assign n14644 = ~n14641 & n14643 ;
  assign n14645 = n14644 ^ n14639 ;
  assign n14646 = n13595 & n14645 ;
  assign n14647 = n14646 ^ n14639 ;
  assign n14669 = n14668 ^ n14647 ;
  assign n14670 = n14669 ^ n12295 ;
  assign n14676 = n14675 ^ n14670 ;
  assign n14628 = n13555 ^ n13170 ;
  assign n14629 = n14628 ^ n13555 ;
  assign n14631 = n14630 ^ n13539 ;
  assign n14632 = n14631 ^ n13555 ;
  assign n14633 = ~n14629 & n14632 ;
  assign n14634 = n14633 ^ n13555 ;
  assign n14635 = n13148 & n14634 ;
  assign n14677 = n14676 ^ n14635 ;
  assign n16242 = n14677 ^ x110 ;
  assign n16243 = n16241 & ~n16242 ;
  assign n16244 = n16243 ^ n16241 ;
  assign n16309 = n16244 ^ n16242 ;
  assign n16310 = n16288 & n16309 ;
  assign n16293 = n16288 ^ n16287 ;
  assign n16294 = n16293 ^ n16245 ;
  assign n16295 = n16244 & ~n16294 ;
  assign n16292 = n16244 & n16288 ;
  assign n16296 = n16295 ^ n16292 ;
  assign n16289 = n16288 ^ n16245 ;
  assign n16290 = n16244 & ~n16289 ;
  assign n16291 = n16290 ^ n16244 ;
  assign n16297 = n16296 ^ n16291 ;
  assign n16311 = n16310 ^ n16297 ;
  assign n16312 = n16311 ^ n16295 ;
  assign n16313 = n16312 ^ n16290 ;
  assign n16306 = n16287 ^ n16241 ;
  assign n16307 = n16242 & ~n16306 ;
  assign n16308 = n16307 ^ n16297 ;
  assign n16314 = n16313 ^ n16308 ;
  assign n16318 = n16314 ^ n16297 ;
  assign n16299 = n16243 ^ n16242 ;
  assign n16301 = ~n16293 & ~n16299 ;
  assign n16317 = n16301 ^ n16293 ;
  assign n16319 = n16318 ^ n16317 ;
  assign n16303 = n16243 & n16288 ;
  assign n16381 = n16319 ^ n16303 ;
  assign n16324 = n16243 & ~n16294 ;
  assign n16380 = n16324 ^ n16243 ;
  assign n16382 = n16381 ^ n16380 ;
  assign n16383 = ~n16337 & ~n16382 ;
  assign n16338 = n16337 ^ n16334 ;
  assign n16300 = ~n16289 & ~n16299 ;
  assign n16377 = n16319 ^ n16300 ;
  assign n16378 = ~n16338 & ~n16377 ;
  assign n16315 = n16314 ^ n16311 ;
  assign n16316 = n16315 ^ n16292 ;
  assign n16320 = n16319 ^ n16316 ;
  assign n16304 = n16303 ^ n16301 ;
  assign n16305 = n16304 ^ n16287 ;
  assign n16321 = n16320 ^ n16305 ;
  assign n16322 = n16321 ^ n16299 ;
  assign n16302 = n16301 ^ n16300 ;
  assign n16323 = n16322 ^ n16302 ;
  assign n16325 = n16324 ^ n16323 ;
  assign n16326 = n16325 ^ n16294 ;
  assign n16327 = n16326 ^ n16313 ;
  assign n16328 = n16327 ^ n16310 ;
  assign n16298 = n16297 ^ n16290 ;
  assign n16329 = n16328 ^ n16298 ;
  assign n16372 = n16329 ^ n16323 ;
  assign n16342 = n16328 ^ n16292 ;
  assign n16343 = n16342 ^ n16309 ;
  assign n16344 = ~n16335 & n16343 ;
  assign n16345 = n16344 ^ n16313 ;
  assign n16371 = n16345 ^ n16307 ;
  assign n16373 = n16372 ^ n16371 ;
  assign n16367 = n16313 ^ n16293 ;
  assign n16368 = n16367 ^ n16323 ;
  assign n16369 = n16368 ^ n16243 ;
  assign n16370 = n16335 & n16369 ;
  assign n16374 = n16373 ^ n16370 ;
  assign n16375 = ~n16334 & ~n16374 ;
  assign n16356 = n16335 ^ n16334 ;
  assign n16330 = n16329 ^ n16321 ;
  assign n16357 = n16330 ^ n16329 ;
  assign n16358 = n16357 ^ n16318 ;
  assign n16359 = n16358 ^ n16329 ;
  assign n16360 = n16359 ^ n16357 ;
  assign n16361 = n16357 ^ n16335 ;
  assign n16362 = n16361 ^ n16357 ;
  assign n16363 = n16360 & n16362 ;
  assign n16364 = n16363 ^ n16357 ;
  assign n16365 = n16356 & n16364 ;
  assign n16347 = n16324 ^ n16300 ;
  assign n16348 = n16347 ^ n16304 ;
  assign n16351 = ~n16334 & n16348 ;
  assign n16352 = n16351 ^ n16304 ;
  assign n16353 = ~n16335 & n16352 ;
  assign n16331 = n16329 ^ n16318 ;
  assign n16332 = n16331 ^ n16309 ;
  assign n16333 = n16332 ^ n16311 ;
  assign n16339 = n16338 ^ n16335 ;
  assign n16340 = n16333 & ~n16339 ;
  assign n16341 = n16340 ^ n16330 ;
  assign n16346 = n16345 ^ n16341 ;
  assign n16354 = n16353 ^ n16346 ;
  assign n16355 = n16354 ^ n13646 ;
  assign n16366 = n16365 ^ n16355 ;
  assign n16376 = n16375 ^ n16366 ;
  assign n16379 = n16378 ^ n16376 ;
  assign n16384 = n16383 ^ n16379 ;
  assign n16385 = n16384 ^ x82 ;
  assign n16386 = n16193 & n16385 ;
  assign n16588 = n16386 ^ n16193 ;
  assign n16024 = n14647 ^ n10783 ;
  assign n15996 = n13543 ^ n13536 ;
  assign n15997 = n13148 & n15996 ;
  assign n15995 = ~n13170 & n13551 ;
  assign n15998 = n15997 ^ n15995 ;
  assign n16020 = n13565 ^ n13545 ;
  assign n16021 = n13171 & n16020 ;
  assign n16006 = n15514 ^ n13557 ;
  assign n16001 = n13555 ^ n13551 ;
  assign n16002 = n16001 ^ n14648 ;
  assign n15999 = n13563 ^ n13559 ;
  assign n16003 = n16002 ^ n15999 ;
  assign n16004 = ~n13148 & n16003 ;
  assign n16000 = n15999 ^ n15514 ;
  assign n16005 = n16004 ^ n16000 ;
  assign n16007 = n16006 ^ n16005 ;
  assign n16010 = n16007 ^ n13557 ;
  assign n16011 = n16010 ^ n16007 ;
  assign n16012 = n16007 ^ n14637 ;
  assign n16013 = n16012 ^ n16007 ;
  assign n16014 = ~n16011 & ~n16013 ;
  assign n16015 = ~n13148 & n16014 ;
  assign n16016 = n16015 ^ n13148 ;
  assign n16008 = n16007 ^ n13148 ;
  assign n16017 = n16016 ^ n16008 ;
  assign n16018 = ~n13595 & n16017 ;
  assign n16019 = n16018 ^ n16005 ;
  assign n16022 = n16021 ^ n16019 ;
  assign n16023 = ~n15998 & ~n16022 ;
  assign n16025 = n16024 ^ n16023 ;
  assign n16445 = n16025 ^ x106 ;
  assign n15681 = ~n14153 & ~n14193 ;
  assign n15672 = n14192 ^ n14146 ;
  assign n15673 = n14202 ^ n14165 ;
  assign n15674 = n15673 ^ n14190 ;
  assign n15675 = n14192 ^ n14190 ;
  assign n15676 = n15675 ^ n14190 ;
  assign n15677 = n15674 & n15676 ;
  assign n15678 = n15677 ^ n14190 ;
  assign n15679 = ~n15672 & ~n15678 ;
  assign n15660 = n14149 ^ n14145 ;
  assign n15661 = n14145 ^ n13975 ;
  assign n15662 = n15661 ^ n14145 ;
  assign n15663 = n15660 & ~n15662 ;
  assign n15664 = n15663 ^ n14145 ;
  assign n15665 = n14010 & ~n15664 ;
  assign n15666 = n15665 ^ n14146 ;
  assign n15667 = n15666 ^ n15495 ;
  assign n15655 = n14160 ^ n14078 ;
  assign n15656 = n14190 & ~n15655 ;
  assign n15657 = n14160 ^ n14044 ;
  assign n15658 = n15657 ^ n14124 ;
  assign n15659 = n15656 & n15658 ;
  assign n15668 = n15667 ^ n15659 ;
  assign n15669 = n15668 ^ n15497 ;
  assign n15670 = n15669 ^ n15492 ;
  assign n15671 = n15670 ^ n11081 ;
  assign n15680 = n15679 ^ n15671 ;
  assign n15682 = n15681 ^ n15680 ;
  assign n15652 = n14141 ^ n14134 ;
  assign n15653 = n15652 ^ n15467 ;
  assign n15654 = n14191 & n15653 ;
  assign n15683 = n15682 ^ n15654 ;
  assign n16446 = n15683 ^ x97 ;
  assign n16447 = ~n16445 & n16446 ;
  assign n16467 = n16447 ^ n16445 ;
  assign n16416 = n13144 ^ n9941 ;
  assign n16402 = n15253 ^ n13070 ;
  assign n16403 = n16402 ^ n13089 ;
  assign n16404 = n13089 ^ n12924 ;
  assign n16405 = n16404 ^ n13089 ;
  assign n16406 = ~n16403 & n16405 ;
  assign n16407 = n16406 ^ n13089 ;
  assign n16408 = ~n13060 & n16407 ;
  assign n16409 = n16408 ^ n13072 ;
  assign n16401 = ~n13064 & n13066 ;
  assign n16410 = n16409 ^ n16401 ;
  assign n16398 = n13098 & ~n13133 ;
  assign n16399 = n16398 ^ n13072 ;
  assign n16400 = n13060 & ~n16399 ;
  assign n16411 = n16410 ^ n16400 ;
  assign n16389 = n13068 ^ n12717 ;
  assign n16412 = n16411 ^ n16389 ;
  assign n16390 = n16389 ^ n16246 ;
  assign n16391 = n16390 ^ n16389 ;
  assign n16392 = n16389 ^ n13060 ;
  assign n16393 = n16392 ^ n16389 ;
  assign n16394 = ~n16391 & n16393 ;
  assign n16395 = n16394 ^ n16389 ;
  assign n16396 = ~n13064 & n16395 ;
  assign n16413 = n16412 ^ n16396 ;
  assign n16414 = ~n13136 & n16413 ;
  assign n16415 = ~n13063 & n16414 ;
  assign n16417 = n16416 ^ n16415 ;
  assign n16418 = n16417 ^ x123 ;
  assign n16430 = n15217 ^ n14348 ;
  assign n16420 = n14372 ^ n14222 ;
  assign n16421 = n16420 ^ n14372 ;
  assign n16422 = ~n15213 & n16421 ;
  assign n16423 = n16422 ^ n14372 ;
  assign n16424 = ~n14256 & ~n16423 ;
  assign n16428 = n16424 ^ n14357 ;
  assign n16425 = n14347 ^ n14335 ;
  assign n16426 = n16425 ^ n14377 ;
  assign n16427 = ~n14222 & ~n16426 ;
  assign n16429 = n16428 ^ n16427 ;
  assign n16431 = n16430 ^ n16429 ;
  assign n16432 = n16431 ^ n16424 ;
  assign n16433 = ~n14257 & n16432 ;
  assign n16434 = n16433 ^ n16429 ;
  assign n16435 = ~n15211 & ~n16434 ;
  assign n16436 = n15244 & n16435 ;
  assign n16437 = ~n15447 & n16436 ;
  assign n16439 = n14222 & n15442 ;
  assign n16440 = n16437 & n16439 ;
  assign n16438 = n16437 ^ n10525 ;
  assign n16441 = n16440 ^ n16438 ;
  assign n16442 = n16441 ^ x80 ;
  assign n16443 = ~n16418 & n16442 ;
  assign n16444 = n16443 ^ n16418 ;
  assign n15923 = n14854 & n14952 ;
  assign n15912 = n14945 ^ n14942 ;
  assign n15913 = n15912 ^ n14938 ;
  assign n15914 = n14855 & n15913 ;
  assign n15915 = n15914 ^ n14856 ;
  assign n15918 = n14950 ^ n14934 ;
  assign n15916 = n14944 ^ n14938 ;
  assign n15917 = n14855 & ~n15916 ;
  assign n15919 = n15918 ^ n15917 ;
  assign n15920 = ~n15915 & ~n15919 ;
  assign n15905 = n14943 ^ n14930 ;
  assign n15906 = n15905 ^ n14961 ;
  assign n15903 = n14939 ^ n14928 ;
  assign n15904 = n15903 ^ n14945 ;
  assign n15907 = n15906 ^ n15904 ;
  assign n15908 = n14853 & n15907 ;
  assign n15909 = n15908 ^ n15904 ;
  assign n15910 = n14854 & n15909 ;
  assign n15891 = n15327 ^ n14926 ;
  assign n15892 = n15891 ^ n15327 ;
  assign n15893 = n15892 ^ n14959 ;
  assign n15894 = n15893 ^ n15892 ;
  assign n15895 = n15892 ^ n14854 ;
  assign n15896 = n15895 ^ n15892 ;
  assign n15897 = n15894 & ~n15896 ;
  assign n15898 = n15897 ^ n15892 ;
  assign n15899 = ~n14977 & n15898 ;
  assign n15900 = n15899 ^ n15891 ;
  assign n15715 = n14928 ^ n14922 ;
  assign n15716 = n15715 ^ n14854 ;
  assign n15717 = n15716 ^ n15715 ;
  assign n15718 = n14981 ^ n14922 ;
  assign n15719 = n15718 ^ n15715 ;
  assign n15720 = n15717 & n15719 ;
  assign n15721 = n15720 ^ n15715 ;
  assign n15722 = n14977 & n15721 ;
  assign n15723 = n15722 ^ n14922 ;
  assign n15901 = n15900 ^ n15723 ;
  assign n15902 = n15901 ^ n11258 ;
  assign n15911 = n15910 ^ n15902 ;
  assign n15921 = n15920 ^ n15911 ;
  assign n15890 = n14855 & ~n14933 ;
  assign n15922 = n15921 ^ n15890 ;
  assign n15924 = n15923 ^ n15922 ;
  assign n16388 = n15924 ^ x82 ;
  assign n15690 = n14565 ^ n14559 ;
  assign n15688 = n14578 ^ n14564 ;
  assign n15689 = n15688 ^ n14542 ;
  assign n15691 = n15690 ^ n15689 ;
  assign n15692 = n14441 & n15691 ;
  assign n15693 = n15692 ^ n15689 ;
  assign n15700 = n15693 ^ n14579 ;
  assign n15698 = n14604 ^ n14572 ;
  assign n15699 = ~n14441 & n15698 ;
  assign n15701 = n15700 ^ n15699 ;
  assign n15696 = n14574 ^ n14558 ;
  assign n15697 = ~n14442 & n15696 ;
  assign n15702 = n15701 ^ n15697 ;
  assign n15703 = n14443 & n15702 ;
  assign n15687 = n14596 ^ n14579 ;
  assign n15694 = n15693 ^ n15687 ;
  assign n15695 = n15694 ^ n15178 ;
  assign n15704 = n15703 ^ n15695 ;
  assign n15705 = n15704 ^ n14528 ;
  assign n15706 = n15705 ^ n11512 ;
  assign n16387 = n15706 ^ x120 ;
  assign n16516 = n16388 ^ n16387 ;
  assign n16515 = n16387 & n16388 ;
  assign n16517 = n16516 ^ n16515 ;
  assign n16539 = n16517 ^ n16388 ;
  assign n16540 = ~n16444 & n16539 ;
  assign n16541 = ~n16467 & n16540 ;
  assign n16542 = n16541 ^ n14518 ;
  assign n16448 = n16447 ^ n16446 ;
  assign n16451 = n16443 & n16448 ;
  assign n16471 = n16451 ^ n16443 ;
  assign n16469 = n16443 & n16447 ;
  assign n16468 = n16443 & ~n16467 ;
  assign n16470 = n16469 ^ n16468 ;
  assign n16472 = n16471 ^ n16470 ;
  assign n16456 = ~n16444 & n16448 ;
  assign n16453 = n16444 ^ n16442 ;
  assign n16454 = n16453 ^ n16418 ;
  assign n16455 = n16448 & n16454 ;
  assign n16457 = n16456 ^ n16455 ;
  assign n16452 = n16451 ^ n16448 ;
  assign n16458 = n16457 ^ n16452 ;
  assign n16473 = n16472 ^ n16458 ;
  assign n16449 = n16448 ^ n16445 ;
  assign n16460 = n16449 & n16454 ;
  assign n16474 = n16473 ^ n16460 ;
  assign n16450 = ~n16444 & n16449 ;
  assign n16459 = n16458 ^ n16450 ;
  assign n16466 = n16459 ^ n16449 ;
  assign n16475 = n16474 ^ n16466 ;
  assign n16478 = ~n16388 & n16475 ;
  assign n16461 = n16460 ^ n16459 ;
  assign n16462 = n16388 & n16461 ;
  assign n16463 = n16462 ^ n16460 ;
  assign n16479 = n16478 ^ n16463 ;
  assign n16480 = n16387 & n16479 ;
  assign n16481 = n16480 ^ n16463 ;
  assign n16527 = n16455 ^ n16450 ;
  assign n16528 = n16527 ^ n16451 ;
  assign n16529 = n16528 ^ n16458 ;
  assign n16482 = n16447 & n16453 ;
  assign n16483 = n16482 ^ n16468 ;
  assign n16525 = n16483 ^ n16451 ;
  assign n16495 = ~n16444 & n16447 ;
  assign n16492 = n16453 & ~n16467 ;
  assign n16524 = n16495 ^ n16492 ;
  assign n16526 = n16525 ^ n16524 ;
  assign n16530 = n16529 ^ n16526 ;
  assign n16531 = n16526 ^ n16388 ;
  assign n16532 = n16531 ^ n16526 ;
  assign n16533 = n16530 & ~n16532 ;
  assign n16534 = n16533 ^ n16526 ;
  assign n16535 = n16387 & n16534 ;
  assign n16493 = n16454 & ~n16467 ;
  assign n16496 = n16495 ^ n16493 ;
  assign n16497 = n16496 ^ n16469 ;
  assign n16504 = n16497 ^ n16492 ;
  assign n16498 = n16497 ^ n16447 ;
  assign n16494 = n16493 ^ n16482 ;
  assign n16499 = n16498 ^ n16494 ;
  assign n16502 = n16499 ^ n16483 ;
  assign n16503 = n16502 ^ n16445 ;
  assign n16505 = n16504 ^ n16503 ;
  assign n16506 = n16505 ^ n16469 ;
  assign n16507 = n16506 ^ n16475 ;
  assign n16508 = n16507 ^ n16482 ;
  assign n16500 = n16499 ^ n16492 ;
  assign n16491 = n16475 ^ n16470 ;
  assign n16501 = n16500 ^ n16491 ;
  assign n16509 = n16508 ^ n16501 ;
  assign n16510 = n16388 & ~n16509 ;
  assign n16511 = n16510 ^ n16508 ;
  assign n16512 = ~n16387 & ~n16511 ;
  assign n16513 = n16512 ^ n16460 ;
  assign n16486 = n16460 ^ n16387 ;
  assign n16487 = n16486 ^ n16460 ;
  assign n16488 = n16483 & n16487 ;
  assign n16489 = n16488 ^ n16460 ;
  assign n16490 = ~n16388 & n16489 ;
  assign n16514 = n16513 ^ n16490 ;
  assign n16519 = n16457 & ~n16516 ;
  assign n16520 = ~n16514 & n16519 ;
  assign n16521 = n16520 ^ n16514 ;
  assign n16536 = n16535 ^ n16521 ;
  assign n16518 = n16517 ^ n16514 ;
  assign n16523 = n16472 & ~n16518 ;
  assign n16537 = n16536 ^ n16523 ;
  assign n16538 = ~n16481 & ~n16537 ;
  assign n16543 = n16542 ^ n16538 ;
  assign n16544 = n16543 ^ x96 ;
  assign n14678 = n14677 ^ x116 ;
  assign n14679 = n14409 ^ x102 ;
  assign n15080 = n14678 & n14679 ;
  assign n15081 = n15080 ^ n14679 ;
  assign n15082 = n15081 ^ n14678 ;
  assign n14802 = n14801 ^ x117 ;
  assign n14833 = n13681 & n13847 ;
  assign n14825 = n13888 ^ n13868 ;
  assign n14826 = n14825 ^ n13680 ;
  assign n14827 = n14826 ^ n13897 ;
  assign n14828 = ~n13861 & ~n14827 ;
  assign n14829 = n14828 ^ n13680 ;
  assign n14830 = n13886 ^ n13861 ;
  assign n14831 = ~n14829 & ~n14830 ;
  assign n14820 = n14819 ^ n13928 ;
  assign n14821 = n14820 ^ n13894 ;
  assign n14810 = n13840 ^ n13835 ;
  assign n14811 = n14810 ^ n13873 ;
  assign n14812 = n13873 ^ n13647 ;
  assign n14813 = n14812 ^ n13873 ;
  assign n14814 = n14811 & n14813 ;
  assign n14815 = n14814 ^ n13873 ;
  assign n14816 = n13842 & ~n14815 ;
  assign n14822 = n14821 ^ n14816 ;
  assign n14808 = n14807 ^ n13833 ;
  assign n14809 = n13680 & n14808 ;
  assign n14823 = n14822 ^ n14809 ;
  assign n14824 = n14823 ^ n13886 ;
  assign n14832 = n14831 ^ n14824 ;
  assign n14834 = n14833 ^ n14832 ;
  assign n14835 = ~n13860 & ~n14834 ;
  assign n14838 = n13835 ^ n13679 ;
  assign n14839 = n14838 ^ n13835 ;
  assign n14840 = n13836 & ~n14839 ;
  assign n14841 = n14840 ^ n13835 ;
  assign n14842 = n13647 & n14841 ;
  assign n14843 = n14835 & ~n14842 ;
  assign n14844 = ~n14806 & n14843 ;
  assign n14845 = ~n14804 & n14844 ;
  assign n14846 = n14845 ^ n12129 ;
  assign n14847 = n14846 ^ x84 ;
  assign n14848 = n14802 & ~n14847 ;
  assign n14852 = n14609 ^ x77 ;
  assign n14996 = n14853 & n14946 ;
  assign n14997 = n14996 ^ n14945 ;
  assign n14998 = n14997 ^ n14931 ;
  assign n14999 = n14998 ^ n14997 ;
  assign n15000 = n14997 ^ n14854 ;
  assign n15001 = n15000 ^ n14997 ;
  assign n15002 = n14999 & n15001 ;
  assign n15003 = n15002 ^ n14997 ;
  assign n15004 = ~n14977 & n15003 ;
  assign n15005 = n15004 ^ n14997 ;
  assign n14988 = n14981 ^ n14959 ;
  assign n14989 = n14959 ^ n14853 ;
  assign n14990 = n14989 ^ n14959 ;
  assign n14991 = n14988 & n14990 ;
  assign n14992 = n14991 ^ n14959 ;
  assign n14993 = n14977 & n14992 ;
  assign n14994 = n14993 ^ n14987 ;
  assign n14964 = n14963 ^ n14922 ;
  assign n14962 = n14961 ^ n14942 ;
  assign n14965 = n14964 ^ n14962 ;
  assign n14957 = n14949 ^ n14926 ;
  assign n14958 = n14957 ^ n14934 ;
  assign n14966 = n14965 ^ n14958 ;
  assign n14967 = n14853 & n14966 ;
  assign n14968 = n14967 ^ n14965 ;
  assign n14995 = n14994 ^ n14968 ;
  assign n15006 = n15005 ^ n14995 ;
  assign n15007 = n15006 ^ n14976 ;
  assign n15008 = n15007 ^ n12083 ;
  assign n14955 = n14941 ^ n14935 ;
  assign n14956 = n14955 ^ n14934 ;
  assign n14969 = n14968 ^ n14956 ;
  assign n14970 = n14854 & n14969 ;
  assign n15009 = n15008 ^ n14970 ;
  assign n14936 = n14935 ^ n14934 ;
  assign n14953 = n14952 ^ n14936 ;
  assign n14954 = n14857 & ~n14953 ;
  assign n15010 = n15009 ^ n14954 ;
  assign n15011 = n15010 ^ x67 ;
  assign n15012 = ~n14852 & n15011 ;
  assign n15015 = n15012 ^ n15011 ;
  assign n15017 = n15015 ^ n14852 ;
  assign n15025 = n15017 ^ n15011 ;
  assign n15026 = n14848 & ~n15025 ;
  assign n14849 = n14848 ^ n14802 ;
  assign n14850 = n14849 ^ n14847 ;
  assign n14851 = n14850 ^ n14802 ;
  assign n15013 = ~n14851 & n15012 ;
  assign n15083 = n15026 ^ n15013 ;
  assign n15084 = ~n15082 & n15083 ;
  assign n15021 = n14848 & n15015 ;
  assign n15016 = ~n14851 & n15015 ;
  assign n15022 = n15021 ^ n15016 ;
  assign n15075 = n15016 ^ n14679 ;
  assign n15076 = n15075 ^ n15016 ;
  assign n15077 = n15022 & ~n15076 ;
  assign n15078 = n15077 ^ n15016 ;
  assign n15079 = n14678 & n15078 ;
  assign n15085 = n15084 ^ n15079 ;
  assign n15023 = n14850 & n15012 ;
  assign n16545 = n15023 & ~n15082 ;
  assign n15027 = n14849 & ~n15025 ;
  assign n15018 = ~n14851 & n15017 ;
  assign n15019 = n15018 ^ n15016 ;
  assign n15014 = n15013 ^ n14851 ;
  assign n15020 = n15019 ^ n15014 ;
  assign n15028 = n15027 ^ n15020 ;
  assign n15029 = n15028 ^ n15026 ;
  assign n15030 = n15029 ^ n15025 ;
  assign n15024 = n14850 & n15017 ;
  assign n15031 = n15030 ^ n15024 ;
  assign n16546 = n15031 ^ n15030 ;
  assign n16547 = n15030 ^ n14678 ;
  assign n16548 = n16547 ^ n15030 ;
  assign n16549 = n16546 & n16548 ;
  assign n16550 = n16549 ^ n15030 ;
  assign n16551 = ~n14679 & n16550 ;
  assign n16552 = n16551 ^ n15030 ;
  assign n16564 = n15029 ^ n15023 ;
  assign n15045 = n14849 & n15017 ;
  assign n15032 = n15031 ^ n14850 ;
  assign n15033 = n15032 ^ n15023 ;
  assign n15034 = n15033 ^ n15015 ;
  assign n15035 = n15034 ^ n15022 ;
  assign n15036 = n15035 ^ n15024 ;
  assign n15046 = n15045 ^ n15036 ;
  assign n15047 = n15046 ^ n15018 ;
  assign n15042 = n15021 ^ n15018 ;
  assign n15043 = n15042 ^ n15027 ;
  assign n15044 = n15043 ^ n15024 ;
  assign n15048 = n15047 ^ n15044 ;
  assign n15040 = n15021 ^ n14848 ;
  assign n15041 = n15040 ^ n14802 ;
  assign n15049 = n15048 ^ n15041 ;
  assign n16565 = n16564 ^ n15049 ;
  assign n16566 = n16565 ^ n15021 ;
  assign n16567 = n16566 ^ n15029 ;
  assign n16568 = n16567 ^ n16565 ;
  assign n16569 = n16565 ^ n14678 ;
  assign n16570 = n16569 ^ n16565 ;
  assign n16571 = ~n16568 & ~n16570 ;
  assign n16572 = n16571 ^ n16565 ;
  assign n16573 = ~n14679 & ~n16572 ;
  assign n16574 = n16573 ^ n15023 ;
  assign n16561 = n15035 ^ n15033 ;
  assign n16560 = n15042 ^ n15028 ;
  assign n16562 = n16561 ^ n16560 ;
  assign n16563 = n15081 & ~n16562 ;
  assign n16575 = n16574 ^ n16563 ;
  assign n14680 = n14679 ^ n14678 ;
  assign n15050 = n15049 ^ n15013 ;
  assign n15039 = n15023 ^ n15012 ;
  assign n15051 = n15050 ^ n15039 ;
  assign n15056 = n15051 ^ n15026 ;
  assign n15057 = n15056 ^ n15040 ;
  assign n15087 = n15057 ^ n15033 ;
  assign n16559 = ~n14680 & n15087 ;
  assign n16576 = n16575 ^ n16559 ;
  assign n16553 = n15019 ^ n15013 ;
  assign n16554 = n16553 ^ n15045 ;
  assign n16555 = n16554 ^ n15051 ;
  assign n16556 = n14679 & n16555 ;
  assign n16557 = n16556 ^ n15019 ;
  assign n16558 = n14678 & n16557 ;
  assign n16577 = n16576 ^ n16558 ;
  assign n15086 = n15030 & ~n15082 ;
  assign n16578 = n16577 ^ n15086 ;
  assign n16579 = ~n16552 & ~n16578 ;
  assign n16580 = ~n16545 & n16579 ;
  assign n16581 = ~n15085 & n16580 ;
  assign n16582 = n16581 ^ n14491 ;
  assign n16583 = n16582 ^ x122 ;
  assign n16584 = n16544 & ~n16583 ;
  assign n16680 = n16584 ^ n16583 ;
  assign n16711 = n16680 ^ n16544 ;
  assign n16721 = n16588 & n16711 ;
  assign n18866 = n16704 & n16721 ;
  assign n19225 = n18866 ^ n14609 ;
  assign n16589 = n16588 ^ n16385 ;
  assign n16716 = ~n16589 & n16711 ;
  assign n16684 = n16584 & ~n16589 ;
  assign n16707 = n16684 ^ n16584 ;
  assign n16705 = n16584 & n16588 ;
  assign n16682 = n16386 & n16584 ;
  assign n16706 = n16705 ^ n16682 ;
  assign n16708 = n16707 ^ n16706 ;
  assign n16717 = n16716 ^ n16708 ;
  assign n16591 = n16589 ^ n16193 ;
  assign n16715 = n16591 & n16711 ;
  assign n16718 = n16717 ^ n16715 ;
  assign n18868 = ~n16638 & n16718 ;
  assign n18869 = n18868 ^ n16715 ;
  assign n18872 = n18869 ^ n16705 ;
  assign n18873 = n18872 ^ n18869 ;
  assign n18874 = ~n16638 & n18873 ;
  assign n18875 = n18874 ^ n18869 ;
  assign n18876 = ~n16678 & n18875 ;
  assign n18877 = n18876 ^ n18869 ;
  assign n16585 = n16584 ^ n16544 ;
  assign n16592 = n16585 & n16591 ;
  assign n16590 = n16585 & ~n16589 ;
  assign n16593 = n16592 ^ n16590 ;
  assign n16754 = n16678 ^ n16592 ;
  assign n16755 = n16754 ^ n16592 ;
  assign n16756 = n16593 & n16755 ;
  assign n16757 = n16756 ^ n16592 ;
  assign n16758 = ~n16638 & n16757 ;
  assign n16681 = n16386 & ~n16680 ;
  assign n16683 = n16682 ^ n16681 ;
  assign n19217 = n16683 ^ n16593 ;
  assign n19211 = n16721 ^ n16705 ;
  assign n19212 = n16721 ^ n16638 ;
  assign n19213 = n19212 ^ n16721 ;
  assign n19214 = n19211 & n19213 ;
  assign n19215 = n19214 ^ n16721 ;
  assign n19216 = n16678 & n19215 ;
  assign n19218 = n19217 ^ n19216 ;
  assign n16586 = n16386 & n16585 ;
  assign n16587 = n16586 ^ n16585 ;
  assign n16594 = n16593 ^ n16587 ;
  assign n19208 = n16684 ^ n16594 ;
  assign n16693 = n16588 & ~n16680 ;
  assign n19204 = n16693 ^ n16586 ;
  assign n16694 = ~n16589 & ~n16680 ;
  assign n16709 = n16708 ^ n16694 ;
  assign n19203 = n16709 ^ n16684 ;
  assign n19205 = n19204 ^ n19203 ;
  assign n16712 = n16386 & n16711 ;
  assign n19206 = n19205 ^ n16712 ;
  assign n19207 = ~n16638 & n19206 ;
  assign n19209 = n19208 ^ n19207 ;
  assign n19210 = ~n16678 & n19209 ;
  assign n19219 = n19218 ^ n19210 ;
  assign n19200 = n16678 & n16705 ;
  assign n19201 = n19200 ^ n16593 ;
  assign n19202 = ~n16638 & n19201 ;
  assign n19220 = n19219 ^ n19202 ;
  assign n16679 = n16678 ^ n16638 ;
  assign n18881 = n16682 ^ n16586 ;
  assign n19191 = n16683 ^ n16638 ;
  assign n19192 = n19191 ^ n16683 ;
  assign n19193 = n18881 & n19192 ;
  assign n19194 = n19193 ^ n16683 ;
  assign n19195 = ~n16679 & n19194 ;
  assign n19221 = n19220 ^ n19195 ;
  assign n19222 = ~n16758 & ~n19221 ;
  assign n16749 = n16679 & n16715 ;
  assign n16695 = n16694 ^ n16693 ;
  assign n16692 = n16681 ^ n16680 ;
  assign n16696 = n16695 ^ n16692 ;
  assign n16743 = n16696 ^ n16693 ;
  assign n16744 = n16693 ^ n16678 ;
  assign n16745 = n16744 ^ n16693 ;
  assign n16746 = ~n16743 & n16745 ;
  assign n16747 = n16746 ^ n16693 ;
  assign n16748 = n16638 & n16747 ;
  assign n16750 = n16749 ^ n16748 ;
  assign n19223 = n19222 ^ n16750 ;
  assign n19224 = ~n18877 & n19223 ;
  assign n19226 = n19225 ^ n19224 ;
  assign n19227 = n19226 ^ x123 ;
  assign n15707 = n15706 ^ x113 ;
  assign n15724 = n14949 ^ n14928 ;
  assign n15725 = n15724 ^ n14924 ;
  assign n15726 = n15725 ^ n15323 ;
  assign n15727 = ~n14856 & ~n15726 ;
  assign n15728 = n15727 ^ n15323 ;
  assign n15730 = n15321 ^ n14854 ;
  assign n15729 = n14938 ^ n14855 ;
  assign n15731 = n15730 ^ n15729 ;
  assign n15732 = n15731 ^ n15321 ;
  assign n15733 = n15728 & ~n15732 ;
  assign n15734 = n15733 ^ n15730 ;
  assign n15735 = n15734 ^ n15723 ;
  assign n15736 = n15735 ^ n14993 ;
  assign n15737 = n15736 ^ n15328 ;
  assign n15738 = n15737 ^ n15005 ;
  assign n15739 = n15738 ^ n14976 ;
  assign n15740 = n15739 ^ n12973 ;
  assign n15708 = n14942 ^ n14855 ;
  assign n15709 = n14941 ^ n14857 ;
  assign n15710 = n14942 ^ n14857 ;
  assign n15711 = n15710 ^ n14857 ;
  assign n15712 = ~n15709 & ~n15711 ;
  assign n15713 = n15712 ^ n14857 ;
  assign n15714 = n15708 & n15713 ;
  assign n15741 = n15740 ^ n15714 ;
  assign n15742 = n15741 ^ x74 ;
  assign n15743 = n15707 & n15742 ;
  assign n15745 = n15141 ^ n15136 ;
  assign n15746 = n14681 & n15745 ;
  assign n15747 = n15746 ^ n15141 ;
  assign n15750 = n15747 ^ n14772 ;
  assign n15749 = n15747 ^ n14761 ;
  assign n15751 = n15750 ^ n15749 ;
  assign n15752 = n15750 ^ n14681 ;
  assign n15753 = n15752 ^ n15750 ;
  assign n15754 = n15751 & ~n15753 ;
  assign n15755 = n15754 ^ n15750 ;
  assign n15756 = n14682 & ~n15755 ;
  assign n15748 = n15747 ^ n12932 ;
  assign n15757 = n15756 ^ n15748 ;
  assign n15758 = n15757 ^ x104 ;
  assign n15759 = n13146 ^ x122 ;
  assign n15760 = ~n15758 & n15759 ;
  assign n15763 = n15760 ^ n15759 ;
  assign n15764 = n15763 ^ n15758 ;
  assign n15778 = n15743 & n15764 ;
  assign n16852 = n15778 ^ n15743 ;
  assign n15822 = n15764 ^ n15759 ;
  assign n15823 = n15743 & ~n15822 ;
  assign n15783 = n15759 ^ n15742 ;
  assign n15801 = n15758 & ~n15783 ;
  assign n15802 = n15801 ^ n15742 ;
  assign n15803 = n15707 & n15802 ;
  assign n15804 = n15803 ^ n15743 ;
  assign n15784 = ~n15707 & n15783 ;
  assign n15786 = n15758 ^ n15742 ;
  assign n15787 = n15786 ^ n15759 ;
  assign n15788 = n15787 ^ n15707 ;
  assign n15789 = n15784 & n15788 ;
  assign n15744 = n15743 ^ n15742 ;
  assign n15762 = n15744 ^ n15707 ;
  assign n15767 = ~n15758 & ~n15762 ;
  assign n15781 = ~n15759 & n15767 ;
  assign n15782 = n15781 ^ n15767 ;
  assign n15790 = n15789 ^ n15782 ;
  assign n15765 = ~n15762 & n15764 ;
  assign n15766 = n15765 ^ n15762 ;
  assign n15768 = n15767 ^ n15766 ;
  assign n15791 = n15790 ^ n15768 ;
  assign n15785 = n15784 ^ n15782 ;
  assign n15792 = n15791 ^ n15785 ;
  assign n15793 = n15792 ^ n15768 ;
  assign n15761 = n15744 & n15760 ;
  assign n15794 = n15793 ^ n15761 ;
  assign n15779 = n15765 ^ n15761 ;
  assign n15780 = n15779 ^ n15778 ;
  assign n15795 = n15794 ^ n15780 ;
  assign n15777 = n15768 ^ n15764 ;
  assign n15796 = n15795 ^ n15777 ;
  assign n15805 = n15804 ^ n15796 ;
  assign n15824 = n15823 ^ n15805 ;
  assign n16853 = n16852 ^ n15824 ;
  assign n16826 = n15796 ^ n15791 ;
  assign n17811 = n16853 ^ n16826 ;
  assign n15806 = n15791 ^ n15744 ;
  assign n15807 = n15806 ^ n15794 ;
  assign n15808 = n15807 ^ n15792 ;
  assign n15809 = n15808 ^ n15805 ;
  assign n15810 = n15809 ^ n15763 ;
  assign n15811 = n15810 ^ n15793 ;
  assign n15775 = n15762 ^ n15742 ;
  assign n15812 = n15811 ^ n15775 ;
  assign n15776 = n15760 & n15775 ;
  assign n15797 = n15796 ^ n15776 ;
  assign n15813 = n15812 ^ n15797 ;
  assign n17821 = n17811 ^ n15813 ;
  assign n15685 = n13938 ^ x107 ;
  assign n15684 = n15683 ^ x81 ;
  assign n17594 = ~n15684 & ~n15809 ;
  assign n17595 = n17594 ^ n15805 ;
  assign n17598 = n17595 ^ n15776 ;
  assign n17599 = n17598 ^ n17595 ;
  assign n17600 = n15684 & n17599 ;
  assign n17601 = n17600 ^ n17595 ;
  assign n17602 = n15685 & ~n17601 ;
  assign n17603 = n17602 ^ n17595 ;
  assign n16835 = n15781 ^ n15776 ;
  assign n16836 = n15781 ^ n15685 ;
  assign n16837 = n16836 ^ n15781 ;
  assign n16838 = n16835 & ~n16837 ;
  assign n16839 = n16838 ^ n15781 ;
  assign n16840 = ~n15684 & n16839 ;
  assign n17820 = n17603 ^ n16840 ;
  assign n17822 = n17821 ^ n17820 ;
  assign n15831 = n15684 & ~n15685 ;
  assign n16844 = n15781 & n15831 ;
  assign n15825 = n15824 ^ n15781 ;
  assign n15826 = n15781 ^ n15684 ;
  assign n15827 = n15826 ^ n15781 ;
  assign n15828 = ~n15825 & ~n15827 ;
  assign n15829 = n15828 ^ n15781 ;
  assign n15830 = n15685 & n15829 ;
  assign n16845 = n16844 ^ n15830 ;
  assign n17823 = n17822 ^ n16845 ;
  assign n15686 = n15685 ^ n15684 ;
  assign n17812 = n17811 ^ n15794 ;
  assign n17813 = n17812 ^ n15795 ;
  assign n17814 = n17813 ^ n17812 ;
  assign n17815 = n17812 ^ n15684 ;
  assign n17816 = n17815 ^ n17812 ;
  assign n17817 = n17814 & ~n17816 ;
  assign n17818 = n17817 ^ n17812 ;
  assign n17819 = n15686 & ~n17818 ;
  assign n17824 = n17823 ^ n17819 ;
  assign n17803 = n15797 ^ n15775 ;
  assign n17804 = n17803 ^ n15684 ;
  assign n17805 = n17804 ^ n17803 ;
  assign n17806 = n17803 ^ n15807 ;
  assign n17807 = n17806 ^ n17803 ;
  assign n17808 = n17805 & ~n17807 ;
  assign n17809 = n17808 ^ n17803 ;
  assign n17810 = n15685 & ~n17809 ;
  assign n17825 = n17824 ^ n17810 ;
  assign n15832 = n15831 ^ n15685 ;
  assign n15833 = n15832 ^ n15684 ;
  assign n15834 = n15782 & n15833 ;
  assign n17826 = n17825 ^ n15834 ;
  assign n15837 = ~n15797 & n15831 ;
  assign n17827 = n17826 ^ n15837 ;
  assign n17828 = n17827 ^ n13710 ;
  assign n17829 = n17828 ^ x64 ;
  assign n17830 = n16637 ^ x90 ;
  assign n17831 = ~n17829 & ~n17830 ;
  assign n17832 = n17831 ^ n17829 ;
  assign n15577 = ~n15464 & n15568 ;
  assign n17179 = n15637 ^ n15590 ;
  assign n17180 = ~n16642 & n17179 ;
  assign n17181 = n17180 ^ n15590 ;
  assign n17182 = ~n15624 & n17181 ;
  assign n17849 = n16648 ^ n15557 ;
  assign n17168 = n15594 ^ n15574 ;
  assign n15596 = n15587 ^ n15573 ;
  assign n17847 = n17168 ^ n15596 ;
  assign n17848 = ~n15462 & ~n17847 ;
  assign n17850 = n17849 ^ n17848 ;
  assign n17851 = ~n15624 & n17850 ;
  assign n17845 = ~n15464 & ~n15591 ;
  assign n17836 = n15585 ^ n15571 ;
  assign n17837 = n17836 ^ n17168 ;
  assign n17838 = n15420 & ~n17837 ;
  assign n17842 = n17838 ^ n15557 ;
  assign n17839 = n17838 ^ n15570 ;
  assign n17834 = n15584 ^ n15563 ;
  assign n17835 = n15420 & n17834 ;
  assign n17840 = n17839 ^ n17835 ;
  assign n17841 = n15462 & n17840 ;
  assign n17843 = n17842 ^ n17841 ;
  assign n17844 = n17843 ^ n16648 ;
  assign n17846 = n17845 ^ n17844 ;
  assign n17852 = n17851 ^ n17846 ;
  assign n17833 = n15463 & n15568 ;
  assign n17853 = n17852 ^ n17833 ;
  assign n17854 = ~n17182 & ~n17853 ;
  assign n17855 = ~n16640 & n17854 ;
  assign n17856 = ~n15621 & n17855 ;
  assign n17857 = ~n15577 & n17856 ;
  assign n17858 = n17857 ^ n13819 ;
  assign n17859 = n17858 ^ x107 ;
  assign n17369 = n15085 ^ n13784 ;
  assign n17370 = n17369 ^ n16545 ;
  assign n17357 = n15026 ^ n15023 ;
  assign n17358 = n15080 & n17357 ;
  assign n17345 = n15027 ^ n15019 ;
  assign n17346 = n17345 ^ n15087 ;
  assign n17347 = ~n14678 & n17346 ;
  assign n17348 = n17347 ^ n15044 ;
  assign n17349 = n17348 ^ n15048 ;
  assign n17350 = n17349 ^ n17348 ;
  assign n17353 = n14678 & n17350 ;
  assign n17354 = n17353 ^ n17348 ;
  assign n17355 = ~n14680 & n17354 ;
  assign n17356 = n17355 ^ n17347 ;
  assign n17359 = n17358 ^ n17356 ;
  assign n17339 = n15020 ^ n14850 ;
  assign n17340 = n17339 ^ n15031 ;
  assign n17341 = n17340 ^ n15049 ;
  assign n17342 = n14678 & ~n17341 ;
  assign n17343 = n17342 ^ n15051 ;
  assign n17344 = ~n14679 & n17343 ;
  assign n17360 = n17359 ^ n17344 ;
  assign n17361 = ~n16552 & ~n17360 ;
  assign n17362 = n15050 ^ n15045 ;
  assign n17363 = n15045 ^ n14678 ;
  assign n17364 = n17363 ^ n15045 ;
  assign n17365 = n17362 & ~n17364 ;
  assign n17366 = n17365 ^ n15045 ;
  assign n17367 = n14680 & n17366 ;
  assign n17368 = n17361 & ~n17367 ;
  assign n17371 = n17370 ^ n17368 ;
  assign n17860 = n17371 ^ x81 ;
  assign n17861 = ~n17859 & n17860 ;
  assign n17862 = n17861 ^ n17860 ;
  assign n17863 = n17862 ^ n17859 ;
  assign n17864 = n17863 ^ n17860 ;
  assign n17865 = ~n17832 & ~n17864 ;
  assign n15862 = n13647 & n13834 ;
  assign n15863 = n15862 ^ n13833 ;
  assign n15881 = n15863 ^ n13887 ;
  assign n15882 = n15881 ^ n13868 ;
  assign n15883 = n15882 ^ n13886 ;
  assign n15884 = n15883 ^ n15863 ;
  assign n15885 = n13647 & ~n15884 ;
  assign n15886 = n15885 ^ n15881 ;
  assign n15887 = n13842 & ~n15886 ;
  assign n15864 = n15102 ^ n13868 ;
  assign n15865 = n13647 & n15864 ;
  assign n15866 = n15865 ^ n13868 ;
  assign n15872 = n15866 ^ n13876 ;
  assign n15873 = n15872 ^ n13883 ;
  assign n15874 = n15873 ^ n13841 ;
  assign n15867 = n15866 ^ n13828 ;
  assign n15868 = n15867 ^ n13847 ;
  assign n15869 = n13878 & n15868 ;
  assign n15870 = n15869 ^ n13847 ;
  assign n15871 = n13842 & n15870 ;
  assign n15875 = n15874 ^ n15871 ;
  assign n15876 = n15875 ^ n15863 ;
  assign n15877 = n15876 ^ n14842 ;
  assign n15878 = n15877 ^ n13411 ;
  assign n15860 = n13888 ^ n13828 ;
  assign n15861 = ~n13842 & ~n15860 ;
  assign n15879 = n15878 ^ n15861 ;
  assign n15858 = n13835 ^ n13825 ;
  assign n15859 = ~n13647 & n15858 ;
  assign n15880 = n15879 ^ n15859 ;
  assign n15888 = n15887 ^ n15880 ;
  assign n15889 = n15888 ^ x112 ;
  assign n15925 = n15924 ^ x98 ;
  assign n15926 = n15889 & ~n15925 ;
  assign n15943 = n14161 ^ n14150 ;
  assign n15944 = n14191 & ~n15943 ;
  assign n15937 = n14157 ^ n14141 ;
  assign n15938 = n15937 ^ n14135 ;
  assign n15939 = n15938 ^ n14177 ;
  assign n15935 = n14170 ^ n14141 ;
  assign n15936 = ~n14010 & ~n15935 ;
  assign n15940 = n15939 ^ n15936 ;
  assign n15941 = n14011 & ~n15940 ;
  assign n15942 = n15941 ^ n14157 ;
  assign n15945 = n15944 ^ n15942 ;
  assign n15951 = ~n14155 & n14192 ;
  assign n15952 = ~n15945 & n15951 ;
  assign n15946 = n15945 ^ n15665 ;
  assign n15934 = n14181 ^ n14178 ;
  assign n15947 = n15946 ^ n15934 ;
  assign n15948 = n15947 ^ n15492 ;
  assign n15949 = n15948 ^ n13370 ;
  assign n15929 = n14166 ^ n14010 ;
  assign n15930 = n15929 ^ n14166 ;
  assign n15931 = n14173 & ~n15930 ;
  assign n15932 = n15931 ^ n14166 ;
  assign n15933 = ~n13975 & n15932 ;
  assign n15950 = n15949 ^ n15933 ;
  assign n15953 = n15952 ^ n15950 ;
  assign n15954 = n15953 ^ x73 ;
  assign n15955 = n15151 ^ x64 ;
  assign n15956 = n15954 & n15955 ;
  assign n15957 = n15956 ^ n15955 ;
  assign n15974 = n15926 & n15957 ;
  assign n16026 = n16025 ^ x66 ;
  assign n15958 = n15957 ^ n15954 ;
  assign n16033 = n15926 & ~n15958 ;
  assign n15973 = ~n15889 & n15957 ;
  assign n15975 = n15974 ^ n15973 ;
  assign n15962 = n15926 ^ n15925 ;
  assign n15963 = n15962 ^ n15889 ;
  assign n15964 = n15963 ^ n15925 ;
  assign n15967 = n15964 ^ n15954 ;
  assign n15984 = n15975 ^ n15967 ;
  assign n15968 = ~n15955 & ~n15967 ;
  assign n15985 = n15984 ^ n15968 ;
  assign n16034 = n16033 ^ n15985 ;
  assign n15857 = n15281 ^ x88 ;
  assign n16035 = n15985 ^ n15857 ;
  assign n16036 = n16035 ^ n15985 ;
  assign n16037 = ~n16034 & ~n16036 ;
  assign n16038 = n16037 ^ n15985 ;
  assign n16039 = n16026 & ~n16038 ;
  assign n15965 = ~n15958 & n15964 ;
  assign n17206 = n15965 ^ n15926 ;
  assign n15976 = n15955 ^ n15954 ;
  assign n15977 = n15976 ^ n15889 ;
  assign n15978 = n15977 ^ n15925 ;
  assign n15979 = n15967 & ~n15978 ;
  assign n16072 = n15979 ^ n15955 ;
  assign n15970 = n15925 ^ n15889 ;
  assign n15982 = n15957 & n15970 ;
  assign n15983 = n15982 ^ n15975 ;
  assign n15986 = n15985 ^ n15983 ;
  assign n15980 = n15979 ^ n15975 ;
  assign n15981 = n15980 ^ n15978 ;
  assign n15987 = n15986 ^ n15981 ;
  assign n15971 = n15970 ^ n15954 ;
  assign n15972 = ~n15955 & n15971 ;
  assign n15988 = n15987 ^ n15972 ;
  assign n16073 = n16072 ^ n15988 ;
  assign n17207 = n17206 ^ n16073 ;
  assign n15989 = n15988 ^ n15968 ;
  assign n15966 = n15965 ^ n15958 ;
  assign n15969 = n15968 ^ n15966 ;
  assign n15990 = n15989 ^ n15969 ;
  assign n17202 = n15990 ^ n15965 ;
  assign n16029 = n15926 & n15956 ;
  assign n16030 = n16029 ^ n15982 ;
  assign n17203 = n17202 ^ n16030 ;
  assign n16063 = n15975 ^ n15957 ;
  assign n16074 = n16073 ^ n16063 ;
  assign n17204 = n17203 ^ n16074 ;
  assign n15959 = n15958 ^ n15955 ;
  assign n15960 = n15926 & n15959 ;
  assign n17205 = n17204 ^ n15960 ;
  assign n17208 = n17207 ^ n17205 ;
  assign n17209 = ~n15857 & ~n17208 ;
  assign n17210 = n17209 ^ n15965 ;
  assign n17211 = ~n16026 & n17210 ;
  assign n17212 = n17211 ^ n15965 ;
  assign n16027 = ~n15857 & ~n16026 ;
  assign n16028 = n16027 ^ n16026 ;
  assign n16064 = n16063 ^ n15983 ;
  assign n16067 = n16064 ^ n16029 ;
  assign n17226 = ~n16028 & n16067 ;
  assign n15961 = n15960 ^ n15959 ;
  assign n15991 = n15990 ^ n15961 ;
  assign n17216 = n15991 ^ n15986 ;
  assign n17213 = n16033 ^ n15980 ;
  assign n17214 = n17213 ^ n16067 ;
  assign n17215 = n15857 & ~n17214 ;
  assign n17217 = n17216 ^ n17215 ;
  assign n17218 = n16026 & n17217 ;
  assign n17219 = n17218 ^ n15991 ;
  assign n16065 = n16027 ^ n15857 ;
  assign n16080 = n16065 ^ n16028 ;
  assign n17220 = n16080 ^ n16073 ;
  assign n16041 = n16033 ^ n15987 ;
  assign n16081 = n16041 ^ n15966 ;
  assign n17221 = n16081 ^ n15960 ;
  assign n17222 = n17221 ^ n16073 ;
  assign n17223 = ~n17220 & n17222 ;
  assign n17224 = n17223 ^ n16073 ;
  assign n17225 = n17219 & n17224 ;
  assign n17227 = n17226 ^ n17225 ;
  assign n17228 = ~n17212 & n17227 ;
  assign n16892 = n16027 & n16029 ;
  assign n17229 = n17228 ^ n16892 ;
  assign n17230 = ~n16039 & n17229 ;
  assign n17231 = ~n15974 & n17230 ;
  assign n17232 = n17231 ^ n13678 ;
  assign n17866 = n17232 ^ x104 ;
  assign n17867 = n16384 ^ x66 ;
  assign n17868 = n17866 & n17867 ;
  assign n17869 = n17868 ^ n17866 ;
  assign n17870 = n17869 ^ n17867 ;
  assign n17871 = n17870 ^ n17866 ;
  assign n17872 = n17865 & n17871 ;
  assign n17874 = n17832 ^ n17830 ;
  assign n17875 = n17863 & ~n17874 ;
  assign n17873 = ~n17832 & n17861 ;
  assign n17876 = n17875 ^ n17873 ;
  assign n17877 = n17869 & n17876 ;
  assign n17878 = ~n17864 & ~n17874 ;
  assign n17887 = n17878 ^ n17874 ;
  assign n17885 = n17861 & ~n17874 ;
  assign n17886 = n17885 ^ n17875 ;
  assign n17888 = n17887 ^ n17886 ;
  assign n17889 = n17888 ^ n17878 ;
  assign n17890 = n17889 ^ n17865 ;
  assign n17891 = n17890 ^ n17886 ;
  assign n17881 = n17864 ^ n17830 ;
  assign n17882 = n17829 & ~n17881 ;
  assign n17880 = n17860 ^ n17859 ;
  assign n17883 = n17882 ^ n17880 ;
  assign n17884 = n17883 ^ n17862 ;
  assign n17892 = n17891 ^ n17884 ;
  assign n17893 = ~n17870 & n17892 ;
  assign n17879 = n17871 & n17878 ;
  assign n17894 = n17893 ^ n17879 ;
  assign n17895 = n17871 ^ n17869 ;
  assign n17936 = n17887 ^ n17882 ;
  assign n17907 = n17831 & n17862 ;
  assign n17906 = n17831 & n17863 ;
  assign n17908 = n17907 ^ n17906 ;
  assign n17909 = n17908 ^ n17892 ;
  assign n17910 = n17909 ^ n17831 ;
  assign n17937 = n17936 ^ n17910 ;
  assign n17938 = n17937 ^ n17908 ;
  assign n17913 = n17859 ^ n17829 ;
  assign n17914 = n17913 ^ n17860 ;
  assign n17915 = ~n17830 & n17914 ;
  assign n17935 = n17915 ^ n17907 ;
  assign n17939 = n17938 ^ n17935 ;
  assign n17940 = n17939 ^ n17936 ;
  assign n17896 = n17874 ^ n17829 ;
  assign n17897 = n17861 & ~n17896 ;
  assign n17934 = n17897 ^ n17896 ;
  assign n17941 = n17940 ^ n17934 ;
  assign n17924 = ~n17832 & n17862 ;
  assign n17954 = n17941 ^ n17924 ;
  assign n17955 = n17895 & ~n17954 ;
  assign n17926 = n17873 ^ n17865 ;
  assign n17932 = n17867 & n17926 ;
  assign n17933 = n17932 ^ n17865 ;
  assign n17942 = n17941 ^ n17933 ;
  assign n17943 = n17942 ^ n17888 ;
  assign n17925 = n17924 ^ n17832 ;
  assign n17927 = n17926 ^ n17925 ;
  assign n17944 = n17943 ^ n17927 ;
  assign n17945 = n17944 ^ n17933 ;
  assign n17946 = n17867 & ~n17945 ;
  assign n17947 = n17946 ^ n17942 ;
  assign n17948 = ~n17895 & ~n17947 ;
  assign n17949 = n17948 ^ n17933 ;
  assign n17931 = ~n17870 & n17907 ;
  assign n17951 = n17949 ^ n17931 ;
  assign n17928 = n17927 ^ n17885 ;
  assign n17929 = ~n17870 & ~n17928 ;
  assign n17922 = n17906 ^ n17897 ;
  assign n17923 = n17869 & n17922 ;
  assign n17930 = n17929 ^ n17923 ;
  assign n17952 = n17951 ^ n17930 ;
  assign n17912 = n17908 ^ n17897 ;
  assign n17916 = n17915 ^ n17912 ;
  assign n17917 = n17915 ^ n17866 ;
  assign n17918 = n17917 ^ n17915 ;
  assign n17919 = n17916 & ~n17918 ;
  assign n17920 = n17919 ^ n17915 ;
  assign n17921 = n17867 & n17920 ;
  assign n17953 = n17952 ^ n17921 ;
  assign n17956 = n17955 ^ n17953 ;
  assign n17911 = n17869 & n17910 ;
  assign n17957 = n17956 ^ n17911 ;
  assign n17899 = n17885 ^ n17865 ;
  assign n17898 = n17897 ^ n17889 ;
  assign n17900 = n17899 ^ n17898 ;
  assign n17901 = n17899 ^ n17866 ;
  assign n17902 = n17901 ^ n17899 ;
  assign n17903 = ~n17900 & ~n17902 ;
  assign n17904 = n17903 ^ n17899 ;
  assign n17905 = ~n17895 & n17904 ;
  assign n17958 = n17957 ^ n17905 ;
  assign n17959 = ~n17894 & ~n17958 ;
  assign n17960 = ~n17877 & n17959 ;
  assign n17961 = ~n17872 & n17960 ;
  assign n17962 = n17961 ^ n13938 ;
  assign n19160 = n17962 ^ x112 ;
  assign n15372 = n15343 ^ n15152 ;
  assign n15373 = n15372 ^ n15154 ;
  assign n15407 = n15406 ^ n15348 ;
  assign n15411 = n15410 ^ n15407 ;
  assign n15412 = n15410 ^ n15132 ;
  assign n15413 = n15412 ^ n15410 ;
  assign n15414 = ~n15411 & ~n15413 ;
  assign n15415 = n15414 ^ n15410 ;
  assign n15416 = ~n15373 & ~n15415 ;
  assign n15417 = n15416 ^ n14009 ;
  assign n15360 = n15152 & n15357 ;
  assign n15350 = n15349 ^ n15348 ;
  assign n15351 = ~n15152 & n15350 ;
  assign n15352 = n15351 ^ n15349 ;
  assign n15361 = n15360 ^ n15352 ;
  assign n15362 = ~n15132 & n15361 ;
  assign n15363 = n15362 ^ n15352 ;
  assign n15394 = n15393 ^ n15392 ;
  assign n15391 = n15390 ^ n15349 ;
  assign n15395 = n15394 ^ n15391 ;
  assign n15396 = ~n15152 & n15395 ;
  assign n15397 = n15396 ^ n15393 ;
  assign n15389 = n15386 ^ n15348 ;
  assign n15398 = n15397 ^ n15389 ;
  assign n15378 = n15357 ^ n15348 ;
  assign n15380 = n15379 ^ n15378 ;
  assign n15387 = n15386 ^ n15380 ;
  assign n15388 = ~n15152 & ~n15387 ;
  assign n15399 = n15398 ^ n15388 ;
  assign n15400 = ~n15132 & ~n15399 ;
  assign n15401 = n15400 ^ n15397 ;
  assign n15377 = ~n15373 & n15376 ;
  assign n15402 = n15401 ^ n15377 ;
  assign n15370 = n15152 & n15367 ;
  assign n15368 = n15367 ^ n15364 ;
  assign n15369 = n15132 & n15368 ;
  assign n15371 = n15370 ^ n15369 ;
  assign n15403 = n15402 ^ n15371 ;
  assign n15404 = ~n15363 & ~n15403 ;
  assign n15405 = ~n15345 & n15404 ;
  assign n15418 = n15417 ^ n15405 ;
  assign n17456 = n15418 ^ x100 ;
  assign n14612 = n14610 ^ n13147 ;
  assign n14618 = n14412 ^ n14220 ;
  assign n14619 = ~n13939 & ~n14618 ;
  assign n14614 = n14613 ^ n14415 ;
  assign n14615 = n14614 ^ n14417 ;
  assign n14434 = n14433 ^ n14415 ;
  assign n14435 = n14434 ^ n14432 ;
  assign n14429 = n14428 ^ n14426 ;
  assign n14430 = n14429 ^ n14423 ;
  assign n14436 = n14435 ^ n14430 ;
  assign n14437 = n14436 ^ n13940 ;
  assign n14616 = n14615 ^ n14437 ;
  assign n14617 = n14616 ^ n14417 ;
  assign n14620 = n14619 ^ n14617 ;
  assign n14621 = n13147 & ~n14620 ;
  assign n14622 = n14621 ^ n14616 ;
  assign n14438 = n14437 ^ n14430 ;
  assign n14439 = ~n13147 & n14438 ;
  assign n14440 = n14439 ^ n14430 ;
  assign n14623 = n14622 ^ n14440 ;
  assign n14624 = ~n14612 & n14623 ;
  assign n14611 = n14610 ^ n14440 ;
  assign n14625 = n14624 ^ n14611 ;
  assign n14626 = n14625 ^ n14123 ;
  assign n17457 = n14626 ^ x101 ;
  assign n16040 = n16026 ^ n15857 ;
  assign n16042 = n16041 ^ n15968 ;
  assign n16043 = ~n16026 & n16042 ;
  assign n16044 = n16043 ^ n15969 ;
  assign n16045 = n16044 ^ n15991 ;
  assign n16046 = n16045 ^ n16044 ;
  assign n16047 = n16044 ^ n15857 ;
  assign n16048 = n16047 ^ n16044 ;
  assign n16049 = ~n16046 & ~n16048 ;
  assign n16050 = n16049 ^ n16044 ;
  assign n16051 = ~n16040 & ~n16050 ;
  assign n16052 = n16051 ^ n16044 ;
  assign n17461 = ~n15857 & ~n16081 ;
  assign n16054 = n16033 ^ n15965 ;
  assign n17460 = ~n16026 & n16054 ;
  assign n17462 = n17461 ^ n17460 ;
  assign n17482 = n16027 & n16064 ;
  assign n17477 = n16026 & ~n16035 ;
  assign n16066 = n15978 ^ n15972 ;
  assign n16068 = n16067 ^ n16066 ;
  assign n16069 = n16068 ^ n15974 ;
  assign n16070 = n16065 & ~n16069 ;
  assign n17476 = n16070 & n16073 ;
  assign n17478 = n17477 ^ n17476 ;
  assign n17479 = n16040 & n17478 ;
  assign n17480 = n17479 ^ n17477 ;
  assign n17481 = n17480 ^ n16035 ;
  assign n17483 = n17482 ^ n17481 ;
  assign n17470 = n16041 ^ n16029 ;
  assign n17471 = ~n16065 & n17470 ;
  assign n17484 = n17483 ^ n17471 ;
  assign n17463 = n17205 ^ n15960 ;
  assign n17464 = n17463 ^ n15960 ;
  assign n17467 = n16026 & n17464 ;
  assign n17468 = n17467 ^ n15960 ;
  assign n17469 = n15857 & n17468 ;
  assign n17485 = n17484 ^ n17469 ;
  assign n17486 = ~n17462 & n17485 ;
  assign n17487 = n16052 & n17486 ;
  assign n17458 = n16892 ^ n14043 ;
  assign n16884 = n16068 ^ n15983 ;
  assign n16885 = ~n16065 & n16884 ;
  assign n17459 = n17458 ^ n16885 ;
  assign n17488 = n17487 ^ n17459 ;
  assign n17489 = n17488 ^ x124 ;
  assign n17490 = n17457 & n17489 ;
  assign n17491 = n17490 ^ n17457 ;
  assign n17550 = n16340 ^ n14119 ;
  assign n16898 = n16296 & ~n16338 ;
  assign n17251 = n16336 ^ n16329 ;
  assign n17252 = n16335 ^ n16290 ;
  assign n17255 = ~n16336 & n17252 ;
  assign n17256 = n17255 ^ n16290 ;
  assign n17257 = n17251 & n17256 ;
  assign n17258 = n17257 ^ n16329 ;
  assign n17250 = n16302 & ~n16339 ;
  assign n17259 = n17258 ^ n17250 ;
  assign n17542 = n17259 ^ n16311 ;
  assign n17236 = n16336 ^ n16333 ;
  assign n17535 = n16338 & ~n17236 ;
  assign n17536 = n17535 ^ n16333 ;
  assign n17537 = n16382 ^ n16302 ;
  assign n17538 = n17537 ^ n16338 ;
  assign n17539 = n17538 ^ n16382 ;
  assign n17540 = n17536 & ~n17539 ;
  assign n17541 = n17540 ^ n17537 ;
  assign n17543 = n17542 ^ n17541 ;
  assign n17528 = n16382 ^ n16335 ;
  assign n17529 = n17528 ^ n16382 ;
  assign n17530 = n16312 & n17529 ;
  assign n17531 = n17530 ^ n16382 ;
  assign n17532 = ~n16334 & ~n17531 ;
  assign n17544 = n17543 ^ n17532 ;
  assign n17519 = n16381 ^ n16296 ;
  assign n17520 = n17519 ^ n16314 ;
  assign n17523 = ~n16334 & ~n17520 ;
  assign n17524 = n17523 ^ n16314 ;
  assign n17525 = ~n16335 & n17524 ;
  assign n17545 = n17544 ^ n17525 ;
  assign n17517 = n16381 ^ n16311 ;
  assign n17518 = ~n16334 & ~n17517 ;
  assign n17546 = n17545 ^ n17518 ;
  assign n17515 = n16325 ^ n16303 ;
  assign n17516 = ~n16337 & ~n17515 ;
  assign n17547 = n17546 ^ n17516 ;
  assign n17260 = n16321 ^ n16319 ;
  assign n17514 = n16336 & ~n17260 ;
  assign n17548 = n17547 ^ n17514 ;
  assign n17549 = ~n16898 & n17548 ;
  assign n17551 = n17550 ^ n17549 ;
  assign n17552 = n17551 ^ x118 ;
  assign n17502 = n16499 ^ n16470 ;
  assign n16794 = n16472 ^ n16456 ;
  assign n17506 = n17502 ^ n16794 ;
  assign n17503 = n17502 ^ n16497 ;
  assign n17504 = n17503 ^ n16528 ;
  assign n17505 = ~n16387 & n17504 ;
  assign n17507 = n17506 ^ n17505 ;
  assign n17508 = ~n16388 & n17507 ;
  assign n17498 = n16794 ^ n16481 ;
  assign n17318 = n16500 ^ n16460 ;
  assign n17319 = ~n16387 & n17318 ;
  assign n17320 = n17319 ^ n16460 ;
  assign n17321 = n17320 ^ n16468 ;
  assign n17322 = n17321 ^ n17320 ;
  assign n17323 = n17320 ^ n16388 ;
  assign n17324 = n17323 ^ n17320 ;
  assign n17325 = n17322 & n17324 ;
  assign n17326 = n17325 ^ n17320 ;
  assign n17327 = ~n16516 & n17326 ;
  assign n17328 = n17327 ^ n17320 ;
  assign n17499 = n17498 ^ n17328 ;
  assign n16781 = n16460 ^ n16458 ;
  assign n16782 = n16781 ^ n16469 ;
  assign n16783 = n16388 & n16782 ;
  assign n16784 = n16783 ^ n16458 ;
  assign n17313 = n16458 ^ n16388 ;
  assign n17314 = n17313 ^ n16458 ;
  assign n17315 = n16784 & n17314 ;
  assign n17316 = n17315 ^ n16458 ;
  assign n17317 = n16387 & n17316 ;
  assign n17500 = n17499 ^ n17317 ;
  assign n16767 = n16505 ^ n16482 ;
  assign n16768 = n16767 ^ n16505 ;
  assign n16769 = n16505 ^ n16388 ;
  assign n16770 = n16769 ^ n16505 ;
  assign n16771 = n16768 & n16770 ;
  assign n16772 = n16771 ^ n16505 ;
  assign n16773 = ~n16516 & ~n16772 ;
  assign n17501 = n17500 ^ n16773 ;
  assign n17509 = n17508 ^ n17501 ;
  assign n17492 = n16494 ^ n16456 ;
  assign n17493 = n16456 ^ n16388 ;
  assign n17494 = n17493 ^ n16456 ;
  assign n17495 = n17492 & n17494 ;
  assign n17496 = n17495 ^ n16456 ;
  assign n17497 = n16516 & n17496 ;
  assign n17510 = n17509 ^ n17497 ;
  assign n17511 = ~n16541 & ~n17510 ;
  assign n17512 = n17511 ^ n14077 ;
  assign n17513 = n17512 ^ x68 ;
  assign n17563 = n17552 ^ n17513 ;
  assign n17564 = n17491 & n17563 ;
  assign n17553 = ~n17513 & n17552 ;
  assign n17554 = n17553 ^ n17513 ;
  assign n17558 = n17491 ^ n17489 ;
  assign n17559 = ~n17554 & ~n17558 ;
  assign n18618 = n17564 ^ n17559 ;
  assign n17555 = n17554 ^ n17552 ;
  assign n17566 = n17491 & n17555 ;
  assign n17562 = ~n17489 & n17553 ;
  assign n17565 = n17564 ^ n17562 ;
  assign n17567 = n17566 ^ n17565 ;
  assign n17568 = n17567 ^ n17558 ;
  assign n17560 = n17555 & ~n17558 ;
  assign n17561 = n17560 ^ n17559 ;
  assign n17569 = n17568 ^ n17561 ;
  assign n19161 = n18618 ^ n17569 ;
  assign n17622 = n17490 & n17553 ;
  assign n17635 = n17622 ^ n17553 ;
  assign n17636 = n17635 ^ n17562 ;
  assign n17556 = n17555 ^ n17513 ;
  assign n17619 = n17490 & n17556 ;
  assign n17662 = n17636 ^ n17619 ;
  assign n19162 = n19161 ^ n17662 ;
  assign n19163 = n19162 ^ n17560 ;
  assign n17653 = n17622 ^ n17619 ;
  assign n17654 = n17653 ^ n17490 ;
  assign n17629 = n17490 & n17555 ;
  assign n17655 = n17654 ^ n17629 ;
  assign n17630 = n17558 ^ n17457 ;
  assign n17632 = n17555 & n17630 ;
  assign n17681 = n17655 ^ n17632 ;
  assign n17620 = n17619 ^ n17556 ;
  assign n17557 = n17491 & n17556 ;
  assign n17570 = n17569 ^ n17557 ;
  assign n17621 = n17620 ^ n17570 ;
  assign n17623 = n17622 ^ n17621 ;
  assign n17637 = n17636 ^ n17623 ;
  assign n17633 = n17632 ^ n17622 ;
  assign n17634 = n17633 ^ n17629 ;
  assign n17638 = n17637 ^ n17634 ;
  assign n17631 = n17630 ^ n17629 ;
  assign n17639 = n17638 ^ n17631 ;
  assign n17682 = n17681 ^ n17639 ;
  assign n17683 = n17682 ^ n17562 ;
  assign n17684 = n17683 ^ n17619 ;
  assign n19164 = n19163 ^ n17684 ;
  assign n19165 = n17456 & n19164 ;
  assign n19166 = n19165 ^ n19162 ;
  assign n17611 = n15834 ^ n13974 ;
  assign n16841 = ~n15686 & ~n15811 ;
  assign n16842 = n16841 ^ n16840 ;
  assign n17606 = n15793 & n15833 ;
  assign n16814 = n15807 ^ n15790 ;
  assign n16815 = n16814 ^ n15813 ;
  assign n17582 = n16815 ^ n15765 ;
  assign n17580 = n15778 ^ n15767 ;
  assign n17581 = n17580 ^ n16826 ;
  assign n17583 = n17582 ^ n17581 ;
  assign n17584 = ~n15685 & ~n17583 ;
  assign n17585 = n17584 ^ n17582 ;
  assign n17604 = n17603 ^ n17585 ;
  assign n17587 = n17585 ^ n15779 ;
  assign n17586 = n17585 ^ n15803 ;
  assign n17588 = n17587 ^ n17586 ;
  assign n17591 = n15685 & n17588 ;
  assign n17592 = n17591 ^ n17587 ;
  assign n17593 = ~n15684 & ~n17592 ;
  assign n17605 = n17604 ^ n17593 ;
  assign n17607 = n17606 ^ n17605 ;
  assign n17579 = ~n15685 & ~n16853 ;
  assign n17608 = n17607 ^ n17579 ;
  assign n17573 = n15824 ^ n15823 ;
  assign n17574 = n15823 ^ n15684 ;
  assign n17575 = n17574 ^ n15823 ;
  assign n17576 = ~n17573 & n17575 ;
  assign n17577 = n17576 ^ n15823 ;
  assign n17578 = ~n15686 & n17577 ;
  assign n17609 = n17608 ^ n17578 ;
  assign n17610 = ~n16842 & ~n17609 ;
  assign n17612 = n17611 ^ n17610 ;
  assign n17613 = n17612 ^ x86 ;
  assign n17624 = ~n17456 & n17613 ;
  assign n17649 = n17624 ^ n17613 ;
  assign n17650 = n17649 ^ n17456 ;
  assign n18608 = n17565 & n17650 ;
  assign n18331 = n17491 & n17624 ;
  assign n18607 = ~n17554 & n18331 ;
  assign n18609 = n18608 ^ n18607 ;
  assign n19175 = n19166 ^ n18609 ;
  assign n17665 = n17613 ^ n17456 ;
  assign n17685 = n17684 ^ n17559 ;
  assign n17679 = n17655 ^ n17513 ;
  assign n17663 = n17662 ^ n17633 ;
  assign n17680 = n17679 ^ n17663 ;
  assign n17686 = n17685 ^ n17680 ;
  assign n17687 = n17456 & n17686 ;
  assign n17688 = n17687 ^ n17655 ;
  assign n17689 = n17665 & n17688 ;
  assign n19176 = n19175 ^ n17689 ;
  assign n17625 = ~n17623 & n17624 ;
  assign n17616 = ~n17570 & ~n17613 ;
  assign n17617 = n17616 ^ n17569 ;
  assign n17618 = n17456 & ~n17617 ;
  assign n17626 = n17625 ^ n17618 ;
  assign n19177 = n19176 ^ n17626 ;
  assign n18332 = n17556 & n18331 ;
  assign n18328 = ~n17613 & n17655 ;
  assign n18329 = n18328 ^ n17560 ;
  assign n18330 = n17665 & n18329 ;
  assign n18333 = n18332 ^ n18330 ;
  assign n19178 = n19177 ^ n18333 ;
  assign n18312 = n17638 ^ n17630 ;
  assign n18313 = n18312 ^ n17636 ;
  assign n18314 = n17636 ^ n17613 ;
  assign n18315 = n18314 ^ n17636 ;
  assign n18316 = ~n18313 & ~n18315 ;
  assign n18317 = n18316 ^ n17636 ;
  assign n18318 = ~n17456 & n18317 ;
  assign n19179 = n19178 ^ n18318 ;
  assign n19180 = n19179 ^ n14219 ;
  assign n19168 = n19166 ^ n17623 ;
  assign n19167 = n19166 ^ n17629 ;
  assign n19169 = n19168 ^ n19167 ;
  assign n19170 = n19168 ^ n17613 ;
  assign n19171 = n19170 ^ n19168 ;
  assign n19172 = ~n19169 & n19171 ;
  assign n19173 = n19172 ^ n19168 ;
  assign n19174 = n17665 & n19173 ;
  assign n19181 = n19180 ^ n19174 ;
  assign n19182 = n19181 ^ x82 ;
  assign n17334 = n16447 & n16540 ;
  assign n16795 = n16794 ^ n16455 ;
  assign n17299 = n16795 ^ n16507 ;
  assign n17297 = n16494 ^ n16470 ;
  assign n17298 = n17297 ^ n16473 ;
  assign n17300 = n17299 ^ n17298 ;
  assign n17301 = ~n16388 & ~n17300 ;
  assign n17302 = n17301 ^ n17299 ;
  assign n16774 = n16527 ^ n16500 ;
  assign n16775 = n16527 ^ n16387 ;
  assign n16776 = n16775 ^ n16527 ;
  assign n16777 = n16774 & n16776 ;
  assign n16778 = n16777 ^ n16527 ;
  assign n16779 = ~n16388 & n16778 ;
  assign n17329 = n17302 ^ n16779 ;
  assign n17330 = n17329 ^ n17328 ;
  assign n16788 = n16496 & n16515 ;
  assign n16787 = n16449 & n16540 ;
  assign n16789 = n16788 ^ n16787 ;
  assign n17331 = n17330 ^ n16789 ;
  assign n17332 = n17331 ^ n17317 ;
  assign n17304 = n17302 ^ n16451 ;
  assign n17303 = n17302 ^ n16527 ;
  assign n17305 = n17304 ^ n17303 ;
  assign n17308 = n16388 & n17305 ;
  assign n17309 = n17308 ^ n17304 ;
  assign n17310 = n16387 & ~n17309 ;
  assign n17333 = n17332 ^ n17310 ;
  assign n17335 = n17334 ^ n17333 ;
  assign n17336 = ~n16541 & n17335 ;
  assign n17337 = n17336 ^ n14255 ;
  assign n17338 = n17337 ^ x120 ;
  assign n17372 = n17371 ^ x65 ;
  assign n17373 = ~n17338 & n17372 ;
  assign n17374 = n17373 ^ n17338 ;
  assign n17233 = n17232 ^ x97 ;
  assign n17261 = n17260 ^ n16243 ;
  assign n17262 = n16334 & n17261 ;
  assign n17263 = n17262 ^ n16381 ;
  assign n17248 = n16347 ^ n16292 ;
  assign n17249 = n16334 & ~n17248 ;
  assign n17268 = n17263 ^ n17249 ;
  assign n17269 = n16356 & ~n17268 ;
  assign n16921 = n16382 ^ n16323 ;
  assign n16922 = n16921 ^ n16298 ;
  assign n16925 = ~n16334 & n16922 ;
  assign n16926 = n16925 ^ n16298 ;
  assign n16927 = n16356 & n16926 ;
  assign n17264 = n17263 ^ n16927 ;
  assign n17265 = n17264 ^ n17259 ;
  assign n17270 = n17269 ^ n17265 ;
  assign n17245 = ~n16328 & ~n16334 ;
  assign n17246 = n17245 ^ n16310 ;
  assign n17247 = n16335 & n17246 ;
  assign n17271 = n17270 ^ n17247 ;
  assign n17234 = n16336 ^ n16314 ;
  assign n17235 = n16338 ^ n16333 ;
  assign n17238 = ~n16336 & n17235 ;
  assign n17239 = n17238 ^ n16333 ;
  assign n17240 = n17234 & ~n17239 ;
  assign n17272 = n17271 ^ n17240 ;
  assign n17273 = ~n16898 & ~n17272 ;
  assign n17274 = ~n16353 & n17273 ;
  assign n17275 = n17274 ^ n14298 ;
  assign n17276 = n17275 ^ x123 ;
  assign n17277 = ~n17233 & n17276 ;
  assign n17279 = n17277 ^ n17233 ;
  assign n17288 = n17279 ^ n17276 ;
  assign n17289 = n17288 ^ n17233 ;
  assign n17171 = n15588 ^ n15585 ;
  assign n17172 = n17171 ^ n15594 ;
  assign n17173 = n17172 ^ n16660 ;
  assign n17174 = ~n15462 & n17173 ;
  assign n17169 = n17168 ^ n15559 ;
  assign n15602 = n15601 ^ n15556 ;
  assign n17170 = n17169 ^ n15602 ;
  assign n17175 = n17174 ^ n17170 ;
  assign n17183 = n17175 ^ n16669 ;
  assign n17184 = n17183 ^ n17182 ;
  assign n15638 = n15637 ^ n15595 ;
  assign n15639 = n15637 ^ n15462 ;
  assign n15640 = n15639 ^ n15637 ;
  assign n15641 = n15638 & ~n15640 ;
  assign n15642 = n15641 ^ n15637 ;
  assign n15643 = ~n15624 & n15642 ;
  assign n17185 = n17184 ^ n15643 ;
  assign n17176 = n17175 ^ n16662 ;
  assign n17164 = n15571 ^ n15558 ;
  assign n17165 = n17164 ^ n15578 ;
  assign n17166 = n17165 ^ n16662 ;
  assign n17167 = n15462 & n17166 ;
  assign n17177 = n17176 ^ n17167 ;
  assign n17178 = n15420 & ~n17177 ;
  assign n17186 = n17185 ^ n17178 ;
  assign n17187 = ~n15577 & n17186 ;
  assign n17188 = n17187 ^ n14323 ;
  assign n17189 = n17188 ^ x106 ;
  assign n17195 = n16179 ^ n14268 ;
  assign n17193 = n14613 ^ n14268 ;
  assign n17191 = n14613 ^ n14434 ;
  assign n17192 = n14610 & n17191 ;
  assign n17194 = n17193 ^ n17192 ;
  assign n17196 = n17195 ^ n17194 ;
  assign n17197 = ~n13147 & ~n17196 ;
  assign n17198 = n17197 ^ n17194 ;
  assign n17190 = n14433 & ~n14610 ;
  assign n17199 = n17198 ^ n17190 ;
  assign n17200 = n17199 ^ x88 ;
  assign n17201 = ~n17189 & ~n17200 ;
  assign n17282 = n17201 ^ n17189 ;
  assign n17382 = n17282 ^ n17200 ;
  assign n17398 = n17289 & ~n17382 ;
  assign n17292 = n17201 & n17288 ;
  assign n17433 = n17398 ^ n17292 ;
  assign n17391 = n17277 & ~n17382 ;
  assign n17284 = ~n17189 & ~n17233 ;
  assign n17283 = ~n17279 & ~n17282 ;
  assign n17285 = n17284 ^ n17283 ;
  assign n17392 = n17391 ^ n17285 ;
  assign n17280 = n17201 & ~n17279 ;
  assign n17390 = n17280 ^ n17277 ;
  assign n17393 = n17392 ^ n17390 ;
  assign n17388 = n17283 ^ n17279 ;
  assign n17383 = ~n17279 & ~n17382 ;
  assign n17384 = n17383 ^ n17280 ;
  assign n17389 = n17388 ^ n17384 ;
  assign n17394 = n17393 ^ n17389 ;
  assign n17376 = n17201 ^ n17200 ;
  assign n17377 = n17288 & ~n17376 ;
  assign n17387 = n17377 ^ n17376 ;
  assign n17395 = n17394 ^ n17387 ;
  assign n17444 = n17433 ^ n17395 ;
  assign n17278 = n17201 & n17277 ;
  assign n17281 = n17280 ^ n17278 ;
  assign n17291 = n17281 ^ n17201 ;
  assign n17293 = n17292 ^ n17291 ;
  assign n17445 = n17444 ^ n17293 ;
  assign n17290 = ~n17189 & n17289 ;
  assign n17294 = n17293 ^ n17290 ;
  assign n17378 = n17377 ^ n17294 ;
  assign n17295 = n17294 ^ n17283 ;
  assign n17286 = n17285 ^ n17281 ;
  assign n17287 = n17286 ^ n17282 ;
  assign n17296 = n17295 ^ n17287 ;
  assign n17379 = n17378 ^ n17296 ;
  assign n17443 = n17379 ^ n17233 ;
  assign n17446 = n17445 ^ n17443 ;
  assign n19116 = n17446 ^ n17378 ;
  assign n19117 = n19116 ^ n17281 ;
  assign n19118 = ~n17374 & ~n19117 ;
  assign n19113 = ~n17338 & n17391 ;
  assign n19106 = n17445 ^ n17392 ;
  assign n19107 = n17392 ^ n17338 ;
  assign n19108 = n19107 ^ n17392 ;
  assign n19109 = n19106 & ~n19108 ;
  assign n19110 = n19109 ^ n17392 ;
  assign n19111 = n17372 & n19110 ;
  assign n17380 = n17374 ^ n17372 ;
  assign n19104 = n17380 & ~n17394 ;
  assign n17385 = n17380 ^ n17373 ;
  assign n17411 = n17393 ^ n17296 ;
  assign n17414 = ~n17372 & ~n17411 ;
  assign n17415 = n17414 ^ n17296 ;
  assign n17416 = ~n17385 & ~n17415 ;
  assign n19105 = n19104 ^ n17416 ;
  assign n19112 = n19111 ^ n19105 ;
  assign n19114 = n19113 ^ n19112 ;
  assign n19102 = n17383 ^ n17286 ;
  assign n19103 = n17385 & n19102 ;
  assign n19115 = n19114 ^ n19103 ;
  assign n19119 = n19118 ^ n19115 ;
  assign n19094 = n17377 ^ n17293 ;
  assign n17417 = n17293 ^ n17283 ;
  assign n18550 = n17417 ^ n17292 ;
  assign n18551 = n18550 ^ n17378 ;
  assign n19095 = n19094 ^ n18551 ;
  assign n19096 = n19095 ^ n19094 ;
  assign n19097 = n19094 ^ n17372 ;
  assign n19098 = n19097 ^ n19094 ;
  assign n19099 = n19096 & ~n19098 ;
  assign n19100 = n19099 ^ n19094 ;
  assign n19101 = n17338 & n19100 ;
  assign n19120 = n19119 ^ n19101 ;
  assign n18567 = n17373 & ~n17389 ;
  assign n19121 = n19120 ^ n18567 ;
  assign n17375 = ~n17296 & ~n17374 ;
  assign n19122 = n19121 ^ n17375 ;
  assign n17441 = n17395 ^ n17372 ;
  assign n17442 = n17441 ^ n17395 ;
  assign n17447 = n17446 ^ n17395 ;
  assign n17450 = n17442 & ~n17447 ;
  assign n17451 = n17450 ^ n17395 ;
  assign n17452 = n17338 & n17451 ;
  assign n19123 = n19122 ^ n17452 ;
  assign n19124 = n19123 ^ n14409 ;
  assign n19125 = n19124 ^ x64 ;
  assign n19230 = n19182 ^ n19125 ;
  assign n16766 = n16192 ^ x91 ;
  assign n16805 = n16784 ^ n16502 ;
  assign n16802 = n16502 ^ n16455 ;
  assign n16803 = n16802 ^ n16474 ;
  assign n16804 = n16388 & n16803 ;
  assign n16806 = n16805 ^ n16804 ;
  assign n16807 = ~n16387 & n16806 ;
  assign n16780 = n16475 ^ n16451 ;
  assign n16798 = n16780 ^ n16504 ;
  assign n16793 = n16504 ^ n16468 ;
  assign n16796 = n16795 ^ n16793 ;
  assign n16797 = ~n16388 & n16796 ;
  assign n16799 = n16798 ^ n16797 ;
  assign n16800 = n16516 & n16799 ;
  assign n16785 = n16784 ^ n16780 ;
  assign n16786 = n16785 ^ n16779 ;
  assign n16790 = n16789 ^ n16786 ;
  assign n16791 = n16790 ^ n16773 ;
  assign n16792 = n16791 ^ n11604 ;
  assign n16801 = n16800 ^ n16792 ;
  assign n16808 = n16807 ^ n16801 ;
  assign n16809 = n16808 ^ x109 ;
  assign n16810 = ~n16766 & ~n16809 ;
  assign n16811 = n16810 ^ n16766 ;
  assign n16812 = n16811 ^ n16809 ;
  assign n16813 = n16812 ^ n16766 ;
  assign n15814 = n15813 ^ n15792 ;
  assign n16856 = n15814 ^ n15791 ;
  assign n16854 = n16853 ^ n15779 ;
  assign n16855 = n16854 ^ n16814 ;
  assign n16857 = n16856 ^ n16855 ;
  assign n16858 = ~n15685 & n16857 ;
  assign n16859 = n16858 ^ n16856 ;
  assign n16860 = n15684 & n16859 ;
  assign n16834 = n15805 ^ n15761 ;
  assign n16843 = n16842 ^ n16834 ;
  assign n16846 = n16845 ^ n16843 ;
  assign n16847 = n16846 ^ n15837 ;
  assign n16848 = n16847 ^ n13324 ;
  assign n16825 = n15805 ^ n15776 ;
  assign n16827 = n16826 ^ n16825 ;
  assign n16828 = n16827 ^ n15805 ;
  assign n16829 = n15805 ^ n15685 ;
  assign n16830 = n16829 ^ n15805 ;
  assign n16831 = n16828 & n16830 ;
  assign n16832 = n16831 ^ n15805 ;
  assign n16833 = n15686 & ~n16832 ;
  assign n16849 = n16848 ^ n16833 ;
  assign n16820 = n15761 ^ n15684 ;
  assign n16821 = n16820 ^ n15761 ;
  assign n16822 = n15823 & ~n16821 ;
  assign n16823 = n16822 ^ n15761 ;
  assign n16824 = ~n15685 & n16823 ;
  assign n16850 = n16849 ^ n16824 ;
  assign n16816 = n16815 ^ n15782 ;
  assign n16817 = ~n15832 & ~n16816 ;
  assign n16851 = n16850 ^ n16817 ;
  assign n16861 = n16860 ^ n16851 ;
  assign n16862 = n16861 ^ x77 ;
  assign n16897 = n16677 ^ x84 ;
  assign n16918 = n16333 ^ n16314 ;
  assign n16919 = ~n16337 & n16918 ;
  assign n16914 = n16329 ^ n16303 ;
  assign n16915 = ~n16356 & n16914 ;
  assign n16909 = n16312 ^ n16301 ;
  assign n16910 = n16909 ^ n16320 ;
  assign n16911 = ~n16335 & ~n16910 ;
  assign n16912 = n16911 ^ n16320 ;
  assign n16913 = ~n16334 & n16912 ;
  assign n16916 = n16915 ^ n16913 ;
  assign n16899 = n16334 ^ n16321 ;
  assign n16900 = n16302 ^ n16299 ;
  assign n16901 = n16900 ^ n16321 ;
  assign n16902 = n16901 ^ n16302 ;
  assign n16903 = n16902 ^ n16324 ;
  assign n16904 = n16335 & ~n16903 ;
  assign n16905 = n16904 ^ n16900 ;
  assign n16906 = n16899 & n16905 ;
  assign n16917 = n16916 ^ n16906 ;
  assign n16920 = n16919 ^ n16917 ;
  assign n16928 = n16920 & ~n16927 ;
  assign n16929 = ~n16898 & n16928 ;
  assign n16930 = ~n16340 & n16929 ;
  assign n16931 = ~n16353 & n16930 ;
  assign n16932 = n16931 ^ n12923 ;
  assign n16933 = n16932 ^ x78 ;
  assign n16934 = n16897 & n16933 ;
  assign n16935 = n16934 ^ n16933 ;
  assign n16953 = ~n16862 & n16935 ;
  assign n15992 = n15991 ^ n15987 ;
  assign n16086 = n16065 ^ n16026 ;
  assign n16889 = ~n15992 & ~n16086 ;
  assign n16886 = n16885 ^ n16028 ;
  assign n16870 = n15968 ^ n15958 ;
  assign n16871 = n16870 ^ n15988 ;
  assign n16872 = n16026 & ~n16871 ;
  assign n16873 = n16872 ^ n15968 ;
  assign n16882 = n16873 ^ n16039 ;
  assign n16875 = n16873 ^ n15980 ;
  assign n16874 = n16873 ^ n16030 ;
  assign n16876 = n16875 ^ n16874 ;
  assign n16879 = n16026 & n16876 ;
  assign n16880 = n16879 ^ n16875 ;
  assign n16881 = ~n16040 & n16880 ;
  assign n16883 = n16882 ^ n16881 ;
  assign n16887 = n16886 ^ n16883 ;
  assign n16055 = n16054 ^ n15985 ;
  assign n16058 = n16026 & ~n16055 ;
  assign n16059 = n16058 ^ n15985 ;
  assign n16060 = n15857 & ~n16059 ;
  assign n16888 = n16887 ^ n16060 ;
  assign n16890 = n16889 ^ n16888 ;
  assign n16863 = n16074 ^ n16028 ;
  assign n16864 = n16065 ^ n16029 ;
  assign n16865 = n16029 ^ n16028 ;
  assign n16866 = n16865 ^ n16029 ;
  assign n16867 = n16864 & n16866 ;
  assign n16868 = n16867 ^ n16029 ;
  assign n16869 = n16863 & ~n16868 ;
  assign n16891 = n16890 ^ n16869 ;
  assign n16893 = n16892 ^ n16891 ;
  assign n16894 = n16893 ^ n13530 ;
  assign n16895 = n16894 ^ x126 ;
  assign n16896 = ~n16862 & ~n16895 ;
  assign n16952 = n16896 & n16935 ;
  assign n16954 = n16953 ^ n16952 ;
  assign n16950 = n16896 ^ n16862 ;
  assign n16951 = n16934 & ~n16950 ;
  assign n16955 = n16954 ^ n16951 ;
  assign n16956 = n16955 ^ n16950 ;
  assign n16938 = n16934 ^ n16897 ;
  assign n16947 = n16896 & n16938 ;
  assign n16939 = n16896 ^ n16895 ;
  assign n16946 = n16938 & ~n16939 ;
  assign n16948 = n16947 ^ n16946 ;
  assign n16940 = n16939 ^ n16862 ;
  assign n16941 = n16938 & ~n16940 ;
  assign n16945 = n16941 ^ n16938 ;
  assign n16949 = n16948 ^ n16945 ;
  assign n16957 = n16956 ^ n16949 ;
  assign n16958 = n16957 ^ n16941 ;
  assign n16936 = n16935 ^ n16897 ;
  assign n16944 = ~n16936 & ~n16939 ;
  assign n16959 = n16958 ^ n16944 ;
  assign n16937 = n16896 & ~n16936 ;
  assign n16942 = n16941 ^ n16937 ;
  assign n16943 = n16942 ^ n16936 ;
  assign n16960 = n16959 ^ n16943 ;
  assign n16961 = ~n16813 & n16960 ;
  assign n16966 = n16946 ^ n16944 ;
  assign n16964 = n16934 & ~n16939 ;
  assign n16965 = n16964 ^ n16939 ;
  assign n16967 = n16966 ^ n16965 ;
  assign n16963 = n16896 & n16934 ;
  assign n16968 = n16967 ^ n16963 ;
  assign n17009 = n16968 ^ n16952 ;
  assign n17010 = n17009 ^ n16952 ;
  assign n17011 = n16952 ^ n16766 ;
  assign n17012 = n17011 ^ n16952 ;
  assign n17013 = ~n17010 & ~n17012 ;
  assign n17014 = n17013 ^ n16952 ;
  assign n17015 = n16809 & n17014 ;
  assign n17016 = n17015 ^ n16952 ;
  assign n16969 = n16968 ^ n16946 ;
  assign n19152 = ~n16811 & ~n16969 ;
  assign n16971 = n16967 ^ n16934 ;
  assign n16970 = n16953 ^ n16933 ;
  assign n16972 = n16971 ^ n16970 ;
  assign n19147 = n16972 ^ n16969 ;
  assign n16992 = n16809 ^ n16766 ;
  assign n18706 = n16949 ^ n16809 ;
  assign n18707 = n18706 ^ n16949 ;
  assign n16974 = n16960 ^ n16941 ;
  assign n16973 = n16972 ^ n16940 ;
  assign n16975 = n16974 ^ n16973 ;
  assign n18708 = n16975 ^ n16949 ;
  assign n18711 = ~n18707 & n18708 ;
  assign n18712 = n18711 ^ n16949 ;
  assign n18713 = ~n16992 & n18712 ;
  assign n19139 = n18713 ^ n16964 ;
  assign n19126 = n16944 ^ n16941 ;
  assign n19127 = n16811 & ~n19126 ;
  assign n19128 = n16958 ^ n16949 ;
  assign n17021 = ~n16813 & n16944 ;
  assign n19129 = n19128 ^ n17021 ;
  assign n19130 = ~n19127 & ~n19129 ;
  assign n19131 = n19130 ^ n16937 ;
  assign n19132 = n19131 ^ n16813 ;
  assign n19133 = n16955 ^ n16811 ;
  assign n19136 = ~n19131 & n19133 ;
  assign n19137 = n19136 ^ n16811 ;
  assign n19138 = ~n19132 & ~n19137 ;
  assign n19140 = n19139 ^ n19138 ;
  assign n19148 = n19147 ^ n19140 ;
  assign n19142 = n16957 ^ n16944 ;
  assign n19143 = n19142 ^ n16964 ;
  assign n18692 = n16972 ^ n16963 ;
  assign n19144 = n19143 ^ n18692 ;
  assign n19145 = ~n16766 & ~n19144 ;
  assign n17008 = n16810 & n16948 ;
  assign n19141 = n19140 ^ n17008 ;
  assign n19146 = n19145 ^ n19141 ;
  assign n19149 = n19148 ^ n19146 ;
  assign n19150 = ~n16809 & ~n19149 ;
  assign n19151 = n19150 ^ n19148 ;
  assign n19153 = n19152 ^ n19151 ;
  assign n19154 = ~n17016 & ~n19153 ;
  assign n17027 = ~n16812 & ~n16958 ;
  assign n19155 = n19154 ^ n17027 ;
  assign n19156 = ~n16961 & n19155 ;
  assign n19157 = n19156 ^ n13613 ;
  assign n19158 = n19157 ^ x73 ;
  assign n19236 = n19158 ^ n19125 ;
  assign n19241 = n19230 & n19236 ;
  assign n19265 = n19160 & n19241 ;
  assign n19231 = n19230 ^ n19160 ;
  assign n19237 = n19160 ^ n19125 ;
  assign n19238 = n19236 & ~n19237 ;
  assign n19239 = n19238 ^ n19160 ;
  assign n19240 = n19231 & ~n19239 ;
  assign n19261 = n19240 ^ n19125 ;
  assign n19159 = ~n19125 & n19158 ;
  assign n19185 = n19159 ^ n19125 ;
  assign n19183 = n19160 & ~n19182 ;
  assign n19186 = n19183 ^ n19182 ;
  assign n19187 = ~n19185 & ~n19186 ;
  assign n19262 = n19261 ^ n19187 ;
  assign n19256 = n19182 ^ n19158 ;
  assign n19244 = ~n19158 & n19160 ;
  assign n19257 = n19244 ^ n19125 ;
  assign n19258 = ~n19256 & n19257 ;
  assign n19248 = n19182 ^ n19160 ;
  assign n19259 = n19258 ^ n19248 ;
  assign n19255 = n19239 ^ n19158 ;
  assign n19260 = n19259 ^ n19255 ;
  assign n19263 = n19262 ^ n19260 ;
  assign n19234 = n19160 ^ n19158 ;
  assign n19243 = n19234 ^ n19230 ;
  assign n19245 = n19244 ^ n19160 ;
  assign n19246 = n19245 ^ n19234 ;
  assign n19247 = n19246 ^ n19160 ;
  assign n19251 = ~n19247 & ~n19248 ;
  assign n19252 = n19251 ^ n19160 ;
  assign n19253 = ~n19243 & n19252 ;
  assign n19254 = n19253 ^ n19244 ;
  assign n19264 = n19263 ^ n19254 ;
  assign n19266 = n19265 ^ n19264 ;
  assign n19232 = n19230 ^ n19159 ;
  assign n19233 = ~n19231 & n19232 ;
  assign n19235 = n19234 ^ n19233 ;
  assign n19267 = n19266 ^ n19235 ;
  assign n19242 = n19241 ^ n19240 ;
  assign n19268 = n19267 ^ n19242 ;
  assign n20748 = n19268 ^ n17199 ;
  assign n15847 = n15824 ^ n15761 ;
  assign n15848 = n15847 ^ n15744 ;
  assign n15849 = n15831 & ~n15848 ;
  assign n15841 = n15789 ^ n15762 ;
  assign n15842 = n15841 ^ n15781 ;
  assign n15843 = ~n15684 & ~n15842 ;
  assign n15835 = n15789 ^ n15788 ;
  assign n15836 = n15835 ^ n15834 ;
  assign n15838 = n15837 ^ n15836 ;
  assign n15839 = n15838 ^ n15834 ;
  assign n15840 = n15839 ^ n15837 ;
  assign n15844 = n15843 ^ n15840 ;
  assign n15845 = n15686 & n15844 ;
  assign n15846 = n15845 ^ n15838 ;
  assign n15850 = n15849 ^ n15846 ;
  assign n15851 = n15850 ^ n15782 ;
  assign n15852 = n15851 ^ n15830 ;
  assign n15853 = n15852 ^ n13059 ;
  assign n15817 = n15782 ^ n15684 ;
  assign n15818 = n15817 ^ n15782 ;
  assign n15819 = ~n15814 & ~n15818 ;
  assign n15820 = n15819 ^ n15782 ;
  assign n15821 = n15685 & n15820 ;
  assign n15854 = n15853 ^ n15821 ;
  assign n15769 = n15768 ^ n15761 ;
  assign n15770 = n15768 ^ n15684 ;
  assign n15771 = n15770 ^ n15768 ;
  assign n15772 = ~n15769 & n15771 ;
  assign n15773 = n15772 ^ n15768 ;
  assign n15774 = ~n15686 & ~n15773 ;
  assign n15855 = n15854 ^ n15774 ;
  assign n17080 = n15855 ^ x125 ;
  assign n17081 = n16932 ^ x116 ;
  assign n17082 = n17080 & ~n17081 ;
  assign n17083 = n17082 ^ n17081 ;
  assign n17073 = n14624 ^ n14622 ;
  assign n17074 = n17073 ^ n12024 ;
  assign n17075 = n17074 ^ x102 ;
  assign n15058 = n15057 ^ n15036 ;
  assign n15054 = n15017 ^ n15016 ;
  assign n15055 = ~n14678 & n15054 ;
  assign n15059 = n15058 ^ n15055 ;
  assign n15052 = n15051 ^ n15028 ;
  assign n15053 = n15052 ^ n15016 ;
  assign n15060 = n15059 ^ n15053 ;
  assign n15061 = n15060 ^ n15059 ;
  assign n15037 = n15036 ^ n15033 ;
  assign n15038 = n15037 ^ n15027 ;
  assign n15062 = n15061 ^ n15038 ;
  assign n15063 = ~n14678 & ~n15062 ;
  assign n15064 = n15063 ^ n15060 ;
  assign n15065 = ~n14679 & ~n15064 ;
  assign n15066 = n15065 ^ n15059 ;
  assign n15092 = n15066 ^ n12392 ;
  assign n15088 = n15082 ^ n14679 ;
  assign n15089 = n15087 & n15088 ;
  assign n15090 = n15089 ^ n15086 ;
  assign n15091 = n15090 ^ n15085 ;
  assign n15093 = n15092 ^ n15091 ;
  assign n15070 = n15013 ^ n14852 ;
  assign n15071 = n15070 ^ n15029 ;
  assign n15072 = n14679 & n15071 ;
  assign n15094 = n15093 ^ n15072 ;
  assign n15069 = n14678 & n15030 ;
  assign n15095 = n15094 ^ n15069 ;
  assign n15067 = ~n15020 & ~n15066 ;
  assign n15068 = ~n14680 & n15067 ;
  assign n15096 = n15095 ^ n15068 ;
  assign n17076 = n15096 ^ x85 ;
  assign n17077 = ~n17075 & n17076 ;
  assign n17092 = n17077 ^ n17075 ;
  assign n17033 = n16808 ^ x75 ;
  assign n17043 = n16596 ^ n15375 ;
  assign n17044 = n17043 ^ n15410 ;
  assign n17045 = n15152 & n17044 ;
  assign n17046 = n17045 ^ n15384 ;
  assign n17047 = n17046 ^ n15367 ;
  assign n17048 = n17047 ^ n15342 ;
  assign n17049 = n17048 ^ n15384 ;
  assign n17050 = n17049 ^ n17047 ;
  assign n17053 = ~n15152 & ~n17050 ;
  assign n17054 = n17053 ^ n17047 ;
  assign n17055 = n15132 & ~n17054 ;
  assign n17056 = n17055 ^ n17045 ;
  assign n17040 = n16595 ^ n15349 ;
  assign n17041 = n17040 ^ n15392 ;
  assign n17042 = ~n15343 & n17041 ;
  assign n17057 = n17056 ^ n17042 ;
  assign n17039 = n15153 & n15374 ;
  assign n17058 = n17057 ^ n17039 ;
  assign n17034 = n15406 ^ n15357 ;
  assign n17035 = n17034 ^ n15406 ;
  assign n17036 = ~n16601 & n17035 ;
  assign n17037 = n17036 ^ n15406 ;
  assign n17038 = n15132 & n17037 ;
  assign n17059 = n17058 ^ n17038 ;
  assign n17060 = n17059 ^ n15344 ;
  assign n17061 = n15374 ^ n15339 ;
  assign n17062 = n15339 ^ n15132 ;
  assign n17063 = n17062 ^ n15339 ;
  assign n17064 = n17061 & ~n17063 ;
  assign n17065 = n17064 ^ n15339 ;
  assign n17066 = n15373 & n17065 ;
  assign n17067 = ~n17060 & ~n17066 ;
  assign n17068 = ~n15363 & n17067 ;
  assign n17069 = ~n15416 & n17068 ;
  assign n17070 = n17069 ^ n12705 ;
  assign n17071 = n17070 ^ x92 ;
  assign n17072 = n17033 & ~n17071 ;
  assign n17087 = n17072 ^ n17071 ;
  assign n17119 = n17087 ^ n17033 ;
  assign n17120 = ~n17092 & n17119 ;
  assign n17078 = n17077 ^ n17076 ;
  assign n17086 = n17078 ^ n17075 ;
  assign n17089 = n17072 ^ n17033 ;
  assign n17090 = n17086 & n17089 ;
  assign n17965 = n17120 ^ n17090 ;
  assign n17966 = ~n17083 & n17965 ;
  assign n17094 = ~n17033 & n17076 ;
  assign n17095 = n17094 ^ n17078 ;
  assign n17079 = n17072 & n17078 ;
  assign n17136 = n17095 ^ n17079 ;
  assign n17100 = ~n17071 & n17077 ;
  assign n17101 = n17100 ^ n17077 ;
  assign n17099 = n17077 & n17089 ;
  assign n17102 = n17101 ^ n17099 ;
  assign n17098 = n17078 & n17089 ;
  assign n17103 = n17102 ^ n17098 ;
  assign n17104 = n17103 ^ n17100 ;
  assign n17137 = n17136 ^ n17104 ;
  assign n17128 = n17102 ^ n17079 ;
  assign n17129 = n17128 ^ n17078 ;
  assign n17126 = n17078 & ~n17087 ;
  assign n17127 = n17126 ^ n17103 ;
  assign n17130 = n17129 ^ n17127 ;
  assign n17982 = n17137 ^ n17130 ;
  assign n17983 = n17982 ^ n17128 ;
  assign n17984 = ~n17080 & n17983 ;
  assign n17093 = n17072 & ~n17092 ;
  assign n17096 = n17095 ^ n17093 ;
  assign n17097 = n17096 ^ n17072 ;
  assign n17105 = n17104 ^ n17097 ;
  assign n17106 = n17105 ^ n17086 ;
  assign n17088 = n17086 & ~n17087 ;
  assign n17091 = n17090 ^ n17088 ;
  assign n17107 = n17106 ^ n17091 ;
  assign n17108 = n17107 ^ n17093 ;
  assign n17980 = n17108 ^ n17105 ;
  assign n17981 = n17082 & n17980 ;
  assign n17985 = n17984 ^ n17981 ;
  assign n17150 = n17083 ^ n17080 ;
  assign n17978 = n17108 ^ n17088 ;
  assign n17979 = n17150 & n17978 ;
  assign n17986 = n17985 ^ n17979 ;
  assign n17085 = n17082 ^ n17080 ;
  assign n17974 = n17126 ^ n17120 ;
  assign n17975 = n17974 ^ n17095 ;
  assign n17976 = n17975 ^ n17108 ;
  assign n17977 = n17085 & ~n17976 ;
  assign n17987 = n17986 ^ n17977 ;
  assign n17967 = n17126 ^ n17105 ;
  assign n17968 = n17967 ^ n17095 ;
  assign n17969 = n17095 ^ n17080 ;
  assign n17970 = n17969 ^ n17095 ;
  assign n17971 = n17968 & ~n17970 ;
  assign n17972 = n17971 ^ n17095 ;
  assign n17973 = ~n17081 & n17972 ;
  assign n17988 = n17987 ^ n17973 ;
  assign n17134 = n17085 ^ n17083 ;
  assign n17116 = ~n17087 & ~n17092 ;
  assign n17157 = n17116 ^ n17092 ;
  assign n17156 = n17120 ^ n17093 ;
  assign n17158 = n17157 ^ n17156 ;
  assign n17159 = n17134 & ~n17158 ;
  assign n17989 = n17988 ^ n17159 ;
  assign n17990 = ~n17966 & ~n17989 ;
  assign n17991 = n17990 ^ n13146 ;
  assign n19228 = n17991 ^ x105 ;
  assign n19184 = n19159 & n19183 ;
  assign n19188 = n19187 ^ n19184 ;
  assign n20745 = n19268 ^ n19188 ;
  assign n20746 = n20745 ^ n19235 ;
  assign n20747 = n19228 & ~n20746 ;
  assign n20749 = n20748 ^ n20747 ;
  assign n20750 = n20749 ^ n17199 ;
  assign n19357 = n19265 ^ n19184 ;
  assign n19358 = n19228 & n19357 ;
  assign n19359 = n19358 ^ n19265 ;
  assign n20738 = n19262 ^ n19228 ;
  assign n20739 = n20738 ^ n19262 ;
  assign n20740 = n19264 ^ n19188 ;
  assign n20741 = n20740 ^ n19262 ;
  assign n20742 = ~n20739 & n20741 ;
  assign n20743 = n20742 ^ n19262 ;
  assign n20744 = ~n19359 & ~n20743 ;
  assign n20751 = n20750 ^ n20744 ;
  assign n20752 = ~n19227 & ~n20751 ;
  assign n20753 = n20752 ^ n20749 ;
  assign n20754 = n20753 ^ x121 ;
  assign n18047 = n17488 ^ x74 ;
  assign n18073 = n15416 ^ n14753 ;
  assign n18070 = n15154 & n15381 ;
  assign n18062 = n17040 ^ n15154 ;
  assign n18063 = n18062 ^ n15409 ;
  assign n18064 = n18063 ^ n15386 ;
  assign n18065 = n15372 & ~n18064 ;
  assign n18066 = n18065 ^ n15154 ;
  assign n18067 = n15406 ^ n15372 ;
  assign n18068 = n18066 & n18067 ;
  assign n18052 = n16618 ^ n15365 ;
  assign n18053 = n18052 ^ n15366 ;
  assign n18054 = n18053 ^ n15365 ;
  assign n18055 = n18054 ^ n15374 ;
  assign n18056 = ~n15132 & ~n18055 ;
  assign n18057 = n18056 ^ n18052 ;
  assign n18050 = n15379 ^ n15355 ;
  assign n18051 = n15152 & ~n18050 ;
  assign n18058 = n18057 ^ n18051 ;
  assign n18059 = ~n16599 & ~n18058 ;
  assign n18060 = n18059 ^ n15132 ;
  assign n18048 = n15391 ^ n15356 ;
  assign n18049 = ~n15132 & n18048 ;
  assign n18061 = n18060 ^ n18049 ;
  assign n18069 = n18068 ^ n18061 ;
  assign n18071 = n18070 ^ n18069 ;
  assign n18072 = ~n17066 & ~n18071 ;
  assign n18074 = n18073 ^ n18072 ;
  assign n18075 = n18074 ^ x89 ;
  assign n18077 = n15045 ^ n15042 ;
  assign n18112 = n17367 ^ n15090 ;
  assign n18079 = n15026 ^ n15025 ;
  assign n18080 = n18079 ^ n15051 ;
  assign n18097 = n18080 ^ n17357 ;
  assign n18082 = n18080 ^ n14678 ;
  assign n18083 = n18082 ^ n15025 ;
  assign n18078 = n15025 ^ n14680 ;
  assign n18081 = n18080 ^ n18078 ;
  assign n18086 = n18081 ^ n18080 ;
  assign n18087 = n18086 ^ n15025 ;
  assign n18088 = ~n18083 & ~n18087 ;
  assign n18089 = n18088 ^ n18081 ;
  assign n18090 = n18088 ^ n18087 ;
  assign n18091 = ~n18079 & ~n18090 ;
  assign n18092 = n18091 ^ n15026 ;
  assign n18093 = n18092 ^ n18079 ;
  assign n18094 = ~n18089 & ~n18093 ;
  assign n18095 = n18094 ^ n18091 ;
  assign n18096 = n18095 ^ n15025 ;
  assign n18098 = n18097 ^ n18096 ;
  assign n18099 = n18098 ^ n17357 ;
  assign n18100 = ~n15088 & n18099 ;
  assign n18101 = n18100 ^ n17357 ;
  assign n18102 = ~n15081 & n18101 ;
  assign n18103 = n18102 ^ n17357 ;
  assign n18104 = n15080 ^ n15018 ;
  assign n18105 = n18104 ^ n18103 ;
  assign n18106 = n16561 ^ n15088 ;
  assign n18107 = ~n15080 & ~n18106 ;
  assign n18108 = n18107 ^ n16561 ;
  assign n18109 = n18105 & ~n18108 ;
  assign n18110 = n18109 ^ n15080 ;
  assign n18111 = ~n18103 & ~n18110 ;
  assign n18113 = n18112 ^ n18111 ;
  assign n18114 = ~n16545 & n18113 ;
  assign n18115 = n15058 ^ n15016 ;
  assign n18116 = n18115 ^ n15050 ;
  assign n18117 = n15050 ^ n14678 ;
  assign n18118 = n18117 ^ n15050 ;
  assign n18119 = n18116 & ~n18118 ;
  assign n18120 = n18119 ^ n15050 ;
  assign n18121 = ~n14679 & n18120 ;
  assign n18122 = n18114 & ~n18121 ;
  assign n18123 = ~n15079 & n18122 ;
  assign n18124 = n15081 & n18123 ;
  assign n18125 = n18077 & n18124 ;
  assign n18126 = n18125 ^ n18123 ;
  assign n18128 = n14680 & n15027 ;
  assign n18129 = n18126 & n18128 ;
  assign n18127 = n18126 ^ n14714 ;
  assign n18130 = n18129 ^ n18127 ;
  assign n18131 = n18130 ^ x98 ;
  assign n18134 = n17337 ^ x99 ;
  assign n18076 = n17612 ^ x80 ;
  assign n18132 = n18131 ^ n18076 ;
  assign n18141 = n18134 ^ n18132 ;
  assign n18142 = n18131 & ~n18141 ;
  assign n18143 = n18142 ^ n18132 ;
  assign n18144 = ~n18075 & ~n18143 ;
  assign n18145 = n18144 ^ n18141 ;
  assign n18135 = n18134 ^ n18076 ;
  assign n18136 = n18131 ^ n18075 ;
  assign n18137 = n18134 & n18136 ;
  assign n18138 = n18137 ^ n18131 ;
  assign n18139 = ~n18135 & ~n18138 ;
  assign n18133 = n18132 ^ n18075 ;
  assign n18140 = n18139 ^ n18133 ;
  assign n18146 = n18145 ^ n18140 ;
  assign n18167 = n17188 ^ x121 ;
  assign n18648 = ~n18146 & ~n18167 ;
  assign n18649 = n18648 ^ n18145 ;
  assign n18642 = n18075 & n18134 ;
  assign n18643 = n18642 ^ n18131 ;
  assign n18644 = n18132 & n18643 ;
  assign n18645 = n18644 ^ n18131 ;
  assign n18646 = n18167 & ~n18645 ;
  assign n18163 = n18134 ^ n18131 ;
  assign n18149 = n18134 ^ n18075 ;
  assign n18156 = ~n18076 & ~n18131 ;
  assign n18157 = ~n18149 & n18156 ;
  assign n18158 = n18157 ^ n18137 ;
  assign n18159 = n18158 ^ n18139 ;
  assign n18160 = n18159 ^ n18149 ;
  assign n18150 = n18149 ^ n18076 ;
  assign n18151 = n18150 ^ n18076 ;
  assign n18152 = ~n18135 & ~n18151 ;
  assign n18153 = n18152 ^ n18076 ;
  assign n18154 = n18141 & n18153 ;
  assign n18155 = n18154 ^ n18076 ;
  assign n18161 = n18160 ^ n18155 ;
  assign n18148 = n18139 ^ n18134 ;
  assign n18162 = n18161 ^ n18148 ;
  assign n18164 = n18163 ^ n18162 ;
  assign n18647 = n18646 ^ n18164 ;
  assign n18650 = n18649 ^ n18647 ;
  assign n18651 = n18047 & ~n18650 ;
  assign n18652 = n18651 ^ n18649 ;
  assign n18653 = n18652 ^ n15546 ;
  assign n18654 = n18653 ^ x86 ;
  assign n16962 = ~n16811 & n16946 ;
  assign n17020 = ~n16813 & n16949 ;
  assign n17022 = n17021 ^ n17020 ;
  assign n16993 = n16951 ^ n16809 ;
  assign n16994 = n16993 ^ n16951 ;
  assign n17001 = n16964 ^ n16952 ;
  assign n17002 = n17001 ^ n16944 ;
  assign n17003 = n17002 ^ n16951 ;
  assign n17004 = n16994 & n17003 ;
  assign n17005 = n17004 ^ n16951 ;
  assign n17006 = ~n16992 & n17005 ;
  assign n18716 = n16810 & n16942 ;
  assign n18699 = n16960 ^ n16957 ;
  assign n18700 = n18699 ^ n17001 ;
  assign n18701 = ~n16809 & ~n18700 ;
  assign n18702 = n18701 ^ n16974 ;
  assign n18714 = n18702 ^ n18692 ;
  assign n18715 = n18714 ^ n18713 ;
  assign n18717 = n18716 ^ n18715 ;
  assign n18703 = n18702 ^ n16969 ;
  assign n18695 = n16957 ^ n16947 ;
  assign n18696 = n18695 ^ n16969 ;
  assign n16983 = n16975 ^ n16954 ;
  assign n16984 = n16983 ^ n16937 ;
  assign n18697 = n18696 ^ n16984 ;
  assign n18698 = n16809 & n18697 ;
  assign n18704 = n18703 ^ n18698 ;
  assign n18705 = ~n16766 & ~n18704 ;
  assign n18718 = n18717 ^ n18705 ;
  assign n18688 = n16957 ^ n16951 ;
  assign n18689 = n18688 ^ n16967 ;
  assign n18690 = n16809 & n18689 ;
  assign n18691 = n18690 ^ n16957 ;
  assign n18693 = n18692 ^ n18691 ;
  assign n18694 = ~n16992 & n18693 ;
  assign n18719 = n18718 ^ n18694 ;
  assign n18720 = ~n17006 & n18719 ;
  assign n18721 = ~n17022 & n18720 ;
  assign n18722 = ~n16962 & n18721 ;
  assign n18723 = n18722 ^ n15543 ;
  assign n18724 = n18723 ^ x76 ;
  assign n18738 = n18654 & n18724 ;
  assign n18739 = n18738 ^ n18654 ;
  assign n18740 = n18739 ^ n18724 ;
  assign n18741 = n18740 ^ n18654 ;
  assign n18319 = ~n17569 & n17650 ;
  assign n18320 = n18319 ^ n17618 ;
  assign n17627 = n17569 ^ n17560 ;
  assign n17628 = n17627 ^ n17621 ;
  assign n17640 = n17639 ^ n17628 ;
  assign n17641 = n17613 & ~n17640 ;
  assign n17642 = n17641 ^ n17621 ;
  assign n17643 = ~n17456 & ~n17642 ;
  assign n18637 = n18320 ^ n17643 ;
  assign n18638 = n18637 ^ n18318 ;
  assign n18639 = n18638 ^ n15502 ;
  assign n18629 = n17682 ^ n17619 ;
  assign n17671 = n17624 ^ n17456 ;
  assign n18621 = n17650 ^ n17489 ;
  assign n18622 = n18621 ^ n17655 ;
  assign n18623 = n18622 ^ n17650 ;
  assign n18626 = ~n17671 & ~n18623 ;
  assign n18627 = n18626 ^ n17650 ;
  assign n18628 = ~n17685 & n18627 ;
  assign n18630 = n17671 & n18628 ;
  assign n18631 = n18629 & n18630 ;
  assign n18632 = n18631 ^ n18628 ;
  assign n18619 = n18618 ^ n17663 ;
  assign n18620 = n17649 & n18619 ;
  assign n18633 = n18632 ^ n18620 ;
  assign n18617 = n17632 & ~n17671 ;
  assign n18634 = n18633 ^ n18617 ;
  assign n18610 = n17619 ^ n17553 ;
  assign n18611 = n18610 ^ n17619 ;
  assign n18614 = n17457 & n18611 ;
  assign n18615 = n18614 ^ n17619 ;
  assign n18616 = n17624 & n18615 ;
  assign n18635 = n18634 ^ n18616 ;
  assign n18636 = ~n18609 & ~n18635 ;
  assign n18640 = n18639 ^ n18636 ;
  assign n18641 = n18640 ^ x69 ;
  assign n18669 = n17869 & ~n17928 ;
  assign n18666 = n17939 ^ n17892 ;
  assign n18667 = n17895 & ~n18666 ;
  assign n18656 = n17924 ^ n17867 ;
  assign n18657 = n17924 ^ n17886 ;
  assign n18658 = n18657 ^ n17891 ;
  assign n18659 = n18658 ^ n18657 ;
  assign n18660 = n18657 ^ n17866 ;
  assign n18661 = n18660 ^ n18657 ;
  assign n18662 = ~n18659 & n18661 ;
  assign n18663 = n18662 ^ n18657 ;
  assign n18664 = n18656 & ~n18663 ;
  assign n18665 = n18664 ^ n17867 ;
  assign n18668 = n18667 ^ n18665 ;
  assign n18670 = n18669 ^ n18668 ;
  assign n18671 = ~n17879 & ~n18670 ;
  assign n18672 = ~n17877 & n18671 ;
  assign n18676 = n17883 ^ n17867 ;
  assign n18673 = n17892 ^ n17831 ;
  assign n18674 = n18673 ^ n17941 ;
  assign n18675 = n17867 & ~n18674 ;
  assign n18677 = n18676 ^ n18675 ;
  assign n18678 = n18675 ^ n17866 ;
  assign n18679 = n18678 ^ n18675 ;
  assign n18680 = n18677 & ~n18679 ;
  assign n18681 = n18680 ^ n18675 ;
  assign n18682 = n18672 & ~n18681 ;
  assign n18683 = ~n17923 & n18682 ;
  assign n18684 = ~n17872 & n18683 ;
  assign n18685 = n18684 ^ n15131 ;
  assign n18686 = n18685 ^ x126 ;
  assign n18742 = n18641 & n18686 ;
  assign n18743 = n18742 ^ n18641 ;
  assign n18744 = n18743 ^ n18686 ;
  assign n18772 = n18741 & ~n18744 ;
  assign n18760 = n18739 & n18743 ;
  assign n18752 = n18741 & n18743 ;
  assign n18761 = n18760 ^ n18752 ;
  assign n18758 = n18738 & n18743 ;
  assign n18759 = n18758 ^ n18743 ;
  assign n18762 = n18761 ^ n18759 ;
  assign n18757 = n18741 & n18742 ;
  assign n18763 = n18762 ^ n18757 ;
  assign n18754 = n18738 & n18742 ;
  assign n18755 = n18754 ^ n18752 ;
  assign n18748 = n18641 & ~n18740 ;
  assign n18756 = n18755 ^ n18748 ;
  assign n18764 = n18763 ^ n18756 ;
  assign n18753 = n18752 ^ n18742 ;
  assign n18765 = n18764 ^ n18753 ;
  assign n18768 = n18765 ^ n18762 ;
  assign n18769 = n18768 ^ n18754 ;
  assign n18773 = n18772 ^ n18769 ;
  assign n18745 = n18744 ^ n18641 ;
  assign n18750 = ~n18740 & n18745 ;
  assign n18749 = n18748 ^ n18740 ;
  assign n18751 = n18750 ^ n18749 ;
  assign n18774 = n18773 ^ n18751 ;
  assign n18771 = n18738 & ~n18744 ;
  assign n18775 = n18774 ^ n18771 ;
  assign n18770 = n18769 ^ n18744 ;
  assign n18776 = n18775 ^ n18770 ;
  assign n18779 = n18776 ^ n18750 ;
  assign n18746 = n18741 & n18745 ;
  assign n18780 = n18779 ^ n18746 ;
  assign n18766 = n18765 ^ n18751 ;
  assign n18735 = n18686 ^ n18654 ;
  assign n18736 = n18641 & n18735 ;
  assign n18655 = n18654 ^ n18641 ;
  assign n18687 = n18686 ^ n18655 ;
  assign n18725 = n18724 ^ n18687 ;
  assign n18726 = n18725 ^ n18641 ;
  assign n18727 = n18726 ^ n18686 ;
  assign n18728 = n18686 ^ n18641 ;
  assign n18731 = ~n18724 & ~n18728 ;
  assign n18732 = n18731 ^ n18641 ;
  assign n18733 = n18727 & ~n18732 ;
  assign n18734 = n18733 ^ n18687 ;
  assign n18737 = n18736 ^ n18734 ;
  assign n18747 = n18746 ^ n18737 ;
  assign n18767 = n18766 ^ n18747 ;
  assign n18777 = n18776 ^ n18767 ;
  assign n18778 = n18777 ^ n18745 ;
  assign n18781 = n18780 ^ n18778 ;
  assign n17420 = n17372 ^ n17338 ;
  assign n18538 = n17447 ^ n17292 ;
  assign n18539 = n18538 ^ n17377 ;
  assign n18540 = n18539 ^ n17338 ;
  assign n18541 = ~n17420 & ~n18540 ;
  assign n18542 = n18541 ^ n17338 ;
  assign n18545 = n17433 ^ n17283 ;
  assign n18546 = n18545 ^ n17278 ;
  assign n18543 = n17283 ^ n17278 ;
  assign n18544 = n18543 ^ n18539 ;
  assign n18547 = n18546 ^ n18544 ;
  assign n18548 = ~n18542 & ~n18547 ;
  assign n18549 = n18548 ^ n18546 ;
  assign n17421 = n17391 ^ n17384 ;
  assign n17422 = n17421 ^ n17391 ;
  assign n17423 = n17391 ^ n17372 ;
  assign n17424 = n17423 ^ n17391 ;
  assign n17425 = n17422 & ~n17424 ;
  assign n17426 = n17425 ^ n17391 ;
  assign n17427 = ~n17420 & n17426 ;
  assign n17428 = n17427 ^ n17391 ;
  assign n18564 = n18549 ^ n17428 ;
  assign n17404 = n17393 ^ n17286 ;
  assign n17405 = n17404 ^ n17389 ;
  assign n17406 = n17389 ^ n17372 ;
  assign n17407 = n17406 ^ n17389 ;
  assign n17408 = ~n17405 & n17407 ;
  assign n17409 = n17408 ^ n17389 ;
  assign n17410 = n17338 & ~n17409 ;
  assign n18565 = n18564 ^ n17410 ;
  assign n18553 = n17200 ^ n17189 ;
  assign n18554 = n18553 ^ n17384 ;
  assign n18555 = n18554 ^ n17291 ;
  assign n18556 = n18555 ^ n17276 ;
  assign n18557 = n18556 ^ n18549 ;
  assign n18552 = n18551 ^ n18549 ;
  assign n18558 = n18557 ^ n18552 ;
  assign n18559 = n18557 ^ n17372 ;
  assign n18560 = n18559 ^ n18557 ;
  assign n18561 = ~n18558 & n18560 ;
  assign n18562 = n18561 ^ n18557 ;
  assign n18563 = ~n17420 & ~n18562 ;
  assign n18566 = n18565 ^ n18563 ;
  assign n18568 = n18567 ^ n18566 ;
  assign n18569 = n18568 ^ n17452 ;
  assign n18570 = n18569 ^ n15461 ;
  assign n18537 = ~n17296 & n17380 ;
  assign n18571 = n18570 ^ n18537 ;
  assign n18572 = n18571 ^ x109 ;
  assign n15097 = n15096 ^ x93 ;
  assign n14627 = n14626 ^ x76 ;
  assign n16103 = n15097 ^ n14627 ;
  assign n15419 = n15418 ^ x94 ;
  assign n15610 = n15601 ^ n15420 ;
  assign n15612 = n15601 ^ n15582 ;
  assign n15611 = n15601 ^ n15573 ;
  assign n15613 = n15612 ^ n15611 ;
  assign n15614 = n15612 ^ n15462 ;
  assign n15615 = n15614 ^ n15612 ;
  assign n15616 = n15613 & n15615 ;
  assign n15617 = n15616 ^ n15612 ;
  assign n15618 = n15610 & n15617 ;
  assign n15619 = n15618 ^ n15420 ;
  assign n15603 = n15602 ^ n15571 ;
  assign n15597 = n15596 ^ n15595 ;
  assign n15604 = n15603 ^ n15597 ;
  assign n15605 = n15597 ^ n15462 ;
  assign n15606 = n15605 ^ n15597 ;
  assign n15607 = ~n15604 & ~n15606 ;
  assign n15608 = n15607 ^ n15597 ;
  assign n15609 = n15420 & n15608 ;
  assign n15620 = n15619 ^ n15609 ;
  assign n15622 = n15621 ^ n15620 ;
  assign n15623 = ~n15577 & n15622 ;
  assign n15625 = n15462 & ~n15589 ;
  assign n15626 = n15625 ^ n15588 ;
  assign n15628 = n15626 ^ n15557 ;
  assign n15627 = n15626 ^ n15592 ;
  assign n15629 = n15628 ^ n15627 ;
  assign n15632 = ~n15462 & ~n15629 ;
  assign n15633 = n15632 ^ n15628 ;
  assign n15634 = n15624 & ~n15633 ;
  assign n15635 = n15634 ^ n15626 ;
  assign n15636 = n15623 & n15635 ;
  assign n15644 = n15636 & ~n15643 ;
  assign n15645 = ~n15576 & n15644 ;
  assign n15646 = n15645 ^ n14918 ;
  assign n15647 = n15646 ^ x69 ;
  assign n15648 = n15419 & ~n15647 ;
  assign n15856 = n15855 ^ x83 ;
  assign n16090 = ~n15992 & ~n16026 ;
  assign n16087 = n16067 & ~n16086 ;
  assign n16082 = n16081 ^ n15989 ;
  assign n16083 = ~n16080 & ~n16082 ;
  assign n16075 = n16074 ^ n15985 ;
  assign n16076 = ~n16027 & ~n16075 ;
  assign n16071 = ~n16064 & n16070 ;
  assign n16077 = n16076 ^ n16071 ;
  assign n16078 = ~n15857 & ~n16077 ;
  assign n16053 = n16052 ^ n16039 ;
  assign n16061 = n16060 ^ n16053 ;
  assign n16062 = n16061 ^ n14879 ;
  assign n16079 = n16078 ^ n16062 ;
  assign n16084 = n16083 ^ n16079 ;
  assign n16031 = n16030 ^ n15965 ;
  assign n16032 = ~n16028 & n16031 ;
  assign n16085 = n16084 ^ n16032 ;
  assign n16088 = n16087 ^ n16085 ;
  assign n15993 = n15992 ^ n15960 ;
  assign n15994 = ~n15857 & ~n15993 ;
  assign n16089 = n16088 ^ n15994 ;
  assign n16091 = n16090 ^ n16089 ;
  assign n16092 = n16091 ^ x117 ;
  assign n16093 = ~n15856 & n16092 ;
  assign n16097 = n16093 ^ n16092 ;
  assign n16138 = n15648 & n16097 ;
  assign n15649 = n15648 ^ n15419 ;
  assign n15650 = n15649 ^ n15647 ;
  assign n15651 = n15650 ^ n15419 ;
  assign n16094 = ~n15651 & n16093 ;
  assign n16132 = n16094 ^ n16093 ;
  assign n16118 = n15648 & n16093 ;
  assign n16108 = n15649 & n16093 ;
  assign n16131 = n16118 ^ n16108 ;
  assign n16133 = n16132 ^ n16131 ;
  assign n16095 = n16093 ^ n15856 ;
  assign n16113 = n16095 ^ n16092 ;
  assign n16130 = n15650 & n16113 ;
  assign n16134 = n16133 ^ n16130 ;
  assign n16163 = n16138 ^ n16134 ;
  assign n16164 = n16138 ^ n15097 ;
  assign n16165 = n16164 ^ n16138 ;
  assign n16166 = n16163 & n16165 ;
  assign n16167 = n16166 ^ n16138 ;
  assign n16168 = n16103 & n16167 ;
  assign n15098 = n14627 & ~n15097 ;
  assign n16098 = ~n15651 & n16097 ;
  assign n16096 = ~n15651 & ~n16095 ;
  assign n16099 = n16098 ^ n16096 ;
  assign n18034 = n16099 ^ n15651 ;
  assign n18035 = n15098 & ~n18034 ;
  assign n16140 = n15648 & n16113 ;
  assign n18004 = n16140 ^ n16108 ;
  assign n18005 = n18004 ^ n16138 ;
  assign n18589 = n15097 & n18005 ;
  assign n15099 = n15098 ^ n15097 ;
  assign n18031 = n16130 ^ n16099 ;
  assign n18032 = ~n15099 & n18031 ;
  assign n16141 = n16140 ^ n16118 ;
  assign n16139 = n16138 ^ n15648 ;
  assign n16142 = n16141 ^ n16139 ;
  assign n16114 = n15649 & n16113 ;
  assign n16143 = n16142 ^ n16114 ;
  assign n18012 = n16143 ^ n16118 ;
  assign n18013 = n15097 & ~n18012 ;
  assign n18014 = n18013 ^ n16118 ;
  assign n18015 = n18014 ^ n14627 ;
  assign n18016 = n18015 ^ n15097 ;
  assign n18017 = n18016 ^ n18014 ;
  assign n16115 = n16114 ^ n16108 ;
  assign n16100 = n16099 ^ n16094 ;
  assign n16101 = n16100 ^ n15651 ;
  assign n16110 = n16101 ^ n16096 ;
  assign n16105 = n16092 ^ n15647 ;
  assign n16106 = n15647 ^ n15419 ;
  assign n16107 = ~n16105 & ~n16106 ;
  assign n16109 = n16108 ^ n16107 ;
  assign n16111 = n16110 ^ n16109 ;
  assign n16112 = n16111 ^ n15649 ;
  assign n16116 = n16115 ^ n16112 ;
  assign n18018 = n16116 ^ n15097 ;
  assign n18019 = n18018 ^ n18014 ;
  assign n18021 = n18019 ^ n16111 ;
  assign n18022 = n18021 ^ n18019 ;
  assign n18025 = n16116 & ~n18022 ;
  assign n18026 = n18018 & n18025 ;
  assign n18027 = n18026 ^ n18018 ;
  assign n18028 = n18027 ^ n18014 ;
  assign n18029 = n18017 & n18028 ;
  assign n18030 = n18029 ^ n18015 ;
  assign n18033 = n18032 ^ n18030 ;
  assign n16102 = n15650 & n16097 ;
  assign n18587 = n18033 ^ n16102 ;
  assign n16150 = n16116 ^ n16111 ;
  assign n16151 = n16150 ^ n16142 ;
  assign n18580 = n16151 ^ n16133 ;
  assign n18583 = n18580 ^ n16118 ;
  assign n17997 = n16134 ^ n16099 ;
  assign n18584 = n18583 ^ n17997 ;
  assign n18585 = n15097 & n18584 ;
  assign n18581 = n18580 ^ n16102 ;
  assign n18582 = n18581 ^ n18033 ;
  assign n18586 = n18585 ^ n18582 ;
  assign n18588 = n18587 ^ n18586 ;
  assign n18590 = n18589 ^ n18588 ;
  assign n18591 = n16103 & n18590 ;
  assign n18592 = n18591 ^ n18586 ;
  assign n18573 = n16102 ^ n14627 ;
  assign n18574 = n18573 ^ n16102 ;
  assign n18577 = n16115 & n18574 ;
  assign n18578 = n18577 ^ n16102 ;
  assign n18579 = ~n15097 & n18578 ;
  assign n18593 = n18592 ^ n18579 ;
  assign n18594 = ~n18035 & ~n18593 ;
  assign n18595 = ~n16168 & n18594 ;
  assign n16129 = n16102 ^ n15650 ;
  assign n16135 = n16134 ^ n16129 ;
  assign n18596 = n16135 ^ n16094 ;
  assign n18597 = n16094 ^ n15097 ;
  assign n18598 = n18597 ^ n16094 ;
  assign n18599 = n18596 & ~n18598 ;
  assign n18600 = n18599 ^ n16094 ;
  assign n18601 = n16103 & n18600 ;
  assign n18602 = n18595 & ~n18601 ;
  assign n18603 = n18602 ^ n15333 ;
  assign n18604 = n18603 ^ x100 ;
  assign n18605 = n18572 & ~n18604 ;
  assign n18606 = n18605 ^ n18604 ;
  assign n19746 = n18606 ^ n18572 ;
  assign n20031 = n18781 & n19746 ;
  assign n20022 = n18604 ^ n18572 ;
  assign n20023 = n18772 ^ n18760 ;
  assign n20024 = n20023 ^ n18772 ;
  assign n20025 = n18772 ^ n18604 ;
  assign n20026 = n20025 ^ n18772 ;
  assign n20027 = n20024 & ~n20026 ;
  assign n20028 = n20027 ^ n18772 ;
  assign n20029 = ~n20022 & n20028 ;
  assign n20030 = n20029 ^ n18772 ;
  assign n20032 = n20031 ^ n20030 ;
  assign n20343 = n18604 & n18737 ;
  assign n20344 = n20343 ^ n18736 ;
  assign n18800 = n18767 ^ n18751 ;
  assign n18811 = n18800 ^ n18776 ;
  assign n18812 = n18605 & ~n18811 ;
  assign n20355 = n20344 ^ n18812 ;
  assign n18784 = n18771 ^ n18746 ;
  assign n20348 = n18784 ^ n18776 ;
  assign n20347 = n18769 ^ n18757 ;
  assign n20349 = n20348 ^ n20347 ;
  assign n20350 = n20349 ^ n20344 ;
  assign n20345 = n20344 ^ n18762 ;
  assign n18801 = n18800 ^ n18757 ;
  assign n18799 = n18760 ^ n18754 ;
  assign n18802 = n18801 ^ n18799 ;
  assign n20346 = n20345 ^ n18802 ;
  assign n20351 = n20350 ^ n20346 ;
  assign n20352 = n18604 & ~n20351 ;
  assign n20353 = n20352 ^ n20350 ;
  assign n20354 = ~n18572 & n20353 ;
  assign n20356 = n20355 ^ n20354 ;
  assign n20357 = ~n20032 & ~n20356 ;
  assign n20358 = n20357 ^ n17188 ;
  assign n20755 = n20358 ^ x74 ;
  assign n20756 = n20754 & n20755 ;
  assign n20757 = n20756 ^ n20754 ;
  assign n18965 = n18649 ^ n18047 ;
  assign n18966 = n18965 ^ n18652 ;
  assign n18967 = n18966 ^ n18647 ;
  assign n18968 = n18967 ^ n14801 ;
  assign n18969 = n18968 ^ x91 ;
  assign n18850 = n17158 ^ n17126 ;
  assign n18840 = n17116 ^ n17105 ;
  assign n18841 = n18840 ^ n17107 ;
  assign n18851 = n18850 ^ n18841 ;
  assign n18852 = n17150 & ~n18851 ;
  assign n18839 = n17098 ^ n17077 ;
  assign n18842 = n18841 ^ n18839 ;
  assign n18416 = n17128 ^ n17090 ;
  assign n18843 = n18842 ^ n18416 ;
  assign n18844 = ~n17081 & n18843 ;
  assign n18835 = n17107 ^ n17088 ;
  assign n18830 = n17157 ^ n17107 ;
  assign n17115 = n17081 ^ n17080 ;
  assign n18831 = n17157 ^ n17081 ;
  assign n18832 = n17115 & n18831 ;
  assign n18833 = n18832 ^ n17081 ;
  assign n18834 = ~n18830 & n18833 ;
  assign n18836 = n18835 ^ n18834 ;
  assign n18838 = n18836 ^ n17104 ;
  assign n18845 = n18844 ^ n18838 ;
  assign n18846 = n17134 & n18845 ;
  assign n18837 = n18836 ^ n17966 ;
  assign n18847 = n18846 ^ n18837 ;
  assign n18848 = n18847 ^ n17126 ;
  assign n18849 = n18848 ^ n16286 ;
  assign n18853 = n18852 ^ n18849 ;
  assign n18823 = n17982 ^ n17079 ;
  assign n18822 = n17158 ^ n17100 ;
  assign n18824 = n18823 ^ n18822 ;
  assign n18825 = n18822 ^ n17081 ;
  assign n18826 = n18825 ^ n18822 ;
  assign n18827 = ~n18824 & n18826 ;
  assign n18828 = n18827 ^ n18822 ;
  assign n18829 = ~n17134 & ~n18828 ;
  assign n18854 = n18853 ^ n18829 ;
  assign n18855 = n18854 ^ x116 ;
  assign n18898 = n16716 ^ n16715 ;
  assign n18899 = n18898 ^ n16592 ;
  assign n18896 = n18881 ^ n16721 ;
  assign n18900 = n18899 ^ n18896 ;
  assign n18901 = n16638 & n18900 ;
  assign n18892 = n16696 ^ n16684 ;
  assign n18893 = n18892 ^ n16694 ;
  assign n18894 = n16704 & ~n18893 ;
  assign n18885 = n16705 ^ n16586 ;
  assign n18884 = n16712 ^ n16594 ;
  assign n18886 = n18885 ^ n18884 ;
  assign n18887 = ~n16678 & n18886 ;
  assign n18861 = n16715 ^ n16590 ;
  assign n18858 = n16681 ^ n16594 ;
  assign n16726 = n16694 ^ n16678 ;
  assign n16727 = n16726 ^ n16694 ;
  assign n16728 = n16695 & n16727 ;
  assign n16729 = n16728 ^ n16694 ;
  assign n16730 = ~n16638 & n16729 ;
  assign n18859 = n18858 ^ n16730 ;
  assign n18862 = n18861 ^ n18859 ;
  assign n18863 = n18862 ^ n16730 ;
  assign n18864 = ~n16678 & n18863 ;
  assign n16759 = n16586 & n16704 ;
  assign n16760 = n16759 ^ n16758 ;
  assign n18860 = n18859 ^ n16760 ;
  assign n18865 = n18864 ^ n18860 ;
  assign n18880 = n18865 ^ n16760 ;
  assign n18882 = n18881 ^ n18880 ;
  assign n18883 = n18882 ^ n16730 ;
  assign n18888 = n18887 ^ n18883 ;
  assign n18889 = n18888 ^ n16696 ;
  assign n18890 = n16679 & ~n18889 ;
  assign n18867 = n18866 ^ n18865 ;
  assign n18878 = n18877 ^ n18867 ;
  assign n18879 = n18878 ^ n16240 ;
  assign n18891 = n18890 ^ n18879 ;
  assign n18895 = n18894 ^ n18891 ;
  assign n18897 = n18896 ^ n18895 ;
  assign n18902 = n18901 ^ n18897 ;
  assign n18903 = n18902 ^ n18895 ;
  assign n18856 = n16679 & n16684 ;
  assign n18857 = n16696 & n18856 ;
  assign n18904 = n18903 ^ n18857 ;
  assign n18905 = n16678 & n18904 ;
  assign n18906 = n18905 ^ n18902 ;
  assign n18907 = n18906 ^ x101 ;
  assign n18908 = n18855 & n18907 ;
  assign n18947 = n18908 ^ n18855 ;
  assign n18924 = n16966 ^ n16935 ;
  assign n18925 = n18924 ^ n16964 ;
  assign n18926 = ~n16809 & n18925 ;
  assign n18927 = n18926 ^ n16966 ;
  assign n18931 = n18927 ^ n17027 ;
  assign n18922 = n16972 ^ n16964 ;
  assign n18923 = n18922 ^ n16983 ;
  assign n18928 = n18927 ^ n18923 ;
  assign n18921 = n16809 & n16970 ;
  assign n18929 = n18928 ^ n18921 ;
  assign n18930 = ~n16766 & ~n18929 ;
  assign n18932 = n18931 ^ n18930 ;
  assign n18933 = n18932 ^ n16949 ;
  assign n18920 = n16809 & n16937 ;
  assign n18934 = n18933 ^ n18920 ;
  assign n18917 = n16975 & n18707 ;
  assign n18918 = n18917 ^ n16949 ;
  assign n18919 = ~n16992 & n18918 ;
  assign n18935 = n18934 ^ n18919 ;
  assign n18936 = n18935 ^ n16947 ;
  assign n18912 = n16947 ^ n16766 ;
  assign n18913 = n18912 ^ n16947 ;
  assign n18914 = n16960 & ~n18913 ;
  assign n18915 = n18914 ^ n16947 ;
  assign n18916 = n16809 & n18915 ;
  assign n18937 = n18936 ^ n18916 ;
  assign n18909 = ~n16992 & ~n18691 ;
  assign n18938 = n18937 ^ n18909 ;
  assign n18939 = ~n18716 & ~n18938 ;
  assign n18940 = ~n16962 & n18939 ;
  assign n18941 = ~n16961 & n18940 ;
  assign n18942 = n18941 ^ n14677 ;
  assign n18943 = n18942 ^ x78 ;
  assign n18944 = n18571 ^ x67 ;
  assign n18945 = ~n18943 & ~n18944 ;
  assign n18949 = n18945 ^ n18943 ;
  assign n18991 = n18949 ^ n18944 ;
  assign n18993 = n18947 & ~n18991 ;
  assign n18976 = n18945 ^ n18944 ;
  assign n18988 = n18908 & ~n18976 ;
  assign n20780 = n18993 ^ n18988 ;
  assign n18952 = n18908 ^ n18907 ;
  assign n18977 = n18952 & ~n18976 ;
  assign n20781 = n20780 ^ n18977 ;
  assign n20782 = n18969 & n20781 ;
  assign n18821 = n18640 ^ x77 ;
  assign n20779 = n18821 & n18977 ;
  assign n20783 = n20782 ^ n20779 ;
  assign n18975 = ~n18821 & ~n18969 ;
  assign n18990 = n18975 ^ n18821 ;
  assign n19023 = n18990 ^ n18969 ;
  assign n18981 = n18947 & ~n18949 ;
  assign n18957 = n18947 ^ n18907 ;
  assign n18958 = n18945 & ~n18957 ;
  assign n18953 = ~n18949 & n18952 ;
  assign n18959 = n18958 ^ n18953 ;
  assign n18950 = n18908 & ~n18949 ;
  assign n18960 = n18959 ^ n18950 ;
  assign n18982 = n18981 ^ n18960 ;
  assign n18980 = n18958 ^ n18949 ;
  assign n18983 = n18982 ^ n18980 ;
  assign n18984 = n18983 ^ n18958 ;
  assign n20775 = n18984 ^ n18957 ;
  assign n20776 = ~n19023 & n20775 ;
  assign n18948 = n18945 & n18947 ;
  assign n18951 = n18950 ^ n18948 ;
  assign n18954 = n18953 ^ n18951 ;
  assign n18946 = n18908 & n18945 ;
  assign n18955 = n18954 ^ n18946 ;
  assign n18956 = n18955 ^ n18945 ;
  assign n20767 = n18956 ^ n18944 ;
  assign n19009 = n18907 ^ n18855 ;
  assign n20768 = n20767 ^ n19009 ;
  assign n20769 = ~n18821 & ~n20768 ;
  assign n20770 = n20769 ^ n18951 ;
  assign n20771 = ~n18969 & n20770 ;
  assign n20772 = n20771 ^ n18951 ;
  assign n19008 = n18969 ^ n18821 ;
  assign n18992 = n18908 & ~n18991 ;
  assign n20760 = n18992 ^ n18984 ;
  assign n18994 = n18981 ^ n18948 ;
  assign n20759 = n18994 ^ n18959 ;
  assign n20761 = n20760 ^ n20759 ;
  assign n20762 = n20760 ^ n18821 ;
  assign n20763 = n20762 ^ n20760 ;
  assign n20764 = ~n20761 & n20763 ;
  assign n20765 = n20764 ^ n20760 ;
  assign n20766 = n19008 & ~n20765 ;
  assign n20773 = n20772 ^ n20766 ;
  assign n18961 = n18960 ^ n18956 ;
  assign n19030 = n18983 ^ n18961 ;
  assign n19048 = ~n19023 & ~n19030 ;
  assign n20774 = n20773 ^ n19048 ;
  assign n20777 = n20776 ^ n20774 ;
  assign n18995 = n18994 ^ n18947 ;
  assign n18996 = n18995 ^ n18993 ;
  assign n18978 = ~n18957 & ~n18976 ;
  assign n18979 = n18978 ^ n18957 ;
  assign n18985 = n18984 ^ n18979 ;
  assign n18997 = n18996 ^ n18985 ;
  assign n18998 = n18997 ^ n18992 ;
  assign n18999 = n18998 ^ n18995 ;
  assign n19000 = n18999 ^ n18991 ;
  assign n19005 = n18975 ^ n18969 ;
  assign n20758 = ~n19000 & ~n19005 ;
  assign n20778 = n20777 ^ n20758 ;
  assign n20784 = n20783 ^ n20778 ;
  assign n19006 = n18997 & ~n19005 ;
  assign n20785 = n20784 ^ n19006 ;
  assign n20786 = n20785 ^ n17275 ;
  assign n20787 = n20786 ^ x120 ;
  assign n18177 = n18142 ^ n18134 ;
  assign n18178 = n18075 & n18177 ;
  assign n18179 = n18178 ^ n18141 ;
  assign n18147 = n18146 ^ n18138 ;
  assign n18165 = n18164 ^ n18147 ;
  assign n18385 = n18179 ^ n18165 ;
  assign n18386 = n18047 & n18385 ;
  assign n18387 = n18386 ^ n18165 ;
  assign n18389 = n18387 ^ n18160 ;
  assign n18388 = n18387 ^ n18155 ;
  assign n18390 = n18389 ^ n18388 ;
  assign n18393 = ~n18047 & n18390 ;
  assign n18394 = n18393 ^ n18389 ;
  assign n18395 = n18167 & ~n18394 ;
  assign n18396 = n18395 ^ n18387 ;
  assign n18397 = ~n18157 & n18396 ;
  assign n18398 = n18397 ^ n15151 ;
  assign n18399 = n18398 ^ x97 ;
  assign n16119 = n16118 ^ n16100 ;
  assign n16117 = n16116 ^ n16108 ;
  assign n16120 = n16119 ^ n16117 ;
  assign n16121 = n16119 ^ n14627 ;
  assign n16122 = n16121 ^ n16119 ;
  assign n16123 = ~n16120 & n16122 ;
  assign n16124 = n16123 ^ n16119 ;
  assign n16125 = ~n15097 & n16124 ;
  assign n16126 = n16125 ^ n16118 ;
  assign n16104 = n16102 & ~n16103 ;
  assign n16127 = n16126 ^ n16104 ;
  assign n16153 = n15419 & ~n16105 ;
  assign n16152 = n16151 ^ n16140 ;
  assign n16154 = n16153 ^ n16152 ;
  assign n16155 = n15097 & n16154 ;
  assign n16156 = n16155 ^ n16153 ;
  assign n16145 = n16134 ^ n16110 ;
  assign n16157 = n16156 ^ n16145 ;
  assign n16147 = n15099 & ~n16138 ;
  assign n16144 = n16143 ^ n16108 ;
  assign n16146 = n16145 ^ n16144 ;
  assign n16148 = n16147 ^ n16146 ;
  assign n16149 = n15097 & n16148 ;
  assign n16158 = n16157 ^ n16149 ;
  assign n16159 = n16103 & ~n16158 ;
  assign n16160 = n16159 ^ n16156 ;
  assign n16128 = n15098 ^ n14627 ;
  assign n16136 = n16135 ^ n16098 ;
  assign n16137 = n16128 & n16136 ;
  assign n16161 = n16160 ^ n16137 ;
  assign n16162 = ~n16127 & ~n16161 ;
  assign n16169 = n16162 & ~n16168 ;
  assign n16172 = n16169 ^ n15924 ;
  assign n15100 = n15099 ^ n14627 ;
  assign n16170 = ~n16101 & n16169 ;
  assign n16171 = n15100 & n16170 ;
  assign n16173 = n16172 ^ n16171 ;
  assign n18400 = n16173 ^ x66 ;
  assign n18401 = n18399 & n18400 ;
  assign n18439 = n18401 ^ n18399 ;
  assign n18345 = n17456 & ~n17638 ;
  assign n18337 = n17630 ^ n17619 ;
  assign n18338 = n18337 ^ n17632 ;
  assign n18339 = n18338 ^ n17671 ;
  assign n18340 = ~n17565 & n18339 ;
  assign n18341 = n18340 ^ n17671 ;
  assign n18342 = n17649 ^ n17565 ;
  assign n18343 = n18341 & n18342 ;
  assign n18322 = n17637 ^ n17565 ;
  assign n17651 = n17559 & n17650 ;
  assign n17644 = n17613 ^ n17513 ;
  assign n17645 = n17491 & n17644 ;
  assign n17646 = n17552 ^ n17456 ;
  assign n17647 = ~n17563 & n17646 ;
  assign n17648 = n17645 & n17647 ;
  assign n17652 = n17651 ^ n17648 ;
  assign n18321 = n18320 ^ n17652 ;
  assign n18323 = n18322 ^ n18321 ;
  assign n18334 = n18333 ^ n18323 ;
  assign n18335 = n18334 ^ n18318 ;
  assign n18336 = n18335 ^ n15953 ;
  assign n18344 = n18343 ^ n18336 ;
  assign n18346 = n18345 ^ n18344 ;
  assign n18303 = n17638 ^ n17637 ;
  assign n18304 = n18303 ^ n17638 ;
  assign n18305 = n18304 ^ n17683 ;
  assign n18306 = n18305 ^ n18303 ;
  assign n18307 = n18303 ^ n17456 ;
  assign n18308 = n18307 ^ n18303 ;
  assign n18309 = n18306 & ~n18308 ;
  assign n18310 = n18309 ^ n18303 ;
  assign n18311 = n17613 & n18310 ;
  assign n18347 = n18346 ^ n18311 ;
  assign n18348 = n18347 ^ x106 ;
  assign n18379 = n17868 & ~n17926 ;
  assign n18372 = n17936 ^ n17876 ;
  assign n18373 = n18372 ^ n17909 ;
  assign n18356 = n17939 ^ n17885 ;
  assign n18374 = n18373 ^ n18356 ;
  assign n18375 = n17867 & n18374 ;
  assign n18370 = n18356 ^ n17876 ;
  assign n18364 = n17892 ^ n17830 ;
  assign n18365 = n18364 ^ n17907 ;
  assign n18366 = n17867 & ~n18365 ;
  assign n18367 = n18366 ^ n17938 ;
  assign n18371 = n18370 ^ n18367 ;
  assign n18376 = n18375 ^ n18371 ;
  assign n18377 = ~n17866 & ~n18376 ;
  assign n18363 = n17949 ^ n17894 ;
  assign n18368 = n18367 ^ n18363 ;
  assign n18369 = n18368 ^ n15888 ;
  assign n18378 = n18377 ^ n18369 ;
  assign n18380 = n18379 ^ n18378 ;
  assign n18355 = n17875 ^ n17869 ;
  assign n18357 = n18356 ^ n17871 ;
  assign n18360 = ~n17875 & n18357 ;
  assign n18361 = n18360 ^ n17871 ;
  assign n18362 = n18355 & n18361 ;
  assign n18381 = n18380 ^ n18362 ;
  assign n18349 = n17922 ^ n17888 ;
  assign n18350 = n17888 ^ n17867 ;
  assign n18351 = n18350 ^ n17888 ;
  assign n18352 = ~n18349 & ~n18351 ;
  assign n18353 = n18352 ^ n17888 ;
  assign n18354 = ~n17866 & ~n18353 ;
  assign n18382 = n18381 ^ n18354 ;
  assign n18383 = n18382 ^ x80 ;
  assign n18384 = n18348 & n18383 ;
  assign n18440 = n18384 ^ n18348 ;
  assign n18454 = n18439 & n18440 ;
  assign n18432 = n17966 ^ n15281 ;
  assign n18433 = n18432 ^ n17981 ;
  assign n18415 = n17088 ^ n17085 ;
  assign n18417 = n18416 ^ n17108 ;
  assign n18418 = n18417 ^ n17083 ;
  assign n18420 = n17085 & n18418 ;
  assign n18421 = n18420 ^ n17083 ;
  assign n18422 = n18415 & n18421 ;
  assign n18423 = n18422 ^ n17088 ;
  assign n18408 = n17974 ^ n17098 ;
  assign n18409 = n18408 ^ n17096 ;
  assign n18410 = n17096 ^ n17080 ;
  assign n18411 = n18410 ^ n17096 ;
  assign n18412 = n18409 & n18411 ;
  assign n18413 = n18412 ^ n17096 ;
  assign n18414 = ~n17081 & n18413 ;
  assign n18424 = n18423 ^ n18414 ;
  assign n17131 = n17130 ^ n17099 ;
  assign n18425 = n17131 ^ n17080 ;
  assign n18426 = n18425 ^ n17131 ;
  assign n18427 = n17081 & ~n17976 ;
  assign n18428 = n18427 ^ n17131 ;
  assign n18429 = ~n18426 & n18428 ;
  assign n18430 = n18429 ^ n17131 ;
  assign n18431 = ~n18424 & ~n18430 ;
  assign n18434 = n18433 ^ n18431 ;
  assign n18435 = n18434 ^ x121 ;
  assign n18402 = n18401 ^ n18400 ;
  assign n18441 = n18440 ^ n18383 ;
  assign n18458 = n18402 & ~n18441 ;
  assign n18459 = n18458 ^ n18402 ;
  assign n18451 = n18402 & n18440 ;
  assign n18405 = n18384 & n18402 ;
  assign n18452 = n18451 ^ n18405 ;
  assign n18460 = n18459 ^ n18452 ;
  assign n18403 = n18402 ^ n18399 ;
  assign n18404 = n18384 & ~n18403 ;
  assign n18461 = n18460 ^ n18404 ;
  assign n18444 = ~n18403 & ~n18441 ;
  assign n18462 = n18461 ^ n18444 ;
  assign n18463 = n18462 ^ n18458 ;
  assign n18464 = n18463 ^ n18399 ;
  assign n18450 = ~n18403 & n18440 ;
  assign n18453 = n18452 ^ n18450 ;
  assign n18465 = n18464 ^ n18453 ;
  assign n18466 = n18465 ^ n18460 ;
  assign n17017 = n17016 ^ n17008 ;
  assign n17007 = n16975 ^ n16951 ;
  assign n17018 = n17017 ^ n17007 ;
  assign n17019 = n17018 ^ n17006 ;
  assign n17023 = n17022 ^ n17019 ;
  assign n16995 = n16972 ^ n16951 ;
  assign n16996 = n16995 ^ n16947 ;
  assign n16997 = n16996 ^ n16951 ;
  assign n16998 = n16994 & ~n16997 ;
  assign n16999 = n16998 ^ n16951 ;
  assign n17000 = ~n16992 & n16999 ;
  assign n17024 = n17023 ^ n17000 ;
  assign n16985 = n16984 ^ n16960 ;
  assign n16986 = n16985 ^ n16959 ;
  assign n16987 = n16959 ^ n16809 ;
  assign n16988 = n16987 ^ n16959 ;
  assign n16989 = ~n16986 & ~n16988 ;
  assign n16990 = n16989 ^ n16959 ;
  assign n16991 = ~n16766 & ~n16990 ;
  assign n17025 = n17024 ^ n16991 ;
  assign n16976 = n16975 ^ n16969 ;
  assign n16977 = n16976 ^ n16975 ;
  assign n16978 = n16975 ^ n16766 ;
  assign n16979 = n16978 ^ n16975 ;
  assign n16980 = ~n16977 & n16979 ;
  assign n16981 = n16980 ^ n16975 ;
  assign n16982 = ~n16809 & n16981 ;
  assign n17026 = n17025 ^ n16982 ;
  assign n17028 = n17027 ^ n17026 ;
  assign n17029 = ~n16962 & ~n17028 ;
  assign n17030 = ~n16961 & n17029 ;
  assign n17031 = n17030 ^ n16025 ;
  assign n18407 = n17031 ^ x99 ;
  assign n18527 = n18460 ^ n18407 ;
  assign n18528 = n18527 ^ n18460 ;
  assign n19800 = ~n18466 & n18528 ;
  assign n19801 = n19800 ^ n18460 ;
  assign n19802 = n18435 & n19801 ;
  assign n18525 = n18435 ^ n18407 ;
  assign n18447 = n18401 & ~n18441 ;
  assign n18526 = n18460 ^ n18447 ;
  assign n18529 = n18526 & n18528 ;
  assign n18530 = n18529 ^ n18460 ;
  assign n18531 = ~n18525 & n18530 ;
  assign n20014 = n19802 ^ n18531 ;
  assign n18442 = n18441 ^ n18348 ;
  assign n18443 = n18439 & n18442 ;
  assign n18457 = n18443 ^ n18442 ;
  assign n18467 = n18466 ^ n18457 ;
  assign n18455 = n18454 ^ n18453 ;
  assign n18449 = n18440 ^ n18405 ;
  assign n18456 = n18455 ^ n18449 ;
  assign n18468 = n18467 ^ n18456 ;
  assign n18448 = n18447 ^ n18401 ;
  assign n18469 = n18468 ^ n18448 ;
  assign n18476 = n18469 ^ n18384 ;
  assign n18406 = n18405 ^ n18404 ;
  assign n18477 = n18476 ^ n18406 ;
  assign n18478 = n18477 ^ n18451 ;
  assign n20001 = ~n18407 & ~n18478 ;
  assign n20000 = n18452 ^ n18444 ;
  assign n20002 = n20001 ^ n20000 ;
  assign n20015 = n20014 ^ n20002 ;
  assign n18436 = ~n18407 & ~n18435 ;
  assign n19804 = n18436 ^ n18435 ;
  assign n19807 = n18443 & ~n19804 ;
  assign n19805 = n18450 ^ n18447 ;
  assign n19806 = ~n19804 & n19805 ;
  assign n19808 = n19807 ^ n19806 ;
  assign n20016 = n20015 ^ n19808 ;
  assign n18479 = ~n18435 & ~n18478 ;
  assign n18480 = n18479 ^ n18451 ;
  assign n18483 = n18480 ^ n18443 ;
  assign n18484 = n18483 ^ n18480 ;
  assign n18485 = n18435 & n18484 ;
  assign n18486 = n18485 ^ n18480 ;
  assign n18487 = ~n18407 & n18486 ;
  assign n18488 = n18487 ^ n18480 ;
  assign n18437 = n18436 ^ n18407 ;
  assign n18471 = n18439 & ~n18441 ;
  assign n18474 = n18471 ^ n18456 ;
  assign n18475 = ~n18437 & n18474 ;
  assign n18489 = n18488 ^ n18475 ;
  assign n20017 = n20016 ^ n18489 ;
  assign n20008 = n18467 ^ n18450 ;
  assign n19778 = n18458 ^ n18406 ;
  assign n20009 = n20008 ^ n19778 ;
  assign n20006 = n18469 ^ n18465 ;
  assign n20005 = n18474 ^ n18458 ;
  assign n20007 = n20006 ^ n20005 ;
  assign n20010 = n20009 ^ n20007 ;
  assign n20011 = ~n18407 & ~n20010 ;
  assign n20003 = n20002 ^ n18467 ;
  assign n20004 = n20003 ^ n19778 ;
  assign n20012 = n20011 ^ n20004 ;
  assign n20013 = ~n18525 & ~n20012 ;
  assign n20018 = n20017 ^ n20013 ;
  assign n20019 = ~n18454 & ~n20018 ;
  assign n20020 = n20019 ^ n17232 ;
  assign n20788 = n20020 ^ x65 ;
  assign n20789 = ~n20787 & ~n20788 ;
  assign n20790 = n20789 ^ n20788 ;
  assign n20815 = n20757 & ~n20790 ;
  assign n20791 = n20790 ^ n20787 ;
  assign n20793 = n20791 ^ n20788 ;
  assign n20794 = n20756 & ~n20793 ;
  assign n20816 = n20815 ^ n20794 ;
  assign n20803 = n20756 & n20789 ;
  assign n20802 = n20757 & n20789 ;
  assign n20804 = n20803 ^ n20802 ;
  assign n20805 = n20804 ^ n20789 ;
  assign n20796 = n20757 ^ n20755 ;
  assign n20800 = n20796 ^ n20754 ;
  assign n20801 = n20789 & n20800 ;
  assign n20806 = n20805 ^ n20801 ;
  assign n20799 = ~n20791 & ~n20796 ;
  assign n20807 = n20806 ^ n20799 ;
  assign n20797 = ~n20790 & ~n20796 ;
  assign n20798 = n20797 ^ n20796 ;
  assign n20808 = n20807 ^ n20798 ;
  assign n20817 = n20816 ^ n20808 ;
  assign n20818 = n20817 ^ n20807 ;
  assign n20810 = n20787 ^ n20755 ;
  assign n20811 = n20788 ^ n20787 ;
  assign n20812 = ~n20810 & ~n20811 ;
  assign n20813 = n20812 ^ n20788 ;
  assign n20814 = n20813 ^ n20757 ;
  assign n20819 = n20818 ^ n20814 ;
  assign n20792 = n20757 & ~n20791 ;
  assign n20820 = n20819 ^ n20792 ;
  assign n20821 = n20820 ^ n20793 ;
  assign n20795 = n20794 ^ n20792 ;
  assign n20809 = n20808 ^ n20795 ;
  assign n20822 = n20821 ^ n20809 ;
  assign n20823 = n20822 ^ n20819 ;
  assign n16174 = n16173 ^ x115 ;
  assign n16733 = n16730 ^ n16705 ;
  assign n16731 = n16721 ^ n16586 ;
  assign n16732 = n16703 & n16731 ;
  assign n16734 = n16733 ^ n16732 ;
  assign n16735 = n16734 ^ n16730 ;
  assign n16722 = n16721 ^ n16682 ;
  assign n16723 = n16678 & n16722 ;
  assign n16736 = n16735 ^ n16723 ;
  assign n16737 = ~n16638 & n16736 ;
  assign n16738 = n16737 ^ n16734 ;
  assign n16719 = n16703 ^ n16678 ;
  assign n16720 = n16718 & ~n16719 ;
  assign n16739 = n16738 ^ n16720 ;
  assign n16710 = n16709 ^ n16590 ;
  assign n16713 = n16712 ^ n16710 ;
  assign n16714 = n16704 & n16713 ;
  assign n16740 = n16739 ^ n16714 ;
  assign n16697 = n16696 ^ n16592 ;
  assign n16700 = n16638 & ~n16697 ;
  assign n16701 = n16700 ^ n16592 ;
  assign n16702 = n16679 & n16701 ;
  assign n16741 = n16740 ^ n16702 ;
  assign n16742 = n16741 ^ n16684 ;
  assign n16751 = n16750 ^ n16742 ;
  assign n16761 = n16760 ^ n16751 ;
  assign n16685 = n16684 ^ n16683 ;
  assign n16686 = n16685 ^ n16684 ;
  assign n16687 = n16684 ^ n16638 ;
  assign n16688 = n16687 ^ n16684 ;
  assign n16689 = n16686 & ~n16688 ;
  assign n16690 = n16689 ^ n16684 ;
  assign n16691 = ~n16679 & n16690 ;
  assign n16762 = n16761 ^ n16691 ;
  assign n16763 = ~n16594 & ~n16762 ;
  assign n16764 = n16763 ^ n15706 ;
  assign n16765 = n16764 ^ x88 ;
  assign n17453 = n17452 ^ n16441 ;
  assign n17432 = n17389 ^ n17278 ;
  assign n17434 = n17433 ^ n17432 ;
  assign n17435 = n17372 & ~n17434 ;
  assign n17436 = n17435 ^ n17417 ;
  assign n17437 = n17338 & n17436 ;
  assign n17418 = n17417 ^ n17416 ;
  assign n17419 = n17418 ^ n17410 ;
  assign n17429 = n17428 ^ n17419 ;
  assign n17399 = n17398 ^ n17377 ;
  assign n17396 = n17395 ^ n17377 ;
  assign n17397 = n17396 ^ n17294 ;
  assign n17400 = n17399 ^ n17397 ;
  assign n17401 = n17372 & n17400 ;
  assign n17402 = n17401 ^ n17399 ;
  assign n17403 = ~n17338 & n17402 ;
  assign n17430 = n17429 ^ n17403 ;
  assign n17386 = n17384 & n17385 ;
  assign n17431 = n17430 ^ n17386 ;
  assign n17438 = n17437 ^ n17431 ;
  assign n17381 = ~n17379 & n17380 ;
  assign n17439 = n17438 ^ n17381 ;
  assign n17440 = ~n17375 & ~n17439 ;
  assign n17454 = n17453 ^ n17440 ;
  assign n17455 = n17454 ^ x113 ;
  assign n17691 = n17567 ^ n17562 ;
  assign n17664 = n17663 ^ n17567 ;
  assign n17677 = n17650 & n17664 ;
  assign n17666 = n17665 ^ n17561 ;
  assign n17672 = n17619 & ~n17671 ;
  assign n17669 = ~n17639 & n17649 ;
  assign n17667 = n17636 ^ n17561 ;
  assign n17668 = n17667 ^ n17629 ;
  assign n17670 = n17669 ^ n17668 ;
  assign n17673 = n17672 ^ n17670 ;
  assign n17674 = ~n17666 & ~n17673 ;
  assign n17675 = n17674 ^ n17665 ;
  assign n17678 = n17677 ^ n17675 ;
  assign n17692 = n17649 & n17678 ;
  assign n17693 = n17691 & n17692 ;
  assign n17690 = n17689 ^ n17678 ;
  assign n17694 = n17693 ^ n17690 ;
  assign n17656 = n17655 ^ n17565 ;
  assign n17659 = ~n17613 & n17656 ;
  assign n17660 = n17659 ^ n17565 ;
  assign n17661 = ~n17456 & n17660 ;
  assign n17695 = n17694 ^ n17661 ;
  assign n17696 = ~n17652 & n17695 ;
  assign n17697 = ~n17643 & n17696 ;
  assign n17698 = ~n17626 & n17697 ;
  assign n17699 = n17698 ^ n15683 ;
  assign n17700 = n17699 ^ x65 ;
  assign n17153 = n17085 & n17107 ;
  assign n17151 = n17127 & n17150 ;
  assign n17146 = n17080 & n17105 ;
  assign n17141 = n17093 ^ n17091 ;
  assign n17132 = n17131 ^ n17100 ;
  assign n17142 = n17141 ^ n17132 ;
  assign n17135 = n17127 ^ n17093 ;
  assign n17138 = n17137 ^ n17135 ;
  assign n17139 = n17138 ^ n17091 ;
  assign n17140 = ~n17081 & n17139 ;
  assign n17143 = n17142 ^ n17140 ;
  assign n17144 = n17134 & n17143 ;
  assign n17133 = n17132 ^ n17120 ;
  assign n17145 = n17144 ^ n17133 ;
  assign n17147 = n17146 ^ n17145 ;
  assign n17117 = n17116 ^ n17081 ;
  assign n17118 = n17117 ^ n17116 ;
  assign n17123 = n17118 & n17120 ;
  assign n17124 = n17123 ^ n17116 ;
  assign n17125 = n17115 & n17124 ;
  assign n17148 = n17147 ^ n17125 ;
  assign n17149 = n17148 ^ n17079 ;
  assign n17152 = n17151 ^ n17149 ;
  assign n17154 = n17153 ^ n17152 ;
  assign n17084 = n17083 ^ n17079 ;
  assign n17109 = n17108 ^ n17085 ;
  assign n17110 = n17108 ^ n17079 ;
  assign n17111 = n17110 ^ n17108 ;
  assign n17112 = ~n17109 & n17111 ;
  assign n17113 = n17112 ^ n17108 ;
  assign n17114 = ~n17084 & n17113 ;
  assign n17155 = n17154 ^ n17114 ;
  assign n17160 = n17159 ^ n17155 ;
  assign n17161 = n17160 ^ n16417 ;
  assign n17162 = n17161 ^ x120 ;
  assign n17032 = n17031 ^ x74 ;
  assign n17714 = n17162 ^ n17032 ;
  assign n17715 = ~n17700 & n17714 ;
  assign n17163 = ~n17032 & n17162 ;
  assign n17719 = n17715 ^ n17163 ;
  assign n17720 = n17719 ^ n17162 ;
  assign n17703 = n17163 & ~n17700 ;
  assign n17718 = n17703 ^ n17032 ;
  assign n17721 = n17720 ^ n17718 ;
  assign n17722 = n17455 & n17721 ;
  assign n17723 = n17722 ^ n17721 ;
  assign n17707 = n17032 & ~n17455 ;
  assign n17724 = n17723 ^ n17707 ;
  assign n17701 = n17455 & ~n17700 ;
  assign n17710 = ~n17162 & n17701 ;
  assign n17711 = ~n17032 & n17710 ;
  assign n17712 = n17711 ^ n17710 ;
  assign n17713 = n17712 ^ n17703 ;
  assign n17716 = n17715 ^ n17713 ;
  assign n17708 = n17162 & n17700 ;
  assign n17709 = n17707 & n17708 ;
  assign n17717 = n17716 ^ n17709 ;
  assign n17725 = n17724 ^ n17717 ;
  assign n17726 = n17725 ^ n17722 ;
  assign n17704 = n17703 ^ n17163 ;
  assign n17702 = n17163 & n17701 ;
  assign n17705 = n17704 ^ n17702 ;
  assign n17706 = n17705 ^ n17163 ;
  assign n17727 = n17726 ^ n17706 ;
  assign n17728 = n16765 & n17727 ;
  assign n17729 = n17728 ^ n17726 ;
  assign n17730 = ~n16174 & n17729 ;
  assign n17733 = n17708 ^ n17700 ;
  assign n17734 = n17733 ^ n17162 ;
  assign n17735 = n17734 ^ n17710 ;
  assign n17736 = n17735 ^ n17716 ;
  assign n17731 = n17710 ^ n17701 ;
  assign n17732 = n17731 ^ n17702 ;
  assign n17737 = n17736 ^ n17732 ;
  assign n17738 = n17736 ^ n16174 ;
  assign n17739 = n17738 ^ n17736 ;
  assign n17740 = ~n17737 & ~n17739 ;
  assign n17741 = n17740 ^ n17736 ;
  assign n17742 = n16765 & ~n17741 ;
  assign n20422 = n17716 ^ n17711 ;
  assign n20423 = ~n16174 & n20422 ;
  assign n20424 = n20423 ^ n17711 ;
  assign n20427 = n20424 ^ n17702 ;
  assign n20428 = n20427 ^ n20424 ;
  assign n20429 = ~n16174 & n20428 ;
  assign n20430 = n20429 ^ n20424 ;
  assign n20431 = ~n16765 & n20430 ;
  assign n20432 = n20431 ^ n20424 ;
  assign n17761 = n16174 & ~n16765 ;
  assign n20404 = n17761 ^ n16765 ;
  assign n20421 = ~n17736 & ~n20404 ;
  assign n20433 = n20432 ^ n20421 ;
  assign n17763 = ~n17455 & n17704 ;
  assign n17764 = n17763 ^ n17704 ;
  assign n17762 = n17736 ^ n17725 ;
  assign n17765 = n17764 ^ n17762 ;
  assign n17766 = n17761 & ~n17765 ;
  assign n17778 = n16765 ^ n16174 ;
  assign n17755 = n17733 ^ n17721 ;
  assign n17756 = n17455 & n17755 ;
  assign n17769 = n17756 ^ n17755 ;
  assign n20407 = n17769 ^ n17763 ;
  assign n17780 = n17723 ^ n17712 ;
  assign n20408 = n20407 ^ n17780 ;
  assign n17757 = n17709 ^ n17708 ;
  assign n17758 = n17757 ^ n17704 ;
  assign n17759 = n17758 ^ n17756 ;
  assign n20409 = n20408 ^ n17759 ;
  assign n20410 = n20409 ^ n20407 ;
  assign n20411 = n20407 ^ n16765 ;
  assign n20412 = n20411 ^ n20407 ;
  assign n20413 = n20410 & ~n20412 ;
  assign n20414 = n20413 ^ n20407 ;
  assign n20415 = n17778 & n20414 ;
  assign n20416 = n20415 ^ n20407 ;
  assign n20405 = n17732 ^ n17723 ;
  assign n20406 = ~n20404 & n20405 ;
  assign n20417 = n20416 ^ n20406 ;
  assign n17748 = n17732 ^ n17709 ;
  assign n20395 = n17748 ^ n17726 ;
  assign n20393 = n17758 ^ n17712 ;
  assign n20392 = n17731 ^ n17455 ;
  assign n20394 = n20393 ^ n20392 ;
  assign n20396 = n20395 ^ n20394 ;
  assign n20399 = n20395 ^ n16174 ;
  assign n20400 = n20399 ^ n20395 ;
  assign n20401 = n20396 & ~n20400 ;
  assign n20402 = n20401 ^ n20395 ;
  assign n20403 = n16765 & n20402 ;
  assign n20418 = n20417 ^ n20403 ;
  assign n20388 = n17709 ^ n17706 ;
  assign n20389 = ~n16765 & n20388 ;
  assign n20390 = n20389 ^ n17709 ;
  assign n20391 = n17778 & n20390 ;
  assign n20419 = n20418 ^ n20391 ;
  assign n20420 = ~n17766 & ~n20419 ;
  assign n20434 = n20433 ^ n20420 ;
  assign n20435 = ~n17742 & n20434 ;
  assign n20436 = ~n17730 & n20435 ;
  assign n20437 = n20436 ^ n17337 ;
  assign n20824 = n20437 ^ x88 ;
  assign n19369 = n19124 ^ x70 ;
  assign n19372 = n18968 ^ x85 ;
  assign n19408 = n17866 & n17924 ;
  assign n19399 = n17885 ^ n17869 ;
  assign n19400 = n17878 ^ n17871 ;
  assign n19403 = ~n17885 & ~n19400 ;
  assign n19404 = n19403 ^ n17871 ;
  assign n19405 = n19399 & n19404 ;
  assign n19396 = n17940 ^ n17926 ;
  assign n19397 = ~n17870 & n19396 ;
  assign n19375 = n17867 ^ n17866 ;
  assign n19376 = n17941 ^ n17937 ;
  assign n19377 = n19376 ^ n17867 ;
  assign n19378 = ~n19375 & ~n19377 ;
  assign n19379 = n19378 ^ n17867 ;
  assign n19380 = n17907 ^ n17892 ;
  assign n19381 = n19380 ^ n17907 ;
  assign n19382 = n19381 ^ n19376 ;
  assign n19383 = n19379 & n19382 ;
  assign n19384 = n19383 ^ n19380 ;
  assign n19393 = n19384 ^ n17930 ;
  assign n19385 = n19384 ^ n19376 ;
  assign n19386 = n19385 ^ n17897 ;
  assign n19387 = n19386 ^ n19384 ;
  assign n19390 = n17867 & n19387 ;
  assign n19391 = n19390 ^ n19384 ;
  assign n19392 = ~n19375 & n19391 ;
  assign n19394 = n19393 ^ n19392 ;
  assign n19374 = n17951 ^ n17869 ;
  assign n19395 = n19394 ^ n19374 ;
  assign n19398 = n19397 ^ n19395 ;
  assign n19406 = n19405 ^ n19398 ;
  assign n19373 = n17867 & n17875 ;
  assign n19407 = n19406 ^ n19373 ;
  assign n19409 = n19408 ^ n19407 ;
  assign n19410 = ~n17872 & ~n19409 ;
  assign n19411 = n19410 ^ n14846 ;
  assign n19412 = n19411 ^ x83 ;
  assign n19413 = ~n19372 & ~n19412 ;
  assign n19441 = n15097 & n16150 ;
  assign n17993 = n16133 ^ n16098 ;
  assign n17994 = n15098 & n17993 ;
  assign n19435 = n17994 ^ n14627 ;
  assign n19428 = n16143 ^ n15099 ;
  assign n19429 = n16141 ^ n16128 ;
  assign n19430 = n16141 ^ n15099 ;
  assign n19431 = n19430 ^ n16141 ;
  assign n19432 = ~n19429 & n19431 ;
  assign n19433 = n19432 ^ n16141 ;
  assign n19434 = ~n19428 & ~n19433 ;
  assign n19436 = n19435 ^ n19434 ;
  assign n19416 = n16147 ^ n16101 ;
  assign n19417 = n16134 ^ n15650 ;
  assign n19418 = n19417 ^ n16128 ;
  assign n19419 = n19416 & n19418 ;
  assign n19420 = n19419 ^ n17993 ;
  assign n19427 = n19420 ^ n18601 ;
  assign n19437 = n19436 ^ n19427 ;
  assign n19438 = n19437 ^ n15010 ;
  assign n19422 = n16138 ^ n16110 ;
  assign n19423 = n19422 ^ n16151 ;
  assign n19424 = ~n15097 & ~n19423 ;
  assign n19415 = n16130 ^ n16110 ;
  assign n19421 = n19420 ^ n19415 ;
  assign n19425 = n19424 ^ n19421 ;
  assign n19426 = n16103 & ~n19425 ;
  assign n19439 = n19438 ^ n19426 ;
  assign n19414 = n15100 & ~n16131 ;
  assign n19440 = n19439 ^ n19414 ;
  assign n19442 = n19441 ^ n19440 ;
  assign n19443 = n19442 ^ x102 ;
  assign n19444 = n19226 ^ x108 ;
  assign n19445 = ~n19443 & n19444 ;
  assign n19456 = n19445 ^ n19444 ;
  assign n19457 = n19456 ^ n19443 ;
  assign n19458 = n19457 ^ n19444 ;
  assign n19505 = n19413 & ~n19458 ;
  assign n19448 = n19413 ^ n19372 ;
  assign n19470 = ~n19448 & n19457 ;
  assign n19450 = n19448 ^ n19412 ;
  assign n19451 = n19450 ^ n19372 ;
  assign n19469 = ~n19451 & n19457 ;
  assign n19471 = n19470 ^ n19469 ;
  assign n19452 = n19445 & ~n19451 ;
  assign n19449 = n19445 & ~n19448 ;
  assign n19453 = n19452 ^ n19449 ;
  assign n19446 = n19413 & n19445 ;
  assign n19447 = n19446 ^ n19445 ;
  assign n19454 = n19453 ^ n19447 ;
  assign n19472 = n19471 ^ n19454 ;
  assign n19462 = n19443 ^ n19412 ;
  assign n19467 = ~n19444 & n19462 ;
  assign n19460 = n19443 ^ n19372 ;
  assign n19461 = n19444 ^ n19412 ;
  assign n19464 = n19443 & ~n19461 ;
  assign n19465 = n19464 ^ n19412 ;
  assign n19466 = n19460 & n19465 ;
  assign n19468 = n19467 ^ n19466 ;
  assign n19473 = n19472 ^ n19468 ;
  assign n19459 = ~n19450 & ~n19458 ;
  assign n19474 = n19473 ^ n19459 ;
  assign n19475 = n19474 ^ n19469 ;
  assign n19476 = n19475 ^ n19467 ;
  assign n19477 = n19476 ^ n19471 ;
  assign n19478 = n19477 ^ n19457 ;
  assign n19506 = n19505 ^ n19478 ;
  assign n19507 = n19506 ^ n19474 ;
  assign n19533 = n19507 ^ n19444 ;
  assign n19534 = n19533 ^ n19477 ;
  assign n19535 = n19534 ^ n19452 ;
  assign n19532 = n19469 ^ n19451 ;
  assign n19536 = n19535 ^ n19532 ;
  assign n19537 = n19536 ^ n19452 ;
  assign n19479 = n19478 ^ n19459 ;
  assign n19455 = n19454 ^ n19450 ;
  assign n19480 = n19479 ^ n19455 ;
  assign n19538 = n19537 ^ n19480 ;
  assign n19370 = n18942 ^ x84 ;
  assign n19539 = n19480 ^ n19370 ;
  assign n19540 = n19539 ^ n19480 ;
  assign n19541 = ~n19538 & ~n19540 ;
  assign n19542 = n19541 ^ n19480 ;
  assign n19543 = n19369 & ~n19542 ;
  assign n19371 = n19370 ^ n19369 ;
  assign n19481 = n19480 ^ n19453 ;
  assign n19482 = n19453 ^ n19370 ;
  assign n19483 = n19482 ^ n19453 ;
  assign n19484 = ~n19481 & ~n19483 ;
  assign n19485 = n19484 ^ n19453 ;
  assign n19486 = ~n19371 & n19485 ;
  assign n20192 = ~n19370 & n19470 ;
  assign n20177 = n19536 ^ n19534 ;
  assign n20178 = n19370 & ~n20177 ;
  assign n20179 = n20178 ^ n19534 ;
  assign n19500 = ~n19448 & n19456 ;
  assign n20182 = n20179 ^ n19500 ;
  assign n20183 = n20182 ^ n20179 ;
  assign n20184 = n19370 & n20183 ;
  assign n20185 = n20184 ^ n20179 ;
  assign n20186 = ~n19369 & ~n20185 ;
  assign n20187 = n20186 ^ n20179 ;
  assign n20148 = n19451 ^ n19449 ;
  assign n20149 = n20148 ^ n19536 ;
  assign n20150 = n20149 ^ n19443 ;
  assign n19487 = n19413 & n19456 ;
  assign n19488 = n19487 ^ n19454 ;
  assign n20147 = n19488 ^ n19473 ;
  assign n20151 = n20150 ^ n20147 ;
  assign n20152 = ~n19370 & n20151 ;
  assign n20153 = n20152 ^ n20150 ;
  assign n20188 = n20187 ^ n20153 ;
  assign n20170 = n19506 ^ n19479 ;
  assign n20171 = n20170 ^ n19478 ;
  assign n20172 = n19478 ^ n19370 ;
  assign n20173 = n20172 ^ n19478 ;
  assign n20174 = n20171 & ~n20173 ;
  assign n20175 = n20174 ^ n19478 ;
  assign n20176 = ~n19371 & n20175 ;
  assign n20189 = n20188 ^ n20176 ;
  assign n20165 = n19459 ^ n19370 ;
  assign n20166 = n20165 ^ n19459 ;
  assign n20167 = n19479 & ~n20166 ;
  assign n20168 = n20167 ^ n19459 ;
  assign n20169 = n19369 & n20168 ;
  assign n20190 = n20189 ^ n20169 ;
  assign n20156 = n20153 ^ n19476 ;
  assign n20154 = n19536 ^ n19446 ;
  assign n20155 = n20154 ^ n20153 ;
  assign n20157 = n20156 ^ n20155 ;
  assign n20158 = n20156 ^ n19369 ;
  assign n20159 = n20158 ^ n20156 ;
  assign n20160 = n20157 & ~n20159 ;
  assign n20161 = n20160 ^ n20156 ;
  assign n20162 = ~n19371 & n20161 ;
  assign n20191 = n20190 ^ n20162 ;
  assign n20193 = n20192 ^ n20191 ;
  assign n20194 = ~n19486 & n20193 ;
  assign n20195 = ~n19543 & n20194 ;
  assign n20196 = n19534 ^ n19476 ;
  assign n20197 = n20196 ^ n19500 ;
  assign n20198 = ~n19370 & ~n20197 ;
  assign n20199 = n20198 ^ n19500 ;
  assign n20200 = n20199 ^ n19480 ;
  assign n20201 = n20200 ^ n20199 ;
  assign n20202 = n20199 ^ n19369 ;
  assign n20203 = n20202 ^ n20199 ;
  assign n20204 = ~n20201 & ~n20203 ;
  assign n20205 = n20204 ^ n20199 ;
  assign n20206 = n19371 & n20205 ;
  assign n20207 = n20206 ^ n20199 ;
  assign n20208 = n20195 & ~n20207 ;
  assign n20209 = n20208 ^ n17371 ;
  assign n20825 = n20209 ^ x98 ;
  assign n20826 = ~n20824 & n20825 ;
  assign n20827 = n20823 & n20826 ;
  assign n20828 = n20825 ^ n20824 ;
  assign n20844 = ~n20791 & n20800 ;
  assign n20845 = ~n20828 & n20844 ;
  assign n20838 = n20799 ^ n20797 ;
  assign n20841 = ~n20824 & n20838 ;
  assign n20842 = n20841 ^ n20797 ;
  assign n20843 = ~n20825 & n20842 ;
  assign n20846 = n20845 ^ n20843 ;
  assign n20864 = ~n20790 & n20800 ;
  assign n20855 = n20822 ^ n20801 ;
  assign n20856 = n20855 ^ n20803 ;
  assign n20848 = n20844 ^ n20802 ;
  assign n20849 = n20848 ^ n20812 ;
  assign n20850 = n20849 ^ n20806 ;
  assign n20853 = n20850 ^ n20822 ;
  assign n20854 = n20853 ^ n20801 ;
  assign n20857 = n20856 ^ n20854 ;
  assign n20852 = n20794 ^ n20756 ;
  assign n20858 = n20857 ^ n20852 ;
  assign n20859 = n20858 ^ n20806 ;
  assign n20872 = n20864 ^ n20859 ;
  assign n20866 = n20815 ^ n20803 ;
  assign n20869 = n20826 ^ n20824 ;
  assign n20870 = n20866 & ~n20869 ;
  assign n20871 = n20870 ^ n20797 ;
  assign n20873 = n20872 ^ n20871 ;
  assign n20876 = n20866 ^ n20858 ;
  assign n20877 = ~n20826 & ~n20876 ;
  assign n20878 = n20873 & n20877 ;
  assign n20865 = n20864 ^ n20792 ;
  assign n20867 = n20866 ^ n20865 ;
  assign n20868 = n20825 & n20867 ;
  assign n20874 = n20873 ^ n20868 ;
  assign n20879 = n20878 ^ n20874 ;
  assign n20880 = ~n20824 & n20879 ;
  assign n20881 = n20880 ^ n20868 ;
  assign n20847 = n20823 ^ n20816 ;
  assign n20851 = n20850 ^ n20847 ;
  assign n20860 = n20859 ^ n20851 ;
  assign n20861 = n20824 & n20860 ;
  assign n20862 = n20861 ^ n20850 ;
  assign n20863 = ~n20825 & n20862 ;
  assign n20882 = n20881 ^ n20863 ;
  assign n20883 = ~n20846 & ~n20882 ;
  assign n20829 = n20826 ^ n20825 ;
  assign n20830 = n20829 ^ n20828 ;
  assign n20831 = n20830 ^ n20828 ;
  assign n20832 = n20824 ^ n20802 ;
  assign n20833 = n20832 ^ n20828 ;
  assign n20834 = n20831 & ~n20833 ;
  assign n20835 = n20834 ^ n20828 ;
  assign n20836 = ~n20801 & ~n20835 ;
  assign n20837 = n20836 ^ n20828 ;
  assign n20884 = n20883 ^ n20837 ;
  assign n20885 = n20799 ^ n20792 ;
  assign n20886 = n20885 ^ n20794 ;
  assign n20887 = ~n20825 & n20886 ;
  assign n20888 = n20887 ^ n20809 ;
  assign n20889 = n20828 & ~n20888 ;
  assign n20890 = n20889 ^ n20808 ;
  assign n20891 = ~n20884 & n20890 ;
  assign n20892 = ~n20827 & n20891 ;
  assign n20893 = n20892 ^ n19124 ;
  assign n20894 = n20893 ^ x101 ;
  assign n18503 = n18477 ^ n18447 ;
  assign n18504 = n18447 ^ n18435 ;
  assign n18505 = n18504 ^ n18447 ;
  assign n18506 = ~n18503 & ~n18505 ;
  assign n18507 = n18506 ^ n18447 ;
  assign n18508 = ~n18407 & n18507 ;
  assign n20337 = ~n18467 & n18525 ;
  assign n20331 = n20007 ^ n18453 ;
  assign n18445 = n18444 ^ n18443 ;
  assign n20332 = n20331 ^ n18445 ;
  assign n20333 = n18407 & n20332 ;
  assign n20329 = n18455 ^ n18444 ;
  assign n20324 = n19778 ^ n18471 ;
  assign n19786 = n18453 ^ n18447 ;
  assign n19787 = n19786 ^ n18474 ;
  assign n20323 = n19787 ^ n18460 ;
  assign n20325 = n20324 ^ n20323 ;
  assign n20326 = ~n18407 & n20325 ;
  assign n20327 = n20326 ^ n20324 ;
  assign n20330 = n20329 ^ n20327 ;
  assign n20334 = n20333 ^ n20330 ;
  assign n20335 = n18435 & n20334 ;
  assign n20328 = n20327 ^ n19806 ;
  assign n20336 = n20335 ^ n20328 ;
  assign n20338 = n20337 ^ n20336 ;
  assign n20339 = ~n18488 & ~n20338 ;
  assign n20340 = ~n18508 & n20339 ;
  assign n20341 = n20340 ^ n17488 ;
  assign n20342 = n20341 ^ x107 ;
  assign n20359 = n20358 ^ x89 ;
  assign n20475 = n19534 ^ n19470 ;
  assign n20476 = n20475 ^ n19536 ;
  assign n20477 = ~n19369 & ~n20476 ;
  assign n20488 = n20477 ^ n20187 ;
  assign n20489 = n20488 ^ n20176 ;
  assign n19489 = n19369 & n19370 ;
  assign n19490 = n19489 ^ n19370 ;
  assign n19491 = n19488 & n19490 ;
  assign n19492 = n19491 ^ n19486 ;
  assign n20490 = n20489 ^ n19492 ;
  assign n20486 = n19473 & n19490 ;
  assign n19521 = n19369 & n19506 ;
  assign n19522 = n19521 ^ n19478 ;
  assign n19523 = n19522 ^ n19446 ;
  assign n19524 = n19523 ^ n19522 ;
  assign n19527 = ~n19369 & n19524 ;
  assign n19528 = n19527 ^ n19522 ;
  assign n19529 = n19371 & n19528 ;
  assign n19530 = n19529 ^ n19522 ;
  assign n20487 = n20486 ^ n19530 ;
  assign n20491 = n20490 ^ n20487 ;
  assign n20492 = n20491 ^ n18130 ;
  assign n20479 = n20154 ^ n19470 ;
  assign n20480 = n20479 ^ n19500 ;
  assign n20481 = n20480 ^ n20477 ;
  assign n20474 = n19487 ^ n19453 ;
  assign n20478 = n20477 ^ n20474 ;
  assign n20482 = n20481 ^ n20478 ;
  assign n20483 = ~n19369 & n20482 ;
  assign n20484 = n20483 ^ n20481 ;
  assign n20485 = ~n19370 & n20484 ;
  assign n20493 = n20492 ^ n20485 ;
  assign n20473 = n19472 & n19489 ;
  assign n20494 = n20493 ^ n20473 ;
  assign n20466 = n19476 ^ n19369 ;
  assign n20467 = n20466 ^ n19476 ;
  assign n20470 = n19474 & n20467 ;
  assign n20471 = n20470 ^ n19476 ;
  assign n20472 = ~n19370 & n20471 ;
  assign n20495 = n20494 ^ n20472 ;
  assign n20496 = n20495 ^ x66 ;
  assign n19549 = n18398 ^ x75 ;
  assign n19551 = n18603 ^ x125 ;
  assign n19566 = n17421 ^ n17395 ;
  assign n19565 = n17404 ^ n17383 ;
  assign n19567 = n19566 ^ n19565 ;
  assign n19568 = n19565 ^ n17372 ;
  assign n19569 = n19568 ^ n19565 ;
  assign n19570 = n19567 & ~n19569 ;
  assign n19571 = n19570 ^ n19565 ;
  assign n19572 = ~n17338 & n19571 ;
  assign n19573 = n19572 ^ n19104 ;
  assign n19563 = n17447 ^ n17283 ;
  assign n19564 = n17373 & ~n19563 ;
  assign n19574 = n19573 ^ n19564 ;
  assign n19562 = ~n17374 & n17433 ;
  assign n19575 = n19574 ^ n19562 ;
  assign n19555 = n17417 ^ n17398 ;
  assign n19552 = n18553 ^ n17233 ;
  assign n19553 = n19552 ^ n17276 ;
  assign n19554 = n19553 ^ n17290 ;
  assign n19556 = n19555 ^ n19554 ;
  assign n19557 = n19554 ^ n17372 ;
  assign n19558 = n19557 ^ n19554 ;
  assign n19559 = ~n19556 & ~n19558 ;
  assign n19560 = n19559 ^ n19554 ;
  assign n19561 = n17338 & ~n19560 ;
  assign n19576 = n19575 ^ n19561 ;
  assign n19577 = n19576 ^ n17381 ;
  assign n19578 = ~n18567 & ~n19577 ;
  assign n19579 = n19578 ^ n17375 ;
  assign n19580 = ~n17294 & n19579 ;
  assign n19581 = n19580 ^ n15248 ;
  assign n19582 = n19581 ^ x124 ;
  assign n19583 = n19551 & n19582 ;
  assign n19614 = n16703 & n16706 ;
  assign n19595 = n16718 ^ n16590 ;
  assign n19596 = n19595 ^ n16592 ;
  assign n19597 = n19596 ^ n16590 ;
  assign n19598 = n19597 ^ n16709 ;
  assign n19599 = ~n16638 & n19598 ;
  assign n19600 = n19599 ^ n19595 ;
  assign n19605 = n19600 ^ n19204 ;
  assign n19591 = n16693 ^ n16592 ;
  assign n19592 = n19591 ^ n18892 ;
  assign n19601 = n19592 ^ n19204 ;
  assign n19602 = n19601 ^ n19600 ;
  assign n19590 = n18884 ^ n16706 ;
  assign n19593 = n19592 ^ n19590 ;
  assign n19594 = ~n16678 & ~n19593 ;
  assign n19603 = n19602 ^ n19594 ;
  assign n19604 = ~n16679 & ~n19603 ;
  assign n19606 = n19605 ^ n19604 ;
  assign n19609 = n16716 ^ n16696 ;
  assign n19610 = n19609 ^ n16593 ;
  assign n19611 = ~n16719 & ~n19610 ;
  assign n19612 = ~n19606 & n19611 ;
  assign n19607 = n19606 ^ n19216 ;
  assign n19613 = n19612 ^ n19607 ;
  assign n19615 = n19614 ^ n19613 ;
  assign n19584 = n18884 ^ n16681 ;
  assign n19585 = n16681 ^ n16638 ;
  assign n19586 = n19585 ^ n16681 ;
  assign n19587 = n19584 & n19586 ;
  assign n19588 = n19587 ^ n16681 ;
  assign n19589 = n16678 & n19588 ;
  assign n19616 = n19615 ^ n19589 ;
  assign n19617 = ~n18866 & ~n19616 ;
  assign n19618 = n19617 ^ n15199 ;
  assign n19619 = n19618 ^ x110 ;
  assign n19620 = n18434 ^ x68 ;
  assign n19621 = n19619 & ~n19620 ;
  assign n19622 = n19621 ^ n19619 ;
  assign n19633 = n19622 ^ n19620 ;
  assign n19637 = n19583 & n19633 ;
  assign n19624 = n19583 ^ n19551 ;
  assign n19634 = n19624 & n19633 ;
  assign n19631 = n19551 & n19621 ;
  assign n19626 = n19583 & n19621 ;
  assign n19632 = n19631 ^ n19626 ;
  assign n19635 = n19634 ^ n19632 ;
  assign n19638 = n19637 ^ n19635 ;
  assign n19625 = n19622 & n19624 ;
  assign n19630 = n19625 ^ n19624 ;
  assign n19636 = n19635 ^ n19630 ;
  assign n19639 = n19638 ^ n19636 ;
  assign n19627 = n19626 ^ n19625 ;
  assign n19623 = n19583 & n19622 ;
  assign n19628 = n19627 ^ n19623 ;
  assign n19629 = n19628 ^ n19551 ;
  assign n19640 = n19639 ^ n19629 ;
  assign n20138 = n19640 ^ n19635 ;
  assign n19548 = n18685 ^ x93 ;
  assign n20139 = n19635 ^ n19548 ;
  assign n20140 = n20139 ^ n19635 ;
  assign n20141 = n20138 & n20140 ;
  assign n20142 = n20141 ^ n19635 ;
  assign n20143 = n19549 & n20142 ;
  assign n20132 = n19627 ^ n19548 ;
  assign n20133 = n20132 ^ n19627 ;
  assign n20134 = n19628 & n20133 ;
  assign n20135 = n20134 ^ n19627 ;
  assign n20136 = ~n19549 & n20135 ;
  assign n19644 = n19624 ^ n19582 ;
  assign n19700 = n19621 & ~n19644 ;
  assign n19687 = ~n19548 & ~n19549 ;
  assign n19688 = n19687 ^ n19549 ;
  assign n19689 = n19688 ^ n19548 ;
  assign n19701 = n19689 ^ n19549 ;
  assign n19702 = n19700 & ~n19701 ;
  assign n19647 = n19583 ^ n19582 ;
  assign n19664 = n19622 & n19647 ;
  assign n19648 = n19621 ^ n19620 ;
  assign n19649 = ~n19644 & ~n19648 ;
  assign n19650 = n19649 ^ n19647 ;
  assign n19645 = n19619 & ~n19644 ;
  assign n19646 = n19645 ^ n19551 ;
  assign n19651 = n19650 ^ n19646 ;
  assign n19652 = n19651 ^ n19637 ;
  assign n19643 = n19634 ^ n19633 ;
  assign n19653 = n19652 ^ n19643 ;
  assign n19662 = n19653 ^ n19649 ;
  assign n19657 = n19640 ^ n19636 ;
  assign n19656 = n19649 ^ n19648 ;
  assign n19658 = n19657 ^ n19656 ;
  assign n19663 = n19662 ^ n19658 ;
  assign n19665 = n19664 ^ n19663 ;
  assign n19666 = n19665 ^ n19650 ;
  assign n19694 = n19666 ^ n19651 ;
  assign n19695 = n19651 ^ n19549 ;
  assign n19696 = n19695 ^ n19651 ;
  assign n19697 = ~n19694 & ~n19696 ;
  assign n19698 = n19697 ^ n19651 ;
  assign n19699 = n19548 & ~n19698 ;
  assign n19703 = n19702 ^ n19699 ;
  assign n19691 = n19632 ^ n19623 ;
  assign n19692 = ~n19689 & n19691 ;
  assign n19690 = n19637 & ~n19689 ;
  assign n19693 = n19692 ^ n19690 ;
  assign n20379 = n19703 ^ n19693 ;
  assign n20362 = n19653 ^ n19645 ;
  assign n20363 = n20362 ^ n19665 ;
  assign n20364 = n19548 & ~n20363 ;
  assign n20365 = n20364 ^ n19665 ;
  assign n20380 = n20379 ^ n20365 ;
  assign n20375 = n19662 ^ n19627 ;
  assign n20376 = ~n19548 & ~n20375 ;
  assign n19705 = n19700 ^ n19644 ;
  assign n19706 = n19705 ^ n19651 ;
  assign n19707 = n19706 ^ n19658 ;
  assign n19708 = ~n19548 & ~n19707 ;
  assign n19709 = n19708 ^ n19706 ;
  assign n20374 = n20365 ^ n19709 ;
  assign n20377 = n20376 ^ n20374 ;
  assign n20378 = n19549 & n20377 ;
  assign n20381 = n20380 ^ n20378 ;
  assign n20371 = n19634 ^ n19626 ;
  assign n20372 = n20371 ^ n19636 ;
  assign n20373 = ~n19688 & n20372 ;
  assign n20382 = n20381 ^ n20373 ;
  assign n19550 = n19549 ^ n19548 ;
  assign n20360 = n19664 ^ n19548 ;
  assign n20361 = n20360 ^ n19664 ;
  assign n20367 = n19664 ^ n19635 ;
  assign n20368 = ~n20361 & n20367 ;
  assign n20369 = n20368 ^ n19664 ;
  assign n20370 = ~n19550 & n20369 ;
  assign n20383 = n20382 ^ n20370 ;
  assign n20384 = ~n20136 & ~n20383 ;
  assign n20385 = ~n20143 & n20384 ;
  assign n20386 = n20385 ^ n18074 ;
  assign n20387 = n20386 ^ x122 ;
  assign n20498 = n20496 ^ n20387 ;
  assign n20438 = n20437 ^ x96 ;
  assign n20525 = ~n20387 & n20438 ;
  assign n17964 = n17699 ^ x114 ;
  assign n17963 = n17962 ^ x104 ;
  assign n18266 = n17964 ^ n17963 ;
  assign n18046 = n16764 ^ x81 ;
  assign n17992 = n17991 ^ x90 ;
  assign n18038 = n16141 ^ n15097 ;
  assign n18039 = n14627 & ~n18038 ;
  assign n18036 = n18035 ^ n18033 ;
  assign n18003 = n16135 ^ n15099 ;
  assign n18006 = n18005 ^ n16128 ;
  assign n18007 = n18005 ^ n16135 ;
  assign n18008 = n18007 ^ n18005 ;
  assign n18009 = ~n18006 & n18008 ;
  assign n18010 = n18009 ^ n18005 ;
  assign n18011 = ~n18003 & ~n18010 ;
  assign n18037 = n18036 ^ n18011 ;
  assign n18040 = n18039 ^ n18037 ;
  assign n17998 = n17997 ^ n16114 ;
  assign n17995 = n16107 ^ n16102 ;
  assign n17999 = n17998 ^ n17995 ;
  assign n18000 = ~n14627 & n17999 ;
  assign n17996 = n17995 ^ n16141 ;
  assign n18001 = n18000 ^ n17996 ;
  assign n18002 = n15097 & ~n18001 ;
  assign n18041 = n18040 ^ n18002 ;
  assign n18042 = ~n17994 & n18041 ;
  assign n18043 = n18042 ^ n15741 ;
  assign n18044 = n18043 ^ x107 ;
  assign n18045 = n17992 & n18044 ;
  assign n18220 = n18045 ^ n18044 ;
  assign n18221 = ~n18046 & n18220 ;
  assign n18166 = n18165 ^ n18157 ;
  assign n18170 = n18166 ^ n18165 ;
  assign n18171 = ~n18155 & ~n18170 ;
  assign n18172 = n18171 ^ n18166 ;
  assign n18173 = n18167 & n18172 ;
  assign n18174 = n18173 ^ n18166 ;
  assign n18175 = n18047 & n18174 ;
  assign n18176 = n18175 ^ n18047 ;
  assign n18180 = ~n18047 & n18179 ;
  assign n18181 = n18180 ^ n18157 ;
  assign n18182 = n18181 ^ n18047 ;
  assign n18183 = n18182 ^ n18180 ;
  assign n18184 = n18180 ^ n18160 ;
  assign n18185 = n18184 ^ n18180 ;
  assign n18186 = ~n18183 & ~n18185 ;
  assign n18187 = n18186 ^ n18180 ;
  assign n18188 = n18167 & n18187 ;
  assign n18189 = n18188 ^ n18180 ;
  assign n18190 = ~n18176 & ~n18189 ;
  assign n18191 = n18190 ^ n15757 ;
  assign n18192 = n18191 ^ x72 ;
  assign n18193 = ~n18046 & n18192 ;
  assign n18194 = n18193 ^ n18046 ;
  assign n18197 = n18045 ^ n17992 ;
  assign n18198 = n18197 ^ n18044 ;
  assign n18200 = n18198 ^ n17992 ;
  assign n18201 = ~n18194 & n18200 ;
  assign n18222 = n18221 ^ n18201 ;
  assign n18204 = n18045 & n18193 ;
  assign n18195 = n18045 & ~n18194 ;
  assign n18218 = n18204 ^ n18195 ;
  assign n18209 = n18194 ^ n18192 ;
  assign n18210 = ~n18198 & n18209 ;
  assign n18211 = n18210 ^ n18198 ;
  assign n18206 = n18193 ^ n18192 ;
  assign n18207 = ~n18198 & n18206 ;
  assign n18199 = ~n18194 & ~n18198 ;
  assign n18208 = n18207 ^ n18199 ;
  assign n18212 = n18211 ^ n18208 ;
  assign n18219 = n18218 ^ n18212 ;
  assign n18223 = n18222 ^ n18219 ;
  assign n18245 = n18223 ^ n18200 ;
  assign n18243 = n18219 ^ n18201 ;
  assign n18214 = n18200 & n18206 ;
  assign n18244 = n18243 ^ n18214 ;
  assign n18246 = n18245 ^ n18244 ;
  assign n18242 = n18197 & n18209 ;
  assign n18247 = n18246 ^ n18242 ;
  assign n18241 = n18210 ^ n18209 ;
  assign n18248 = n18247 ^ n18241 ;
  assign n18286 = n18248 ^ n18214 ;
  assign n18287 = n18248 ^ n17964 ;
  assign n18288 = n18287 ^ n18248 ;
  assign n18289 = n18286 & ~n18288 ;
  assign n18290 = n18289 ^ n18248 ;
  assign n18291 = n18266 & n18290 ;
  assign n18249 = n18248 ^ n18045 ;
  assign n18250 = n18249 ^ n18218 ;
  assign n18202 = n18201 ^ n18199 ;
  assign n18196 = n18195 ^ n18194 ;
  assign n18203 = n18202 ^ n18196 ;
  assign n20446 = n18250 ^ n18203 ;
  assign n20454 = n20446 ^ n18223 ;
  assign n18261 = n18242 ^ n18207 ;
  assign n20442 = n18261 ^ n18212 ;
  assign n18217 = n18196 ^ n18046 ;
  assign n18224 = n18223 ^ n18217 ;
  assign n20441 = n18224 ^ n18208 ;
  assign n20443 = n20442 ^ n20441 ;
  assign n20444 = n17964 & n20443 ;
  assign n20445 = n20444 ^ n20442 ;
  assign n20453 = n20445 ^ n18210 ;
  assign n20455 = n20454 ^ n20453 ;
  assign n20450 = n18218 ^ n18210 ;
  assign n18251 = n18250 ^ n18208 ;
  assign n18205 = n18204 ^ n18203 ;
  assign n18213 = n18212 ^ n18205 ;
  assign n18270 = n18251 ^ n18213 ;
  assign n18271 = n18270 ^ n18244 ;
  assign n18269 = n18192 ^ n18046 ;
  assign n18272 = n18271 ^ n18269 ;
  assign n18273 = n18272 ^ n18246 ;
  assign n20076 = n18273 ^ n18207 ;
  assign n20077 = n20076 ^ n18210 ;
  assign n20078 = n20077 ^ n18223 ;
  assign n20451 = n20450 ^ n20078 ;
  assign n20452 = n17963 & ~n20451 ;
  assign n20456 = n20455 ^ n20452 ;
  assign n20457 = ~n18266 & ~n20456 ;
  assign n20447 = n20446 ^ n20445 ;
  assign n19840 = n18202 ^ n18201 ;
  assign n19841 = n18201 ^ n17964 ;
  assign n19842 = n19841 ^ n18201 ;
  assign n19843 = n19840 & n19842 ;
  assign n19844 = n19843 ^ n18201 ;
  assign n19845 = ~n18266 & n19844 ;
  assign n19846 = n19845 ^ n18201 ;
  assign n20448 = n20447 ^ n19846 ;
  assign n18292 = n18248 ^ n18222 ;
  assign n18293 = n18222 ^ n17964 ;
  assign n18294 = n18293 ^ n18222 ;
  assign n18295 = n18292 & ~n18294 ;
  assign n18296 = n18295 ^ n18222 ;
  assign n18297 = n17963 & n18296 ;
  assign n20449 = n20448 ^ n18297 ;
  assign n20458 = n20457 ^ n20449 ;
  assign n18265 = n17963 & ~n17964 ;
  assign n18267 = n18266 ^ n18265 ;
  assign n18268 = n18267 ^ n17963 ;
  assign n19853 = n18247 & ~n18268 ;
  assign n20459 = n20458 ^ n19853 ;
  assign n20440 = ~n17963 & n18272 ;
  assign n20460 = n20459 ^ n20440 ;
  assign n20461 = ~n18291 & ~n20460 ;
  assign n20462 = n20461 ^ n17612 ;
  assign n20463 = n20462 ^ x113 ;
  assign n20526 = n20525 ^ n20463 ;
  assign n20527 = ~n20498 & n20526 ;
  assign n20504 = n20496 ^ n20438 ;
  assign n20528 = n20527 ^ n20504 ;
  assign n20499 = n20438 & n20498 ;
  assign n20524 = n20499 ^ n20387 ;
  assign n20529 = n20528 ^ n20524 ;
  assign n20530 = n20529 ^ n20504 ;
  assign n20464 = n20463 ^ n20387 ;
  assign n20439 = n20438 ^ n20387 ;
  assign n20465 = n20464 ^ n20439 ;
  assign n20516 = ~n20463 & ~n20496 ;
  assign n20517 = n20516 ^ n20463 ;
  assign n20518 = n20498 & ~n20517 ;
  assign n20519 = n20518 ^ n20387 ;
  assign n20520 = n20465 & ~n20519 ;
  assign n20521 = n20520 ^ n20516 ;
  assign n20522 = n20521 ^ n20387 ;
  assign n20523 = n20522 ^ n20463 ;
  assign n20531 = n20530 ^ n20523 ;
  assign n20532 = n20531 ^ n20530 ;
  assign n20507 = n20463 ^ n20438 ;
  assign n20533 = n20525 ^ n20507 ;
  assign n20534 = ~n20496 & n20533 ;
  assign n20537 = ~n20532 & ~n20534 ;
  assign n20538 = n20537 ^ n20530 ;
  assign n20539 = n20359 & n20538 ;
  assign n20540 = n20539 ^ n20530 ;
  assign n20508 = n20496 & n20507 ;
  assign n20509 = n20508 ^ n20438 ;
  assign n20510 = n20387 & n20509 ;
  assign n20505 = n20504 ^ n20463 ;
  assign n20511 = n20510 ^ n20505 ;
  assign n20506 = n20505 ^ n20499 ;
  assign n20512 = n20511 ^ n20506 ;
  assign n20497 = n20496 ^ n20464 ;
  assign n20500 = n20499 ^ n20497 ;
  assign n20501 = n20500 ^ n20439 ;
  assign n20502 = ~n20465 & ~n20501 ;
  assign n20503 = n20502 ^ n20497 ;
  assign n20513 = n20512 ^ n20503 ;
  assign n20514 = ~n20359 & ~n20513 ;
  assign n20515 = n20514 ^ n20511 ;
  assign n20541 = n20540 ^ n20515 ;
  assign n20542 = n20342 & n20541 ;
  assign n20543 = n20542 ^ n20342 ;
  assign n20544 = n20543 ^ n20540 ;
  assign n20545 = n20544 ^ n18968 ;
  assign n20546 = n20545 ^ x116 ;
  assign n20144 = n20143 ^ n16637 ;
  assign n20119 = n19700 ^ n19653 ;
  assign n20120 = n20119 ^ n19623 ;
  assign n20121 = n19623 ^ n19549 ;
  assign n20122 = n20121 ^ n19623 ;
  assign n20123 = ~n20120 & ~n20122 ;
  assign n20124 = n20123 ^ n19623 ;
  assign n20125 = ~n19548 & n20124 ;
  assign n20126 = n20125 ^ n19699 ;
  assign n20106 = n19645 ^ n19628 ;
  assign n20104 = n19666 ^ n19636 ;
  assign n20096 = n19700 ^ n19657 ;
  assign n20097 = n20096 ^ n19652 ;
  assign n20098 = n20097 ^ n19657 ;
  assign n20099 = n19657 ^ n19548 ;
  assign n20100 = n20099 ^ n19657 ;
  assign n20101 = ~n20098 & n20100 ;
  assign n20102 = n20101 ^ n19657 ;
  assign n20103 = ~n19549 & n20102 ;
  assign n20105 = n20104 ^ n20103 ;
  assign n20107 = n20106 ^ n20105 ;
  assign n20108 = n20107 ^ n20103 ;
  assign n20109 = n19548 & n20108 ;
  assign n20110 = n20109 ^ n20105 ;
  assign n20127 = n20126 ^ n20110 ;
  assign n19711 = n19708 ^ n19658 ;
  assign n19712 = n19711 ^ n19664 ;
  assign n19713 = n19712 ^ n19711 ;
  assign n19716 = n19548 & n19713 ;
  assign n19717 = n19716 ^ n19711 ;
  assign n19718 = ~n19549 & ~n19717 ;
  assign n19719 = n19718 ^ n19711 ;
  assign n19704 = ~n19653 & ~n19701 ;
  assign n19720 = n19719 ^ n19704 ;
  assign n20128 = n20127 ^ n19720 ;
  assign n20111 = n20110 ^ n20103 ;
  assign n20114 = n20111 ^ n19706 ;
  assign n20115 = n20114 ^ n20111 ;
  assign n20116 = ~n19548 & n20115 ;
  assign n20117 = n20116 ^ n20111 ;
  assign n20118 = ~n19549 & n20117 ;
  assign n20129 = n20128 ^ n20118 ;
  assign n20137 = n20129 & ~n20136 ;
  assign n20145 = n20144 ^ n20137 ;
  assign n20547 = n20145 ^ x112 ;
  assign n18816 = n18765 ^ n18758 ;
  assign n18817 = n18605 & n18816 ;
  assign n18818 = n18817 ^ n16677 ;
  assign n18782 = n18781 ^ n18606 ;
  assign n18783 = n18605 ^ n18572 ;
  assign n18785 = n18784 ^ n18783 ;
  assign n18786 = n18784 ^ n18606 ;
  assign n18787 = n18786 ^ n18784 ;
  assign n18788 = ~n18785 & n18787 ;
  assign n18789 = n18788 ^ n18784 ;
  assign n18790 = ~n18782 & n18789 ;
  assign n18791 = n18790 ^ n18781 ;
  assign n18793 = n18755 ^ n18746 ;
  assign n18792 = n18751 ^ n18736 ;
  assign n18794 = n18793 ^ n18792 ;
  assign n18795 = ~n18572 & ~n18794 ;
  assign n18796 = n18795 ^ n18793 ;
  assign n18813 = n18812 ^ n18796 ;
  assign n18798 = n18771 ^ n18752 ;
  assign n18803 = n18802 ^ n18798 ;
  assign n18804 = n18803 ^ n18796 ;
  assign n18797 = n18796 ^ n18734 ;
  assign n18805 = n18804 ^ n18797 ;
  assign n18806 = n18804 ^ n18572 ;
  assign n18807 = n18806 ^ n18804 ;
  assign n18808 = ~n18805 & ~n18807 ;
  assign n18809 = n18808 ^ n18804 ;
  assign n18810 = n18604 & ~n18809 ;
  assign n18814 = n18813 ^ n18810 ;
  assign n18815 = ~n18791 & ~n18814 ;
  assign n18819 = n18818 ^ n18815 ;
  assign n20548 = n18819 ^ x105 ;
  assign n20549 = n20547 & n20548 ;
  assign n20550 = n20549 ^ n20548 ;
  assign n17751 = n16174 & n17748 ;
  assign n17743 = n17726 ^ n17702 ;
  assign n17744 = n16174 & n17743 ;
  assign n17745 = n17744 ^ n17726 ;
  assign n17752 = n17751 ^ n17745 ;
  assign n17753 = ~n16765 & n17752 ;
  assign n17754 = n17753 ^ n17745 ;
  assign n20569 = n20396 ^ n17705 ;
  assign n17779 = n17769 ^ n17764 ;
  assign n17781 = n17780 ^ n17779 ;
  assign n17760 = n17759 ^ n17716 ;
  assign n17782 = n17781 ^ n17760 ;
  assign n20570 = n20569 ^ n17782 ;
  assign n20571 = n16174 & ~n20570 ;
  assign n20572 = n20571 ^ n17759 ;
  assign n20573 = ~n16765 & n20572 ;
  assign n20567 = n16174 & n17779 ;
  assign n20554 = n17715 ^ n17703 ;
  assign n20555 = n20554 ^ n17780 ;
  assign n20556 = n17780 ^ n16765 ;
  assign n20557 = n17778 & n20556 ;
  assign n20558 = n20557 ^ n16765 ;
  assign n20559 = n20555 & n20558 ;
  assign n20560 = n20559 ^ n17780 ;
  assign n20561 = n20560 ^ n17725 ;
  assign n20562 = n20561 ^ n17709 ;
  assign n20565 = n20562 ^ n20432 ;
  assign n20551 = n17758 ^ n17731 ;
  assign n20552 = n20551 ^ n17755 ;
  assign n20553 = n16765 & n20552 ;
  assign n20563 = n20562 ^ n20553 ;
  assign n20564 = n17778 & n20563 ;
  assign n20566 = n20565 ^ n20564 ;
  assign n20568 = n20567 ^ n20566 ;
  assign n20574 = n20573 ^ n20568 ;
  assign n20575 = ~n17754 & ~n20574 ;
  assign n20576 = ~n20421 & n20575 ;
  assign n20577 = n20576 ^ n16543 ;
  assign n20578 = n20577 ^ x64 ;
  assign n19229 = n19228 ^ n19227 ;
  assign n19269 = n19268 ^ n19261 ;
  assign n19270 = ~n19227 & ~n19269 ;
  assign n19271 = n19270 ^ n19261 ;
  assign n19272 = n19271 ^ n19235 ;
  assign n19273 = n19272 ^ n19267 ;
  assign n19274 = n19273 ^ n19272 ;
  assign n19277 = n19227 & n19274 ;
  assign n19278 = n19277 ^ n19272 ;
  assign n19279 = n19229 & n19278 ;
  assign n19280 = n19279 ^ n19271 ;
  assign n19281 = ~n19188 & ~n19280 ;
  assign n19282 = n19281 ^ n16192 ;
  assign n20605 = n19282 ^ x81 ;
  assign n20650 = ~n20578 & ~n20605 ;
  assign n20583 = n19474 ^ n19446 ;
  assign n20584 = n20583 ^ n19488 ;
  assign n20581 = n19466 ^ n19462 ;
  assign n20582 = n19369 & n20581 ;
  assign n20585 = n20584 ^ n20582 ;
  assign n20597 = n20585 ^ n20487 ;
  assign n20598 = n20597 ^ n20169 ;
  assign n20579 = n19488 ^ n19478 ;
  assign n20580 = n20579 ^ n19535 ;
  assign n20586 = n20585 ^ n20580 ;
  assign n20587 = n20586 ^ n20585 ;
  assign n20588 = n20587 ^ n19477 ;
  assign n20589 = n20588 ^ n20587 ;
  assign n20590 = n20587 ^ n19537 ;
  assign n20591 = n20590 ^ n20587 ;
  assign n20592 = ~n20589 & ~n20591 ;
  assign n20593 = n20592 ^ n20587 ;
  assign n20594 = ~n19369 & n20593 ;
  assign n20595 = n20594 ^ n20586 ;
  assign n20596 = n19370 & ~n20595 ;
  assign n20599 = n20598 ^ n20596 ;
  assign n20600 = ~n20207 & ~n20599 ;
  assign n20601 = n20600 ^ n16582 ;
  assign n20602 = n20601 ^ x90 ;
  assign n20603 = ~n20578 & n20602 ;
  assign n20604 = n20603 ^ n20578 ;
  assign n19949 = n19030 ^ n18994 ;
  assign n19957 = n18988 ^ n18821 ;
  assign n19959 = n18988 ^ n18960 ;
  assign n19958 = n18988 ^ n18981 ;
  assign n19960 = n19959 ^ n19958 ;
  assign n19961 = n19959 ^ n18969 ;
  assign n19962 = n19961 ^ n19959 ;
  assign n19963 = n19960 & n19962 ;
  assign n19964 = n19963 ^ n19959 ;
  assign n19965 = n19957 & ~n19964 ;
  assign n19966 = n19965 ^ n18821 ;
  assign n19024 = n18992 ^ n18977 ;
  assign n19025 = n19024 ^ n18978 ;
  assign n19950 = n19025 ^ n18988 ;
  assign n19951 = n19950 ^ n18955 ;
  assign n19954 = ~n18969 & n19951 ;
  assign n19955 = n19954 ^ n18955 ;
  assign n19956 = ~n18821 & n19955 ;
  assign n19967 = n19966 ^ n19956 ;
  assign n19968 = n19967 ^ n19048 ;
  assign n19969 = n19008 ^ n18995 ;
  assign n19970 = n19969 ^ n18995 ;
  assign n19972 = n18821 & n18998 ;
  assign n19973 = n19972 ^ n18995 ;
  assign n19974 = ~n19970 & n19973 ;
  assign n19975 = n19974 ^ n18995 ;
  assign n19976 = ~n19968 & n19975 ;
  assign n19977 = n19976 ^ n19968 ;
  assign n19978 = n18969 & ~n19977 ;
  assign n19979 = n18977 ^ n18821 ;
  assign n19980 = n19979 ^ n18977 ;
  assign n19983 = ~n19000 & ~n19980 ;
  assign n19984 = n19983 ^ n18977 ;
  assign n19985 = n19978 & n19984 ;
  assign n19986 = n19985 ^ n19977 ;
  assign n19987 = n18975 & ~n19986 ;
  assign n19988 = ~n19949 & n19987 ;
  assign n19989 = n19988 ^ n19986 ;
  assign n19001 = n19000 ^ n18978 ;
  assign n18989 = n18988 ^ n18983 ;
  assign n19990 = n18989 ^ n18977 ;
  assign n19991 = n19990 ^ n18994 ;
  assign n19993 = n19991 ^ n19005 ;
  assign n19994 = n19001 & ~n19993 ;
  assign n19995 = n19994 ^ n19005 ;
  assign n19992 = n19991 ^ n19001 ;
  assign n19996 = n19995 ^ n19992 ;
  assign n19997 = ~n19989 & ~n19996 ;
  assign n19998 = n19997 ^ n16384 ;
  assign n20606 = n19998 ^ x115 ;
  assign n20607 = ~n20605 & n20606 ;
  assign n20608 = n20607 ^ n20605 ;
  assign n20634 = ~n20604 & ~n20608 ;
  assign n20622 = n20603 & n20607 ;
  assign n20635 = n20634 ^ n20622 ;
  assign n20651 = n20650 ^ n20635 ;
  assign n20618 = n20578 & ~n20606 ;
  assign n20619 = n20602 ^ n20578 ;
  assign n20620 = n20618 & ~n20619 ;
  assign n20631 = n20620 ^ n20619 ;
  assign n20632 = ~n20605 & ~n20631 ;
  assign n20633 = n20632 ^ n20607 ;
  assign n20636 = n20635 ^ n20633 ;
  assign n20609 = n20608 ^ n20606 ;
  assign n20611 = n20604 ^ n20602 ;
  assign n20628 = n20609 & n20611 ;
  assign n20612 = n20609 ^ n20605 ;
  assign n20626 = ~n20604 & n20612 ;
  assign n20629 = n20628 ^ n20626 ;
  assign n20613 = n20611 & n20612 ;
  assign n20630 = n20629 ^ n20613 ;
  assign n20637 = n20636 ^ n20630 ;
  assign n20627 = n20626 ^ n20611 ;
  assign n20638 = n20637 ^ n20627 ;
  assign n20641 = n20638 ^ n20622 ;
  assign n20642 = n20641 ^ n20634 ;
  assign n20616 = n20603 ^ n20602 ;
  assign n20617 = n20609 & n20616 ;
  assign n20621 = n20620 ^ n20617 ;
  assign n20623 = n20622 ^ n20621 ;
  assign n20640 = n20623 ^ n20608 ;
  assign n20643 = n20642 ^ n20640 ;
  assign n20652 = n20651 ^ n20643 ;
  assign n20653 = n20652 ^ n20641 ;
  assign n20639 = n20638 ^ n20636 ;
  assign n20649 = n20639 ^ n20607 ;
  assign n20654 = n20653 ^ n20649 ;
  assign n20655 = n20654 ^ n20643 ;
  assign n20615 = n20603 & n20609 ;
  assign n20656 = n20655 ^ n20615 ;
  assign n20647 = n20602 & n20606 ;
  assign n20648 = n20647 ^ n20603 ;
  assign n20657 = n20656 ^ n20648 ;
  assign n20719 = n20657 ^ n20638 ;
  assign n20720 = n20550 & n20719 ;
  assign n20721 = n20720 ^ n19226 ;
  assign n20713 = n20654 ^ n20617 ;
  assign n20714 = n20617 ^ n20548 ;
  assign n20715 = n20714 ^ n20617 ;
  assign n20716 = ~n20713 & n20715 ;
  assign n20717 = n20716 ^ n20617 ;
  assign n20718 = ~n20547 & n20717 ;
  assign n20722 = n20721 ^ n20718 ;
  assign n20686 = n20549 ^ n20547 ;
  assign n20687 = n20621 & n20686 ;
  assign n20658 = n20657 ^ n20629 ;
  assign n20659 = n20658 ^ n20617 ;
  assign n20644 = n20643 ^ n20639 ;
  assign n20645 = n20644 ^ n20632 ;
  assign n20624 = n20623 ^ n20615 ;
  assign n20610 = ~n20604 & n20609 ;
  assign n20614 = n20613 ^ n20610 ;
  assign n20625 = n20624 ^ n20614 ;
  assign n20646 = n20645 ^ n20625 ;
  assign n20660 = n20659 ^ n20646 ;
  assign n20672 = n20660 ^ n20628 ;
  assign n20671 = n20657 ^ n20655 ;
  assign n20673 = n20672 ^ n20671 ;
  assign n20674 = n20547 & n20673 ;
  assign n20675 = n20674 ^ n20656 ;
  assign n20663 = n20652 ^ n20617 ;
  assign n20684 = n20675 ^ n20663 ;
  assign n20676 = n20675 ^ n20614 ;
  assign n20677 = n20676 ^ n20657 ;
  assign n20678 = n20677 ^ n20675 ;
  assign n20681 = n20547 & n20678 ;
  assign n20682 = n20681 ^ n20675 ;
  assign n20683 = n20548 & n20682 ;
  assign n20685 = n20684 ^ n20683 ;
  assign n20688 = n20687 ^ n20685 ;
  assign n20664 = n20663 ^ n20637 ;
  assign n20665 = n20664 ^ n20663 ;
  assign n20666 = n20663 ^ n20547 ;
  assign n20667 = n20666 ^ n20663 ;
  assign n20668 = n20665 & ~n20667 ;
  assign n20669 = n20668 ^ n20663 ;
  assign n20670 = ~n20548 & ~n20669 ;
  assign n20689 = n20688 ^ n20670 ;
  assign n20690 = n20548 ^ n20547 ;
  assign n20691 = n20636 ^ n20634 ;
  assign n20692 = n20636 ^ n20548 ;
  assign n20693 = n20692 ^ n20636 ;
  assign n20694 = n20691 & n20693 ;
  assign n20695 = n20694 ^ n20636 ;
  assign n20696 = n20690 & n20695 ;
  assign n20697 = n20689 & ~n20696 ;
  assign n20661 = n20660 ^ n20610 ;
  assign n20662 = n20550 & n20661 ;
  assign n20698 = n20697 ^ n20662 ;
  assign n20701 = n20639 & ~n20693 ;
  assign n20702 = n20701 ^ n20636 ;
  assign n20703 = n20547 & n20702 ;
  assign n20704 = n20698 & ~n20703 ;
  assign n20705 = n20641 ^ n20548 ;
  assign n20706 = n20705 ^ n20641 ;
  assign n20709 = ~n20653 & ~n20706 ;
  assign n20710 = n20709 ^ n20641 ;
  assign n20711 = n20547 & n20710 ;
  assign n20712 = n20704 & ~n20711 ;
  assign n20723 = n20722 ^ n20712 ;
  assign n20724 = n20723 ^ x76 ;
  assign n20725 = ~n20546 & ~n20724 ;
  assign n20726 = n20725 ^ n20546 ;
  assign n19340 = n19230 ^ n19158 ;
  assign n19341 = n19340 ^ n19260 ;
  assign n19348 = n19341 ^ n19265 ;
  assign n19344 = n19254 ^ n19182 ;
  assign n19345 = n19344 ^ n19160 ;
  assign n19346 = n19345 ^ n19125 ;
  assign n19347 = n19346 ^ n19184 ;
  assign n19349 = n19348 ^ n19347 ;
  assign n19350 = ~n19228 & n19349 ;
  assign n19351 = n19350 ^ n19347 ;
  assign n19352 = n19351 ^ n19259 ;
  assign n19353 = n19352 ^ n19351 ;
  assign n19337 = n19182 ^ n19159 ;
  assign n19338 = ~n19160 & n19337 ;
  assign n19339 = n19338 ^ n19236 ;
  assign n19354 = n19353 ^ n19339 ;
  assign n19355 = n19228 & ~n19354 ;
  assign n19356 = n19355 ^ n19352 ;
  assign n19360 = n19359 ^ n19356 ;
  assign n19361 = n19229 & ~n19360 ;
  assign n19362 = n19361 ^ n19339 ;
  assign n19342 = n19341 ^ n19339 ;
  assign n19343 = ~n19228 & n19342 ;
  assign n19363 = n19362 ^ n19343 ;
  assign n19365 = ~n19227 & n19359 ;
  assign n19366 = ~n19363 & n19365 ;
  assign n19364 = n19363 ^ n14626 ;
  assign n19367 = n19366 ^ n19364 ;
  assign n19368 = n19367 ^ x75 ;
  assign n19510 = n19470 ^ n19452 ;
  assign n19511 = n19510 ^ n19474 ;
  assign n19512 = n19511 ^ n19506 ;
  assign n19513 = ~n19369 & n19512 ;
  assign n19503 = n19454 ^ n19444 ;
  assign n19504 = ~n19369 & ~n19503 ;
  assign n19508 = n19507 ^ n19504 ;
  assign n19509 = n19508 ^ n19475 ;
  assign n19514 = n19513 ^ n19509 ;
  assign n19515 = n19370 & n19514 ;
  assign n19516 = n19515 ^ n19508 ;
  assign n19501 = n19489 ^ n19369 ;
  assign n19502 = n19500 & n19501 ;
  assign n19517 = n19516 ^ n19502 ;
  assign n19518 = n19517 ^ n19449 ;
  assign n19495 = n19449 ^ n19369 ;
  assign n19496 = n19495 ^ n19449 ;
  assign n19497 = n19487 & n19496 ;
  assign n19498 = n19497 ^ n19449 ;
  assign n19499 = n19370 & n19498 ;
  assign n19519 = n19518 ^ n19499 ;
  assign n19520 = ~n19492 & ~n19519 ;
  assign n19531 = n19520 & ~n19530 ;
  assign n19544 = n19531 & ~n19543 ;
  assign n19545 = n19544 ^ n15096 ;
  assign n19546 = n19545 ^ x124 ;
  assign n19909 = n19368 & n19546 ;
  assign n19911 = n19909 ^ n19368 ;
  assign n19910 = n19909 ^ n19546 ;
  assign n19912 = n19911 ^ n19910 ;
  assign n19721 = n19720 ^ n19703 ;
  assign n19661 = n19634 ^ n19625 ;
  assign n19667 = n19666 ^ n19661 ;
  assign n19642 = n19620 ^ n19619 ;
  assign n19654 = n19653 ^ n19642 ;
  assign n19641 = n19640 ^ n19632 ;
  assign n19655 = n19654 ^ n19641 ;
  assign n19659 = n19658 ^ n19655 ;
  assign n19660 = ~n19548 & n19659 ;
  assign n19668 = n19667 ^ n19660 ;
  assign n19722 = n19721 ^ n19668 ;
  assign n19723 = n19722 ^ n19693 ;
  assign n19676 = n19664 ^ n19625 ;
  assign n19677 = ~n19549 & n19676 ;
  assign n19678 = n19677 ^ n19625 ;
  assign n19681 = n19678 ^ n19662 ;
  assign n19682 = n19681 ^ n19678 ;
  assign n19683 = ~n19549 & ~n19682 ;
  assign n19684 = n19683 ^ n19678 ;
  assign n19685 = n19548 & n19684 ;
  assign n19686 = n19685 ^ n19678 ;
  assign n19724 = n19723 ^ n19686 ;
  assign n19725 = n19724 ^ n15418 ;
  assign n19669 = n19668 ^ n19639 ;
  assign n19670 = n19669 ^ n19657 ;
  assign n19671 = n19670 ^ n19664 ;
  assign n19672 = n19671 ^ n19668 ;
  assign n19673 = ~n19548 & n19672 ;
  assign n19674 = n19673 ^ n19669 ;
  assign n19675 = n19550 & n19674 ;
  assign n19726 = n19725 ^ n19675 ;
  assign n19727 = n19726 ^ x125 ;
  assign n18262 = n17964 & n18261 ;
  assign n19847 = n18262 ^ n18203 ;
  assign n19848 = ~n18266 & ~n19847 ;
  assign n19849 = n19848 ^ n18203 ;
  assign n19830 = ~n17964 & ~n18271 ;
  assign n19817 = n18248 & n18265 ;
  assign n19818 = n19817 ^ n18214 ;
  assign n19819 = n19818 ^ n18272 ;
  assign n19820 = n19819 ^ n18210 ;
  assign n19821 = n19820 ^ n18267 ;
  assign n19822 = n18265 ^ n18218 ;
  assign n19825 = ~n19820 & ~n19822 ;
  assign n19826 = n19825 ^ n18265 ;
  assign n19827 = n19821 & n19826 ;
  assign n19828 = n19827 ^ n18267 ;
  assign n19829 = n19828 ^ n18244 ;
  assign n19831 = n19830 ^ n19829 ;
  assign n19850 = n19849 ^ n19831 ;
  assign n19851 = n19850 ^ n19846 ;
  assign n19832 = n19831 ^ n19828 ;
  assign n19833 = n19832 ^ n17963 ;
  assign n19834 = n19833 ^ n19832 ;
  assign n18225 = n18224 ^ n18222 ;
  assign n19835 = n19832 ^ n18225 ;
  assign n19836 = n19835 ^ n19832 ;
  assign n19837 = n19834 & ~n19836 ;
  assign n19838 = n19837 ^ n19832 ;
  assign n19839 = n18266 & ~n19838 ;
  assign n19852 = n19851 ^ n19839 ;
  assign n19854 = n19853 ^ n19852 ;
  assign n19855 = ~n18291 & ~n19854 ;
  assign n19856 = n19855 ^ n15855 ;
  assign n19857 = n19856 ^ x118 ;
  assign n19858 = ~n19727 & n19857 ;
  assign n19728 = ~n18604 & n18780 ;
  assign n19729 = n19728 ^ n18746 ;
  assign n19730 = n19729 ^ n18757 ;
  assign n19731 = n19730 ^ n18758 ;
  assign n19732 = n19731 ^ n19729 ;
  assign n19735 = n18604 & n19732 ;
  assign n19736 = n19735 ^ n19729 ;
  assign n19737 = ~n18572 & n19736 ;
  assign n19738 = n19737 ^ n19729 ;
  assign n19747 = n18772 ^ n18748 ;
  assign n19753 = n19747 ^ n18765 ;
  assign n19750 = n18761 ^ n18757 ;
  assign n19751 = n19750 ^ n19747 ;
  assign n19752 = n18572 & n19751 ;
  assign n19754 = n19753 ^ n19752 ;
  assign n19755 = ~n18767 & ~n19754 ;
  assign n19756 = ~n18604 & ~n19755 ;
  assign n19748 = n19747 ^ n18777 ;
  assign n19749 = n19746 & n19748 ;
  assign n19757 = n19756 ^ n19749 ;
  assign n19741 = n18771 ^ n18604 ;
  assign n19742 = n19741 ^ n18771 ;
  assign n19743 = ~n18775 & n19742 ;
  assign n19744 = n19743 ^ n18771 ;
  assign n19745 = n18572 & n19744 ;
  assign n19758 = n19757 ^ n19745 ;
  assign n19759 = n18760 ^ n18750 ;
  assign n19760 = n18760 ^ n18572 ;
  assign n19761 = n19760 ^ n18760 ;
  assign n19762 = n19759 & ~n19761 ;
  assign n19763 = n19762 ^ n18760 ;
  assign n19764 = n18604 & n19763 ;
  assign n19765 = ~n19758 & ~n19764 ;
  assign n19766 = ~n19738 & n19765 ;
  assign n19767 = ~n18791 & n19766 ;
  assign n19768 = n19767 ^ n15646 ;
  assign n19769 = n19768 ^ x100 ;
  assign n19777 = n18465 ^ n18463 ;
  assign n19779 = n19778 ^ n19777 ;
  assign n19780 = n19779 ^ n18463 ;
  assign n19781 = n18463 ^ n18407 ;
  assign n19782 = n19781 ^ n18463 ;
  assign n19783 = ~n19780 & ~n19782 ;
  assign n19784 = n19783 ^ n18463 ;
  assign n19785 = ~n18456 & ~n19784 ;
  assign n19788 = n19787 ^ n19785 ;
  assign n19789 = n19788 ^ n18477 ;
  assign n19790 = n19789 ^ n19785 ;
  assign n19791 = n19785 ^ n18407 ;
  assign n19792 = n19791 ^ n19785 ;
  assign n19793 = ~n19790 & n19792 ;
  assign n19794 = n19793 ^ n19785 ;
  assign n19795 = n18435 & ~n19794 ;
  assign n19796 = n19795 ^ n19785 ;
  assign n19772 = n18467 ^ n18454 ;
  assign n19770 = n18451 ^ n18406 ;
  assign n18470 = n18469 ^ n18454 ;
  assign n18472 = n18471 ^ n18470 ;
  assign n19771 = n19770 ^ n18472 ;
  assign n19773 = n19772 ^ n19771 ;
  assign n19774 = n18435 & n19773 ;
  assign n19775 = n19774 ^ n19772 ;
  assign n19776 = ~n18407 & ~n19775 ;
  assign n19797 = n19796 ^ n19776 ;
  assign n19803 = n19797 & ~n19802 ;
  assign n19809 = n19808 ^ n19803 ;
  assign n19810 = ~n18508 & n19809 ;
  assign n19811 = n19810 ^ n16091 ;
  assign n19812 = n19811 ^ x85 ;
  assign n19813 = n19769 & ~n19812 ;
  assign n19866 = n19813 ^ n19812 ;
  assign n19920 = n19858 & ~n19866 ;
  assign n19814 = n19813 ^ n19769 ;
  assign n19815 = n19814 ^ n19812 ;
  assign n19859 = n19858 ^ n19727 ;
  assign n19896 = n19815 & ~n19859 ;
  assign n19921 = n19920 ^ n19896 ;
  assign n19913 = n19814 & n19858 ;
  assign n19940 = n19921 ^ n19913 ;
  assign n19938 = n19812 ^ n19727 ;
  assign n19889 = n19857 ^ n19727 ;
  assign n19890 = n19857 ^ n19769 ;
  assign n19891 = n19857 ^ n19812 ;
  assign n19892 = n19891 ^ n19857 ;
  assign n19893 = ~n19890 & n19892 ;
  assign n19894 = n19893 ^ n19857 ;
  assign n19895 = ~n19889 & ~n19894 ;
  assign n19939 = n19938 ^ n19895 ;
  assign n19941 = n19940 ^ n19939 ;
  assign n19924 = n19814 & ~n19859 ;
  assign n19874 = n19813 & ~n19859 ;
  assign n19925 = n19924 ^ n19874 ;
  assign n19897 = n19896 ^ n19859 ;
  assign n19926 = n19925 ^ n19897 ;
  assign n19942 = n19941 ^ n19926 ;
  assign n19860 = n19859 ^ n19857 ;
  assign n19869 = n19813 & n19860 ;
  assign n19943 = n19942 ^ n19869 ;
  assign n19944 = ~n19546 & n19943 ;
  assign n19945 = n19944 ^ n19939 ;
  assign n19946 = ~n19912 & ~n19945 ;
  assign n19861 = n19860 ^ n19727 ;
  assign n19872 = n19813 & n19861 ;
  assign n19876 = n19872 ^ n19869 ;
  assign n19875 = n19874 ^ n19813 ;
  assign n19877 = n19876 ^ n19875 ;
  assign n19922 = n19921 ^ n19877 ;
  assign n19914 = n19913 ^ n19896 ;
  assign n19919 = n19914 ^ n19858 ;
  assign n19923 = n19922 ^ n19919 ;
  assign n19927 = n19926 ^ n19923 ;
  assign n19898 = n19897 ^ n19895 ;
  assign n19864 = n19815 & n19860 ;
  assign n19899 = n19898 ^ n19864 ;
  assign n19900 = n19899 ^ n19872 ;
  assign n19816 = n19727 & n19815 ;
  assign n19862 = n19861 ^ n19816 ;
  assign n19901 = n19900 ^ n19862 ;
  assign n19902 = n19901 ^ n19869 ;
  assign n19928 = n19927 ^ n19902 ;
  assign n19929 = ~n19546 & n19928 ;
  assign n19915 = n19912 & n19914 ;
  assign n19867 = n19860 & ~n19866 ;
  assign n19903 = n19902 ^ n19867 ;
  assign n19904 = n19867 ^ n19368 ;
  assign n19905 = n19904 ^ n19867 ;
  assign n19906 = ~n19903 & ~n19905 ;
  assign n19907 = n19906 ^ n19867 ;
  assign n19908 = n19546 & n19907 ;
  assign n19916 = n19915 ^ n19908 ;
  assign n19917 = n19916 ^ n19442 ;
  assign n19547 = n19546 ^ n19368 ;
  assign n19865 = n19864 ^ n19816 ;
  assign n19868 = n19867 ^ n19865 ;
  assign n19870 = n19869 ^ n19868 ;
  assign n19863 = n19862 ^ n19727 ;
  assign n19871 = n19870 ^ n19863 ;
  assign n19873 = n19872 ^ n19871 ;
  assign n19878 = n19877 ^ n19873 ;
  assign n19879 = ~n19546 & n19878 ;
  assign n19880 = n19879 ^ n19877 ;
  assign n19881 = n19880 ^ n19874 ;
  assign n19882 = n19881 ^ n19880 ;
  assign n19883 = n19880 ^ n19368 ;
  assign n19884 = n19883 ^ n19880 ;
  assign n19885 = n19882 & n19884 ;
  assign n19886 = n19885 ^ n19880 ;
  assign n19887 = ~n19547 & n19886 ;
  assign n19888 = n19887 ^ n19880 ;
  assign n19918 = n19917 ^ n19888 ;
  assign n19930 = n19929 ^ n19918 ;
  assign n19933 = n19930 ^ n19442 ;
  assign n19934 = n19933 ^ n19888 ;
  assign n19931 = n19898 ^ n19868 ;
  assign n19932 = n19931 ^ n19916 ;
  assign n19935 = n19934 ^ n19932 ;
  assign n19936 = ~n19368 & ~n19935 ;
  assign n19937 = n19936 ^ n19930 ;
  assign n19947 = n19946 ^ n19937 ;
  assign n19948 = n19947 ^ x70 ;
  assign n20057 = n18817 ^ n17858 ;
  assign n20039 = n18771 ^ n18765 ;
  assign n20040 = n20039 ^ n18767 ;
  assign n20041 = n18604 & n20040 ;
  assign n20042 = n20041 ^ n18800 ;
  assign n20043 = ~n18572 & ~n20042 ;
  assign n20044 = n20043 ^ n18756 ;
  assign n20034 = n18756 ^ n18604 ;
  assign n20035 = n20034 ^ n18756 ;
  assign n20036 = n18763 & ~n20035 ;
  assign n20037 = n20036 ^ n18756 ;
  assign n20038 = n20022 & n20037 ;
  assign n20045 = n20044 ^ n20038 ;
  assign n20046 = n18746 ^ n18604 ;
  assign n20047 = n20046 ^ n18746 ;
  assign n20048 = n18572 & n18777 ;
  assign n20049 = n20048 ^ n18746 ;
  assign n20050 = n20047 & n20049 ;
  assign n20051 = n20050 ^ n18746 ;
  assign n20052 = ~n20045 & n20051 ;
  assign n20053 = n20052 ^ n20045 ;
  assign n20054 = ~n19764 & ~n20053 ;
  assign n20055 = ~n20032 & n20054 ;
  assign n20056 = ~n19738 & n20055 ;
  assign n20058 = n20057 ^ n20056 ;
  assign n20059 = n20058 ^ x104 ;
  assign n20091 = n19853 ^ n17828 ;
  assign n20063 = n17963 & n19818 ;
  assign n20061 = n18266 & n18273 ;
  assign n20060 = n18250 ^ n18214 ;
  assign n20062 = n20061 ^ n20060 ;
  assign n20064 = n20063 ^ n20062 ;
  assign n20065 = n20064 ^ n17963 ;
  assign n20068 = n18199 ^ n18195 ;
  assign n20069 = n20068 ^ n17964 ;
  assign n20070 = ~n20064 & n20069 ;
  assign n20071 = n20070 ^ n17964 ;
  assign n20072 = ~n20065 & ~n20071 ;
  assign n20073 = n20072 ^ n17963 ;
  assign n20080 = n18192 ^ n18044 ;
  assign n18239 = n18212 ^ n18195 ;
  assign n20079 = n18239 ^ n18222 ;
  assign n20081 = n20080 ^ n20079 ;
  assign n20082 = n20081 ^ n20078 ;
  assign n20083 = n17964 & n20082 ;
  assign n20084 = n20083 ^ n20079 ;
  assign n20085 = n20084 ^ n18212 ;
  assign n20074 = n18204 ^ n18193 ;
  assign n20075 = ~n17964 & n20074 ;
  assign n20086 = n20085 ^ n20075 ;
  assign n20087 = ~n17963 & n20086 ;
  assign n20088 = n20087 ^ n20084 ;
  assign n20089 = n20073 & n20088 ;
  assign n20090 = n19849 & n20089 ;
  assign n20092 = n20091 ^ n20090 ;
  assign n20093 = n20092 ^ x97 ;
  assign n20146 = n20145 ^ x123 ;
  assign n20210 = n20209 ^ x114 ;
  assign n20211 = ~n20146 & ~n20210 ;
  assign n20222 = n20093 & n20211 ;
  assign n20232 = n20059 & n20222 ;
  assign n20094 = n20059 & ~n20093 ;
  assign n20228 = n20094 ^ n20059 ;
  assign n20233 = n20232 ^ n20228 ;
  assign n20212 = n20211 ^ n20210 ;
  assign n20230 = ~n20212 & n20228 ;
  assign n20213 = n20212 ^ n20146 ;
  assign n20229 = ~n20213 & n20228 ;
  assign n20231 = n20230 ^ n20229 ;
  assign n20234 = n20233 ^ n20231 ;
  assign n20095 = n20094 ^ n20093 ;
  assign n20217 = n20211 ^ n20146 ;
  assign n20226 = ~n20095 & ~n20217 ;
  assign n20248 = n20234 ^ n20226 ;
  assign n20214 = ~n20095 & ~n20213 ;
  assign n20249 = n20248 ^ n20214 ;
  assign n20220 = ~n20095 & n20211 ;
  assign n20235 = n20234 ^ n20220 ;
  assign n20247 = n20235 ^ n20095 ;
  assign n20250 = n20249 ^ n20247 ;
  assign n20218 = n20095 ^ n20059 ;
  assign n20241 = n20210 & n20218 ;
  assign n20219 = ~n20217 & n20218 ;
  assign n20242 = n20241 ^ n20219 ;
  assign n20251 = n20250 ^ n20242 ;
  assign n20245 = n20241 ^ n20218 ;
  assign n20238 = n20232 ^ n20222 ;
  assign n20246 = n20245 ^ n20238 ;
  assign n20252 = n20251 ^ n20246 ;
  assign n19999 = n19998 ^ x99 ;
  assign n20021 = n20020 ^ x72 ;
  assign n20284 = n19999 & ~n20021 ;
  assign n20285 = n20284 ^ n20021 ;
  assign n20286 = n20285 ^ n19999 ;
  assign n20300 = n20286 ^ n20021 ;
  assign n20312 = ~n20252 & n20300 ;
  assign n20221 = n20220 ^ n20211 ;
  assign n20223 = n20222 ^ n20221 ;
  assign n20301 = n20223 & n20300 ;
  assign n20227 = n20226 ^ n20222 ;
  assign n20236 = n20235 ^ n20227 ;
  assign n20224 = n20223 ^ n20219 ;
  assign n20225 = n20224 ^ n20146 ;
  assign n20237 = n20236 ^ n20225 ;
  assign n20297 = n20237 ^ n20232 ;
  assign n20298 = n20297 ^ n20226 ;
  assign n20295 = n20230 & ~n20285 ;
  assign n20270 = n20021 ^ n19999 ;
  assign n20289 = n20238 ^ n20224 ;
  assign n20290 = n20238 ^ n19999 ;
  assign n20291 = n20290 ^ n20238 ;
  assign n20292 = n20289 & ~n20291 ;
  assign n20293 = n20292 ^ n20238 ;
  assign n20294 = n20270 & n20293 ;
  assign n20296 = n20295 ^ n20294 ;
  assign n20299 = n20298 ^ n20296 ;
  assign n20302 = n20301 ^ n20299 ;
  assign n20243 = n20242 ^ n20230 ;
  assign n20244 = n20243 ^ n20212 ;
  assign n20253 = n20252 ^ n20244 ;
  assign n20309 = n20302 ^ n20253 ;
  assign n20304 = n20253 ^ n20242 ;
  assign n20305 = n20304 ^ n20229 ;
  assign n20306 = ~n20021 & n20305 ;
  assign n20303 = n20302 ^ n20296 ;
  assign n20307 = n20306 ^ n20303 ;
  assign n20308 = ~n19999 & ~n20307 ;
  assign n20310 = n20309 ^ n20308 ;
  assign n20287 = n20238 ^ n20234 ;
  assign n20288 = n20286 & n20287 ;
  assign n20311 = n20310 ^ n20288 ;
  assign n20313 = n20312 ^ n20311 ;
  assign n20239 = n20238 ^ n20220 ;
  assign n20240 = n20239 ^ n20237 ;
  assign n20254 = n20253 ^ n20240 ;
  assign n20278 = n20254 ^ n20253 ;
  assign n20279 = n20253 ^ n20021 ;
  assign n20280 = n20279 ^ n20253 ;
  assign n20281 = ~n20278 & ~n20280 ;
  assign n20282 = n20281 ^ n20253 ;
  assign n20283 = ~n20270 & n20282 ;
  assign n20314 = n20313 ^ n20283 ;
  assign n20315 = n20314 ^ n20214 ;
  assign n20271 = n20230 ^ n19999 ;
  assign n20272 = n20271 ^ n20230 ;
  assign n20275 = n20231 & ~n20272 ;
  assign n20276 = n20275 ^ n20230 ;
  assign n20277 = n20270 & n20276 ;
  assign n20316 = n20315 ^ n20277 ;
  assign n20264 = n20229 ^ n20226 ;
  assign n20265 = n20229 ^ n19999 ;
  assign n20266 = n20265 ^ n20229 ;
  assign n20267 = n20264 & ~n20266 ;
  assign n20268 = n20267 ^ n20229 ;
  assign n20269 = ~n20021 & n20268 ;
  assign n20317 = n20316 ^ n20269 ;
  assign n20318 = n20317 ^ n19411 ;
  assign n20215 = n20214 ^ n20021 ;
  assign n20216 = n20215 ^ n20214 ;
  assign n20255 = n20239 ^ n20223 ;
  assign n20256 = n20255 ^ n20094 ;
  assign n20257 = n20256 ^ n20254 ;
  assign n20258 = n20257 ^ n20246 ;
  assign n20261 = n20216 & ~n20258 ;
  assign n20262 = n20261 ^ n20214 ;
  assign n20263 = ~n19999 & n20262 ;
  assign n20319 = n20318 ^ n20263 ;
  assign n20320 = n20319 ^ x118 ;
  assign n20321 = n19948 & ~n20320 ;
  assign n20322 = n20321 ^ n19948 ;
  assign n20731 = n20322 ^ n20320 ;
  assign n20907 = ~n20726 & n20731 ;
  assign n20727 = n20726 ^ n20724 ;
  assign n20900 = ~n20727 & n20731 ;
  assign n20908 = n20907 ^ n20900 ;
  assign n20905 = n20321 & ~n20727 ;
  assign n20732 = n20731 ^ n19948 ;
  assign n20904 = ~n20726 & ~n20732 ;
  assign n20906 = n20905 ^ n20904 ;
  assign n20909 = n20908 ^ n20906 ;
  assign n20902 = n20546 ^ n19948 ;
  assign n20903 = n20724 & n20902 ;
  assign n20910 = n20909 ^ n20903 ;
  assign n20901 = n20900 ^ n20724 ;
  assign n20911 = n20910 ^ n20901 ;
  assign n20728 = n20727 ^ n20546 ;
  assign n20729 = n20322 & ~n20728 ;
  assign n20915 = n20911 ^ n20729 ;
  assign n20913 = n20322 & n20725 ;
  assign n20914 = n20913 ^ n20322 ;
  assign n20916 = n20915 ^ n20914 ;
  assign n20923 = n20916 ^ n20900 ;
  assign n20922 = n20906 ^ n20724 ;
  assign n20924 = n20923 ^ n20922 ;
  assign n20920 = n20320 ^ n19948 ;
  assign n20921 = n20920 ^ n20546 ;
  assign n20925 = n20924 ^ n20921 ;
  assign n20733 = ~n20728 & ~n20732 ;
  assign n20730 = n20321 & n20725 ;
  assign n20734 = n20733 ^ n20730 ;
  assign n20735 = n20734 ^ n20729 ;
  assign n20926 = n20925 ^ n20735 ;
  assign n20927 = n20926 ^ n20731 ;
  assign n20928 = n20927 ^ n20908 ;
  assign n20964 = n20928 ^ n20730 ;
  assign n20944 = n20905 ^ n20726 ;
  assign n20945 = n20944 ^ n20910 ;
  assign n20965 = n20964 ^ n20945 ;
  assign n20931 = n20926 ^ n20733 ;
  assign n20932 = n20931 ^ n20913 ;
  assign n20966 = n20965 ^ n20932 ;
  assign n17790 = n17763 ^ n17711 ;
  assign n17791 = n17790 ^ n16765 ;
  assign n17792 = n17791 ^ n17790 ;
  assign n17793 = n17790 ^ n17709 ;
  assign n17794 = n17793 ^ n17790 ;
  assign n17795 = n17792 & n17794 ;
  assign n17796 = n17795 ^ n17790 ;
  assign n17797 = n16174 & n17796 ;
  assign n17784 = n17760 ^ n16765 ;
  assign n17785 = n17784 ^ n17760 ;
  assign n17786 = n17781 & n17785 ;
  assign n17787 = n17786 ^ n17760 ;
  assign n17788 = n17778 & n17787 ;
  assign n17770 = n17769 ^ n17703 ;
  assign n17771 = n17770 ^ n17723 ;
  assign n17772 = n17723 ^ n16174 ;
  assign n17773 = n17772 ^ n17723 ;
  assign n17774 = n17771 & ~n17773 ;
  assign n17775 = n17774 ^ n17723 ;
  assign n17776 = ~n16765 & n17775 ;
  assign n17767 = n17766 ^ n17760 ;
  assign n17768 = n17767 ^ n17754 ;
  assign n17777 = n17776 ^ n17768 ;
  assign n17789 = n17788 ^ n17777 ;
  assign n17798 = n17797 ^ n17789 ;
  assign n17799 = ~n17742 & ~n17798 ;
  assign n17800 = ~n17730 & n17799 ;
  assign n17801 = n17800 ^ n16808 ;
  assign n17802 = n17801 ^ x77 ;
  assign n18298 = n18297 ^ n18291 ;
  assign n18274 = n18273 ^ n18203 ;
  assign n18275 = ~n18268 & ~n18274 ;
  assign n18263 = n18262 ^ n18250 ;
  assign n18226 = n18225 ^ n18201 ;
  assign n18236 = n18226 ^ n18212 ;
  assign n18215 = n18214 ^ n18213 ;
  assign n18216 = n18215 ^ n18212 ;
  assign n18227 = n18226 ^ n18216 ;
  assign n18230 = ~n18215 & n18227 ;
  assign n18237 = n18236 ^ n18230 ;
  assign n18228 = n18227 ^ n18226 ;
  assign n18232 = n18230 ^ n18228 ;
  assign n18233 = n17964 & ~n18232 ;
  assign n18234 = n18233 ^ n18226 ;
  assign n18235 = ~n17963 & ~n18234 ;
  assign n18238 = n18237 ^ n18235 ;
  assign n18252 = n18251 ^ n18199 ;
  assign n18253 = n18252 ^ n18247 ;
  assign n18240 = n18239 ^ n18225 ;
  assign n18254 = n18253 ^ n18240 ;
  assign n18255 = n18253 ^ n17964 ;
  assign n18256 = n18255 ^ n18253 ;
  assign n18257 = n18254 & ~n18256 ;
  assign n18258 = n18257 ^ n18253 ;
  assign n18259 = n17963 & n18258 ;
  assign n18260 = ~n18238 & ~n18259 ;
  assign n18264 = n18263 ^ n18260 ;
  assign n18276 = n18275 ^ n18264 ;
  assign n18299 = n18298 ^ n18276 ;
  assign n18300 = n18299 ^ n16861 ;
  assign n18277 = n18276 ^ n18263 ;
  assign n18279 = n18242 ^ n18199 ;
  assign n18278 = n18239 ^ n18224 ;
  assign n18280 = n18279 ^ n18278 ;
  assign n18281 = ~n17964 & n18280 ;
  assign n18282 = n18281 ^ n18278 ;
  assign n18283 = n18277 & n18282 ;
  assign n18284 = n18283 ^ n18263 ;
  assign n18285 = n17963 & n18284 ;
  assign n18301 = n18300 ^ n18285 ;
  assign n18302 = n18301 ^ x108 ;
  assign n18491 = n18461 ^ n18450 ;
  assign n18473 = n18468 ^ n18443 ;
  assign n18492 = n18491 ^ n18473 ;
  assign n18493 = n18435 & ~n18492 ;
  assign n18490 = n18489 ^ n18473 ;
  assign n18494 = n18493 ^ n18490 ;
  assign n18509 = n18508 ^ n18494 ;
  assign n18495 = n18494 ^ n18489 ;
  assign n18496 = n18495 ^ n18472 ;
  assign n18497 = n18496 ^ n18495 ;
  assign n18500 = ~n18435 & ~n18497 ;
  assign n18501 = n18500 ^ n18495 ;
  assign n18502 = ~n18407 & ~n18501 ;
  assign n18510 = n18509 ^ n18502 ;
  assign n18446 = n18436 & n18445 ;
  assign n18511 = n18510 ^ n18446 ;
  assign n18438 = n18406 & ~n18437 ;
  assign n18512 = n18511 ^ n18438 ;
  assign n18516 = n18458 ^ n18450 ;
  assign n18517 = n18516 ^ n18465 ;
  assign n18514 = n18472 ^ n18465 ;
  assign n18515 = n18435 & n18514 ;
  assign n18518 = n18517 ^ n18515 ;
  assign n18521 = n18407 & ~n18518 ;
  assign n18513 = n18472 ^ n18451 ;
  assign n18519 = n18518 ^ n18513 ;
  assign n18520 = n18435 & n18519 ;
  assign n18522 = n18521 ^ n18520 ;
  assign n18523 = n18522 ^ n18451 ;
  assign n18524 = n18512 & ~n18523 ;
  assign n18532 = n18524 & ~n18531 ;
  assign n18533 = n18532 ^ n16894 ;
  assign n18534 = n18533 ^ x94 ;
  assign n18535 = n18302 & ~n18534 ;
  assign n18536 = n18535 ^ n18534 ;
  assign n18820 = n18819 ^ x83 ;
  assign n19049 = n19048 ^ n16932 ;
  assign n19026 = n19025 ^ n18993 ;
  assign n19027 = ~n19023 & n19026 ;
  assign n19010 = n19009 ^ n18943 ;
  assign n19011 = n19010 ^ n18944 ;
  assign n19012 = ~n18969 & ~n19011 ;
  assign n19015 = n18943 ^ n18907 ;
  assign n19016 = n19015 ^ n18943 ;
  assign n19017 = n18944 & n19016 ;
  assign n19018 = n19017 ^ n18943 ;
  assign n19019 = n19012 & ~n19018 ;
  assign n19002 = n19001 ^ n18996 ;
  assign n19003 = ~n18990 & ~n19002 ;
  assign n19004 = n19003 ^ n18989 ;
  assign n19020 = n19019 ^ n19004 ;
  assign n19021 = ~n19008 & ~n19020 ;
  assign n19007 = n19006 ^ n19004 ;
  assign n19022 = n19021 ^ n19007 ;
  assign n19028 = n19027 ^ n19022 ;
  assign n18986 = n18985 ^ n18977 ;
  assign n18987 = n18975 & n18986 ;
  assign n19029 = n19028 ^ n18987 ;
  assign n19031 = n19030 ^ n18948 ;
  assign n19032 = n19031 ^ n18950 ;
  assign n19033 = n19032 ^ n18948 ;
  assign n19034 = n18948 ^ n18821 ;
  assign n19035 = n19034 ^ n18948 ;
  assign n19036 = ~n19033 & ~n19035 ;
  assign n19037 = n19036 ^ n18948 ;
  assign n19038 = n19008 & n19037 ;
  assign n19039 = n19029 & ~n19038 ;
  assign n18962 = n18961 ^ n18950 ;
  assign n18970 = n18969 ^ n18953 ;
  assign n18971 = n18970 ^ n18953 ;
  assign n18972 = n18962 & ~n18971 ;
  assign n18973 = n18972 ^ n18953 ;
  assign n18974 = n18821 & n18973 ;
  assign n19040 = n19039 ^ n18974 ;
  assign n19041 = n19001 ^ n18946 ;
  assign n19042 = n18946 ^ n18821 ;
  assign n19043 = n19042 ^ n18946 ;
  assign n19044 = ~n19041 & ~n19043 ;
  assign n19045 = n19044 ^ n18946 ;
  assign n19046 = ~n19008 & n19045 ;
  assign n19047 = n19040 & ~n19046 ;
  assign n19050 = n19049 ^ n19047 ;
  assign n19051 = n19050 ^ x109 ;
  assign n19052 = ~n18820 & n19051 ;
  assign n19070 = ~n18536 & n19052 ;
  assign n19053 = n19052 ^ n19051 ;
  assign n19055 = n18535 ^ n18302 ;
  assign n19057 = n19055 ^ n18534 ;
  assign n19058 = n19053 & n19057 ;
  assign n19056 = n19052 & n19055 ;
  assign n19059 = n19058 ^ n19056 ;
  assign n19054 = ~n18536 & n19053 ;
  assign n19060 = n19059 ^ n19054 ;
  assign n19085 = n19070 ^ n19060 ;
  assign n19066 = n19053 ^ n18820 ;
  assign n19082 = ~n18536 & n19066 ;
  assign n19083 = n19082 ^ n19059 ;
  assign n19084 = n19083 ^ n18536 ;
  assign n19086 = n19085 ^ n19084 ;
  assign n19067 = n18535 & n19066 ;
  assign n19087 = n19086 ^ n19067 ;
  assign n19064 = n19052 ^ n18820 ;
  assign n19081 = n19055 & ~n19064 ;
  assign n19088 = n19087 ^ n19081 ;
  assign n19065 = n18535 & ~n19064 ;
  assign n19068 = n19067 ^ n19065 ;
  assign n19080 = n19068 ^ n19064 ;
  assign n19089 = n19088 ^ n19080 ;
  assign n19079 = n19056 ^ n19054 ;
  assign n19090 = n19089 ^ n19079 ;
  assign n19283 = n19282 ^ x126 ;
  assign n19284 = n19090 & n19283 ;
  assign n19285 = n19284 ^ n19089 ;
  assign n19091 = n19090 ^ n19057 ;
  assign n19062 = n18535 & n19052 ;
  assign n19063 = n19062 ^ n18535 ;
  assign n19069 = n19068 ^ n19063 ;
  assign n19073 = n19069 ^ n19060 ;
  assign n19072 = n19056 ^ n19053 ;
  assign n19074 = n19073 ^ n19072 ;
  assign n19075 = n19074 ^ n19062 ;
  assign n19071 = n19070 ^ n19069 ;
  assign n19076 = n19075 ^ n19071 ;
  assign n19061 = n19060 ^ n19051 ;
  assign n19077 = n19076 ^ n19061 ;
  assign n19078 = n19077 ^ n19060 ;
  assign n19092 = n19091 ^ n19078 ;
  assign n19093 = n19092 ^ n19087 ;
  assign n19286 = n19285 ^ n19093 ;
  assign n19287 = n19286 ^ n19062 ;
  assign n19288 = n19287 ^ n19087 ;
  assign n19289 = n19288 ^ n19286 ;
  assign n19290 = n19286 ^ n19283 ;
  assign n19291 = n19290 ^ n19286 ;
  assign n19292 = ~n19289 & n19291 ;
  assign n19293 = n19292 ^ n19286 ;
  assign n19294 = ~n17802 & ~n19293 ;
  assign n19295 = n19294 ^ n19285 ;
  assign n19309 = n19283 ^ n17802 ;
  assign n19324 = n19082 ^ n19065 ;
  assign n19325 = n19309 & n19324 ;
  assign n19319 = ~n17802 & ~n19283 ;
  assign n19320 = n19319 ^ n19309 ;
  assign n19321 = n19089 ^ n19069 ;
  assign n19322 = ~n19320 & n19321 ;
  assign n19296 = n19088 ^ n19076 ;
  assign n19297 = ~n17802 & ~n19296 ;
  assign n19298 = n19297 ^ n19088 ;
  assign n19311 = n19298 ^ n19056 ;
  assign n19310 = n19298 ^ n19085 ;
  assign n19312 = n19311 ^ n19310 ;
  assign n19313 = n19311 ^ n17802 ;
  assign n19314 = n19313 ^ n19311 ;
  assign n19315 = n19312 & n19314 ;
  assign n19316 = n19315 ^ n19311 ;
  assign n19317 = n19309 & ~n19316 ;
  assign n19299 = n19055 & n19066 ;
  assign n19300 = n19299 ^ n17802 ;
  assign n19301 = n19300 ^ n19299 ;
  assign n19302 = n19077 ^ n19074 ;
  assign n19303 = n19302 ^ n19070 ;
  assign n19304 = n19303 ^ n19299 ;
  assign n19305 = ~n19301 & n19304 ;
  assign n19306 = n19305 ^ n19299 ;
  assign n19307 = n19283 & n19306 ;
  assign n19308 = n19307 ^ n19298 ;
  assign n19318 = n19317 ^ n19308 ;
  assign n19323 = n19322 ^ n19318 ;
  assign n19326 = n19325 ^ n19323 ;
  assign n19327 = ~n19295 & n19326 ;
  assign n19328 = n19299 ^ n19089 ;
  assign n19329 = n19089 ^ n17802 ;
  assign n19330 = n19329 ^ n19089 ;
  assign n19331 = n19328 & n19330 ;
  assign n19332 = n19331 ^ n19089 ;
  assign n19333 = ~n19283 & n19332 ;
  assign n19334 = n19327 & ~n19333 ;
  assign n19335 = n19334 ^ n18942 ;
  assign n19336 = n19335 ^ x83 ;
  assign n20967 = n20932 ^ n19336 ;
  assign n20968 = n20967 ^ n20932 ;
  assign n20969 = ~n20966 & n20968 ;
  assign n20970 = n20969 ^ n20932 ;
  assign n20971 = ~n20894 & n20970 ;
  assign n20933 = n20932 ^ n20725 ;
  assign n20934 = n20933 ^ n20734 ;
  assign n20935 = n20934 ^ n20928 ;
  assign n20958 = ~n19336 & n20894 ;
  assign n20962 = n20935 & n20958 ;
  assign n20959 = n20958 ^ n20894 ;
  assign n20960 = n20923 & n20959 ;
  assign n20942 = n20911 ^ n20906 ;
  assign n20947 = n20942 ^ n20726 ;
  assign n20917 = n20916 ^ n20905 ;
  assign n20912 = n20911 ^ n20907 ;
  assign n20918 = n20917 ^ n20912 ;
  assign n20948 = n20947 ^ n20918 ;
  assign n20949 = n20948 ^ n20900 ;
  assign n20946 = n20945 ^ n20905 ;
  assign n20950 = n20949 ^ n20946 ;
  assign n20936 = n20935 ^ n20926 ;
  assign n20929 = n20928 ^ n20729 ;
  assign n20919 = n20733 ^ n20728 ;
  assign n20930 = n20929 ^ n20919 ;
  assign n20937 = n20936 ^ n20930 ;
  assign n20938 = n20937 ^ n20918 ;
  assign n20939 = ~n20894 & ~n20938 ;
  assign n20940 = n20939 ^ n20937 ;
  assign n20951 = n20950 ^ n20940 ;
  assign n20943 = n20942 ^ n20913 ;
  assign n20952 = n20951 ^ n20943 ;
  assign n20953 = n20952 ^ n20940 ;
  assign n20954 = n20894 & n20953 ;
  assign n20955 = n20954 ^ n20951 ;
  assign n20956 = ~n19336 & ~n20955 ;
  assign n20736 = n20735 ^ n20734 ;
  assign n20737 = n20736 ^ n20734 ;
  assign n20897 = n20737 & ~n20894 ;
  assign n20898 = n20897 ^ n20734 ;
  assign n20899 = ~n19336 & n20898 ;
  assign n20941 = n20940 ^ n20899 ;
  assign n20957 = n20956 ^ n20941 ;
  assign n20961 = n20960 ^ n20957 ;
  assign n20963 = n20962 ^ n20961 ;
  assign n20972 = n20971 ^ n20963 ;
  assign n20978 = n20904 & n20959 ;
  assign n20975 = n20894 & n20915 ;
  assign n20976 = n20975 ^ n20729 ;
  assign n20977 = n19336 & n20976 ;
  assign n20979 = n20978 ^ n20977 ;
  assign n20980 = n20972 & ~n20979 ;
  assign n20981 = n20980 ^ n20209 ;
  assign n20982 = n19726 ^ x68 ;
  assign n20983 = n20462 ^ x117 ;
  assign n20984 = ~n20982 & ~n20983 ;
  assign n20985 = n20984 ^ n20982 ;
  assign n21049 = n17769 ^ n17702 ;
  assign n21048 = n20390 ^ n17790 ;
  assign n21050 = n21049 ^ n21048 ;
  assign n21051 = n21050 ^ n20390 ;
  assign n21052 = n16765 & n21051 ;
  assign n21053 = n21052 ^ n21048 ;
  assign n21054 = ~n17778 & n21053 ;
  assign n21045 = n17705 & n17761 ;
  assign n21039 = n17736 ^ n17717 ;
  assign n21040 = n21039 ^ n17755 ;
  assign n21041 = n16765 & ~n21040 ;
  assign n21037 = n17729 ^ n17717 ;
  assign n21025 = n17732 ^ n17722 ;
  assign n21026 = n21025 ^ n16765 ;
  assign n21027 = n17778 ^ n16765 ;
  assign n21028 = n21026 & ~n21027 ;
  assign n21029 = n21028 ^ n16765 ;
  assign n21030 = n17780 ^ n17748 ;
  assign n21031 = n21030 ^ n17780 ;
  assign n21032 = n21031 ^ n21025 ;
  assign n21033 = ~n21029 & n21032 ;
  assign n21034 = n21033 ^ n21030 ;
  assign n21038 = n21037 ^ n21034 ;
  assign n21042 = n21041 ^ n21038 ;
  assign n21043 = ~n16174 & n21042 ;
  assign n21035 = n20390 ^ n17756 ;
  assign n21036 = n21035 ^ n21034 ;
  assign n21044 = n21043 ^ n21036 ;
  assign n21046 = n21045 ^ n21044 ;
  assign n21020 = n17756 ^ n16765 ;
  assign n21021 = n21020 ^ n17756 ;
  assign n21022 = n20393 & n21021 ;
  assign n21023 = n21022 ^ n17756 ;
  assign n21024 = n17778 & n21023 ;
  assign n21047 = n21046 ^ n21024 ;
  assign n21055 = n21054 ^ n21047 ;
  assign n21056 = ~n20421 & ~n21055 ;
  assign n21057 = ~n17742 & n21056 ;
  assign n21058 = n21057 ^ n17512 ;
  assign n21059 = n21058 ^ x67 ;
  assign n21060 = n20341 ^ x92 ;
  assign n21061 = n21059 & n21060 ;
  assign n21079 = n21061 ^ n21060 ;
  assign n20986 = n19367 ^ x69 ;
  assign n21006 = n19006 ^ n18969 ;
  assign n20998 = n18997 ^ n18959 ;
  assign n20999 = n20998 ^ n20780 ;
  assign n20997 = n18984 ^ n18962 ;
  assign n21000 = n20999 ^ n20997 ;
  assign n21001 = n20999 ^ n18969 ;
  assign n21002 = n21001 ^ n20999 ;
  assign n21003 = n21000 & ~n21002 ;
  assign n21004 = n21003 ^ n20999 ;
  assign n21005 = ~n18821 & ~n21004 ;
  assign n21007 = n21006 ^ n21005 ;
  assign n20995 = n19023 ^ n19001 ;
  assign n20996 = ~n19995 & n20995 ;
  assign n21008 = n21007 ^ n20996 ;
  assign n20994 = ~n18969 & n18992 ;
  assign n21009 = n21008 ^ n20994 ;
  assign n20993 = n18962 & n19008 ;
  assign n21010 = n21009 ^ n20993 ;
  assign n20987 = n18996 ^ n18981 ;
  assign n20988 = n18981 ^ n18821 ;
  assign n20989 = n20988 ^ n18981 ;
  assign n20990 = n20987 & ~n20989 ;
  assign n20991 = n20990 ^ n18981 ;
  assign n20992 = ~n18969 & n20991 ;
  assign n21011 = n21010 ^ n20992 ;
  assign n21012 = ~n19046 & ~n21011 ;
  assign n21013 = n21012 ^ n17551 ;
  assign n21014 = n21013 ^ x86 ;
  assign n21015 = n20986 & ~n21014 ;
  assign n21086 = n21015 ^ n20986 ;
  assign n21089 = n21079 & n21086 ;
  assign n21083 = n21015 & n21079 ;
  assign n21090 = n21089 ^ n21083 ;
  assign n21016 = n21015 ^ n21014 ;
  assign n21080 = ~n21016 & n21079 ;
  assign n21088 = n21080 ^ n21079 ;
  assign n21091 = n21090 ^ n21088 ;
  assign n21092 = n21091 ^ n21089 ;
  assign n21087 = n21061 & n21086 ;
  assign n21093 = n21092 ^ n21087 ;
  assign n21017 = n21016 ^ n20986 ;
  assign n21082 = n21017 & n21061 ;
  assign n21084 = n21083 ^ n21082 ;
  assign n21078 = n21015 & n21061 ;
  assign n21081 = n21080 ^ n21078 ;
  assign n21085 = n21084 ^ n21081 ;
  assign n21094 = n21093 ^ n21085 ;
  assign n21095 = n21094 ^ n21060 ;
  assign n21099 = n21095 ^ n21078 ;
  assign n21062 = n21061 ^ n21059 ;
  assign n21072 = n21015 & n21062 ;
  assign n21098 = n21089 ^ n21072 ;
  assign n21100 = n21099 ^ n21098 ;
  assign n21096 = n21095 ^ n21090 ;
  assign n21097 = n21096 ^ n21015 ;
  assign n21101 = n21100 ^ n21097 ;
  assign n21070 = n21017 & n21062 ;
  assign n21102 = n21101 ^ n21070 ;
  assign n21068 = ~n21016 & n21062 ;
  assign n21103 = n21102 ^ n21068 ;
  assign n21104 = n21103 ^ n21060 ;
  assign n21065 = ~n21016 & ~n21060 ;
  assign n21069 = n21068 ^ n21065 ;
  assign n21071 = n21070 ^ n21069 ;
  assign n21073 = n21072 ^ n21071 ;
  assign n21063 = n21062 ^ n21060 ;
  assign n21066 = n21065 ^ n21063 ;
  assign n21067 = n21066 ^ n21060 ;
  assign n21074 = n21073 ^ n21067 ;
  assign n21064 = n21017 & ~n21063 ;
  assign n21075 = n21074 ^ n21064 ;
  assign n21076 = n21075 ^ n21069 ;
  assign n21077 = n21076 ^ n21072 ;
  assign n21105 = n21104 ^ n21077 ;
  assign n21106 = ~n20985 & ~n21105 ;
  assign n21149 = ~n20985 & n21091 ;
  assign n21114 = n20985 ^ n20983 ;
  assign n21146 = ~n21066 & ~n21114 ;
  assign n21136 = n20983 ^ n20982 ;
  assign n21141 = n21099 ^ n21084 ;
  assign n21137 = n21098 ^ n20983 ;
  assign n21138 = ~n21136 & n21137 ;
  assign n21139 = n21138 ^ n20983 ;
  assign n21140 = n21100 & ~n21139 ;
  assign n21142 = n21141 ^ n21140 ;
  assign n21131 = n21079 ^ n21015 ;
  assign n21132 = n21131 ^ n21070 ;
  assign n21133 = ~n20983 & n21132 ;
  assign n21143 = n21142 ^ n21133 ;
  assign n21144 = n21136 & n21143 ;
  assign n21124 = n21080 ^ n21068 ;
  assign n21125 = n21080 ^ n20982 ;
  assign n21126 = n21125 ^ n21080 ;
  assign n21127 = n21124 & ~n21126 ;
  assign n21128 = n21127 ^ n21080 ;
  assign n21129 = n20983 & n21128 ;
  assign n21130 = n21129 ^ n21074 ;
  assign n21134 = n21133 ^ n21130 ;
  assign n21117 = n21095 ^ n21087 ;
  assign n21118 = n21117 ^ n21105 ;
  assign n21119 = n21105 ^ n20983 ;
  assign n21120 = n21119 ^ n21105 ;
  assign n21121 = ~n21118 & n21120 ;
  assign n21122 = n21121 ^ n21105 ;
  assign n21123 = n20982 & ~n21122 ;
  assign n21135 = n21134 ^ n21123 ;
  assign n21145 = n21144 ^ n21135 ;
  assign n21147 = n21146 ^ n21145 ;
  assign n21115 = n21114 ^ n20982 ;
  assign n21116 = n21076 & ~n21115 ;
  assign n21148 = n21147 ^ n21116 ;
  assign n21150 = n21149 ^ n21148 ;
  assign n21107 = n21074 ^ n20983 ;
  assign n21108 = n21107 ^ n21074 ;
  assign n21111 = n21083 & n21108 ;
  assign n21112 = n21111 ^ n21074 ;
  assign n21113 = n20982 & n21112 ;
  assign n21151 = n21150 ^ n21113 ;
  assign n21152 = ~n21106 & ~n21151 ;
  assign n21153 = n21152 ^ n17699 ;
  assign n21154 = n21153 ^ x82 ;
  assign n21182 = n20230 ^ n20214 ;
  assign n21183 = n20286 & n21182 ;
  assign n21168 = ~n20285 & ~n20287 ;
  assign n21178 = n20094 & n20217 ;
  assign n21179 = n21168 & n21178 ;
  assign n21174 = ~n20257 & n20284 ;
  assign n21175 = n21174 ^ n20277 ;
  assign n21170 = n20297 ^ n20220 ;
  assign n21171 = n21170 ^ n20304 ;
  assign n21172 = n20300 & ~n21171 ;
  assign n21165 = n20250 ^ n20229 ;
  assign n21166 = n20300 & ~n21165 ;
  assign n21167 = n21166 ^ n20285 ;
  assign n21169 = n21168 ^ n21167 ;
  assign n21173 = n21172 ^ n21169 ;
  assign n21176 = n21175 ^ n21173 ;
  assign n21177 = n21176 ^ n20294 ;
  assign n21180 = n21179 ^ n21177 ;
  assign n21155 = n20232 ^ n20226 ;
  assign n21156 = n21155 ^ n20246 ;
  assign n21157 = n21156 ^ n20232 ;
  assign n21158 = n21157 ^ n20224 ;
  assign n21159 = n21158 ^ n21156 ;
  assign n21160 = n21156 ^ n20021 ;
  assign n21161 = n21160 ^ n21156 ;
  assign n21162 = n21159 & ~n21161 ;
  assign n21163 = n21162 ^ n21156 ;
  assign n21164 = n20270 & n21163 ;
  assign n21181 = n21180 ^ n21164 ;
  assign n21184 = n21183 ^ n21181 ;
  assign n21185 = n20250 ^ n20219 ;
  assign n21186 = n21185 ^ n20241 ;
  assign n21187 = n21186 ^ n20219 ;
  assign n21188 = n20219 ^ n19999 ;
  assign n21189 = n21188 ^ n20219 ;
  assign n21190 = ~n21187 & ~n21189 ;
  assign n21191 = n21190 ^ n20219 ;
  assign n21192 = ~n20270 & n21191 ;
  assign n21193 = n21184 & ~n21192 ;
  assign n21194 = ~n20269 & n21193 ;
  assign n21195 = n21194 ^ n17962 ;
  assign n21196 = n21195 ^ x72 ;
  assign n21197 = ~n21154 & n21196 ;
  assign n21198 = n21197 ^ n21196 ;
  assign n21200 = n19856 ^ x93 ;
  assign n21201 = n19050 ^ x84 ;
  assign n21296 = n21200 & ~n21201 ;
  assign n21297 = n21296 ^ n21201 ;
  assign n21233 = n19549 & n19709 ;
  assign n21211 = n19657 ^ n19627 ;
  assign n21210 = n20372 ^ n19637 ;
  assign n21212 = n21211 ^ n21210 ;
  assign n21213 = n21210 ^ n19548 ;
  assign n21215 = n19549 & n21213 ;
  assign n21216 = n21215 ^ n19548 ;
  assign n21217 = n21212 & n21216 ;
  assign n21218 = n21217 ^ n21210 ;
  assign n21227 = n21218 ^ n19719 ;
  assign n21219 = n21218 ^ n20371 ;
  assign n21220 = n21219 ^ n19653 ;
  assign n21221 = n21220 ^ n21218 ;
  assign n21222 = n21218 ^ n19548 ;
  assign n21223 = n21222 ^ n21218 ;
  assign n21224 = ~n21221 & n21223 ;
  assign n21225 = n21224 ^ n21218 ;
  assign n21226 = n19549 & n21225 ;
  assign n21228 = n21227 ^ n21226 ;
  assign n21209 = n19666 & n19687 ;
  assign n21229 = n21228 ^ n21209 ;
  assign n21202 = n19700 ^ n19548 ;
  assign n21203 = n21202 ^ n19700 ;
  assign n21204 = n19651 ^ n19641 ;
  assign n21205 = n21204 ^ n19700 ;
  assign n21206 = ~n21203 & ~n21205 ;
  assign n21207 = n21206 ^ n19700 ;
  assign n21208 = n19550 & n21207 ;
  assign n21230 = n21229 ^ n21208 ;
  assign n21231 = ~n19692 & n21230 ;
  assign n21232 = n21231 ^ n20125 ;
  assign n21234 = n21233 ^ n21232 ;
  assign n21235 = ~n19686 & n21234 ;
  assign n21236 = n21235 ^ n17070 ;
  assign n21237 = n21236 ^ x91 ;
  assign n21239 = ~n19227 & n19356 ;
  assign n21238 = n19351 ^ n17074 ;
  assign n21240 = n21239 ^ n21238 ;
  assign n21241 = n21240 ^ x70 ;
  assign n21242 = ~n21237 & ~n21241 ;
  assign n21243 = n21242 ^ n21241 ;
  assign n21246 = n17801 ^ x110 ;
  assign n21247 = n19545 ^ x116 ;
  assign n21248 = ~n21246 & n21247 ;
  assign n21259 = n21248 ^ n21246 ;
  assign n21260 = n21259 ^ n21247 ;
  assign n21275 = ~n21243 & n21260 ;
  assign n21244 = n21243 ^ n21237 ;
  assign n21245 = n21244 ^ n21241 ;
  assign n21272 = ~n21245 & n21260 ;
  assign n21267 = n21246 ^ n21241 ;
  assign n21268 = n21267 ^ n21247 ;
  assign n21269 = ~n21259 & n21268 ;
  assign n21270 = n21269 ^ n21259 ;
  assign n21266 = n21242 & ~n21259 ;
  assign n21271 = n21270 ^ n21266 ;
  assign n21273 = n21272 ^ n21271 ;
  assign n21301 = n21275 ^ n21273 ;
  assign n21261 = n21260 ^ n21246 ;
  assign n21262 = ~n21244 & n21261 ;
  assign n21251 = n21241 ^ n21237 ;
  assign n21252 = n21247 ^ n21241 ;
  assign n21253 = n21252 ^ n21247 ;
  assign n21254 = n21247 ^ n21246 ;
  assign n21255 = n21254 ^ n21247 ;
  assign n21256 = ~n21253 & n21255 ;
  assign n21257 = n21256 ^ n21247 ;
  assign n21258 = ~n21251 & n21257 ;
  assign n21263 = n21262 ^ n21258 ;
  assign n21264 = ~n21246 & n21263 ;
  assign n21299 = n21264 ^ n21263 ;
  assign n21300 = n21299 ^ n21271 ;
  assign n21302 = n21301 ^ n21300 ;
  assign n21334 = n21302 ^ n21260 ;
  assign n21335 = ~n21297 & n21334 ;
  assign n21305 = n21301 ^ n21245 ;
  assign n21249 = ~n21245 & n21248 ;
  assign n21250 = n21249 ^ n21248 ;
  assign n21265 = n21264 ^ n21250 ;
  assign n21279 = n21275 ^ n21265 ;
  assign n21280 = n21279 ^ n21262 ;
  assign n21277 = n21237 & n21254 ;
  assign n21278 = n21277 ^ n21244 ;
  assign n21281 = n21280 ^ n21278 ;
  assign n21282 = n21281 ^ n21269 ;
  assign n21283 = n21282 ^ n21271 ;
  assign n21276 = n21275 ^ n21249 ;
  assign n21284 = n21283 ^ n21276 ;
  assign n21306 = n21305 ^ n21284 ;
  assign n21333 = ~n21297 & n21306 ;
  assign n21336 = n21335 ^ n21333 ;
  assign n21327 = n21299 ^ n21201 ;
  assign n21328 = n21327 ^ n21299 ;
  assign n21304 = n21281 ^ n21272 ;
  assign n21307 = n21306 ^ n21304 ;
  assign n21308 = n21307 ^ n21271 ;
  assign n21303 = n21280 ^ n21249 ;
  assign n21309 = n21308 ^ n21303 ;
  assign n21287 = n21284 ^ n21268 ;
  assign n21310 = n21309 ^ n21287 ;
  assign n21311 = n21310 ^ n21302 ;
  assign n21312 = n21311 ^ n21264 ;
  assign n21329 = n21312 ^ n21299 ;
  assign n21330 = ~n21328 & n21329 ;
  assign n21331 = n21330 ^ n21299 ;
  assign n21332 = ~n21200 & n21331 ;
  assign n21337 = n21336 ^ n21332 ;
  assign n21338 = n21337 ^ n17991 ;
  assign n21313 = n21312 ^ n21266 ;
  assign n21298 = n21263 ^ n21242 ;
  assign n21314 = n21313 ^ n21298 ;
  assign n21315 = n21314 ^ n21249 ;
  assign n21316 = ~n21297 & n21315 ;
  assign n21285 = n21284 ^ n21269 ;
  assign n21286 = ~n21201 & ~n21285 ;
  assign n21288 = n21287 ^ n21286 ;
  assign n21317 = n21316 ^ n21288 ;
  assign n21289 = n21268 ^ n21258 ;
  assign n21290 = n21289 ^ n21288 ;
  assign n21274 = n21273 ^ n21265 ;
  assign n21291 = n21290 ^ n21274 ;
  assign n21292 = n21291 ^ n21288 ;
  assign n21293 = ~n21201 & ~n21292 ;
  assign n21294 = n21293 ^ n21290 ;
  assign n21295 = ~n21200 & ~n21294 ;
  assign n21318 = n21317 ^ n21295 ;
  assign n21319 = n21201 ^ n21200 ;
  assign n21320 = n21314 ^ n21304 ;
  assign n21321 = n21304 ^ n21201 ;
  assign n21322 = n21321 ^ n21304 ;
  assign n21323 = ~n21320 & n21322 ;
  assign n21324 = n21323 ^ n21304 ;
  assign n21325 = n21319 & ~n21324 ;
  assign n21326 = n21318 & ~n21325 ;
  assign n21339 = n21338 ^ n21326 ;
  assign n21340 = n21339 ^ x123 ;
  assign n21402 = n19874 ^ n19868 ;
  assign n21403 = n21402 ^ n19874 ;
  assign n21404 = n19874 ^ n19368 ;
  assign n21405 = n21404 ^ n19874 ;
  assign n21406 = n21403 & ~n21405 ;
  assign n21407 = n21406 ^ n19874 ;
  assign n21408 = ~n19547 & n21407 ;
  assign n21409 = n21408 ^ n19874 ;
  assign n21432 = n19913 ^ n19873 ;
  assign n21433 = n21432 ^ n19899 ;
  assign n21434 = n21433 ^ n19873 ;
  assign n21435 = n19873 ^ n19368 ;
  assign n21436 = n21435 ^ n19873 ;
  assign n21437 = ~n21434 & n21436 ;
  assign n21438 = n21437 ^ n19873 ;
  assign n21439 = n19547 & n21438 ;
  assign n21440 = n21439 ^ n19873 ;
  assign n21425 = n19940 ^ n19901 ;
  assign n21423 = n19924 ^ n19877 ;
  assign n21424 = n21423 ^ n19914 ;
  assign n21426 = n21425 ^ n21424 ;
  assign n21427 = n21424 ^ n19546 ;
  assign n21428 = n21427 ^ n21424 ;
  assign n21429 = ~n21426 & n21428 ;
  assign n21430 = n21429 ^ n21424 ;
  assign n21431 = ~n19912 & n21430 ;
  assign n21441 = n21440 ^ n21431 ;
  assign n21442 = n21441 ^ n19926 ;
  assign n21417 = n19923 ^ n19920 ;
  assign n21418 = n19920 ^ n19546 ;
  assign n21419 = n21418 ^ n19920 ;
  assign n21420 = n21417 & n21419 ;
  assign n21421 = n21420 ^ n19920 ;
  assign n21422 = n19912 & n21421 ;
  assign n21443 = n21442 ^ n21422 ;
  assign n21410 = n19926 ^ n19910 ;
  assign n21411 = n19911 ^ n19816 ;
  assign n21414 = n19926 & ~n21411 ;
  assign n21415 = n21414 ^ n19911 ;
  assign n21416 = ~n21410 & ~n21415 ;
  assign n21444 = n21443 ^ n21416 ;
  assign n21445 = ~n21409 & n21444 ;
  assign n21446 = ~n19908 & n21445 ;
  assign n21447 = ~n19888 & n21446 ;
  assign n21448 = n21447 ^ n18043 ;
  assign n21449 = n21448 ^ x104 ;
  assign n21450 = ~n21340 & n21449 ;
  assign n21451 = n21450 ^ n21449 ;
  assign n21352 = n20626 ^ n20613 ;
  assign n21353 = n21352 ^ n20655 ;
  assign n21354 = n20547 & n21353 ;
  assign n21362 = n21354 ^ n20625 ;
  assign n21361 = n20650 ^ n20647 ;
  assign n21363 = n21362 ^ n21361 ;
  assign n21364 = n21363 ^ n21354 ;
  assign n21365 = ~n20547 & n21364 ;
  assign n21366 = n21365 ^ n21362 ;
  assign n21367 = ~n20548 & n21366 ;
  assign n21356 = n20617 & n20686 ;
  assign n21355 = n20550 & n20615 ;
  assign n21357 = n21356 ^ n21355 ;
  assign n21358 = n21357 ^ n21354 ;
  assign n21348 = n20636 ^ n20617 ;
  assign n21349 = ~n20715 & n21348 ;
  assign n21350 = n21349 ^ n20617 ;
  assign n21351 = ~n20690 & n21350 ;
  assign n21359 = n21358 ^ n21351 ;
  assign n21360 = n21359 ^ n20711 ;
  assign n21368 = n21367 ^ n21360 ;
  assign n21343 = n20657 ^ n20615 ;
  assign n21344 = n21343 ^ n20613 ;
  assign n21345 = n21344 ^ n20642 ;
  assign n21341 = n20658 ^ n20602 ;
  assign n21342 = n21341 ^ n20624 ;
  assign n21346 = n21345 ^ n21342 ;
  assign n21347 = n20550 & ~n21346 ;
  assign n21369 = n21368 ^ n21347 ;
  assign n21370 = n21369 ^ n20628 ;
  assign n21371 = n21370 ^ n20720 ;
  assign n21372 = n21371 ^ n16764 ;
  assign n21373 = n21372 ^ x114 ;
  assign n21388 = n20523 ^ n20439 ;
  assign n21389 = n21388 ^ n20528 ;
  assign n21382 = n20534 ^ n20438 ;
  assign n21383 = n21382 ^ n20521 ;
  assign n21381 = n20534 ^ n20525 ;
  assign n21384 = n21383 ^ n21381 ;
  assign n21385 = n21384 ^ n20521 ;
  assign n21386 = n20464 & n21385 ;
  assign n21387 = n21386 ^ n21383 ;
  assign n21390 = n21389 ^ n21387 ;
  assign n21391 = n21390 ^ n20528 ;
  assign n21392 = n20359 & ~n21391 ;
  assign n21393 = n21392 ^ n21390 ;
  assign n21374 = n20518 ^ n20509 ;
  assign n21375 = n21374 ^ n20530 ;
  assign n21376 = n21375 ^ n20505 ;
  assign n21377 = n21376 ^ n20503 ;
  assign n21378 = n20359 & n21377 ;
  assign n21379 = n21378 ^ n21376 ;
  assign n21380 = n21379 ^ n18191 ;
  assign n21394 = n21393 ^ n21380 ;
  assign n21395 = n21394 ^ n18191 ;
  assign n21396 = n20342 & ~n21395 ;
  assign n21397 = n21396 ^ n21380 ;
  assign n21398 = n21397 ^ x105 ;
  assign n21399 = ~n21373 & n21398 ;
  assign n21452 = n21399 ^ n21373 ;
  assign n21465 = n21452 ^ n21398 ;
  assign n21466 = n21451 & n21465 ;
  assign n21467 = n21466 ^ n21451 ;
  assign n21456 = n21451 ^ n21340 ;
  assign n21458 = ~n21373 & n21456 ;
  assign n21400 = n21340 & n21399 ;
  assign n21459 = n21458 ^ n21400 ;
  assign n21457 = ~n21452 & n21456 ;
  assign n21460 = n21459 ^ n21457 ;
  assign n21454 = n21450 & ~n21452 ;
  assign n21461 = n21460 ^ n21454 ;
  assign n21453 = n21451 & ~n21452 ;
  assign n21455 = n21454 ^ n21453 ;
  assign n21462 = n21461 ^ n21455 ;
  assign n21468 = n21467 ^ n21462 ;
  assign n21469 = n21198 & n21468 ;
  assign n21470 = n21450 & n21465 ;
  assign n21471 = n21154 & n21470 ;
  assign n21472 = n21196 ^ n21154 ;
  assign n21501 = n21457 ^ n21452 ;
  assign n21502 = n21501 ^ n21455 ;
  assign n21474 = n21450 ^ n21340 ;
  assign n21475 = n21465 & ~n21474 ;
  assign n21476 = n21475 ^ n21466 ;
  assign n21477 = n21476 ^ n21465 ;
  assign n21478 = n21477 ^ n21470 ;
  assign n21489 = n21478 ^ n21460 ;
  assign n21484 = n21398 ^ n21373 ;
  assign n21486 = n21449 ^ n21373 ;
  assign n21487 = n21486 ^ n21340 ;
  assign n21488 = n21484 & n21487 ;
  assign n21490 = n21489 ^ n21488 ;
  assign n21485 = n21484 ^ n21470 ;
  assign n21491 = n21490 ^ n21485 ;
  assign n21492 = n21491 ^ n21457 ;
  assign n21493 = n21492 ^ n21373 ;
  assign n21494 = n21493 ^ n21461 ;
  assign n21482 = n21398 ^ n21340 ;
  assign n21483 = n21482 ^ n21449 ;
  assign n21495 = n21494 ^ n21483 ;
  assign n21473 = n21458 ^ n21456 ;
  assign n21479 = n21478 ^ n21473 ;
  assign n21480 = n21479 ^ n21476 ;
  assign n21496 = n21495 ^ n21480 ;
  assign n21514 = n21502 ^ n21496 ;
  assign n21515 = n21514 ^ n21400 ;
  assign n21513 = n21457 ^ n21373 ;
  assign n21516 = n21515 ^ n21513 ;
  assign n21517 = ~n21154 & n21516 ;
  assign n21511 = n21475 ^ n21473 ;
  assign n21497 = n21496 ^ n21468 ;
  assign n21498 = n21497 ^ n21478 ;
  assign n21499 = n21498 ^ n21470 ;
  assign n21481 = n21480 ^ n21373 ;
  assign n21500 = n21499 ^ n21481 ;
  assign n21503 = n21502 ^ n21466 ;
  assign n21504 = n21503 ^ n21497 ;
  assign n21505 = n21502 ^ n21196 ;
  assign n21506 = n21472 & n21505 ;
  assign n21507 = n21506 ^ n21196 ;
  assign n21508 = ~n21504 & ~n21507 ;
  assign n21509 = n21508 ^ n21502 ;
  assign n21510 = ~n21500 & n21509 ;
  assign n21512 = n21511 ^ n21510 ;
  assign n21518 = n21517 ^ n21512 ;
  assign n21519 = n21472 & ~n21518 ;
  assign n21520 = n21519 ^ n21510 ;
  assign n21521 = ~n21471 & n21520 ;
  assign n21522 = ~n21469 & n21521 ;
  assign n21199 = n21198 ^ n21154 ;
  assign n21401 = n21400 ^ n21399 ;
  assign n21463 = n21462 ^ n21401 ;
  assign n21464 = n21199 & n21463 ;
  assign n21523 = n21522 ^ n21464 ;
  assign n21524 = n21472 ^ n21458 ;
  assign n21526 = n21461 ^ n21458 ;
  assign n21525 = n21461 ^ n21196 ;
  assign n21527 = n21526 ^ n21525 ;
  assign n21528 = n21526 ^ n21462 ;
  assign n21529 = n21528 ^ n21526 ;
  assign n21530 = ~n21527 & n21529 ;
  assign n21531 = n21530 ^ n21526 ;
  assign n21532 = ~n21524 & n21531 ;
  assign n21533 = n21532 ^ n21458 ;
  assign n21534 = n21523 & ~n21533 ;
  assign n21535 = n21534 ^ n20462 ;
  assign n21536 = n21535 ^ x93 ;
  assign n21546 = n19999 & n20227 ;
  assign n21554 = n21546 ^ n20258 ;
  assign n21552 = n20224 & ~n20285 ;
  assign n21553 = n21552 ^ n21166 ;
  assign n21555 = n21554 ^ n21553 ;
  assign n21548 = n20242 ^ n20214 ;
  assign n21549 = ~n19999 & n21548 ;
  assign n21544 = n20235 ^ n20214 ;
  assign n21545 = n21544 ^ n20253 ;
  assign n21547 = n21546 ^ n21545 ;
  assign n21550 = n21549 ^ n21547 ;
  assign n21551 = n20270 & n21550 ;
  assign n21556 = n21555 ^ n21551 ;
  assign n21539 = n20258 ^ n20021 ;
  assign n21540 = n21539 ^ n20258 ;
  assign n21541 = ~n20297 & ~n21540 ;
  assign n21542 = n21541 ^ n20258 ;
  assign n21543 = ~n19999 & ~n21542 ;
  assign n21557 = n21556 ^ n21543 ;
  assign n21558 = ~n21183 & n21557 ;
  assign n21559 = ~n21192 & n21558 ;
  assign n21560 = ~n20296 & n21559 ;
  assign n21561 = ~n20269 & n21560 ;
  assign n21562 = n21561 ^ n18685 ;
  assign n21563 = n21562 ^ x124 ;
  assign n21564 = n21392 ^ n21387 ;
  assign n21565 = n21564 ^ n21379 ;
  assign n21566 = n21379 ^ n20342 ;
  assign n21567 = n21566 ^ n21379 ;
  assign n21568 = ~n21565 & ~n21567 ;
  assign n21569 = n21568 ^ n21379 ;
  assign n21570 = n21389 & ~n21569 ;
  assign n21571 = n21570 ^ n18398 ;
  assign n21572 = n21571 ^ x110 ;
  assign n21721 = n21563 & n21572 ;
  assign n21722 = n21721 ^ n21572 ;
  assign n21723 = n21722 ^ n21563 ;
  assign n21590 = n19910 ^ n19871 ;
  assign n21591 = n19920 ^ n19911 ;
  assign n21592 = n19911 ^ n19871 ;
  assign n21593 = n21592 ^ n19911 ;
  assign n21594 = ~n21591 & ~n21593 ;
  assign n21595 = n21594 ^ n19911 ;
  assign n21596 = n21590 & ~n21595 ;
  assign n21588 = ~n19546 & n19870 ;
  assign n21577 = n19924 ^ n19921 ;
  assign n21578 = n21577 ^ n19923 ;
  assign n21583 = n21578 ^ n19900 ;
  assign n21579 = n19901 ^ n19864 ;
  assign n21580 = n21579 ^ n21578 ;
  assign n21573 = n19869 ^ n19813 ;
  assign n21574 = n21573 ^ n19899 ;
  assign n21575 = n21574 ^ n19895 ;
  assign n21576 = n21575 ^ n19870 ;
  assign n21581 = n21580 ^ n21576 ;
  assign n21582 = ~n19546 & n21581 ;
  assign n21584 = n21583 ^ n21582 ;
  assign n21585 = ~n19912 & ~n21584 ;
  assign n21586 = n21585 ^ n19871 ;
  assign n21587 = n21586 ^ n21422 ;
  assign n21589 = n21588 ^ n21587 ;
  assign n21597 = n21596 ^ n21589 ;
  assign n21598 = ~n21409 & ~n21597 ;
  assign n21599 = ~n19916 & n21598 ;
  assign n21600 = n21599 ^ n18603 ;
  assign n21601 = n21600 ^ x93 ;
  assign n21610 = n20820 ^ n20799 ;
  assign n21611 = n21610 ^ n20848 ;
  assign n21612 = n20825 & ~n21611 ;
  assign n21613 = n21612 ^ n20848 ;
  assign n21620 = n21613 ^ n20864 ;
  assign n21621 = n21620 ^ n20837 ;
  assign n21615 = n20858 ^ n20808 ;
  assign n21616 = n21615 ^ n20866 ;
  assign n21617 = n20825 & ~n21616 ;
  assign n21609 = n20866 ^ n20806 ;
  assign n21614 = n21613 ^ n21609 ;
  assign n21618 = n21617 ^ n21614 ;
  assign n21619 = n20828 & n21618 ;
  assign n21622 = n21621 ^ n21619 ;
  assign n21602 = n20864 ^ n20853 ;
  assign n21603 = n20869 ^ n20829 ;
  assign n21604 = n21603 ^ n20826 ;
  assign n21605 = n20853 ^ n20826 ;
  assign n21606 = n21604 & ~n21605 ;
  assign n21607 = n21606 ^ n20826 ;
  assign n21608 = ~n21602 & n21607 ;
  assign n21623 = n21622 ^ n21608 ;
  assign n21624 = n20844 ^ n20803 ;
  assign n21625 = n21624 ^ n20853 ;
  assign n21626 = n20853 ^ n20824 ;
  assign n21627 = n21626 ^ n20853 ;
  assign n21628 = ~n21625 & ~n21627 ;
  assign n21629 = n21628 ^ n20853 ;
  assign n21630 = n20825 & ~n21629 ;
  assign n21631 = n21623 & ~n21630 ;
  assign n21632 = n20820 ^ n20794 ;
  assign n21635 = ~n20824 & ~n21632 ;
  assign n21636 = n21635 ^ n20820 ;
  assign n21637 = ~n20825 & ~n21636 ;
  assign n21638 = n21631 & ~n21637 ;
  assign n21639 = n21638 ^ n20870 ;
  assign n21640 = ~n20792 & n21639 ;
  assign n21641 = n21640 ^ n19581 ;
  assign n21642 = n21641 ^ x92 ;
  assign n21643 = ~n21601 & ~n21642 ;
  assign n21724 = n21643 ^ n21642 ;
  assign n21725 = n21724 ^ n21601 ;
  assign n21726 = n21725 ^ n21642 ;
  assign n21644 = n21296 ^ n21200 ;
  assign n21663 = n21289 ^ n21277 ;
  assign n21661 = n21271 ^ n21243 ;
  assign n21662 = n21661 ^ n21279 ;
  assign n21664 = n21663 ^ n21662 ;
  assign n21665 = n21644 & n21664 ;
  assign n21657 = n21299 ^ n21265 ;
  assign n21654 = n21264 ^ n21254 ;
  assign n21655 = n21654 ^ n21237 ;
  assign n21656 = ~n21201 & n21655 ;
  assign n21658 = n21657 ^ n21656 ;
  assign n21659 = n21319 & n21658 ;
  assign n21660 = n21659 ^ n21657 ;
  assign n21666 = n21665 ^ n21660 ;
  assign n21647 = n21311 ^ n21262 ;
  assign n21648 = n21647 ^ n21287 ;
  assign n21649 = n21287 ^ n21201 ;
  assign n21650 = n21649 ^ n21287 ;
  assign n21651 = ~n21648 & ~n21650 ;
  assign n21652 = n21651 ^ n21287 ;
  assign n21653 = ~n21200 & ~n21652 ;
  assign n21667 = n21666 ^ n21653 ;
  assign n21646 = n21283 & ~n21297 ;
  assign n21668 = n21667 ^ n21646 ;
  assign n21669 = n21668 ^ n21335 ;
  assign n21670 = n21669 ^ n21333 ;
  assign n21671 = n21670 ^ n18434 ;
  assign n21645 = n21312 & n21644 ;
  assign n21672 = n21671 ^ n21645 ;
  assign n21673 = n21672 ^ x67 ;
  assign n21688 = n20629 ^ n20610 ;
  assign n21689 = n20549 & n21688 ;
  assign n21675 = n20548 & ~n20645 ;
  assign n21676 = n21675 ^ n20632 ;
  assign n21685 = n21676 ^ n20703 ;
  assign n21678 = n21676 ^ n20658 ;
  assign n21677 = n21676 ^ n20624 ;
  assign n21679 = n21678 ^ n21677 ;
  assign n21680 = n21678 ^ n20547 ;
  assign n21681 = n21680 ^ n21678 ;
  assign n21682 = n21679 & n21681 ;
  assign n21683 = n21682 ^ n21678 ;
  assign n21684 = ~n20690 & n21683 ;
  assign n21686 = n21685 ^ n21684 ;
  assign n21687 = ~n20718 & ~n21686 ;
  assign n21690 = n21689 ^ n21687 ;
  assign n21674 = n20550 & n20613 ;
  assign n21691 = n21690 ^ n21674 ;
  assign n21696 = n20642 ^ n20547 ;
  assign n21697 = n21696 ^ n20642 ;
  assign n21698 = n21345 & n21697 ;
  assign n21699 = n21698 ^ n20642 ;
  assign n21700 = ~n20548 & n21699 ;
  assign n21701 = n21691 & n21700 ;
  assign n21692 = n21691 ^ n21357 ;
  assign n21702 = n21701 ^ n21692 ;
  assign n21703 = ~n21351 & n21702 ;
  assign n21704 = ~n20662 & n21703 ;
  assign n21705 = n21704 ^ n19618 ;
  assign n21706 = n21705 ^ x78 ;
  assign n21707 = ~n21673 & n21706 ;
  assign n21727 = n21707 ^ n21673 ;
  assign n21728 = ~n21726 & ~n21727 ;
  assign n21729 = ~n21723 & n21728 ;
  assign n21708 = n21707 ^ n21706 ;
  assign n21709 = n21708 ^ n21673 ;
  assign n21710 = n21643 & n21709 ;
  assign n21711 = n21710 ^ n21572 ;
  assign n21712 = n21711 ^ n21710 ;
  assign n21713 = n21706 ^ n21673 ;
  assign n21714 = n21643 & ~n21713 ;
  assign n21715 = n21714 ^ n21710 ;
  assign n21718 = n21712 & n21715 ;
  assign n21719 = n21718 ^ n21710 ;
  assign n21720 = ~n21563 & n21719 ;
  assign n21730 = n21729 ^ n21720 ;
  assign n21731 = n21723 ^ n21572 ;
  assign n21732 = n21728 & n21731 ;
  assign n21737 = n21708 & ~n21725 ;
  assign n21736 = ~n21725 & ~n21727 ;
  assign n21738 = n21737 ^ n21736 ;
  assign n21734 = n21707 & ~n21725 ;
  assign n21735 = n21734 ^ n21725 ;
  assign n21739 = n21738 ^ n21735 ;
  assign n21733 = ~n21724 & ~n21727 ;
  assign n21740 = n21739 ^ n21733 ;
  assign n21741 = n21740 ^ n21737 ;
  assign n21742 = ~n21723 & ~n21741 ;
  assign n21743 = n21734 ^ n21710 ;
  assign n21744 = n21710 ^ n21563 ;
  assign n21745 = n21744 ^ n21710 ;
  assign n21746 = n21743 & n21745 ;
  assign n21747 = n21746 ^ n21710 ;
  assign n21748 = n21572 & n21747 ;
  assign n21782 = n21715 ^ n21643 ;
  assign n21767 = n21708 & ~n21726 ;
  assign n21783 = n21782 ^ n21767 ;
  assign n21784 = n21783 ^ n21728 ;
  assign n21785 = n21728 ^ n21572 ;
  assign n21786 = n21785 ^ n21728 ;
  assign n21787 = n21784 & ~n21786 ;
  assign n21788 = n21787 ^ n21728 ;
  assign n21789 = ~n21563 & n21788 ;
  assign n21749 = n21708 & ~n21724 ;
  assign n21761 = n21749 ^ n21739 ;
  assign n21762 = n21761 ^ n21724 ;
  assign n21759 = n21709 & ~n21724 ;
  assign n21760 = n21759 ^ n21740 ;
  assign n21763 = n21762 ^ n21760 ;
  assign n21764 = n21643 & ~n21706 ;
  assign n21765 = n21764 ^ n21715 ;
  assign n21751 = n21707 & ~n21726 ;
  assign n21768 = n21765 ^ n21751 ;
  assign n21773 = n21768 ^ n21759 ;
  assign n21769 = n21768 ^ n21767 ;
  assign n21770 = n21769 ^ n21728 ;
  assign n21766 = n21765 ^ n21726 ;
  assign n21771 = n21770 ^ n21766 ;
  assign n21772 = n21771 ^ n21733 ;
  assign n21774 = n21773 ^ n21772 ;
  assign n21775 = n21772 ^ n21572 ;
  assign n21776 = n21775 ^ n21772 ;
  assign n21777 = ~n21774 & ~n21776 ;
  assign n21778 = n21777 ^ n21772 ;
  assign n21779 = n21763 & n21778 ;
  assign n21780 = n21563 & ~n21779 ;
  assign n21750 = n21749 ^ n21722 ;
  assign n21752 = n21751 ^ n21731 ;
  assign n21755 = ~n21749 & ~n21752 ;
  assign n21756 = n21755 ^ n21731 ;
  assign n21757 = n21750 & n21756 ;
  assign n21758 = n21757 ^ n21722 ;
  assign n21781 = n21780 ^ n21758 ;
  assign n21790 = n21789 ^ n21781 ;
  assign n21791 = n21790 ^ n21734 ;
  assign n21793 = n21791 ^ n21790 ;
  assign n21794 = n21790 ^ n21572 ;
  assign n21795 = n21794 ^ n21790 ;
  assign n21796 = n21790 ^ n21780 ;
  assign n21797 = n21796 ^ n21790 ;
  assign n21798 = ~n21795 & ~n21797 ;
  assign n21799 = n21793 & n21798 ;
  assign n21800 = n21799 ^ n21793 ;
  assign n21801 = n21800 ^ n21791 ;
  assign n21802 = ~n21748 & ~n21801 ;
  assign n21803 = n21783 ^ n21771 ;
  assign n21804 = n21771 ^ n21572 ;
  assign n21805 = n21804 ^ n21771 ;
  assign n21806 = ~n21803 & n21805 ;
  assign n21807 = n21806 ^ n21771 ;
  assign n21808 = n21563 & ~n21807 ;
  assign n21809 = n21802 & ~n21808 ;
  assign n21810 = ~n21742 & n21809 ;
  assign n21811 = ~n21732 & n21810 ;
  assign n21812 = ~n21730 & n21811 ;
  assign n21814 = n21759 ^ n21736 ;
  assign n21813 = n21737 ^ n21733 ;
  assign n21815 = n21814 ^ n21813 ;
  assign n21816 = n21814 ^ n21563 ;
  assign n21817 = n21816 ^ n21814 ;
  assign n21818 = n21815 & ~n21817 ;
  assign n21819 = n21818 ^ n21814 ;
  assign n21820 = n21572 & n21819 ;
  assign n21821 = n21812 & ~n21820 ;
  assign n21822 = n21821 ^ n19726 ;
  assign n21823 = n21822 ^ x75 ;
  assign n22649 = ~n21536 & ~n21823 ;
  assign n22650 = n22649 ^ n21823 ;
  assign n22563 = n20723 ^ x120 ;
  assign n22551 = n21339 ^ x73 ;
  assign n22106 = n19299 & n19319 ;
  assign n22508 = n19068 ^ n19054 ;
  assign n22509 = ~n19089 & n19309 ;
  assign n22510 = n19283 & n22509 ;
  assign n22511 = n22508 & n22510 ;
  assign n22512 = n22511 ^ n22509 ;
  assign n22513 = n22512 ^ n19309 ;
  assign n22514 = n22513 ^ n19083 ;
  assign n22502 = n19062 ^ n19058 ;
  assign n22107 = n19077 ^ n19069 ;
  assign n22503 = n22502 ^ n22107 ;
  assign n22501 = n19092 ^ n19086 ;
  assign n22504 = n22503 ^ n22501 ;
  assign n22505 = ~n19283 & ~n22504 ;
  assign n22506 = n22505 ^ n19083 ;
  assign n22507 = ~n17802 & n22506 ;
  assign n22515 = n22514 ^ n22507 ;
  assign n22516 = n19081 ^ n17802 ;
  assign n22517 = n22516 ^ n19081 ;
  assign n22520 = n19075 & ~n19283 ;
  assign n22521 = n22520 ^ n19081 ;
  assign n22522 = n22517 & n22521 ;
  assign n22523 = n22522 ^ n19081 ;
  assign n22524 = ~n22515 & ~n22523 ;
  assign n22136 = n19087 ^ n19075 ;
  assign n22137 = n22136 ^ n19087 ;
  assign n22138 = n19283 & n22137 ;
  assign n22139 = n22138 ^ n19087 ;
  assign n22140 = n17802 & ~n22139 ;
  assign n22525 = n22524 ^ n22140 ;
  assign n22526 = ~n19307 & n22525 ;
  assign n22527 = ~n22106 & n22526 ;
  assign n22528 = n22527 ^ n19157 ;
  assign n22529 = n22528 ^ x106 ;
  assign n22497 = n21195 ^ x80 ;
  assign n22534 = n22529 ^ n22497 ;
  assign n22500 = n20893 ^ x97 ;
  assign n22576 = n22534 ^ n22500 ;
  assign n22577 = n22576 ^ n22534 ;
  assign n22579 = ~n22529 & ~n22577 ;
  assign n22580 = n22579 ^ n22534 ;
  assign n21953 = n21091 ^ n21072 ;
  assign n21954 = ~n20983 & n21953 ;
  assign n21955 = n21954 ^ n21091 ;
  assign n21956 = n20982 & n21955 ;
  assign n21948 = n20984 & n21083 ;
  assign n22480 = n21091 ^ n21062 ;
  assign n22481 = n22480 ^ n21069 ;
  assign n22482 = n22481 ^ n21064 ;
  assign n22483 = ~n20983 & n22482 ;
  assign n22484 = n22483 ^ n21073 ;
  assign n22485 = ~n20982 & n22484 ;
  assign n22486 = n22485 ^ n21106 ;
  assign n22479 = n21081 & ~n21136 ;
  assign n22487 = n22486 ^ n22479 ;
  assign n22476 = n21092 ^ n21074 ;
  assign n21957 = n21101 ^ n21069 ;
  assign n22477 = n22476 ^ n21957 ;
  assign n22478 = ~n21115 & n22477 ;
  assign n22488 = n22487 ^ n22478 ;
  assign n22489 = n22488 ^ n21082 ;
  assign n21985 = n21117 ^ n21103 ;
  assign n21986 = n21103 ^ n20983 ;
  assign n21987 = n21986 ^ n21103 ;
  assign n21988 = n21985 & ~n21987 ;
  assign n21989 = n21988 ^ n21103 ;
  assign n21990 = n20982 & n21989 ;
  assign n22490 = n22489 ^ n21990 ;
  assign n22475 = ~n20985 & n21096 ;
  assign n22491 = n22490 ^ n22475 ;
  assign n22468 = n21082 ^ n21075 ;
  assign n22469 = n22468 ^ n21082 ;
  assign n22470 = n21082 ^ n20983 ;
  assign n22471 = n22470 ^ n21082 ;
  assign n22472 = n22469 & n22471 ;
  assign n22473 = n22472 ^ n21082 ;
  assign n22474 = n20982 & n22473 ;
  assign n22492 = n22491 ^ n22474 ;
  assign n22493 = ~n21948 & ~n22492 ;
  assign n22494 = ~n21956 & n22493 ;
  assign n22495 = n22494 ^ n19181 ;
  assign n22496 = n22495 ^ x115 ;
  assign n22581 = n22534 ^ n22496 ;
  assign n22582 = n22581 ^ n22500 ;
  assign n22583 = n22582 ^ n22529 ;
  assign n22584 = ~n22580 & ~n22583 ;
  assign n22585 = n22584 ^ n22534 ;
  assign n22549 = n22497 ^ n22496 ;
  assign n22564 = n22549 ^ n22500 ;
  assign n22566 = n22549 ^ n22497 ;
  assign n22569 = ~n22534 & ~n22566 ;
  assign n22570 = n22569 ^ n22497 ;
  assign n22571 = n22564 & ~n22570 ;
  assign n22572 = n22571 ^ n22500 ;
  assign n22586 = n22585 ^ n22572 ;
  assign n22498 = n22496 & ~n22497 ;
  assign n22499 = n22498 ^ n22496 ;
  assign n22532 = n22500 ^ n22496 ;
  assign n22530 = n22529 ^ n22500 ;
  assign n22533 = n22532 ^ n22530 ;
  assign n22537 = n22530 ^ n22529 ;
  assign n22538 = n22534 & ~n22537 ;
  assign n22539 = n22538 ^ n22529 ;
  assign n22540 = n22533 & n22539 ;
  assign n22541 = n22540 ^ n22532 ;
  assign n22542 = n22498 & n22541 ;
  assign n22531 = n22500 & n22530 ;
  assign n22543 = n22542 ^ n22531 ;
  assign n22544 = n22543 ^ n22500 ;
  assign n22545 = n22544 ^ n22529 ;
  assign n22546 = n22545 ^ n22543 ;
  assign n22547 = ~n22499 & ~n22546 ;
  assign n22548 = n22547 ^ n22544 ;
  assign n22575 = n22548 ^ n22497 ;
  assign n22587 = n22586 ^ n22575 ;
  assign n22574 = n22532 ^ n22529 ;
  assign n22588 = n22587 ^ n22574 ;
  assign n22565 = n22564 ^ n22543 ;
  assign n22573 = n22572 ^ n22565 ;
  assign n22589 = n22588 ^ n22573 ;
  assign n22590 = n22551 & ~n22589 ;
  assign n22591 = n22590 ^ n22588 ;
  assign n22552 = n22530 ^ n22496 ;
  assign n22553 = n22552 ^ n22548 ;
  assign n22554 = n22553 ^ n22496 ;
  assign n22555 = n22554 ^ n22531 ;
  assign n22556 = n22555 ^ n22553 ;
  assign n22557 = n22553 ^ n22497 ;
  assign n22558 = n22557 ^ n22553 ;
  assign n22559 = n22556 & ~n22558 ;
  assign n22560 = n22559 ^ n22553 ;
  assign n22561 = n22551 & ~n22560 ;
  assign n22550 = n22549 ^ n22548 ;
  assign n22562 = n22561 ^ n22550 ;
  assign n22592 = n22591 ^ n22562 ;
  assign n22593 = ~n22563 & n22592 ;
  assign n22594 = n22593 ^ n22563 ;
  assign n22595 = n22594 ^ n22562 ;
  assign n22596 = n22595 ^ n19367 ;
  assign n22597 = n22596 ^ x108 ;
  assign n21947 = n20545 ^ x126 ;
  assign n21852 = n20547 & ~n20652 ;
  assign n21851 = n20548 & n20623 ;
  assign n21853 = n21852 ^ n21851 ;
  assign n21827 = n20634 ^ n20602 ;
  assign n21828 = n21827 ^ n20658 ;
  assign n21829 = ~n20548 & ~n21828 ;
  assign n21830 = n21829 ^ n20643 ;
  assign n21831 = ~n20690 & ~n21830 ;
  assign n21832 = ~n20635 & ~n20659 ;
  assign n21833 = n20672 ^ n20614 ;
  assign n21834 = n20548 & n21833 ;
  assign n21835 = n21834 ^ n20549 ;
  assign n21836 = n21835 ^ n20547 ;
  assign n21837 = n21836 ^ n21834 ;
  assign n21838 = n21832 & n21837 ;
  assign n21839 = n21838 ^ n21835 ;
  assign n21840 = n21839 ^ n20547 ;
  assign n21841 = n21840 ^ n21839 ;
  assign n21842 = n21840 ^ n20613 ;
  assign n21843 = n21842 ^ n21840 ;
  assign n21844 = n21840 ^ n21834 ;
  assign n21845 = n21844 ^ n21840 ;
  assign n21846 = ~n21843 & n21845 ;
  assign n21847 = ~n21841 & n21846 ;
  assign n21848 = n21847 ^ n21841 ;
  assign n21849 = n21848 ^ n21839 ;
  assign n21850 = ~n21831 & ~n21849 ;
  assign n21854 = n21853 ^ n21850 ;
  assign n21855 = n21854 ^ n21355 ;
  assign n21856 = ~n20696 & n21855 ;
  assign n21825 = n20720 ^ n18906 ;
  assign n21826 = n21825 ^ n20718 ;
  assign n21857 = n21856 ^ n21826 ;
  assign n21858 = n21857 ^ x69 ;
  assign n21905 = n21335 ^ n18854 ;
  assign n21887 = n21300 ^ n21282 ;
  assign n21888 = n21887 ^ n21275 ;
  assign n21885 = n21304 ^ n21279 ;
  assign n21886 = n21885 ^ n21647 ;
  assign n21889 = n21888 ^ n21886 ;
  assign n21890 = ~n21200 & ~n21889 ;
  assign n21891 = n21890 ^ n21888 ;
  assign n21892 = n21201 & n21891 ;
  assign n21864 = n21662 ^ n21265 ;
  assign n21865 = n21864 ^ n21314 ;
  assign n21866 = n21314 ^ n21201 ;
  assign n21867 = n21319 ^ n21201 ;
  assign n21868 = ~n21866 & ~n21867 ;
  assign n21869 = n21868 ^ n21201 ;
  assign n21870 = n21865 & ~n21869 ;
  assign n21871 = n21870 ^ n21314 ;
  assign n21872 = n21871 ^ n21249 ;
  assign n21873 = n21872 ^ n21306 ;
  assign n21882 = n21873 ^ n21316 ;
  assign n21874 = n21873 ^ n21311 ;
  assign n21875 = n21874 ^ n21275 ;
  assign n21876 = n21875 ^ n21873 ;
  assign n21877 = n21873 ^ n21201 ;
  assign n21878 = n21877 ^ n21873 ;
  assign n21879 = n21876 & ~n21878 ;
  assign n21880 = n21879 ^ n21873 ;
  assign n21881 = ~n21200 & n21880 ;
  assign n21883 = n21882 ^ n21881 ;
  assign n21863 = n21296 & n21334 ;
  assign n21884 = n21883 ^ n21863 ;
  assign n21893 = n21892 ^ n21884 ;
  assign n21894 = ~n21325 & ~n21893 ;
  assign n21859 = n21281 ^ n21266 ;
  assign n21860 = ~n21200 & ~n21859 ;
  assign n21861 = n21860 ^ n21266 ;
  assign n21862 = ~n21201 & n21861 ;
  assign n21895 = n21894 ^ n21862 ;
  assign n21896 = ~n21646 & n21895 ;
  assign n21899 = n21266 ^ n21200 ;
  assign n21900 = n21899 ^ n21266 ;
  assign n21901 = n21313 & n21900 ;
  assign n21902 = n21901 ^ n21266 ;
  assign n21903 = n21201 & n21902 ;
  assign n21904 = n21896 & ~n21903 ;
  assign n21906 = n21905 ^ n21904 ;
  assign n21907 = n21906 ^ x84 ;
  assign n21908 = n21858 & n21907 ;
  assign n21939 = n21908 ^ n21858 ;
  assign n21940 = n21939 ^ n21907 ;
  assign n21909 = n19335 ^ x109 ;
  assign n21921 = n20815 ^ n20802 ;
  assign n21922 = n20826 & n21921 ;
  assign n21916 = n20890 ^ n20802 ;
  assign n21917 = n21916 ^ n21630 ;
  assign n21918 = n21917 ^ n21637 ;
  assign n21911 = n20788 ^ n20754 ;
  assign n21912 = n21911 ^ n20755 ;
  assign n21913 = n21912 ^ n20787 ;
  assign n21914 = ~n20813 & n21913 ;
  assign n21915 = ~n20828 & n21914 ;
  assign n21919 = n21918 ^ n21915 ;
  assign n21910 = ~n20819 & ~n20869 ;
  assign n21920 = n21919 ^ n21910 ;
  assign n21923 = n21922 ^ n21920 ;
  assign n21924 = n20864 ^ n20807 ;
  assign n21925 = n21924 ^ n20818 ;
  assign n21926 = n21925 ^ n21924 ;
  assign n21927 = n21924 ^ n20825 ;
  assign n21928 = n21927 ^ n21924 ;
  assign n21929 = ~n21926 & ~n21928 ;
  assign n21930 = n21929 ^ n21924 ;
  assign n21931 = n20828 & n21930 ;
  assign n21932 = n21923 & ~n21931 ;
  assign n21933 = n21932 ^ n18571 ;
  assign n21934 = n21933 ^ x102 ;
  assign n21935 = ~n21909 & n21934 ;
  assign n22002 = n21935 ^ n21934 ;
  assign n22019 = ~n21940 & n22002 ;
  assign n21936 = n21935 ^ n21909 ;
  assign n21937 = n21936 ^ n21934 ;
  assign n21943 = n21940 ^ n21858 ;
  assign n21944 = n21937 & n21943 ;
  assign n21945 = n21944 ^ n21937 ;
  assign n21941 = n21937 & ~n21940 ;
  assign n21938 = n21908 & n21937 ;
  assign n21942 = n21941 ^ n21938 ;
  assign n21946 = n21945 ^ n21942 ;
  assign n22045 = n22019 ^ n21946 ;
  assign n22035 = ~n21936 & n21943 ;
  assign n22017 = n21943 & n22002 ;
  assign n22043 = n22035 ^ n22017 ;
  assign n22042 = n21908 & n21935 ;
  assign n22044 = n22043 ^ n22042 ;
  assign n22046 = n22045 ^ n22044 ;
  assign n22047 = n21947 & n22046 ;
  assign n22032 = n21935 & n21939 ;
  assign n22031 = n21908 & ~n21936 ;
  assign n22033 = n22032 ^ n22031 ;
  assign n22052 = n22047 ^ n22033 ;
  assign n21950 = ~n20982 & n21089 ;
  assign n21949 = ~n20983 & n21080 ;
  assign n21951 = n21950 ^ n21949 ;
  assign n21958 = n21091 ^ n21077 ;
  assign n21959 = n21958 ^ n21957 ;
  assign n21960 = n20983 & n21959 ;
  assign n21961 = n21960 ^ n21077 ;
  assign n21978 = n21961 ^ n21106 ;
  assign n21979 = n21978 ^ n21123 ;
  assign n21971 = n21083 ^ n21071 ;
  assign n21969 = n21087 ^ n21082 ;
  assign n21970 = n21969 ^ n21078 ;
  assign n21972 = n21971 ^ n21970 ;
  assign n21973 = n21970 ^ n20983 ;
  assign n21974 = n21973 ^ n21970 ;
  assign n21975 = n21972 & ~n21974 ;
  assign n21976 = n21975 ^ n21970 ;
  assign n21977 = n21136 & n21976 ;
  assign n21980 = n21979 ^ n21977 ;
  assign n21964 = n21961 ^ n21089 ;
  assign n21965 = n21964 ^ n21961 ;
  assign n21966 = n20983 & n21965 ;
  assign n21967 = n21966 ^ n21961 ;
  assign n21968 = n20982 & n21967 ;
  assign n21981 = n21980 ^ n21968 ;
  assign n21982 = ~n21956 & ~n21981 ;
  assign n21952 = n21072 & ~n21114 ;
  assign n21983 = n21982 ^ n21952 ;
  assign n21984 = ~n21951 & n21983 ;
  assign n21991 = n21984 & ~n21990 ;
  assign n21992 = ~n21948 & n21991 ;
  assign n21994 = n20984 & n21095 ;
  assign n21995 = n21992 & n21994 ;
  assign n21993 = n21992 ^ n18640 ;
  assign n21996 = n21995 ^ n21993 ;
  assign n21997 = n21996 ^ x108 ;
  assign n22048 = n21935 & ~n21940 ;
  assign n22003 = n21939 & n22002 ;
  assign n22018 = n22017 ^ n22003 ;
  assign n22020 = n22019 ^ n22018 ;
  assign n22021 = n22020 ^ n22002 ;
  assign n22022 = n22021 ^ n21944 ;
  assign n22049 = n22048 ^ n22022 ;
  assign n22050 = n22049 ^ n22047 ;
  assign n22051 = n21997 & n22050 ;
  assign n22053 = n22052 ^ n22051 ;
  assign n21998 = n21947 & ~n21997 ;
  assign n22013 = n21998 ^ n21997 ;
  assign n22014 = n22013 ^ n21947 ;
  assign n22015 = n22014 ^ n21998 ;
  assign n22039 = n21941 & n21997 ;
  assign n22038 = n22033 ^ n21941 ;
  assign n22040 = n22039 ^ n22038 ;
  assign n22041 = ~n22015 & n22040 ;
  assign n22054 = n22053 ^ n22041 ;
  assign n22001 = n21935 & n21943 ;
  assign n22034 = n22033 ^ n22001 ;
  assign n22036 = n22035 ^ n22034 ;
  assign n22037 = ~n22013 & n22036 ;
  assign n22055 = n22054 ^ n22037 ;
  assign n22056 = n22055 ^ n22003 ;
  assign n22029 = n22017 ^ n21941 ;
  assign n22030 = n22014 & n22029 ;
  assign n22057 = n22056 ^ n22030 ;
  assign n22016 = ~n21936 & n21939 ;
  assign n22023 = n22022 ^ n22016 ;
  assign n22024 = n22022 ^ n21997 ;
  assign n22025 = n22024 ^ n22022 ;
  assign n22026 = n22023 & n22025 ;
  assign n22027 = n22026 ^ n22022 ;
  assign n22028 = ~n22015 & n22027 ;
  assign n22058 = n22057 ^ n22028 ;
  assign n22005 = ~n21936 & ~n21940 ;
  assign n22004 = n22003 ^ n22001 ;
  assign n22006 = n22005 ^ n22004 ;
  assign n22007 = n22006 ^ n22003 ;
  assign n22008 = n22003 ^ n21997 ;
  assign n22009 = n22008 ^ n22003 ;
  assign n22010 = n22007 & n22009 ;
  assign n22011 = n22010 ^ n22003 ;
  assign n22012 = n21947 & n22011 ;
  assign n22059 = n22058 ^ n22012 ;
  assign n21999 = n21998 ^ n21947 ;
  assign n22000 = n21946 & n21999 ;
  assign n22060 = n22059 ^ n22000 ;
  assign n22063 = n21997 ^ n21941 ;
  assign n22064 = n22063 ^ n21941 ;
  assign n22065 = n21942 & n22064 ;
  assign n22066 = n22065 ^ n21941 ;
  assign n22067 = n21947 & n22066 ;
  assign n22068 = ~n22060 & ~n22067 ;
  assign n22069 = n22068 ^ n21013 ;
  assign n22070 = n22069 ^ x125 ;
  assign n22300 = n21672 ^ x89 ;
  assign n22122 = n17802 & n19073 ;
  assign n22123 = n22122 ^ n19081 ;
  assign n22124 = n22123 ^ n19092 ;
  assign n22125 = n19309 & n22124 ;
  assign n22112 = n19065 ^ n17802 ;
  assign n22114 = n19071 ^ n19059 ;
  assign n22115 = ~n19283 & n22114 ;
  assign n22113 = n19078 ^ n19065 ;
  assign n22116 = n22115 ^ n22113 ;
  assign n22117 = ~n22112 & ~n22116 ;
  assign n22118 = n22117 ^ n17802 ;
  assign n22119 = n22118 ^ n19092 ;
  assign n22108 = n22107 ^ n19299 ;
  assign n22109 = n19301 & n22108 ;
  assign n22110 = n22109 ^ n19299 ;
  assign n22111 = n19283 & n22110 ;
  assign n22120 = n22119 ^ n22111 ;
  assign n22126 = n22125 ^ n22120 ;
  assign n22127 = n19082 ^ n19081 ;
  assign n22128 = n19082 ^ n17802 ;
  assign n22129 = n22128 ^ n19082 ;
  assign n22130 = n22127 & n22129 ;
  assign n22131 = n22130 ^ n19082 ;
  assign n22132 = n19283 & n22131 ;
  assign n22133 = n22126 & ~n22132 ;
  assign n22141 = n22133 & ~n22140 ;
  assign n22142 = ~n22106 & n22141 ;
  assign n22143 = ~n19333 & n22142 ;
  assign n22144 = n22143 ^ n17031 ;
  assign n22301 = n22144 ^ x96 ;
  assign n22448 = ~n22300 & ~n22301 ;
  assign n22449 = n22448 ^ n22300 ;
  assign n22450 = n22449 ^ n22301 ;
  assign n22093 = n19868 & n19910 ;
  assign n22089 = n19902 ^ n19899 ;
  assign n22090 = n19909 & n22089 ;
  assign n22083 = n19867 ^ n19546 ;
  assign n22084 = n22083 ^ n19899 ;
  assign n22085 = ~n19368 & ~n22084 ;
  assign n22079 = n19925 ^ n19913 ;
  assign n22073 = n19926 ^ n19871 ;
  assign n22074 = n22073 ^ n19925 ;
  assign n22075 = n22073 ^ n19368 ;
  assign n22076 = ~n19547 & ~n22075 ;
  assign n22077 = n22076 ^ n19368 ;
  assign n22078 = ~n22074 & ~n22077 ;
  assign n22080 = n22079 ^ n22078 ;
  assign n22081 = n22080 ^ n19923 ;
  assign n22072 = n19922 ^ n19871 ;
  assign n22082 = n22081 ^ n22072 ;
  assign n22086 = n22085 ^ n22082 ;
  assign n22087 = ~n19912 & n22086 ;
  assign n22088 = n22087 ^ n22081 ;
  assign n22091 = n22090 ^ n22088 ;
  assign n22071 = n19876 & n19912 ;
  assign n22092 = n22091 ^ n22071 ;
  assign n22094 = n22093 ^ n22092 ;
  assign n22100 = n22094 ^ n16173 ;
  assign n22095 = ~n19546 & ~n22094 ;
  assign n22096 = n19874 ^ n19816 ;
  assign n22097 = n21405 & n22096 ;
  assign n22098 = n22097 ^ n19874 ;
  assign n22099 = n22095 & n22098 ;
  assign n22101 = n22100 ^ n22099 ;
  assign n22303 = n22101 ^ x99 ;
  assign n22304 = n21571 ^ x65 ;
  assign n22305 = n22303 & ~n22304 ;
  assign n22386 = n22305 ^ n22304 ;
  assign n22389 = n22386 ^ n22303 ;
  assign n22323 = n21089 ^ n21070 ;
  assign n22324 = ~n20985 & n22323 ;
  assign n22317 = n21074 ^ n21068 ;
  assign n22320 = n22317 ^ n21948 ;
  assign n22313 = n21096 ^ n21078 ;
  assign n22314 = n22313 ^ n21102 ;
  assign n22315 = n22314 ^ n21064 ;
  assign n22316 = ~n20983 & n22315 ;
  assign n22318 = n22317 ^ n22316 ;
  assign n22319 = n21136 & n22318 ;
  assign n22321 = n22320 ^ n22319 ;
  assign n22308 = n21093 ^ n20983 ;
  assign n22309 = n22308 ^ n21093 ;
  assign n22310 = n21094 & n22309 ;
  assign n22311 = n22310 ^ n21093 ;
  assign n22312 = ~n20982 & n22311 ;
  assign n22322 = n22321 ^ n22312 ;
  assign n22325 = n22324 ^ n22322 ;
  assign n22326 = n21072 ^ n21069 ;
  assign n22327 = n22326 ^ n21105 ;
  assign n22328 = n22327 ^ n21969 ;
  assign n22329 = n20983 & ~n22328 ;
  assign n22330 = n22329 ^ n21069 ;
  assign n22331 = ~n21136 & n22330 ;
  assign n22332 = ~n22325 & ~n22331 ;
  assign n22333 = ~n21129 & n22332 ;
  assign n22334 = n21955 ^ n21101 ;
  assign n22335 = n21101 ^ n20982 ;
  assign n22336 = n22335 ^ n21101 ;
  assign n22337 = n22334 & n22336 ;
  assign n22338 = n22337 ^ n21101 ;
  assign n22339 = n22333 & ~n22338 ;
  assign n22340 = n22339 ^ n18347 ;
  assign n22341 = n22340 ^ x74 ;
  assign n22349 = n20146 ^ n20059 ;
  assign n22350 = n22349 ^ n20210 ;
  assign n22351 = n22350 ^ n20241 ;
  assign n22352 = n19999 & ~n22351 ;
  assign n22347 = n20253 ^ n20220 ;
  assign n22348 = n22347 ^ n21182 ;
  assign n22353 = n22352 ^ n22348 ;
  assign n22354 = n22353 ^ n20226 ;
  assign n22355 = n22354 ^ n20255 ;
  assign n22356 = n22355 ^ n22353 ;
  assign n22359 = n19999 & n22356 ;
  assign n22360 = n22359 ^ n22353 ;
  assign n22361 = n20021 & n22360 ;
  assign n22362 = n22361 ^ n22353 ;
  assign n22344 = n20237 ^ n20219 ;
  assign n22345 = n22344 ^ n20222 ;
  assign n22346 = n20286 & ~n22345 ;
  assign n22363 = n22362 ^ n22346 ;
  assign n22364 = n22363 ^ n20214 ;
  assign n22365 = n22364 ^ n21175 ;
  assign n22366 = n22365 ^ n21553 ;
  assign n22367 = n22366 ^ n18382 ;
  assign n22343 = n20243 & n20300 ;
  assign n22368 = n22367 ^ n22343 ;
  assign n22371 = n22368 ^ n20250 ;
  assign n22369 = n22368 ^ n20214 ;
  assign n22342 = ~n19999 & n20248 ;
  assign n22370 = n22369 ^ n22342 ;
  assign n22372 = n22371 ^ n22370 ;
  assign n22373 = n22372 ^ n22347 ;
  assign n22374 = n22373 ^ n20250 ;
  assign n22375 = n22374 ^ n22372 ;
  assign n22378 = n20021 & ~n22375 ;
  assign n22379 = n22378 ^ n22372 ;
  assign n22380 = n20270 & ~n22379 ;
  assign n22381 = n22380 ^ n22370 ;
  assign n22382 = n22381 ^ x113 ;
  assign n22383 = n22341 & n22382 ;
  assign n22397 = n22383 ^ n22341 ;
  assign n22398 = n22397 ^ n22382 ;
  assign n22453 = n22389 & ~n22398 ;
  assign n22384 = n22383 ^ n22382 ;
  assign n22406 = n22389 ^ n22304 ;
  assign n22407 = n22384 & n22406 ;
  assign n22408 = n22407 ^ n22384 ;
  assign n22404 = n22384 & ~n22386 ;
  assign n22385 = n22305 & n22384 ;
  assign n22405 = n22404 ^ n22385 ;
  assign n22409 = n22408 ^ n22405 ;
  assign n22392 = n22383 ^ n22303 ;
  assign n22393 = n22304 & n22392 ;
  assign n22394 = n22393 ^ n22304 ;
  assign n22390 = n22383 & n22389 ;
  assign n22391 = n22390 ^ n22389 ;
  assign n22395 = n22394 ^ n22391 ;
  assign n22410 = n22409 ^ n22395 ;
  assign n22457 = n22453 ^ n22410 ;
  assign n22458 = n22457 ^ n22394 ;
  assign n22399 = n22305 & ~n22398 ;
  assign n22400 = n22399 ^ n22390 ;
  assign n22446 = n22400 ^ n22395 ;
  assign n22429 = n22382 ^ n22341 ;
  assign n22430 = n22304 ^ n22303 ;
  assign n22432 = n22382 & n22430 ;
  assign n22433 = n22432 ^ n22303 ;
  assign n22434 = ~n22429 & n22433 ;
  assign n22447 = n22446 ^ n22434 ;
  assign n22459 = n22458 ^ n22447 ;
  assign n22460 = ~n22450 & n22459 ;
  assign n22402 = ~n22386 & ~n22398 ;
  assign n22456 = n22402 & n22448 ;
  assign n22461 = n22460 ^ n22456 ;
  assign n22454 = n22453 ^ n22407 ;
  assign n22455 = ~n22449 & n22454 ;
  assign n22462 = n22461 ^ n22455 ;
  assign n22427 = n22382 ^ n22303 ;
  assign n22387 = n22383 & ~n22386 ;
  assign n22416 = n22387 ^ n22386 ;
  assign n22424 = n22416 ^ n22385 ;
  assign n22428 = n22427 ^ n22424 ;
  assign n22435 = n22434 ^ n22428 ;
  assign n22436 = n22301 & ~n22435 ;
  assign n22415 = n22404 ^ n22402 ;
  assign n22417 = n22416 ^ n22415 ;
  assign n22418 = n22417 ^ n22390 ;
  assign n22419 = n22418 ^ n22398 ;
  assign n22412 = n22383 ^ n22305 ;
  assign n22388 = n22387 ^ n22385 ;
  assign n22396 = n22395 ^ n22388 ;
  assign n22401 = n22400 ^ n22396 ;
  assign n22413 = n22412 ^ n22401 ;
  assign n22414 = n22413 ^ n22387 ;
  assign n22420 = n22419 ^ n22414 ;
  assign n22421 = ~n22300 & ~n22420 ;
  assign n22411 = n22410 ^ n22390 ;
  assign n22422 = n22421 ^ n22411 ;
  assign n22423 = ~n22301 & n22422 ;
  assign n22425 = n22424 ^ n22423 ;
  assign n22437 = n22436 ^ n22425 ;
  assign n22463 = n22462 ^ n22437 ;
  assign n22451 = n22450 ^ n22300 ;
  assign n22452 = n22447 & ~n22451 ;
  assign n22464 = n22463 ^ n22452 ;
  assign n22465 = n22464 ^ n20341 ;
  assign n22302 = n22301 ^ n22300 ;
  assign n22438 = n22437 ^ n22423 ;
  assign n22403 = n22402 ^ n22401 ;
  assign n22439 = n22438 ^ n22403 ;
  assign n22440 = n22439 ^ n22438 ;
  assign n22441 = n22438 ^ n22300 ;
  assign n22442 = n22441 ^ n22438 ;
  assign n22443 = n22440 & n22442 ;
  assign n22444 = n22443 ^ n22438 ;
  assign n22445 = ~n22302 & ~n22444 ;
  assign n22466 = n22465 ^ n22445 ;
  assign n22467 = n22466 ^ x68 ;
  assign n22614 = n22070 & ~n22467 ;
  assign n22615 = n22597 & n22614 ;
  assign n22664 = n22615 ^ n22614 ;
  assign n22598 = n22467 & n22597 ;
  assign n22632 = n22598 ^ n22467 ;
  assign n22103 = n21372 ^ x121 ;
  assign n22102 = n22101 ^ x112 ;
  assign n22104 = n22103 ^ n22102 ;
  assign n22105 = n21153 ^ x98 ;
  assign n22145 = n22144 ^ x107 ;
  assign n22146 = ~n22105 & ~n22145 ;
  assign n22161 = n20804 & ~n20824 ;
  assign n22158 = n20859 ^ n20820 ;
  assign n22159 = ~n20828 & ~n22158 ;
  assign n22155 = n20846 ^ n20827 ;
  assign n22156 = n22155 ^ n21931 ;
  assign n22157 = n22156 ^ n17454 ;
  assign n22160 = n22159 ^ n22157 ;
  assign n22162 = n22161 ^ n22160 ;
  assign n22154 = n20826 & n20850 ;
  assign n22163 = n22162 ^ n22154 ;
  assign n22149 = n20856 ^ n20825 ;
  assign n22150 = n22149 ^ n20856 ;
  assign n22151 = n20857 & ~n22150 ;
  assign n22152 = n22151 ^ n20856 ;
  assign n22153 = n20824 & ~n22152 ;
  assign n22164 = n22163 ^ n22153 ;
  assign n22165 = n22164 ^ x81 ;
  assign n22166 = n21662 ^ n21314 ;
  assign n22167 = n22166 ^ n21311 ;
  assign n22191 = n22167 ^ n21333 ;
  assign n22179 = n21200 & n21309 ;
  assign n22180 = n22179 ^ n21303 ;
  assign n22192 = n22191 ^ n22180 ;
  assign n22193 = n22192 ^ n21332 ;
  assign n22194 = n22193 ^ n21903 ;
  assign n22195 = n22194 ^ n17161 ;
  assign n22181 = n22180 ^ n21301 ;
  assign n22182 = n22181 ^ n21861 ;
  assign n22183 = n22182 ^ n21300 ;
  assign n22184 = n22183 ^ n21301 ;
  assign n22185 = n22184 ^ n22182 ;
  assign n22188 = ~n21200 & n22185 ;
  assign n22189 = n22188 ^ n22182 ;
  assign n22190 = ~n21201 & ~n22189 ;
  assign n22196 = n22195 ^ n22190 ;
  assign n22176 = n21303 ^ n21275 ;
  assign n22177 = n22176 ^ n21314 ;
  assign n22178 = n21296 & n22177 ;
  assign n22197 = n22196 ^ n22178 ;
  assign n22168 = n22167 ^ n21334 ;
  assign n22169 = n22168 ^ n21282 ;
  assign n22170 = n22169 ^ n22167 ;
  assign n22171 = n22167 ^ n21201 ;
  assign n22172 = n22171 ^ n22167 ;
  assign n22173 = ~n22170 & n22172 ;
  assign n22174 = n22173 ^ n22167 ;
  assign n22175 = n21319 & n22174 ;
  assign n22198 = n22197 ^ n22175 ;
  assign n22199 = n22198 ^ x88 ;
  assign n22200 = n22165 & ~n22199 ;
  assign n22201 = n22200 ^ n22165 ;
  assign n22202 = n22201 ^ n22199 ;
  assign n22203 = n22202 ^ n22165 ;
  assign n22204 = n22146 & ~n22203 ;
  assign n22220 = n22102 & n22204 ;
  assign n22206 = n22146 ^ n22145 ;
  assign n22209 = n22206 ^ n22105 ;
  assign n22213 = ~n22203 & ~n22209 ;
  assign n22212 = n22200 & ~n22209 ;
  assign n22214 = n22213 ^ n22212 ;
  assign n22210 = n22202 & ~n22209 ;
  assign n22211 = n22210 ^ n22209 ;
  assign n22215 = n22214 ^ n22211 ;
  assign n22207 = n22202 & ~n22206 ;
  assign n22205 = n22146 & n22201 ;
  assign n22208 = n22207 ^ n22205 ;
  assign n22216 = n22215 ^ n22208 ;
  assign n22217 = ~n22102 & ~n22216 ;
  assign n22218 = n22217 ^ n22215 ;
  assign n22219 = n22218 ^ n22204 ;
  assign n22221 = n22220 ^ n22219 ;
  assign n22222 = ~n22104 & ~n22221 ;
  assign n22223 = n22222 ^ n22218 ;
  assign n22234 = n22146 & n22200 ;
  assign n22235 = n22102 & ~n22103 ;
  assign n22236 = n22234 & n22235 ;
  assign n22224 = n22209 ^ n22145 ;
  assign n22225 = n22202 & ~n22224 ;
  assign n22226 = n22225 ^ n22207 ;
  assign n22229 = n22207 ^ n22102 ;
  assign n22230 = n22229 ^ n22207 ;
  assign n22231 = n22226 & ~n22230 ;
  assign n22232 = n22231 ^ n22207 ;
  assign n22233 = ~n22103 & n22232 ;
  assign n22237 = n22236 ^ n22233 ;
  assign n22269 = n22225 ^ n22204 ;
  assign n22270 = n22269 ^ n22203 ;
  assign n22241 = ~n22203 & ~n22224 ;
  assign n22242 = n22241 ^ n22212 ;
  assign n22243 = n22242 ^ n22225 ;
  assign n22244 = n22243 ^ n22214 ;
  assign n22271 = n22270 ^ n22244 ;
  assign n22238 = n22201 & ~n22224 ;
  assign n22278 = n22271 ^ n22238 ;
  assign n22276 = n22225 ^ n22212 ;
  assign n22246 = n22201 & ~n22206 ;
  assign n22277 = n22276 ^ n22246 ;
  assign n22279 = n22278 ^ n22277 ;
  assign n22280 = n22102 & ~n22279 ;
  assign n22281 = n22280 ^ n22246 ;
  assign n22282 = n22104 & n22281 ;
  assign n22272 = n22271 ^ n22234 ;
  assign n22273 = ~n22104 & ~n22272 ;
  assign n22283 = n22282 ^ n22273 ;
  assign n22268 = n22242 ^ n22215 ;
  assign n22274 = ~n22102 & ~n22273 ;
  assign n22275 = ~n22268 & n22274 ;
  assign n22284 = n22283 ^ n22275 ;
  assign n22253 = n22226 ^ n22202 ;
  assign n22254 = n22253 ^ n22210 ;
  assign n22285 = n22284 ^ n22254 ;
  assign n22256 = ~n22102 & ~n22103 ;
  assign n22257 = n22256 ^ n22102 ;
  assign n22255 = n22254 ^ n22103 ;
  assign n22258 = n22257 ^ n22255 ;
  assign n22260 = n22225 ^ n22213 ;
  assign n22259 = n22200 & ~n22206 ;
  assign n22261 = n22260 ^ n22259 ;
  assign n22262 = n22261 ^ n22257 ;
  assign n22263 = n22257 ^ n22254 ;
  assign n22264 = n22263 ^ n22257 ;
  assign n22265 = n22262 & ~n22264 ;
  assign n22266 = n22265 ^ n22257 ;
  assign n22267 = ~n22258 & n22266 ;
  assign n22286 = n22285 ^ n22267 ;
  assign n22239 = n22238 ^ n22213 ;
  assign n22240 = n22239 ^ n22224 ;
  assign n22245 = n22244 ^ n22240 ;
  assign n22247 = n22246 ^ n22245 ;
  assign n22248 = n22246 ^ n22103 ;
  assign n22249 = n22248 ^ n22246 ;
  assign n22250 = ~n22247 & n22249 ;
  assign n22251 = n22250 ^ n22246 ;
  assign n22252 = ~n22102 & n22251 ;
  assign n22287 = n22286 ^ n22252 ;
  assign n22288 = n22245 ^ n22210 ;
  assign n22289 = n22288 ^ n22204 ;
  assign n22290 = n22204 ^ n22103 ;
  assign n22291 = n22290 ^ n22204 ;
  assign n22292 = ~n22289 & n22291 ;
  assign n22293 = n22292 ^ n22204 ;
  assign n22294 = n22102 & n22293 ;
  assign n22295 = ~n22287 & ~n22294 ;
  assign n22296 = ~n22237 & n22295 ;
  assign n22297 = n22223 & n22296 ;
  assign n22298 = n22297 ^ n21058 ;
  assign n22299 = n22298 ^ x110 ;
  assign n22603 = n22299 & ~n22597 ;
  assign n22604 = n22467 & n22603 ;
  assign n22633 = n22632 ^ n22604 ;
  assign n22631 = n22603 ^ n22597 ;
  assign n22634 = n22633 ^ n22631 ;
  assign n22642 = n22634 ^ n22467 ;
  assign n22619 = n22299 & n22615 ;
  assign n22620 = n22619 ^ n22615 ;
  assign n22617 = n22614 ^ n22467 ;
  assign n22618 = n22603 & ~n22617 ;
  assign n22621 = n22620 ^ n22618 ;
  assign n22622 = n22621 ^ n22619 ;
  assign n22613 = n22598 ^ n22597 ;
  assign n22616 = n22615 ^ n22613 ;
  assign n22623 = n22622 ^ n22616 ;
  assign n22643 = n22642 ^ n22623 ;
  assign n22665 = n22664 ^ n22643 ;
  assign n22666 = n22665 ^ n22620 ;
  assign n22667 = n22666 ^ n22643 ;
  assign n22660 = n22299 ^ n22070 ;
  assign n22661 = n22660 ^ n22597 ;
  assign n22662 = ~n22467 & n22661 ;
  assign n22663 = n22662 ^ n22642 ;
  assign n22668 = n22667 ^ n22663 ;
  assign n22705 = ~n22650 & n22668 ;
  assign n22599 = n22299 & n22598 ;
  assign n22600 = n22599 ^ n22598 ;
  assign n22601 = ~n22070 & n22600 ;
  assign n22602 = n22601 ^ n22600 ;
  assign n22651 = n22650 ^ n21536 ;
  assign n22704 = n22602 & ~n22651 ;
  assign n22706 = n22705 ^ n22704 ;
  assign n22637 = n22070 & n22599 ;
  assign n22692 = n22643 ^ n22637 ;
  assign n22693 = n22643 ^ n21823 ;
  assign n22694 = n22693 ^ n22643 ;
  assign n22695 = n22692 & ~n22694 ;
  assign n22696 = n22695 ^ n22643 ;
  assign n22697 = ~n21536 & n22696 ;
  assign n22638 = n22637 ^ n22599 ;
  assign n22605 = ~n22070 & n22604 ;
  assign n22639 = n22638 ^ n22605 ;
  assign n22640 = n22639 ^ n22601 ;
  assign n22636 = n22617 ^ n22070 ;
  assign n22641 = n22640 ^ n22636 ;
  assign n22655 = n22641 ^ n22633 ;
  assign n22679 = n22655 ^ n22637 ;
  assign n22676 = n22665 ^ n22634 ;
  assign n22677 = n22676 ^ n22620 ;
  assign n21824 = n21823 ^ n21536 ;
  assign n22669 = n22668 ^ n22616 ;
  assign n22659 = n22641 ^ n22601 ;
  assign n22670 = n22669 ^ n22659 ;
  assign n22671 = n22659 ^ n21536 ;
  assign n22672 = n22671 ^ n22659 ;
  assign n22673 = n22670 & ~n22672 ;
  assign n22674 = n22673 ^ n22659 ;
  assign n22675 = n21824 & n22674 ;
  assign n22678 = n22677 ^ n22675 ;
  assign n22680 = n22679 ^ n22678 ;
  assign n22681 = n22680 ^ n22675 ;
  assign n22682 = n21536 & ~n22681 ;
  assign n22683 = n22682 ^ n22678 ;
  assign n22698 = n22697 ^ n22683 ;
  assign n22684 = n22683 ^ n22675 ;
  assign n22653 = n22605 ^ n22604 ;
  assign n22685 = n22684 ^ n22653 ;
  assign n22686 = n22685 ^ n22684 ;
  assign n22687 = n22684 ^ n21823 ;
  assign n22688 = n22687 ^ n22684 ;
  assign n22689 = n22686 & ~n22688 ;
  assign n22690 = n22689 ^ n22684 ;
  assign n22691 = ~n21824 & ~n22690 ;
  assign n22699 = n22698 ^ n22691 ;
  assign n22652 = n22651 ^ n21823 ;
  assign n22656 = n22655 ^ n22602 ;
  assign n22654 = n22653 ^ n22638 ;
  assign n22657 = n22656 ^ n22654 ;
  assign n22658 = ~n22652 & n22657 ;
  assign n22700 = n22699 ^ n22658 ;
  assign n22644 = n22643 ^ n22641 ;
  assign n22630 = n22619 ^ n22605 ;
  assign n22635 = n22634 ^ n22630 ;
  assign n22645 = n22644 ^ n22635 ;
  assign n22646 = n21536 & ~n22645 ;
  assign n22647 = n22646 ^ n22644 ;
  assign n22648 = ~n21824 & n22647 ;
  assign n22701 = n22700 ^ n22648 ;
  assign n22702 = n22701 ^ n22616 ;
  assign n22625 = n22616 ^ n21536 ;
  assign n22626 = n22625 ^ n22616 ;
  assign n22627 = n22622 & n22626 ;
  assign n22628 = n22627 ^ n22616 ;
  assign n22629 = n21824 & n22628 ;
  assign n22703 = n22702 ^ n22629 ;
  assign n22707 = n22706 ^ n22703 ;
  assign n22606 = n22605 ^ n22602 ;
  assign n22607 = n22606 ^ n22601 ;
  assign n22608 = n22601 ^ n21536 ;
  assign n22609 = n22608 ^ n22601 ;
  assign n22610 = n22607 & ~n22609 ;
  assign n22611 = n22610 ^ n22601 ;
  assign n22612 = ~n21824 & n22611 ;
  assign n22708 = n22707 ^ n22612 ;
  assign n22709 = n22708 ^ n21153 ;
  assign n22998 = n20981 ^ x74 ;
  assign n22956 = n22458 ^ n22404 ;
  assign n22957 = ~n22449 & n22956 ;
  assign n22953 = ~n22451 & n22457 ;
  assign n22950 = ~n22407 & n22450 ;
  assign n22951 = n22393 & ~n22950 ;
  assign n22944 = n22414 ^ n22399 ;
  assign n22945 = n22944 ^ n22402 ;
  assign n22946 = ~n22449 & n22945 ;
  assign n22942 = n22413 & ~n22451 ;
  assign n22943 = n22942 ^ n22456 ;
  assign n22947 = n22946 ^ n22943 ;
  assign n22937 = n22417 ^ n22301 ;
  assign n22938 = n22937 ^ n22417 ;
  assign n22939 = ~n22418 & n22938 ;
  assign n22940 = n22939 ^ n22417 ;
  assign n22941 = n22302 & ~n22940 ;
  assign n22948 = n22947 ^ n22941 ;
  assign n22949 = n22948 ^ n20020 ;
  assign n22952 = n22951 ^ n22949 ;
  assign n22954 = n22953 ^ n22952 ;
  assign n22927 = n22447 ^ n22410 ;
  assign n22929 = n22927 ^ n22413 ;
  assign n22916 = n22405 ^ n22402 ;
  assign n22930 = n22929 ^ n22916 ;
  assign n22931 = n22930 ^ n22427 ;
  assign n22932 = n22931 ^ n22403 ;
  assign n22928 = n22927 ^ n22417 ;
  assign n22933 = n22932 ^ n22928 ;
  assign n22934 = n22448 & ~n22933 ;
  assign n22955 = n22954 ^ n22934 ;
  assign n22958 = n22957 ^ n22955 ;
  assign n22926 = n22388 & ~n22451 ;
  assign n22959 = n22958 ^ n22926 ;
  assign n22917 = n22416 ^ n22392 ;
  assign n22918 = n22917 ^ n22394 ;
  assign n22919 = n22918 ^ n22916 ;
  assign n22920 = n22919 ^ n22918 ;
  assign n22921 = n22918 ^ n22300 ;
  assign n22922 = n22921 ^ n22918 ;
  assign n22923 = n22920 & n22922 ;
  assign n22924 = n22923 ^ n22918 ;
  assign n22925 = ~n22302 & n22924 ;
  assign n22960 = n22959 ^ n22925 ;
  assign n22961 = n22960 ^ x106 ;
  assign n22535 = n22534 ^ n22529 ;
  assign n22967 = n22549 ^ n22529 ;
  assign n22968 = ~n22535 & n22967 ;
  assign n22969 = n22968 ^ n22529 ;
  assign n22970 = n22530 & ~n22969 ;
  assign n22971 = n22970 ^ n22549 ;
  assign n22973 = ~n22563 & n22971 ;
  assign n22972 = n22971 ^ n22563 ;
  assign n22974 = n22973 ^ n22972 ;
  assign n22975 = n22974 ^ n22541 ;
  assign n22983 = n22975 ^ n20753 ;
  assign n22962 = n22543 ^ n22541 ;
  assign n22963 = n22962 ^ n22587 ;
  assign n22966 = n22963 ^ n22585 ;
  assign n22976 = n22975 ^ n22966 ;
  assign n22965 = n22572 ^ n22541 ;
  assign n22977 = n22976 ^ n22965 ;
  assign n22980 = ~n22563 & n22977 ;
  assign n22981 = n22980 ^ n22976 ;
  assign n22982 = n22551 & ~n22981 ;
  assign n22984 = n22983 ^ n22982 ;
  assign n22964 = ~n22563 & ~n22963 ;
  assign n22985 = n22984 ^ n22964 ;
  assign n22986 = n22985 ^ x97 ;
  assign n22987 = n22961 & n22986 ;
  assign n23008 = n22987 ^ n22961 ;
  assign n23009 = n23008 ^ n22986 ;
  assign n22760 = n19302 ^ n19067 ;
  assign n22761 = n22760 ^ n19324 ;
  assign n22762 = n19283 & n22761 ;
  assign n22763 = n22762 ^ n19087 ;
  assign n22764 = n17802 & ~n22763 ;
  assign n22765 = n22764 ^ n19087 ;
  assign n22756 = n22501 ^ n19081 ;
  assign n22757 = ~n19283 & ~n22756 ;
  assign n22758 = n22757 ^ n19081 ;
  assign n22759 = n19309 & n22758 ;
  assign n22766 = n22765 ^ n22759 ;
  assign n22767 = n22766 ^ n19073 ;
  assign n22747 = n22502 ^ n19071 ;
  assign n22746 = n22502 ^ n19302 ;
  assign n22748 = n22747 ^ n22746 ;
  assign n22749 = n22746 ^ n19283 ;
  assign n22750 = n22749 ^ n22746 ;
  assign n22751 = n22748 & ~n22750 ;
  assign n22752 = n22751 ^ n22746 ;
  assign n22753 = n19309 & n22752 ;
  assign n22754 = n22753 ^ n19073 ;
  assign n22755 = ~n19319 & n22754 ;
  assign n22768 = n22767 ^ n22755 ;
  assign n22769 = ~n22132 & n22768 ;
  assign n22770 = n22769 ^ n22106 ;
  assign n22771 = ~n19333 & n22770 ;
  assign n22774 = n22771 ^ n18723 ;
  assign n22772 = n17802 & n19285 ;
  assign n22773 = n22771 & n22772 ;
  assign n22775 = n22774 ^ n22773 ;
  assign n22776 = n22775 ^ x75 ;
  assign n22777 = n21996 ^ x100 ;
  assign n22778 = n22776 & n22777 ;
  assign n22779 = n22778 ^ n22776 ;
  assign n22780 = n21562 ^ x94 ;
  assign n22782 = n20542 ^ n20515 ;
  assign n22783 = n22782 ^ n18653 ;
  assign n22784 = n22783 ^ x117 ;
  assign n22785 = n22780 & ~n22784 ;
  assign n22791 = n22785 ^ n22780 ;
  assign n22792 = n22791 ^ n22784 ;
  assign n22806 = n22779 & n22792 ;
  assign n22807 = n22806 ^ n22779 ;
  assign n22829 = n22807 ^ n22791 ;
  assign n22819 = n22784 ^ n22776 ;
  assign n22812 = n22780 ^ n22776 ;
  assign n22820 = ~n22776 & ~n22812 ;
  assign n22821 = n22820 ^ n22778 ;
  assign n22822 = n22819 & ~n22821 ;
  assign n22830 = n22829 ^ n22822 ;
  assign n22795 = n22779 ^ n22777 ;
  assign n22796 = n22795 ^ n22776 ;
  assign n22798 = n22785 ^ n22784 ;
  assign n22799 = n22796 & ~n22798 ;
  assign n22866 = n22830 ^ n22799 ;
  assign n22788 = n21933 ^ x77 ;
  assign n22745 = n21600 ^ x68 ;
  assign n22793 = n22792 ^ n22785 ;
  assign n22818 = n22793 ^ n22777 ;
  assign n22823 = n22822 ^ n22818 ;
  assign n22816 = n22778 & n22785 ;
  assign n22800 = n22799 ^ n22796 ;
  assign n22797 = n22780 & n22796 ;
  assign n22801 = n22800 ^ n22797 ;
  assign n22817 = n22816 ^ n22801 ;
  assign n22824 = n22823 ^ n22817 ;
  assign n22814 = n22792 & ~n22795 ;
  assign n22813 = n22812 ^ n22777 ;
  assign n22815 = n22814 ^ n22813 ;
  assign n22825 = n22824 ^ n22815 ;
  assign n22786 = n22779 & n22785 ;
  assign n22781 = n22779 & n22780 ;
  assign n22787 = n22786 ^ n22781 ;
  assign n22828 = n22825 ^ n22787 ;
  assign n22831 = n22830 ^ n22828 ;
  assign n22810 = n22785 & n22796 ;
  assign n22811 = n22810 ^ n22797 ;
  assign n22826 = n22825 ^ n22811 ;
  assign n22827 = n22826 ^ n22791 ;
  assign n22832 = n22831 ^ n22827 ;
  assign n22809 = ~n22795 & ~n22798 ;
  assign n22833 = n22832 ^ n22809 ;
  assign n22808 = n22807 ^ n22781 ;
  assign n22834 = n22833 ^ n22808 ;
  assign n22789 = n22745 & n22788 ;
  assign n22790 = n22789 ^ n22788 ;
  assign n22794 = n22777 & n22793 ;
  assign n22802 = n22794 & ~n22801 ;
  assign n22803 = ~n22790 & n22802 ;
  assign n22804 = n22803 ^ n22794 ;
  assign n22805 = n22804 ^ n22787 ;
  assign n22835 = n22834 ^ n22805 ;
  assign n22836 = n22835 ^ n22804 ;
  assign n22837 = n22804 ^ n22788 ;
  assign n22838 = n22837 ^ n22804 ;
  assign n22839 = n22836 & ~n22838 ;
  assign n22840 = n22839 ^ n22804 ;
  assign n22841 = n22745 & n22840 ;
  assign n22842 = n22841 ^ n22804 ;
  assign n22846 = n22814 ^ n22786 ;
  assign n22844 = n22816 ^ n22806 ;
  assign n22843 = n22811 ^ n22808 ;
  assign n22845 = n22844 ^ n22843 ;
  assign n22847 = n22846 ^ n22845 ;
  assign n22848 = ~n22788 & n22847 ;
  assign n22849 = n22848 ^ n22808 ;
  assign n22850 = n22849 ^ n22823 ;
  assign n22851 = n22850 ^ n22824 ;
  assign n22852 = n22851 ^ n22850 ;
  assign n22855 = ~n22788 & n22852 ;
  assign n22856 = n22855 ^ n22850 ;
  assign n22857 = n22745 & n22856 ;
  assign n22858 = n22857 ^ n22849 ;
  assign n22859 = ~n22842 & ~n22858 ;
  assign n22867 = ~n22788 & n22859 ;
  assign n22868 = n22866 & n22867 ;
  assign n22862 = n22814 ^ n22787 ;
  assign n22863 = n22790 & n22862 ;
  assign n22861 = n22790 & n22809 ;
  assign n22864 = n22863 ^ n22861 ;
  assign n22860 = n22859 ^ n20358 ;
  assign n22865 = n22864 ^ n22860 ;
  assign n22869 = n22868 ^ n22865 ;
  assign n22870 = n22869 ^ x115 ;
  assign n22908 = n22032 ^ n22005 ;
  assign n22909 = n21998 & n22908 ;
  assign n22907 = ~n22013 & n22048 ;
  assign n22910 = n22909 ^ n22907 ;
  assign n22871 = ~n22013 & n22016 ;
  assign n22872 = n22871 ^ n22030 ;
  assign n22900 = n22045 ^ n22022 ;
  assign n22901 = n22900 ^ n22033 ;
  assign n22902 = ~n22013 & n22901 ;
  assign n22890 = n22048 ^ n22005 ;
  assign n22888 = n21908 & n21909 ;
  assign n22889 = n22888 ^ n22042 ;
  assign n22891 = n22890 ^ n22889 ;
  assign n22892 = n22891 ^ n21998 ;
  assign n22893 = n22014 & ~n22892 ;
  assign n22894 = n22893 ^ n21998 ;
  assign n22879 = n22019 ^ n21944 ;
  assign n22880 = ~n21998 & ~n22879 ;
  assign n22881 = n22880 ^ n22017 ;
  assign n22882 = n21947 & ~n22881 ;
  assign n22896 = n22882 ^ n22014 ;
  assign n22895 = n22882 ^ n22035 ;
  assign n22897 = n22896 ^ n22895 ;
  assign n22898 = n22894 & n22897 ;
  assign n22899 = n22898 ^ n22896 ;
  assign n22903 = n22902 ^ n22899 ;
  assign n22875 = n22003 ^ n21938 ;
  assign n22876 = n22875 ^ n22001 ;
  assign n22877 = n22876 ^ n22045 ;
  assign n22878 = n22877 ^ n22001 ;
  assign n22885 = ~n22878 & n22882 ;
  assign n22886 = n22885 ^ n22001 ;
  assign n22887 = n21998 & n22886 ;
  assign n22904 = n22903 ^ n22887 ;
  assign n22873 = n22034 ^ n22005 ;
  assign n22874 = n21999 & n22873 ;
  assign n22905 = n22904 ^ n22874 ;
  assign n22906 = ~n22872 & ~n22905 ;
  assign n22911 = n22910 ^ n22906 ;
  assign n22912 = n22911 ^ n22000 ;
  assign n22913 = n22912 ^ n20786 ;
  assign n22914 = n22913 ^ x96 ;
  assign n22915 = n22870 & n22914 ;
  assign n22991 = n22915 ^ n22914 ;
  assign n23013 = n22991 ^ n22870 ;
  assign n23014 = ~n23009 & ~n23013 ;
  assign n23072 = n22998 & n23014 ;
  assign n23039 = n22987 & ~n23013 ;
  assign n23038 = n22915 & n22987 ;
  assign n23040 = n23039 ^ n23038 ;
  assign n23036 = n22987 & n22991 ;
  assign n23037 = n23036 ^ n22987 ;
  assign n23041 = n23040 ^ n23037 ;
  assign n22738 = n22256 & n22259 ;
  assign n22711 = n22271 ^ n22254 ;
  assign n22735 = n22256 & ~n22711 ;
  assign n22726 = n22205 ^ n22204 ;
  assign n22727 = n22726 ^ n22210 ;
  assign n22728 = n22210 ^ n22102 ;
  assign n22729 = n22728 ^ n22210 ;
  assign n22730 = n22727 & n22729 ;
  assign n22731 = n22730 ^ n22210 ;
  assign n22732 = n22104 & n22731 ;
  assign n22733 = n22732 ^ n22220 ;
  assign n22721 = n22242 ^ n22234 ;
  assign n22722 = n22721 ^ n22278 ;
  assign n22723 = ~n22102 & ~n22722 ;
  assign n22734 = n22733 ^ n22723 ;
  assign n22736 = n22735 ^ n22734 ;
  assign n22737 = n22736 ^ n22237 ;
  assign n22739 = n22738 ^ n22737 ;
  assign n22720 = n22288 ^ n22215 ;
  assign n22724 = n22723 ^ n22720 ;
  assign n22725 = ~n22104 & n22724 ;
  assign n22740 = n22739 ^ n22725 ;
  assign n22712 = n22711 ^ n22241 ;
  assign n22713 = n22712 ^ n22246 ;
  assign n22710 = n22261 ^ n22245 ;
  assign n22714 = n22713 ^ n22710 ;
  assign n22715 = n22710 ^ n22103 ;
  assign n22716 = n22715 ^ n22710 ;
  assign n22717 = n22714 & n22716 ;
  assign n22718 = n22717 ^ n22710 ;
  assign n22719 = n22102 & ~n22718 ;
  assign n22741 = n22740 ^ n22719 ;
  assign n22742 = n22223 & ~n22741 ;
  assign n22743 = n22742 ^ n20437 ;
  assign n22744 = n22743 ^ x64 ;
  assign n23004 = n22998 ^ n22744 ;
  assign n23005 = ~n22998 & n23004 ;
  assign n23068 = n23041 ^ n23005 ;
  assign n22993 = n22915 ^ n22870 ;
  assign n23020 = n22993 & n23008 ;
  assign n23006 = n23005 ^ n22744 ;
  assign n23007 = n23006 ^ n22998 ;
  assign n23069 = n23020 ^ n23007 ;
  assign n23070 = n23068 & n23069 ;
  assign n23019 = n22991 & n23008 ;
  assign n23061 = n23006 & n23019 ;
  assign n23027 = n23008 & ~n23013 ;
  assign n23028 = n23027 ^ n23008 ;
  assign n23021 = n23020 ^ n23019 ;
  assign n23029 = n23028 ^ n23021 ;
  assign n23059 = n23036 ^ n23029 ;
  assign n23060 = n23005 & n23059 ;
  assign n23062 = n23061 ^ n23060 ;
  assign n23012 = n22991 & ~n23009 ;
  assign n23015 = n23014 ^ n23012 ;
  assign n23010 = n22915 & ~n23009 ;
  assign n23011 = n23010 ^ n23009 ;
  assign n23016 = n23015 ^ n23011 ;
  assign n23056 = n23005 & ~n23016 ;
  assign n23055 = n23004 & n23012 ;
  assign n23057 = n23056 ^ n23055 ;
  assign n22988 = n22987 ^ n22986 ;
  assign n22994 = n22988 & n22993 ;
  assign n22992 = n22988 & n22991 ;
  assign n22995 = n22994 ^ n22992 ;
  assign n22989 = n22915 & n22988 ;
  assign n22990 = n22989 ^ n22988 ;
  assign n22996 = n22995 ^ n22990 ;
  assign n22997 = n22996 ^ n22992 ;
  assign n23022 = n23005 ^ n22998 ;
  assign n23052 = n22997 & ~n23022 ;
  assign n23042 = n23041 ^ n23027 ;
  assign n23043 = n23042 ^ n23040 ;
  assign n23046 = n23043 ^ n22744 ;
  assign n23047 = n23046 ^ n23043 ;
  assign n23048 = n23039 & n23047 ;
  assign n23049 = n23048 ^ n23043 ;
  assign n23050 = ~n23004 & n23049 ;
  assign n23051 = n23050 ^ n23040 ;
  assign n23053 = n23052 ^ n23051 ;
  assign n23024 = n23010 ^ n22989 ;
  assign n23054 = n23053 ^ n23024 ;
  assign n23058 = n23057 ^ n23054 ;
  assign n23063 = n23062 ^ n23058 ;
  assign n23025 = n23024 ^ n22744 ;
  assign n23026 = n23025 ^ n23024 ;
  assign n23030 = n23029 ^ n22994 ;
  assign n23033 = ~n23026 & n23030 ;
  assign n23034 = n23033 ^ n23024 ;
  assign n23035 = n23004 & n23034 ;
  assign n23064 = n23063 ^ n23035 ;
  assign n23023 = n23021 & ~n23022 ;
  assign n23065 = n23064 ^ n23023 ;
  assign n23017 = n23007 & ~n23016 ;
  assign n23001 = n22997 & ~n22998 ;
  assign n23002 = n23001 ^ n22992 ;
  assign n23003 = n22744 & n23002 ;
  assign n23018 = n23017 ^ n23003 ;
  assign n23066 = n23065 ^ n23018 ;
  assign n23067 = n23066 ^ n20893 ;
  assign n23071 = n23070 ^ n23067 ;
  assign n23073 = n23072 ^ n23071 ;
  assign n23092 = n21473 ^ n21470 ;
  assign n23093 = n23092 ^ n21514 ;
  assign n23094 = n21197 & ~n23093 ;
  assign n23089 = ~n21472 & ~n21494 ;
  assign n23082 = n21465 ^ n21373 ;
  assign n23083 = n23082 ^ n21468 ;
  assign n23084 = n23083 ^ n21470 ;
  assign n23085 = ~n21154 & n23084 ;
  assign n23086 = n23085 ^ n21499 ;
  assign n23087 = ~n21196 & n23086 ;
  assign n23079 = n21197 & n21500 ;
  assign n23078 = n21199 & n21492 ;
  assign n23080 = n23079 ^ n23078 ;
  assign n23077 = n21469 ^ n19856 ;
  assign n23081 = n23080 ^ n23077 ;
  assign n23088 = n23087 ^ n23081 ;
  assign n23090 = n23089 ^ n23088 ;
  assign n23075 = n21500 ^ n21476 ;
  assign n23076 = n21198 & n23075 ;
  assign n23091 = n23090 ^ n23076 ;
  assign n23095 = n23094 ^ n23091 ;
  assign n23074 = n21461 & n21472 ;
  assign n23096 = n23095 ^ n23074 ;
  assign n23125 = ~n23016 & ~n23022 ;
  assign n23123 = n23039 ^ n23020 ;
  assign n23124 = n23006 & n23123 ;
  assign n23126 = n23125 ^ n23124 ;
  assign n23127 = n23126 ^ n23057 ;
  assign n23122 = n23007 & n23059 ;
  assign n23128 = n23127 ^ n23122 ;
  assign n23129 = n23128 ^ n23042 ;
  assign n23111 = n22744 & n23015 ;
  assign n23112 = n23111 ^ n23014 ;
  assign n23113 = n23112 ^ n22744 ;
  assign n23114 = n23113 ^ n23112 ;
  assign n23115 = n23112 ^ n22992 ;
  assign n23116 = n23115 ^ n23112 ;
  assign n23117 = n23114 & n23116 ;
  assign n23118 = n23117 ^ n23112 ;
  assign n23119 = n23004 & n23118 ;
  assign n23120 = n23119 ^ n23112 ;
  assign n23110 = n23060 ^ n23017 ;
  assign n23121 = n23120 ^ n23110 ;
  assign n23130 = n23129 ^ n23121 ;
  assign n23103 = n23036 ^ n23014 ;
  assign n23104 = n23103 ^ n22994 ;
  assign n23107 = n22998 & n23104 ;
  assign n23108 = n23107 ^ n22994 ;
  assign n23109 = n22744 & n23108 ;
  assign n23131 = n23130 ^ n23109 ;
  assign n23099 = n23040 ^ n22989 ;
  assign n23100 = ~n22744 & n23099 ;
  assign n23098 = n23042 ^ n22996 ;
  assign n23101 = n23100 ^ n23098 ;
  assign n23102 = ~n23004 & n23101 ;
  assign n23132 = n23131 ^ n23102 ;
  assign n23133 = n23132 ^ n23023 ;
  assign n23134 = n23133 ^ n21933 ;
  assign n23097 = n22998 & n23024 ;
  assign n23135 = n23134 ^ n23097 ;
  assign n23146 = n22789 ^ n22745 ;
  assign n23147 = n23146 ^ n22788 ;
  assign n23169 = n22832 & ~n23147 ;
  assign n23138 = n22801 ^ n22781 ;
  assign n23139 = n23138 ^ n22825 ;
  assign n23140 = n23139 ^ n22833 ;
  assign n23141 = n22745 & n23140 ;
  assign n23137 = n22830 ^ n22786 ;
  assign n23142 = n23141 ^ n23137 ;
  assign n23143 = n22788 & n23142 ;
  assign n23170 = n23169 ^ n23143 ;
  assign n23151 = n22778 & n22792 ;
  assign n23148 = n22809 ^ n22786 ;
  assign n23149 = n23148 ^ n22801 ;
  assign n23150 = ~n23147 & n23149 ;
  assign n23152 = n23151 ^ n23150 ;
  assign n23171 = n23170 ^ n23152 ;
  assign n23161 = n22825 ^ n22810 ;
  assign n23162 = n23161 ^ n22797 ;
  assign n23163 = n23162 ^ n22810 ;
  assign n23164 = n22810 ^ n22788 ;
  assign n23165 = n23164 ^ n22810 ;
  assign n23166 = n23163 & n23165 ;
  assign n23167 = n23166 ^ n22810 ;
  assign n23168 = ~n22745 & n23167 ;
  assign n23172 = n23171 ^ n23168 ;
  assign n23173 = n23172 ^ n22864 ;
  assign n23174 = n23173 ^ n18819 ;
  assign n23154 = n23151 ^ n22788 ;
  assign n23155 = n23154 ^ n23151 ;
  assign n23156 = n23151 ^ n22823 ;
  assign n23157 = n23156 ^ n23151 ;
  assign n23158 = ~n23155 & n23157 ;
  assign n23159 = n23158 ^ n23151 ;
  assign n23160 = n22745 & n23159 ;
  assign n23175 = n23174 ^ n23160 ;
  assign n23136 = n22788 ^ n22745 ;
  assign n23145 = n22844 & ~n23136 ;
  assign n23176 = n23175 ^ n23145 ;
  assign n23177 = n23096 ^ x69 ;
  assign n23200 = n21997 & n22042 ;
  assign n23197 = n22873 ^ n21946 ;
  assign n23198 = n22014 & n23197 ;
  assign n23179 = n22880 ^ n22003 ;
  assign n23182 = n22022 ^ n21946 ;
  assign n23183 = ~n21999 & ~n23182 ;
  assign n23184 = ~n23179 & n23183 ;
  assign n23178 = n22031 ^ n22001 ;
  assign n23180 = n23179 ^ n23178 ;
  assign n23185 = n23184 ^ n23180 ;
  assign n23188 = n23185 ^ n22875 ;
  assign n23189 = n23188 ^ n22043 ;
  assign n23190 = n23189 ^ n23185 ;
  assign n23191 = n23185 ^ n21997 ;
  assign n23192 = n23191 ^ n23185 ;
  assign n23193 = n23190 & ~n23192 ;
  assign n23194 = n23193 ^ n23185 ;
  assign n23195 = ~n21947 & ~n23194 ;
  assign n23186 = n22872 ^ n22028 ;
  assign n23187 = n23186 ^ n23185 ;
  assign n23196 = n23195 ^ n23187 ;
  assign n23199 = n23198 ^ n23196 ;
  assign n23201 = n23200 ^ n23199 ;
  assign n23202 = ~n22907 & n23201 ;
  assign n23203 = ~n22909 & n23202 ;
  assign n23204 = ~n22067 & n23203 ;
  assign n23205 = n23204 ^ n19050 ;
  assign n23206 = n23205 ^ x91 ;
  assign n23207 = n23177 & n23206 ;
  assign n23208 = n23207 ^ n23206 ;
  assign n23209 = n23208 ^ n23177 ;
  assign n23210 = n21751 ^ n21710 ;
  assign n23211 = ~n21563 & n23210 ;
  assign n23212 = n23211 ^ n21710 ;
  assign n23215 = n23212 ^ n21814 ;
  assign n23216 = n23215 ^ n23212 ;
  assign n23217 = ~n21563 & n23216 ;
  assign n23218 = n23217 ^ n23212 ;
  assign n23219 = n21572 & n23218 ;
  assign n23220 = n23219 ^ n23212 ;
  assign n23231 = n21763 ^ n21739 ;
  assign n23232 = n23231 ^ n21783 ;
  assign n23233 = n21563 & n23232 ;
  assign n23234 = n23233 ^ n21783 ;
  assign n23224 = n21768 ^ n21728 ;
  assign n23226 = n21767 ^ n21732 ;
  assign n23225 = n21751 ^ n21714 ;
  assign n23227 = n23226 ^ n23225 ;
  assign n23228 = ~n21721 & n23227 ;
  assign n23229 = ~n23224 & n23228 ;
  assign n23230 = n23229 ^ n23227 ;
  assign n23235 = n23234 ^ n23230 ;
  assign n23236 = n23235 ^ n23234 ;
  assign n23221 = n21771 ^ n21763 ;
  assign n23222 = n23221 ^ n21734 ;
  assign n23223 = ~n21572 & n23222 ;
  assign n23237 = n23236 ^ n23223 ;
  assign n23238 = ~n21563 & n23237 ;
  assign n23239 = n23238 ^ n23235 ;
  assign n23240 = n23239 ^ n23234 ;
  assign n23241 = n21761 ^ n21563 ;
  assign n23242 = n23241 ^ n21761 ;
  assign n23245 = n21813 & n23242 ;
  assign n23246 = n23245 ^ n21761 ;
  assign n23247 = ~n23240 & ~n23246 ;
  assign n23248 = n23247 ^ n23234 ;
  assign n23249 = ~n21572 & n23248 ;
  assign n23250 = n23249 ^ n23239 ;
  assign n23251 = ~n23220 & ~n23250 ;
  assign n23252 = ~n21730 & n23251 ;
  assign n23253 = ~n21820 & n23252 ;
  assign n23254 = n23253 ^ n21236 ;
  assign n23255 = n23254 ^ x67 ;
  assign n23261 = n20930 ^ n20913 ;
  assign n23273 = n23261 ^ n20729 ;
  assign n23274 = n23273 ^ n20934 ;
  assign n23267 = n20546 ^ n20320 ;
  assign n23268 = n20724 & n23267 ;
  assign n23266 = n20937 ^ n20924 ;
  assign n23269 = n23268 ^ n23266 ;
  assign n23270 = n19336 & ~n23269 ;
  assign n23271 = n23270 ^ n23268 ;
  assign n23272 = n23271 ^ n20945 ;
  assign n23275 = n23274 ^ n23272 ;
  assign n23276 = n23275 ^ n23271 ;
  assign n23279 = n19336 & n23276 ;
  assign n23280 = n23279 ^ n23271 ;
  assign n23281 = n20894 & n23280 ;
  assign n23282 = n23281 ^ n23271 ;
  assign n23259 = n20911 ^ n20731 ;
  assign n23260 = n23259 ^ n20934 ;
  assign n23262 = n23261 ^ n23260 ;
  assign n23263 = n20894 & ~n23262 ;
  assign n23264 = n23263 ^ n20936 ;
  assign n23265 = ~n19336 & n23264 ;
  assign n23283 = n23282 ^ n23265 ;
  assign n23284 = ~n20899 & ~n23283 ;
  assign n23257 = ~n20949 & n20959 ;
  assign n23256 = n20729 & n20958 ;
  assign n23258 = n23257 ^ n23256 ;
  assign n23285 = n23284 ^ n23258 ;
  assign n23286 = ~n20978 & n23285 ;
  assign n23287 = n23286 ^ n19545 ;
  assign n23288 = n23287 ^ x92 ;
  assign n23289 = ~n23255 & n23288 ;
  assign n23292 = n22593 ^ n22591 ;
  assign n23293 = n23292 ^ n21240 ;
  assign n23294 = n23293 ^ x109 ;
  assign n23328 = n22738 ^ n17801 ;
  assign n23315 = ~n22104 & n22239 ;
  assign n23298 = n22225 ^ n22205 ;
  assign n23296 = n22246 ^ n22234 ;
  assign n23295 = n22712 ^ n22259 ;
  assign n23297 = n23296 ^ n23295 ;
  assign n23299 = n23298 ^ n23297 ;
  assign n23300 = n22103 & ~n23299 ;
  assign n23301 = n23300 ^ n23296 ;
  assign n23310 = n23301 ^ n22233 ;
  assign n23311 = n23310 ^ n22294 ;
  assign n23312 = n23311 ^ n22733 ;
  assign n23313 = n23312 ^ n22735 ;
  assign n23303 = n23301 ^ n22207 ;
  assign n23302 = n23301 ^ n22268 ;
  assign n23304 = n23303 ^ n23302 ;
  assign n23307 = ~n22103 & ~n23304 ;
  assign n23308 = n23307 ^ n23303 ;
  assign n23309 = n22102 & n23308 ;
  assign n23314 = n23313 ^ n23309 ;
  assign n23316 = n23315 ^ n23314 ;
  assign n23317 = n22102 & n22720 ;
  assign n23318 = n23317 ^ n22215 ;
  assign n23319 = n23318 ^ n23296 ;
  assign n23320 = n23319 ^ n23318 ;
  assign n23323 = n22102 & n23320 ;
  assign n23324 = n23323 ^ n23318 ;
  assign n23325 = ~n22104 & ~n23324 ;
  assign n23326 = n23325 ^ n23318 ;
  assign n23327 = ~n23316 & n23326 ;
  assign n23329 = n23328 ^ n23327 ;
  assign n23330 = n23329 ^ x86 ;
  assign n23331 = n23294 & n23330 ;
  assign n23341 = n23289 & n23331 ;
  assign n23290 = n23289 ^ n23288 ;
  assign n23291 = n23290 ^ n23255 ;
  assign n23340 = n23291 & n23331 ;
  assign n23342 = n23341 ^ n23340 ;
  assign n23338 = n23290 & n23331 ;
  assign n23339 = n23338 ^ n23331 ;
  assign n23343 = n23342 ^ n23339 ;
  assign n23332 = n23331 ^ n23294 ;
  assign n23333 = n23332 ^ n23330 ;
  assign n23335 = n23289 ^ n23255 ;
  assign n23337 = ~n23333 & ~n23335 ;
  assign n23344 = n23343 ^ n23337 ;
  assign n23345 = n23344 ^ n23335 ;
  assign n23336 = n23332 & ~n23335 ;
  assign n23346 = n23345 ^ n23336 ;
  assign n23334 = n23291 & ~n23333 ;
  assign n23347 = n23346 ^ n23334 ;
  assign n23348 = n23347 ^ n23343 ;
  assign n23349 = ~n23209 & ~n23348 ;
  assign n23398 = n23207 ^ n23177 ;
  assign n23361 = n23333 ^ n23294 ;
  assign n23362 = n23289 & n23361 ;
  assign n23399 = n23398 ^ n23362 ;
  assign n23356 = n23290 & ~n23333 ;
  assign n23368 = n23356 ^ n23341 ;
  assign n23369 = n23368 ^ n23362 ;
  assign n23358 = n23337 ^ n23334 ;
  assign n23357 = n23356 ^ n23333 ;
  assign n23359 = n23358 ^ n23357 ;
  assign n23370 = n23369 ^ n23359 ;
  assign n23367 = n23356 ^ n23289 ;
  assign n23371 = n23370 ^ n23367 ;
  assign n23372 = n23371 ^ n23368 ;
  assign n23373 = n23372 ^ n23338 ;
  assign n23365 = n23290 & n23361 ;
  assign n23366 = n23365 ^ n23359 ;
  assign n23374 = n23373 ^ n23366 ;
  assign n23364 = n23362 ^ n23288 ;
  assign n23375 = n23374 ^ n23364 ;
  assign n23397 = n23375 ^ n23344 ;
  assign n23400 = n23399 ^ n23397 ;
  assign n23376 = n23371 ^ n23365 ;
  assign n23401 = n23376 ^ n23208 ;
  assign n23404 = n23398 & n23401 ;
  assign n23405 = n23404 ^ n23208 ;
  assign n23406 = n23400 & n23405 ;
  assign n23407 = n23406 ^ n23206 ;
  assign n23352 = n23291 & n23332 ;
  assign n23390 = n23366 ^ n23352 ;
  assign n23388 = n23340 ^ n23291 ;
  assign n23389 = n23388 ^ n23352 ;
  assign n23391 = n23390 ^ n23389 ;
  assign n23392 = n23390 ^ n23206 ;
  assign n23393 = n23392 ^ n23390 ;
  assign n23394 = n23391 & n23393 ;
  assign n23395 = n23394 ^ n23390 ;
  assign n23396 = ~n23177 & n23395 ;
  assign n23408 = n23407 ^ n23396 ;
  assign n23380 = n23356 ^ n23338 ;
  assign n23409 = n23408 ^ n23380 ;
  assign n23377 = n23376 ^ n23375 ;
  assign n23353 = n23352 ^ n23334 ;
  assign n23354 = n23353 ^ n23343 ;
  assign n23350 = n23288 ^ n23255 ;
  assign n23351 = n23350 ^ n23330 ;
  assign n23355 = n23354 ^ n23351 ;
  assign n23360 = n23359 ^ n23355 ;
  assign n23363 = n23362 ^ n23360 ;
  assign n23378 = n23377 ^ n23363 ;
  assign n23379 = n23378 ^ n23351 ;
  assign n23381 = n23380 ^ n23379 ;
  assign n23382 = n23381 ^ n23380 ;
  assign n23383 = n23380 ^ n23206 ;
  assign n23384 = n23383 ^ n23380 ;
  assign n23385 = ~n23382 & n23384 ;
  assign n23386 = n23385 ^ n23380 ;
  assign n23387 = n23177 & n23386 ;
  assign n23410 = n23409 ^ n23387 ;
  assign n23411 = ~n23349 & n23410 ;
  assign n23412 = n23388 ^ n23334 ;
  assign n23413 = n23398 & n23412 ;
  assign n23414 = n23411 & ~n23413 ;
  assign n23415 = n23414 ^ n21672 ;
  assign n23441 = n23148 ^ n22820 ;
  assign n23417 = n22831 ^ n22810 ;
  assign n23442 = n23441 ^ n23417 ;
  assign n23443 = n23146 & ~n23442 ;
  assign n23428 = n22799 ^ n22789 ;
  assign n23429 = n23147 ^ n22801 ;
  assign n23430 = n22801 ^ n22789 ;
  assign n23431 = n23430 ^ n22801 ;
  assign n23432 = n23429 & ~n23431 ;
  assign n23433 = n23432 ^ n22801 ;
  assign n23434 = n23428 & n23433 ;
  assign n23435 = n23434 ^ n22799 ;
  assign n23436 = n23435 ^ n23150 ;
  assign n23437 = n23436 ^ n23417 ;
  assign n23438 = n23437 ^ n20058 ;
  assign n23419 = n22793 ^ n22776 ;
  assign n23420 = n23419 ^ n22777 ;
  assign n23418 = n23417 ^ n22781 ;
  assign n23421 = n23420 ^ n23418 ;
  assign n23422 = n23421 ^ n23417 ;
  assign n23423 = n23417 ^ n22788 ;
  assign n23424 = n23423 ^ n23417 ;
  assign n23425 = n23422 & n23424 ;
  assign n23426 = n23425 ^ n23417 ;
  assign n23427 = n23136 & n23426 ;
  assign n23439 = n23438 ^ n23427 ;
  assign n23416 = n22789 & n22846 ;
  assign n23440 = n23439 ^ n23416 ;
  assign n23444 = n23443 ^ n23440 ;
  assign n23446 = ~n23209 & n23336 ;
  assign n23457 = n23388 ^ n23353 ;
  assign n23458 = n23206 & n23457 ;
  assign n23462 = n23458 ^ n23206 ;
  assign n23456 = n23352 ^ n23347 ;
  assign n23459 = n23458 ^ n23456 ;
  assign n23454 = n23342 ^ n23334 ;
  assign n23455 = ~n23206 & ~n23454 ;
  assign n23460 = n23459 ^ n23455 ;
  assign n23461 = ~n23177 & ~n23460 ;
  assign n23463 = n23462 ^ n23461 ;
  assign n23450 = n23354 ^ n23208 ;
  assign n23451 = n23398 & ~n23450 ;
  assign n23452 = n23451 ^ n23208 ;
  assign n23453 = n23399 & n23452 ;
  assign n23464 = n23463 ^ n23453 ;
  assign n23465 = n23464 ^ n23366 ;
  assign n23449 = n23207 & n23336 ;
  assign n23466 = n23465 ^ n23449 ;
  assign n23447 = n23206 ^ n23177 ;
  assign n23448 = n23374 & n23447 ;
  assign n23467 = n23466 ^ n23448 ;
  assign n23468 = ~n23446 & ~n23467 ;
  assign n23445 = n23207 & n23397 ;
  assign n23469 = n23468 ^ n23445 ;
  assign n23470 = n23375 ^ n23340 ;
  assign n23471 = n23340 ^ n23206 ;
  assign n23472 = n23471 ^ n23340 ;
  assign n23473 = n23470 & ~n23472 ;
  assign n23474 = n23473 ^ n23340 ;
  assign n23475 = ~n23447 & n23474 ;
  assign n23476 = n23469 & ~n23475 ;
  assign n23477 = n23476 ^ n22198 ;
  assign n23511 = n21814 ^ n21737 ;
  assign n23512 = n21721 & n23511 ;
  assign n23494 = n21764 ^ n21762 ;
  assign n23495 = n23494 ^ n21751 ;
  assign n23496 = n23495 ^ n21771 ;
  assign n23497 = n21563 & ~n23496 ;
  assign n23498 = n23497 ^ n21762 ;
  assign n23508 = n23498 ^ n20386 ;
  assign n23509 = n23508 ^ n21748 ;
  assign n23492 = n21572 ^ n21563 ;
  assign n23499 = n21782 ^ n21728 ;
  assign n23500 = n23499 ^ n21714 ;
  assign n23501 = n23500 ^ n23498 ;
  assign n23493 = n21770 ^ n21762 ;
  assign n23502 = n23501 ^ n23493 ;
  assign n23503 = n23501 ^ n21563 ;
  assign n23504 = n23503 ^ n23501 ;
  assign n23505 = n23502 & ~n23504 ;
  assign n23506 = n23505 ^ n23501 ;
  assign n23507 = ~n23492 & n23506 ;
  assign n23510 = n23509 ^ n23507 ;
  assign n23513 = n23512 ^ n23510 ;
  assign n23484 = n21763 ^ n21761 ;
  assign n23485 = n23484 ^ n21736 ;
  assign n23486 = n23485 ^ n21763 ;
  assign n23487 = n21763 ^ n21563 ;
  assign n23488 = n23487 ^ n21763 ;
  assign n23489 = ~n23486 & n23488 ;
  assign n23490 = n23489 ^ n21763 ;
  assign n23491 = ~n21572 & ~n23490 ;
  assign n23514 = n23513 ^ n23491 ;
  assign n23478 = n21769 ^ n21760 ;
  assign n23479 = n21760 ^ n21572 ;
  assign n23480 = n23479 ^ n21760 ;
  assign n23481 = ~n23478 & n23480 ;
  assign n23482 = n23481 ^ n21760 ;
  assign n23483 = ~n21563 & ~n23482 ;
  assign n23515 = n23514 ^ n23483 ;
  assign n23529 = n23176 ^ x126 ;
  assign n23543 = n21199 ^ n21196 ;
  assign n23544 = n21470 ^ n21468 ;
  assign n23545 = ~n23543 & n23544 ;
  assign n23546 = n23545 ^ n21471 ;
  assign n23536 = n23075 ^ n21492 ;
  assign n23537 = n21154 & n23536 ;
  assign n23538 = n23537 ^ n21492 ;
  assign n23547 = n23546 ^ n23538 ;
  assign n23542 = n21197 & n21461 ;
  assign n23548 = n23547 ^ n23542 ;
  assign n23539 = n23538 ^ n21480 ;
  assign n23533 = n21502 ^ n21476 ;
  assign n23534 = n23533 ^ n21473 ;
  assign n23535 = ~n21154 & ~n23534 ;
  assign n23540 = n23539 ^ n23535 ;
  assign n23541 = ~n21472 & n23540 ;
  assign n23549 = n23548 ^ n23541 ;
  assign n23531 = n21473 ^ n21465 ;
  assign n23532 = n21197 & n23531 ;
  assign n23550 = n23549 ^ n23532 ;
  assign n23530 = n21198 & ~n21515 ;
  assign n23551 = n23550 ^ n23530 ;
  assign n23552 = n21468 ^ n21453 ;
  assign n23553 = n23552 ^ n21526 ;
  assign n23554 = n21526 ^ n21154 ;
  assign n23555 = n23554 ^ n21526 ;
  assign n23556 = n23553 & n23555 ;
  assign n23557 = n23556 ^ n21526 ;
  assign n23558 = ~n21196 & n23557 ;
  assign n23559 = ~n23551 & ~n23558 ;
  assign n23560 = ~n23078 & n23559 ;
  assign n23561 = n23560 ^ n18301 ;
  assign n23562 = n23561 ^ x84 ;
  assign n23563 = ~n23529 & n23562 ;
  assign n23564 = n23205 ^ x85 ;
  assign n23584 = n22932 ^ n22409 ;
  assign n23579 = n22405 ^ n22395 ;
  assign n23578 = n22417 ^ n22399 ;
  assign n23580 = n23579 ^ n23578 ;
  assign n23581 = n22301 & ~n23580 ;
  assign n23565 = n22932 ^ n22918 ;
  assign n23574 = n23565 ^ n22404 ;
  assign n23566 = n22414 ^ n22405 ;
  assign n23567 = n23566 ^ n23565 ;
  assign n23568 = n23567 ^ n23566 ;
  assign n23569 = n23566 ^ n22301 ;
  assign n23570 = n23569 ^ n23566 ;
  assign n23571 = n23568 & ~n23570 ;
  assign n23572 = n23571 ^ n23566 ;
  assign n23573 = n22300 & n23572 ;
  assign n23575 = ~n22301 & n23573 ;
  assign n23576 = ~n23574 & n23575 ;
  assign n23577 = n23576 ^ n23573 ;
  assign n23582 = n23581 ^ n23577 ;
  assign n23583 = n23582 ^ n23576 ;
  assign n23585 = n23584 ^ n23583 ;
  assign n23586 = n23585 ^ n23573 ;
  assign n23587 = ~n22302 & n23586 ;
  assign n23588 = n23587 ^ n23582 ;
  assign n23597 = n23588 ^ n22462 ;
  assign n23589 = ~n22301 & ~n23588 ;
  assign n23590 = n22454 ^ n22395 ;
  assign n23591 = n23590 ^ n22401 ;
  assign n23592 = n22401 ^ n22300 ;
  assign n23593 = n23592 ^ n22401 ;
  assign n23594 = n23591 & n23593 ;
  assign n23595 = n23594 ^ n22401 ;
  assign n23596 = n23589 & n23595 ;
  assign n23598 = n23597 ^ n23596 ;
  assign n23599 = ~n22452 & ~n23598 ;
  assign n23600 = ~n22941 & n23599 ;
  assign n23601 = n23600 ^ n18533 ;
  assign n23602 = n23601 ^ x70 ;
  assign n23603 = ~n23564 & n23602 ;
  assign n23606 = n23603 ^ n23564 ;
  assign n23611 = n23563 & ~n23606 ;
  assign n23605 = n23563 ^ n23529 ;
  assign n23609 = n23605 ^ n23562 ;
  assign n23678 = n23611 ^ n23609 ;
  assign n23516 = n22973 ^ n22541 ;
  assign n23518 = n23516 ^ n22572 ;
  assign n23517 = n23516 ^ n22585 ;
  assign n23519 = n23518 ^ n23517 ;
  assign n23522 = ~n22563 & n23519 ;
  assign n23523 = n23522 ^ n23518 ;
  assign n23524 = n22551 & ~n23523 ;
  assign n23525 = n23524 ^ n23516 ;
  assign n23526 = n22963 & ~n23525 ;
  assign n23527 = n23526 ^ n19282 ;
  assign n23528 = n23527 ^ x102 ;
  assign n23622 = n23329 ^ x116 ;
  assign n23636 = n23528 & n23622 ;
  assign n23637 = n23636 ^ n23622 ;
  assign n23638 = n23637 ^ n23528 ;
  assign n23679 = n23638 ^ n23602 ;
  assign n23680 = n23679 ^ n23638 ;
  assign n23683 = ~n23636 & ~n23680 ;
  assign n23684 = n23683 ^ n23638 ;
  assign n23685 = ~n23564 & ~n23684 ;
  assign n23686 = n23678 & ~n23685 ;
  assign n23640 = n23603 ^ n23602 ;
  assign n23644 = n23563 & n23640 ;
  assign n23610 = ~n23606 & n23609 ;
  assign n23612 = n23611 ^ n23610 ;
  assign n23607 = ~n23605 & ~n23606 ;
  assign n23608 = n23607 ^ n23606 ;
  assign n23613 = n23612 ^ n23608 ;
  assign n23659 = n23644 ^ n23613 ;
  assign n23641 = n23606 ^ n23602 ;
  assign n23675 = n23659 ^ n23641 ;
  assign n23676 = ~n23638 & ~n23675 ;
  assign n23665 = n23609 & n23641 ;
  assign n23666 = n23665 ^ n23641 ;
  assign n23642 = n23562 & n23641 ;
  assign n23667 = n23666 ^ n23642 ;
  assign n23672 = n23622 & n23667 ;
  assign n23639 = n23638 ^ n23622 ;
  assign n23660 = n23659 ^ n23611 ;
  assign n23618 = n23603 & n23609 ;
  assign n23604 = n23563 & n23603 ;
  assign n23619 = n23618 ^ n23604 ;
  assign n23661 = n23660 ^ n23619 ;
  assign n23662 = n23661 ^ n23642 ;
  assign n23657 = n23618 ^ n23563 ;
  assign n23658 = n23657 ^ n23613 ;
  assign n23663 = n23662 ^ n23658 ;
  assign n23664 = n23663 ^ n23641 ;
  assign n23668 = n23667 ^ n23664 ;
  assign n23669 = n23639 & n23668 ;
  assign n23615 = n23609 ^ n23529 ;
  assign n23616 = n23603 & n23615 ;
  assign n23617 = n23616 ^ n23603 ;
  assign n23620 = n23619 ^ n23617 ;
  assign n23654 = n23620 & n23637 ;
  assign n23653 = n23616 & n23639 ;
  assign n23655 = n23654 ^ n23653 ;
  assign n23648 = n23609 & n23640 ;
  assign n23647 = ~n23605 & n23640 ;
  assign n23649 = n23648 ^ n23647 ;
  assign n23643 = n23642 ^ n23640 ;
  assign n23645 = n23644 ^ n23643 ;
  assign n23646 = ~n23639 & n23645 ;
  assign n23650 = n23649 ^ n23646 ;
  assign n23628 = n23619 ^ n23528 ;
  assign n23629 = n23628 ^ n23619 ;
  assign n23630 = n23619 ^ n23607 ;
  assign n23631 = n23630 ^ n23619 ;
  assign n23632 = ~n23629 & n23631 ;
  assign n23633 = n23632 ^ n23619 ;
  assign n23634 = ~n23622 & n23633 ;
  assign n23635 = n23634 ^ n23619 ;
  assign n23651 = n23650 ^ n23635 ;
  assign n23614 = n23613 ^ n23604 ;
  assign n23621 = n23620 ^ n23614 ;
  assign n23625 = ~n23621 & ~n23622 ;
  assign n23626 = n23625 ^ n23620 ;
  assign n23627 = n23528 & n23626 ;
  assign n23652 = n23651 ^ n23627 ;
  assign n23656 = n23655 ^ n23652 ;
  assign n23670 = n23669 ^ n23656 ;
  assign n23671 = n23670 ^ n22528 ;
  assign n23673 = n23672 ^ n23671 ;
  assign n23674 = n23673 ^ n23609 ;
  assign n23677 = n23676 ^ n23674 ;
  assign n23687 = n23686 ^ n23677 ;
  assign n23718 = n22943 ^ n22452 ;
  assign n23701 = n22390 ^ n22385 ;
  assign n23702 = n23701 ^ n23584 ;
  assign n23703 = n22451 & ~n23702 ;
  assign n23704 = n22458 ^ n22409 ;
  assign n23705 = n23704 ^ n22458 ;
  assign n23706 = n22950 ^ n22458 ;
  assign n23707 = n23706 ^ n22458 ;
  assign n23708 = ~n23705 & n23707 ;
  assign n23709 = n23708 ^ n22458 ;
  assign n23710 = ~n23703 & ~n23709 ;
  assign n23719 = n23718 ^ n23710 ;
  assign n23711 = n23710 ^ n22930 ;
  assign n23712 = n23711 ^ n22390 ;
  assign n23713 = n23712 ^ n23590 ;
  assign n23714 = n23713 ^ n23710 ;
  assign n23715 = ~n22301 & n23714 ;
  assign n23716 = n23715 ^ n23711 ;
  assign n23717 = ~n22300 & n23716 ;
  assign n23720 = n23719 ^ n23717 ;
  assign n23700 = ~n22302 & ~n23578 ;
  assign n23721 = n23720 ^ n23700 ;
  assign n23695 = n22404 ^ n22300 ;
  assign n23696 = n23695 ^ n22404 ;
  assign n23697 = n22415 & n23696 ;
  assign n23698 = n23697 ^ n22404 ;
  assign n23699 = ~n22301 & n23698 ;
  assign n23722 = n23721 ^ n23699 ;
  assign n23688 = n22918 ^ n22301 ;
  assign n23689 = n23688 ^ n22918 ;
  assign n23692 = n22387 & n23689 ;
  assign n23693 = n23692 ^ n22918 ;
  assign n23694 = n22300 & n23693 ;
  assign n23723 = n23722 ^ n23694 ;
  assign n23724 = ~n22941 & ~n23723 ;
  assign n23725 = n23724 ^ n19811 ;
  assign n23813 = n23527 ^ x122 ;
  assign n23830 = n22042 ^ n22016 ;
  assign n23826 = n22035 ^ n22016 ;
  assign n23827 = n23826 ^ n21946 ;
  assign n23828 = n23827 ^ n22032 ;
  assign n23829 = n21997 & n23828 ;
  assign n23831 = n23830 ^ n23829 ;
  assign n23832 = n22015 & n23831 ;
  assign n23821 = n21858 & n21909 ;
  assign n23822 = ~n21997 & n23821 ;
  assign n23816 = n22888 ^ n22048 ;
  assign n23817 = n23816 ^ n23178 ;
  assign n23818 = n21997 & n23817 ;
  assign n23819 = n23818 ^ n22888 ;
  assign n23820 = n23819 ^ n22022 ;
  assign n23823 = n23822 ^ n23820 ;
  assign n23824 = ~n21947 & n23823 ;
  assign n23825 = n23824 ^ n23819 ;
  assign n23833 = n23832 ^ n23825 ;
  assign n23834 = n23833 ^ n22000 ;
  assign n23835 = n23834 ^ n22909 ;
  assign n23814 = n23178 ^ n22005 ;
  assign n23815 = ~n22013 & n23814 ;
  assign n23836 = n23835 ^ n23815 ;
  assign n23837 = ~n22039 & ~n23836 ;
  assign n23838 = n22019 ^ n21997 ;
  assign n23839 = n23838 ^ n21947 ;
  assign n23840 = n23839 ^ n22019 ;
  assign n23841 = n22020 ^ n22019 ;
  assign n23842 = n21947 & n23841 ;
  assign n23843 = n23842 ^ n22019 ;
  assign n23844 = ~n23840 & n23843 ;
  assign n23845 = n23844 ^ n22019 ;
  assign n23846 = n23837 & n23845 ;
  assign n23847 = n23846 ^ n23837 ;
  assign n23848 = ~n22907 & n23847 ;
  assign n23849 = ~n22067 & n23848 ;
  assign n23850 = n23849 ^ n19998 ;
  assign n23851 = n23850 ^ x120 ;
  assign n23852 = n23813 & ~n23851 ;
  assign n23853 = n23852 ^ n23813 ;
  assign n23773 = n22278 ^ n22252 ;
  assign n23774 = n23773 ^ n23326 ;
  assign n23766 = n23298 ^ n22244 ;
  assign n23767 = n23766 ^ n22269 ;
  assign n23768 = n22269 ^ n22103 ;
  assign n23769 = n23768 ^ n22269 ;
  assign n23770 = n23767 & ~n23769 ;
  assign n23771 = n23770 ^ n22269 ;
  assign n23772 = ~n22102 & n23771 ;
  assign n23775 = n23774 ^ n23772 ;
  assign n23776 = n23775 ^ n22738 ;
  assign n23777 = n23776 ^ n22223 ;
  assign n23778 = n23777 ^ n20577 ;
  assign n23764 = n22243 ^ n22210 ;
  assign n23765 = ~n22104 & n23764 ;
  assign n23779 = n23778 ^ n23765 ;
  assign n23759 = n22239 ^ n22204 ;
  assign n23760 = n23759 ^ n23296 ;
  assign n23761 = n22102 & n23760 ;
  assign n23762 = n23761 ^ n22278 ;
  assign n23763 = ~n22103 & ~n23762 ;
  assign n23780 = n23779 ^ n23763 ;
  assign n23781 = n23780 ^ x105 ;
  assign n23809 = n20979 ^ n20601 ;
  assign n23782 = n20894 ^ n19336 ;
  assign n23798 = n20935 ^ n20733 ;
  assign n23795 = n20931 ^ n20904 ;
  assign n23796 = n23795 ^ n20964 ;
  assign n23797 = n23796 ^ n20949 ;
  assign n23799 = n23798 ^ n23797 ;
  assign n23800 = n23797 ^ n19336 ;
  assign n23801 = n23800 ^ n23797 ;
  assign n23802 = ~n23799 & n23801 ;
  assign n23803 = n23802 ^ n23797 ;
  assign n23804 = n23782 & ~n23803 ;
  assign n23788 = n20929 ^ n20909 ;
  assign n23789 = n23788 ^ n20903 ;
  assign n23790 = n20903 ^ n19336 ;
  assign n23791 = n23790 ^ n20903 ;
  assign n23792 = n23789 & ~n23791 ;
  assign n23793 = n23792 ^ n20903 ;
  assign n23794 = ~n20894 & n23793 ;
  assign n23805 = n23804 ^ n23794 ;
  assign n23784 = n20926 ^ n20730 ;
  assign n23785 = n23784 ^ n20946 ;
  assign n23786 = n20959 & ~n23785 ;
  assign n23806 = n23805 ^ n23786 ;
  assign n23783 = ~n23261 & ~n23782 ;
  assign n23807 = n23806 ^ n23783 ;
  assign n23808 = ~n23256 & ~n23807 ;
  assign n23810 = n23809 ^ n23808 ;
  assign n23811 = n23810 ^ x66 ;
  assign n23812 = n23781 & n23811 ;
  assign n23857 = n23812 ^ n23811 ;
  assign n23866 = n23857 ^ n23781 ;
  assign n23867 = n23866 ^ n23811 ;
  assign n23869 = n23853 & n23867 ;
  assign n23753 = n21742 ^ n20145 ;
  assign n23754 = n23753 ^ n21808 ;
  assign n23749 = n23220 ^ n21758 ;
  assign n23736 = n21764 ^ n21740 ;
  assign n23734 = n21749 ^ n21714 ;
  assign n23726 = n21738 ^ n21734 ;
  assign n23727 = n23726 ^ n23499 ;
  assign n23728 = n23727 ^ n21738 ;
  assign n23729 = n21738 ^ n21572 ;
  assign n23730 = n23729 ^ n21738 ;
  assign n23731 = n23728 & ~n23730 ;
  assign n23732 = n23731 ^ n21738 ;
  assign n23733 = n21563 & n23732 ;
  assign n23735 = n23734 ^ n23733 ;
  assign n23737 = n23736 ^ n23735 ;
  assign n23738 = n23737 ^ n23733 ;
  assign n23739 = n21563 & ~n23738 ;
  assign n23740 = n23739 ^ n23735 ;
  assign n23750 = n23749 ^ n23740 ;
  assign n23741 = n23740 ^ n23733 ;
  assign n23742 = n23741 ^ n23221 ;
  assign n23743 = n23742 ^ n23741 ;
  assign n23744 = n23741 ^ n21563 ;
  assign n23745 = n23744 ^ n23741 ;
  assign n23746 = n23743 & ~n23745 ;
  assign n23747 = n23746 ^ n23741 ;
  assign n23748 = n23492 & n23747 ;
  assign n23751 = n23750 ^ n23748 ;
  assign n23752 = ~n21720 & ~n23751 ;
  assign n23755 = n23754 ^ n23752 ;
  assign n23756 = n23755 ^ x88 ;
  assign n23757 = n23176 ^ x81 ;
  assign n23887 = ~n23756 & ~n23757 ;
  assign n23933 = n23869 & n23887 ;
  assign n23854 = n23853 ^ n23851 ;
  assign n23871 = n23854 ^ n23813 ;
  assign n23872 = ~n23866 & ~n23871 ;
  assign n23858 = n23852 & n23857 ;
  assign n23856 = n23812 & n23853 ;
  assign n23859 = n23858 ^ n23856 ;
  assign n23926 = n23872 ^ n23859 ;
  assign n23927 = ~n23756 & n23926 ;
  assign n23879 = n23858 ^ n23857 ;
  assign n23877 = n23857 & ~n23871 ;
  assign n23876 = n23853 & n23857 ;
  assign n23878 = n23877 ^ n23876 ;
  assign n23880 = n23879 ^ n23878 ;
  assign n23855 = n23812 & n23854 ;
  assign n23881 = n23880 ^ n23855 ;
  assign n23873 = ~n23813 & ~n23866 ;
  assign n23874 = n23873 ^ n23872 ;
  assign n23875 = n23874 ^ n23854 ;
  assign n23882 = n23881 ^ n23875 ;
  assign n23885 = n23882 ^ n23877 ;
  assign n23886 = n23885 ^ n23874 ;
  assign n23888 = n23887 ^ n23757 ;
  assign n23889 = ~n23886 & n23888 ;
  assign n23891 = n23880 ^ n23873 ;
  assign n23890 = n23885 & n23887 ;
  assign n23892 = n23891 ^ n23890 ;
  assign n23893 = ~n23889 & n23892 ;
  assign n23883 = n23882 ^ n23867 ;
  assign n23868 = n23852 & n23867 ;
  assign n23870 = n23869 ^ n23868 ;
  assign n23884 = n23883 ^ n23870 ;
  assign n23894 = n23893 ^ n23884 ;
  assign n23928 = n23927 ^ n23894 ;
  assign n23930 = n23928 ^ n23880 ;
  assign n23931 = n23757 & n23930 ;
  assign n23913 = n23812 & ~n23871 ;
  assign n23895 = n23852 & ~n23866 ;
  assign n23896 = n23895 ^ n23856 ;
  assign n23921 = n23913 ^ n23896 ;
  assign n23922 = n23887 & n23921 ;
  assign n23914 = n23913 ^ n23870 ;
  assign n23915 = n23914 ^ n23870 ;
  assign n23916 = n23870 ^ n23756 ;
  assign n23917 = n23916 ^ n23870 ;
  assign n23918 = n23915 & ~n23917 ;
  assign n23919 = n23918 ^ n23870 ;
  assign n23920 = n23757 & n23919 ;
  assign n23923 = n23922 ^ n23920 ;
  assign n23897 = n23896 ^ n23868 ;
  assign n23898 = n23897 ^ n23852 ;
  assign n23899 = n23898 ^ n23859 ;
  assign n23900 = n23899 ^ n23756 ;
  assign n23901 = n23895 ^ n23866 ;
  assign n23902 = n23901 ^ n23873 ;
  assign n23907 = n23902 ^ n23899 ;
  assign n23904 = n23874 ^ n23855 ;
  assign n23903 = n23902 ^ n23878 ;
  assign n23905 = n23904 ^ n23903 ;
  assign n23906 = n23757 & ~n23905 ;
  assign n23908 = n23907 ^ n23906 ;
  assign n23909 = n23900 & n23908 ;
  assign n23910 = n23909 ^ n23756 ;
  assign n23911 = n23910 ^ n23894 ;
  assign n23758 = n23757 ^ n23756 ;
  assign n23860 = n23859 ^ n23855 ;
  assign n23861 = n23859 ^ n23757 ;
  assign n23862 = n23861 ^ n23859 ;
  assign n23863 = n23860 & n23862 ;
  assign n23864 = n23863 ^ n23859 ;
  assign n23865 = n23758 & n23864 ;
  assign n23912 = n23911 ^ n23865 ;
  assign n23924 = n23923 ^ n23912 ;
  assign n23925 = n23924 ^ n21857 ;
  assign n23932 = n23931 ^ n23925 ;
  assign n23934 = n23933 ^ n23932 ;
  assign n23951 = n23880 ^ n23757 ;
  assign n23952 = n23951 ^ n23880 ;
  assign n23955 = n23881 & ~n23952 ;
  assign n23956 = n23955 ^ n23880 ;
  assign n23957 = ~n23758 & n23956 ;
  assign n23944 = n23882 ^ n23872 ;
  assign n23945 = n23944 ^ n23904 ;
  assign n23946 = ~n23757 & n23945 ;
  assign n23947 = n23946 ^ n23904 ;
  assign n23958 = n23957 ^ n23947 ;
  assign n23943 = n23921 ^ n23885 ;
  assign n23948 = n23947 ^ n23943 ;
  assign n23939 = n23885 ^ n23852 ;
  assign n23940 = n23939 ^ n23884 ;
  assign n23941 = n23940 ^ n23921 ;
  assign n23942 = ~n23757 & n23941 ;
  assign n23949 = n23948 ^ n23942 ;
  assign n23950 = n23756 & n23949 ;
  assign n23959 = n23958 ^ n23950 ;
  assign n23960 = n23877 ^ n23757 ;
  assign n23961 = n23960 ^ n23877 ;
  assign n23964 = n23878 & ~n23961 ;
  assign n23965 = n23964 ^ n23877 ;
  assign n23966 = n23758 & n23965 ;
  assign n23967 = ~n23959 & ~n23966 ;
  assign n23968 = n23899 ^ n23876 ;
  assign n23969 = n23968 ^ n23904 ;
  assign n23970 = n23904 ^ n23757 ;
  assign n23971 = n23970 ^ n23904 ;
  assign n23972 = n23969 & n23971 ;
  assign n23973 = n23972 ^ n23904 ;
  assign n23974 = n23758 & n23973 ;
  assign n23975 = n23967 & ~n23974 ;
  assign n23936 = n23902 ^ n23858 ;
  assign n23937 = n23887 & ~n23936 ;
  assign n23935 = n23923 ^ n21705 ;
  assign n23938 = n23937 ^ n23935 ;
  assign n23976 = n23975 ^ n23938 ;
  assign n24009 = n21198 & n21470 ;
  assign n24006 = ~n21196 & ~n21502 ;
  assign n23988 = n21479 ^ n21196 ;
  assign n23991 = n21154 & ~n21476 ;
  assign n23992 = n23991 ^ n21496 ;
  assign n23995 = n23988 ^ n21479 ;
  assign n23996 = ~n23992 & ~n23995 ;
  assign n23997 = n23996 ^ n21154 ;
  assign n23998 = ~n23988 & n23997 ;
  assign n23999 = n23998 ^ n21196 ;
  assign n23987 = n21457 & ~n23543 ;
  assign n24000 = n23999 ^ n23987 ;
  assign n24003 = n24000 ^ n23080 ;
  assign n23986 = n21491 ^ n21453 ;
  assign n24001 = ~n21472 & n24000 ;
  assign n24002 = n23986 & n24001 ;
  assign n24004 = n24003 ^ n24002 ;
  assign n23984 = n21475 ^ n21458 ;
  assign n23985 = n21198 & n23984 ;
  assign n24005 = n24004 ^ n23985 ;
  assign n24007 = n24006 ^ n24005 ;
  assign n23979 = n21460 ^ n21196 ;
  assign n23980 = n23979 ^ n21460 ;
  assign n23981 = n21490 & n23980 ;
  assign n23982 = n23981 ^ n21460 ;
  assign n23983 = n21472 & n23982 ;
  assign n24008 = n24007 ^ n23983 ;
  assign n24010 = n24009 ^ n24008 ;
  assign n24011 = ~n23545 & n24010 ;
  assign n24012 = ~n21469 & n24011 ;
  assign n24013 = ~n23542 & n24012 ;
  assign n24014 = n24013 ^ n20092 ;
  assign n24036 = n23027 ^ n22989 ;
  assign n24037 = n24036 ^ n23030 ;
  assign n24038 = n22744 & n24037 ;
  assign n24025 = n23038 ^ n23036 ;
  assign n24024 = n23010 ^ n22995 ;
  assign n24026 = n24025 ^ n24024 ;
  assign n24017 = n23041 ^ n23019 ;
  assign n24018 = n24017 ^ n23038 ;
  assign n24023 = n24018 ^ n23029 ;
  assign n24027 = n24026 ^ n24023 ;
  assign n24028 = ~n22744 & n24027 ;
  assign n24029 = n24028 ^ n24023 ;
  assign n24039 = n24038 ^ n24029 ;
  assign n24040 = n22998 & n24039 ;
  assign n24015 = n23005 ^ n22996 ;
  assign n24016 = n24015 ^ n23103 ;
  assign n24019 = n24018 ^ n24016 ;
  assign n24020 = ~n23010 & ~n24019 ;
  assign n24021 = n24020 ^ n23005 ;
  assign n24031 = n23124 ^ n23010 ;
  assign n24022 = n23124 ^ n23007 ;
  assign n24030 = n24029 ^ n24022 ;
  assign n24032 = n24031 ^ n24030 ;
  assign n24033 = n24032 ^ n24029 ;
  assign n24034 = n24021 & n24033 ;
  assign n24035 = n24034 ^ n24030 ;
  assign n24041 = n24040 ^ n24035 ;
  assign n24042 = n24041 ^ n23056 ;
  assign n24043 = n24042 ^ n23120 ;
  assign n24044 = ~n23023 & ~n24043 ;
  assign n24045 = ~n23018 & n24044 ;
  assign n24046 = n24045 ^ n22164 ;
  assign n24066 = n20924 & n20958 ;
  assign n24059 = n20964 ^ n20904 ;
  assign n24060 = ~n20894 & n24059 ;
  assign n24056 = n20931 ^ n20917 ;
  assign n24050 = n20935 ^ n20730 ;
  assign n24048 = n20946 ^ n20908 ;
  assign n24049 = n24048 ^ n23274 ;
  assign n24051 = n24050 ^ n24049 ;
  assign n24052 = n19336 & n24051 ;
  assign n24053 = n24052 ^ n24050 ;
  assign n24057 = n24056 ^ n24053 ;
  assign n24054 = n24053 ^ n23258 ;
  assign n24058 = n24057 ^ n24054 ;
  assign n24061 = n24060 ^ n24058 ;
  assign n24062 = ~n20913 & ~n24061 ;
  assign n24063 = n24062 ^ n24054 ;
  assign n24064 = ~n23782 & ~n24063 ;
  assign n24047 = n20978 ^ n20495 ;
  assign n24055 = n24054 ^ n24047 ;
  assign n24065 = n24064 ^ n24055 ;
  assign n24067 = n24066 ^ n24065 ;
  assign n24094 = n22653 ^ n22601 ;
  assign n24095 = n22649 & n24094 ;
  assign n24079 = n22705 ^ n22651 ;
  assign n24080 = n22668 ^ n22619 ;
  assign n24081 = n24080 ^ n22666 ;
  assign n24082 = ~n24079 & n24081 ;
  assign n24077 = n22668 ^ n22621 ;
  assign n24078 = ~n22652 & n24077 ;
  assign n24083 = n24082 ^ n24078 ;
  assign n24075 = n22676 ^ n22643 ;
  assign n24074 = n22637 ^ n22633 ;
  assign n24076 = n24075 ^ n24074 ;
  assign n24084 = n24083 ^ n24076 ;
  assign n24085 = n24084 ^ n24083 ;
  assign n24086 = n24085 ^ n22662 ;
  assign n24087 = n24086 ^ n24085 ;
  assign n24090 = ~n21536 & n24087 ;
  assign n24091 = n24090 ^ n24085 ;
  assign n24092 = ~n21824 & ~n24091 ;
  assign n24093 = n24092 ^ n24084 ;
  assign n24096 = n24095 ^ n24093 ;
  assign n24068 = n22641 ^ n22605 ;
  assign n24069 = n22605 ^ n21823 ;
  assign n24070 = n24069 ^ n22605 ;
  assign n24071 = n24068 & n24070 ;
  assign n24072 = n24071 ^ n22605 ;
  assign n24073 = n21536 & n24072 ;
  assign n24097 = n24096 ^ n24073 ;
  assign n24100 = n22656 ^ n21823 ;
  assign n24101 = n24100 ^ n22656 ;
  assign n24102 = n22657 & n24101 ;
  assign n24103 = n24102 ^ n22656 ;
  assign n24104 = n21536 & n24103 ;
  assign n24105 = n24097 & ~n24104 ;
  assign n24106 = ~n22612 & n24105 ;
  assign n24107 = n24106 ^ n22495 ;
  assign n24138 = n23420 ^ n22797 ;
  assign n24139 = n23146 & n24138 ;
  assign n24134 = n22863 ^ n22788 ;
  assign n24124 = n22806 ^ n22787 ;
  assign n24125 = n24124 ^ n22834 ;
  assign n24126 = n22834 ^ n22788 ;
  assign n24127 = n23136 & ~n24126 ;
  assign n24128 = n24127 ^ n22788 ;
  assign n24129 = n24125 & ~n24128 ;
  assign n24130 = n24129 ^ n22834 ;
  assign n24131 = n24130 ^ n22786 ;
  assign n24135 = n24134 ^ n24131 ;
  assign n24136 = n24135 ^ n23169 ;
  assign n24116 = n22785 ^ n22776 ;
  assign n24117 = n24116 ^ n22777 ;
  assign n24118 = n24117 ^ n22785 ;
  assign n24121 = n22793 & n24118 ;
  assign n24122 = n24121 ^ n22785 ;
  assign n24123 = ~n22745 & ~n24122 ;
  assign n24132 = n24131 ^ n24123 ;
  assign n24133 = n23136 & ~n24132 ;
  assign n24137 = n24136 ^ n24133 ;
  assign n24140 = n24139 ^ n24137 ;
  assign n24115 = n22789 & n22830 ;
  assign n24141 = n24140 ^ n24115 ;
  assign n24108 = n23147 ^ n22811 ;
  assign n24109 = n22808 ^ n22789 ;
  assign n24112 = ~n23147 & ~n24109 ;
  assign n24113 = n24112 ^ n22789 ;
  assign n24114 = ~n24108 & n24113 ;
  assign n24142 = n24141 ^ n24114 ;
  assign n24143 = ~n23435 & n24142 ;
  assign n24144 = ~n23168 & n24143 ;
  assign n24145 = n24144 ^ n19768 ;
  assign n24155 = n23377 ^ n23341 ;
  assign n24147 = n23330 ^ n23294 ;
  assign n24148 = n24147 ^ n23288 ;
  assign n24149 = n24148 ^ n23294 ;
  assign n24152 = ~n23350 & ~n24149 ;
  assign n24153 = n24152 ^ n23294 ;
  assign n24154 = ~n23177 & n24153 ;
  assign n24156 = n24155 ^ n24154 ;
  assign n24157 = n23206 & ~n24156 ;
  assign n24165 = n23359 ^ n23206 ;
  assign n24167 = n23362 ^ n23338 ;
  assign n24170 = n24167 ^ n23359 ;
  assign n24166 = n23371 ^ n23342 ;
  assign n24168 = n24167 ^ n24166 ;
  assign n24169 = n23177 & ~n24168 ;
  assign n24171 = n24170 ^ n24169 ;
  assign n24172 = n24165 & n24171 ;
  assign n24173 = n24172 ^ n23206 ;
  assign n24164 = n23358 & n23398 ;
  assign n24174 = n24173 ^ n24164 ;
  assign n24158 = n23370 ^ n23347 ;
  assign n24159 = n23347 ^ n23177 ;
  assign n24160 = n24159 ^ n23347 ;
  assign n24161 = n24158 & ~n24160 ;
  assign n24162 = n24161 ^ n23347 ;
  assign n24163 = n23206 & ~n24162 ;
  assign n24175 = n24174 ^ n24163 ;
  assign n24176 = ~n23449 & n24175 ;
  assign n24177 = ~n23475 & n24176 ;
  assign n24178 = ~n24157 & n24177 ;
  assign n24179 = ~n23446 & n24178 ;
  assign n24180 = ~n23413 & n24179 ;
  assign n24183 = n24180 ^ n21906 ;
  assign n24146 = n23457 ^ n23347 ;
  assign n24181 = ~n23209 & n24180 ;
  assign n24182 = ~n24146 & n24181 ;
  assign n24184 = n24183 ^ n24182 ;
  assign n24193 = n24024 ^ n23014 ;
  assign n24194 = n24193 ^ n23007 ;
  assign n24196 = ~n23020 & ~n24194 ;
  assign n24197 = n24196 ^ n23007 ;
  assign n24199 = n23100 ^ n23005 ;
  assign n24198 = n23100 ^ n23020 ;
  assign n24200 = n24199 ^ n24198 ;
  assign n24201 = n24197 & n24200 ;
  assign n24202 = n24201 ^ n24199 ;
  assign n24203 = n24202 ^ n23052 ;
  assign n24189 = n23100 ^ n22994 ;
  assign n24186 = n23038 ^ n23010 ;
  assign n24190 = n24189 ^ n24186 ;
  assign n24185 = n24018 ^ n23012 ;
  assign n24187 = n24186 ^ n24185 ;
  assign n24188 = ~n22744 & n24187 ;
  assign n24191 = n24190 ^ n24188 ;
  assign n24192 = ~n23004 & n24191 ;
  assign n24204 = n24203 ^ n24192 ;
  assign n24205 = n24204 ^ n23122 ;
  assign n24206 = n24205 ^ n23062 ;
  assign n24207 = n24206 ^ n23126 ;
  assign n24208 = n24207 ^ n23018 ;
  assign n24209 = ~n22996 & ~n24208 ;
  assign n24210 = n24209 ^ n21641 ;
  assign n24211 = n23620 & n23639 ;
  assign n24226 = n23649 ^ n23644 ;
  assign n24235 = n24226 ^ n23640 ;
  assign n24236 = n24235 ^ n23607 ;
  assign n24237 = n24236 ^ n23644 ;
  assign n24233 = n24226 ^ n23665 ;
  assign n24220 = n23663 ^ n23647 ;
  assign n24221 = n24220 ^ n23667 ;
  assign n24227 = n24226 ^ n24221 ;
  assign n24229 = n24221 ^ n23528 ;
  assign n24230 = n23622 & ~n24229 ;
  assign n24231 = n24230 ^ n23528 ;
  assign n24232 = n24227 & n24231 ;
  assign n24234 = n24233 ^ n24232 ;
  assign n24238 = n24237 ^ n24234 ;
  assign n24239 = n24238 ^ n23613 ;
  assign n24240 = n24239 ^ n24234 ;
  assign n24241 = n24234 ^ n23528 ;
  assign n24242 = n24241 ^ n24234 ;
  assign n24243 = ~n24240 & n24242 ;
  assign n24244 = n24243 ^ n24234 ;
  assign n24245 = n23622 & n24244 ;
  assign n24246 = n24245 ^ n24234 ;
  assign n24212 = n23622 ^ n23528 ;
  assign n24225 = n23611 & n24212 ;
  assign n24247 = n24246 ^ n24225 ;
  assign n24222 = n24221 ^ n23644 ;
  assign n24223 = n23637 & n24222 ;
  assign n24219 = n23615 & n23685 ;
  assign n24224 = n24223 ^ n24219 ;
  assign n24248 = n24247 ^ n24224 ;
  assign n24249 = n24248 ^ n23653 ;
  assign n24250 = n24249 ^ n23635 ;
  assign n24213 = n23668 ^ n23612 ;
  assign n24216 = n23622 & n24213 ;
  assign n24217 = n24216 ^ n23612 ;
  assign n24218 = ~n24212 & n24217 ;
  assign n24251 = n24250 ^ n24218 ;
  assign n24252 = ~n24211 & ~n24251 ;
  assign n24253 = n24252 ^ n22144 ;
  assign n24254 = n22960 ^ x113 ;
  assign n24255 = n23850 ^ x104 ;
  assign n24256 = n24254 & ~n24255 ;
  assign n24257 = n24256 ^ n24254 ;
  assign n24258 = n24257 ^ n24255 ;
  assign n24259 = n24258 ^ n24254 ;
  assign n24260 = n23444 ^ x80 ;
  assign n24261 = n20981 ^ x90 ;
  assign n24262 = n24260 & ~n24261 ;
  assign n24263 = n24262 ^ n24261 ;
  assign n24269 = n24263 ^ n24260 ;
  assign n24270 = n24269 ^ n24261 ;
  assign n24264 = n23755 ^ x99 ;
  assign n24265 = n24014 ^ x73 ;
  assign n24266 = n24264 & ~n24265 ;
  assign n24273 = n24266 ^ n24265 ;
  assign n24284 = n24270 & ~n24273 ;
  assign n24274 = n24273 ^ n24264 ;
  assign n24275 = ~n24263 & n24274 ;
  assign n24288 = n24284 ^ n24275 ;
  assign n24287 = n24262 & n24274 ;
  assign n24289 = n24288 ^ n24287 ;
  assign n24286 = n24270 & n24274 ;
  assign n24290 = n24289 ^ n24286 ;
  assign n24285 = n24284 ^ n24274 ;
  assign n24291 = n24290 ^ n24285 ;
  assign n24292 = n24291 ^ n24269 ;
  assign n24282 = n24269 & ~n24273 ;
  assign n24281 = n24266 & n24269 ;
  assign n24283 = n24282 ^ n24281 ;
  assign n24293 = n24292 ^ n24283 ;
  assign n24278 = ~n24260 & n24264 ;
  assign n24271 = n24266 & n24270 ;
  assign n24267 = n24266 ^ n24264 ;
  assign n24268 = ~n24263 & n24267 ;
  assign n24272 = n24271 ^ n24268 ;
  assign n24279 = n24278 ^ n24272 ;
  assign n24280 = n24279 ^ n24266 ;
  assign n24294 = n24293 ^ n24280 ;
  assign n24295 = n24294 ^ n24281 ;
  assign n24277 = n24271 ^ n24266 ;
  assign n24296 = n24295 ^ n24277 ;
  assign n24297 = n24296 ^ n24271 ;
  assign n24298 = n24297 ^ n24263 ;
  assign n24276 = n24275 ^ n24272 ;
  assign n24299 = n24298 ^ n24276 ;
  assign n24300 = n24299 ^ n24286 ;
  assign n24301 = ~n24259 & ~n24300 ;
  assign n24353 = n24296 ^ n24293 ;
  assign n24360 = n24353 ^ n24294 ;
  assign n24361 = n24258 & n24360 ;
  assign n24338 = n24255 ^ n24254 ;
  assign n24308 = n24299 ^ n24284 ;
  assign n24354 = n24353 ^ n24308 ;
  assign n24355 = n24353 ^ n24255 ;
  assign n24356 = n24355 ^ n24353 ;
  assign n24357 = ~n24354 & n24356 ;
  assign n24358 = n24357 ^ n24353 ;
  assign n24359 = n24338 & n24358 ;
  assign n24362 = n24361 ^ n24359 ;
  assign n24307 = n24282 ^ n24273 ;
  assign n24309 = n24308 ^ n24307 ;
  assign n24310 = n24309 ^ n24291 ;
  assign n24311 = n24310 ^ n24276 ;
  assign n24304 = n24294 ^ n24268 ;
  assign n24303 = n24267 & n24270 ;
  assign n24305 = n24304 ^ n24303 ;
  assign n24306 = n24305 ^ n24291 ;
  assign n24312 = n24311 ^ n24306 ;
  assign n24302 = n24290 ^ n24260 ;
  assign n24313 = n24312 ^ n24302 ;
  assign n24314 = n24257 & n24313 ;
  assign n24324 = ~n24259 & n24304 ;
  assign n24322 = n24281 ^ n24275 ;
  assign n24323 = n24322 ^ n24271 ;
  assign n24325 = n24324 ^ n24323 ;
  assign n24326 = n24325 ^ n24257 ;
  assign n24327 = n24300 ^ n24294 ;
  assign n24328 = n24327 ^ n24259 ;
  assign n24331 = ~n24325 & ~n24328 ;
  assign n24332 = n24331 ^ n24259 ;
  assign n24333 = n24326 & ~n24332 ;
  assign n24334 = n24333 ^ n24257 ;
  assign n24320 = n24303 ^ n24287 ;
  assign n24321 = n24258 & n24320 ;
  assign n24335 = n24334 ^ n24321 ;
  assign n24316 = n24282 ^ n24275 ;
  assign n24317 = n24316 ^ n24286 ;
  assign n24315 = n24313 ^ n24309 ;
  assign n24318 = n24317 ^ n24315 ;
  assign n24319 = n24256 & n24318 ;
  assign n24336 = n24335 ^ n24319 ;
  assign n24337 = ~n24314 & ~n24336 ;
  assign n24339 = n24284 ^ n24282 ;
  assign n24340 = n24284 ^ n24255 ;
  assign n24341 = n24340 ^ n24284 ;
  assign n24342 = n24339 & n24341 ;
  assign n24343 = n24342 ^ n24284 ;
  assign n24344 = ~n24338 & n24343 ;
  assign n24345 = n24337 & ~n24344 ;
  assign n24346 = n24303 ^ n24291 ;
  assign n24347 = n24291 ^ n24255 ;
  assign n24348 = n24347 ^ n24291 ;
  assign n24349 = n24346 & ~n24348 ;
  assign n24350 = n24349 ^ n24291 ;
  assign n24351 = n24338 & n24350 ;
  assign n24352 = n24345 & ~n24351 ;
  assign n24363 = n24362 ^ n24352 ;
  assign n24364 = ~n24301 & n24363 ;
  assign n24365 = n24364 ^ n21195 ;
  assign n24387 = ~n23615 & ~n23637 ;
  assign n24388 = n24221 & n24387 ;
  assign n24384 = n23648 ^ n23610 ;
  assign n24385 = n24384 ^ n24221 ;
  assign n24375 = n24237 ^ n23648 ;
  assign n24376 = n24375 ^ n23658 ;
  assign n24377 = ~n23622 & ~n24376 ;
  assign n24378 = n24377 ^ n23661 ;
  assign n24383 = n24378 ^ n23607 ;
  assign n24386 = n24385 ^ n24383 ;
  assign n24389 = n24388 ^ n24386 ;
  assign n24381 = n23616 ^ n23607 ;
  assign n24382 = n23622 & n24381 ;
  assign n24390 = n24389 ^ n24382 ;
  assign n24391 = n24212 & ~n24390 ;
  assign n24374 = n23655 ^ n23610 ;
  assign n24379 = n24378 ^ n24374 ;
  assign n24370 = n23619 ^ n23612 ;
  assign n24371 = ~n23622 & n24370 ;
  assign n24372 = n24371 ^ n23612 ;
  assign n24373 = ~n23528 & n24372 ;
  assign n24380 = n24379 ^ n24373 ;
  assign n24392 = n24391 ^ n24380 ;
  assign n24393 = n24392 ^ n24211 ;
  assign n24394 = n24393 ^ n23669 ;
  assign n24395 = n24394 ^ n19335 ;
  assign n24366 = n24235 ^ n24220 ;
  assign n24367 = ~n23622 & n24366 ;
  assign n24368 = n24367 ^ n24220 ;
  assign n24369 = n23528 & n24368 ;
  assign n24396 = n24395 ^ n24369 ;
  assign n24397 = n22596 ^ x118 ;
  assign n24398 = n23287 ^ x100 ;
  assign n24471 = n24397 & ~n24398 ;
  assign n24472 = n24471 ^ n24397 ;
  assign n24403 = n23096 ^ x94 ;
  assign n24404 = n21822 ^ x101 ;
  assign n24405 = n24403 & ~n24404 ;
  assign n24406 = n24405 ^ n24403 ;
  assign n24407 = n24406 ^ n24404 ;
  assign n24400 = n23725 ^ x124 ;
  assign n24401 = n24145 ^ x76 ;
  assign n24402 = ~n24400 & n24401 ;
  assign n24425 = n24402 ^ n24400 ;
  assign n24426 = n24407 & ~n24425 ;
  assign n24420 = n24402 & n24406 ;
  assign n24496 = n24426 ^ n24420 ;
  assign n24497 = n24472 & n24496 ;
  assign n24399 = n24398 ^ n24397 ;
  assign n24409 = n24402 ^ n24401 ;
  assign n24422 = n24407 & n24409 ;
  assign n24483 = n24422 ^ n24406 ;
  assign n24410 = n24409 ^ n24400 ;
  assign n24411 = n24406 & n24410 ;
  assign n24427 = n24426 ^ n24411 ;
  assign n24408 = n24402 & n24407 ;
  assign n24428 = n24427 ^ n24408 ;
  assign n24419 = n24400 & n24404 ;
  assign n24424 = n24419 ^ n24407 ;
  assign n24429 = n24428 ^ n24424 ;
  assign n24423 = n24422 ^ n24420 ;
  assign n24430 = n24429 ^ n24423 ;
  assign n24431 = n24430 ^ n24411 ;
  assign n24484 = n24483 ^ n24431 ;
  assign n24421 = n24420 ^ n24419 ;
  assign n24432 = n24431 ^ n24421 ;
  assign n24433 = n24432 ^ n24429 ;
  assign n24485 = n24484 ^ n24433 ;
  assign n24486 = n24485 ^ n24397 ;
  assign n24487 = n24486 ^ n24485 ;
  assign n24435 = n24407 ^ n24403 ;
  assign n24439 = n24409 & ~n24435 ;
  assign n24438 = n24402 & ~n24435 ;
  assign n24440 = n24439 ^ n24438 ;
  assign n24436 = n24410 & ~n24435 ;
  assign n24437 = n24436 ^ n24435 ;
  assign n24441 = n24440 ^ n24437 ;
  assign n24488 = n24484 ^ n24441 ;
  assign n24489 = n24488 ^ n24485 ;
  assign n24490 = ~n24487 & ~n24489 ;
  assign n24491 = n24490 ^ n24485 ;
  assign n24492 = ~n24399 & n24491 ;
  assign n24493 = n24492 ^ n24484 ;
  assign n24494 = n24493 ^ n21600 ;
  assign n24452 = n24429 ^ n24422 ;
  assign n24451 = n24439 ^ n24409 ;
  assign n24453 = n24452 ^ n24451 ;
  assign n24454 = n24453 ^ n24436 ;
  assign n24456 = n24453 ^ n24438 ;
  assign n24455 = n24405 & ~n24425 ;
  assign n24457 = n24456 ^ n24455 ;
  assign n24458 = n24398 & ~n24457 ;
  assign n24459 = n24458 ^ n24457 ;
  assign n24460 = n24459 ^ n24397 ;
  assign n24461 = n24460 ^ n24459 ;
  assign n24464 = n24459 ^ n24439 ;
  assign n24465 = n24464 ^ n24459 ;
  assign n24466 = n24458 & ~n24465 ;
  assign n24467 = ~n24461 & n24466 ;
  assign n24468 = n24467 ^ n24461 ;
  assign n24469 = n24468 ^ n24460 ;
  assign n24470 = ~n24454 & ~n24469 ;
  assign n24473 = n24472 ^ n24398 ;
  assign n24474 = n24456 & n24472 ;
  assign n24475 = n24474 ^ n24439 ;
  assign n24443 = n24405 & n24410 ;
  assign n24476 = n24475 ^ n24443 ;
  assign n24477 = ~n24473 & ~n24476 ;
  assign n24478 = n24477 ^ n24397 ;
  assign n24479 = n24399 ^ n24397 ;
  assign n24480 = ~n24478 & n24479 ;
  assign n24481 = n24480 ^ n24397 ;
  assign n24482 = ~n24470 & n24481 ;
  assign n24495 = n24494 ^ n24482 ;
  assign n24498 = n24497 ^ n24495 ;
  assign n24444 = n24443 ^ n24441 ;
  assign n24445 = n24444 ^ n24438 ;
  assign n24446 = n24445 ^ n24402 ;
  assign n24434 = n24433 ^ n24420 ;
  assign n24442 = n24441 ^ n24434 ;
  assign n24447 = n24446 ^ n24442 ;
  assign n24448 = ~n24397 & n24447 ;
  assign n24449 = n24448 ^ n24423 ;
  assign n24450 = ~n24398 & n24449 ;
  assign n24499 = n24498 ^ n24450 ;
  assign n24412 = n24411 ^ n24408 ;
  assign n24413 = n24412 ^ n24411 ;
  assign n24414 = n24411 ^ n24397 ;
  assign n24415 = n24414 ^ n24411 ;
  assign n24416 = n24413 & ~n24415 ;
  assign n24417 = n24416 ^ n24411 ;
  assign n24418 = n24399 & n24417 ;
  assign n24500 = n24499 ^ n24418 ;
  assign n24536 = n24452 & n24471 ;
  assign n24532 = n24477 ^ n24455 ;
  assign n24512 = n24474 ^ n24399 ;
  assign n24514 = n24402 & n24405 ;
  assign n24515 = n24514 ^ n24436 ;
  assign n24513 = n24475 ^ n24411 ;
  assign n24516 = n24515 ^ n24513 ;
  assign n24517 = ~n24471 & ~n24516 ;
  assign n24518 = n24512 & ~n24517 ;
  assign n24533 = ~n24436 & n24518 ;
  assign n24534 = n24532 & n24533 ;
  assign n24529 = n24493 ^ n24426 ;
  assign n24527 = n24420 & n24473 ;
  assign n24519 = n24441 ^ n24411 ;
  assign n24520 = n24519 ^ n24442 ;
  assign n24521 = n24520 ^ n24519 ;
  assign n24522 = n24519 ^ n24397 ;
  assign n24523 = n24522 ^ n24519 ;
  assign n24524 = ~n24521 & ~n24523 ;
  assign n24525 = n24524 ^ n24519 ;
  assign n24526 = ~n24399 & ~n24525 ;
  assign n24528 = n24527 ^ n24526 ;
  assign n24530 = n24529 ^ n24528 ;
  assign n24531 = n24530 ^ n24518 ;
  assign n24535 = n24534 ^ n24531 ;
  assign n24537 = n24536 ^ n24535 ;
  assign n24504 = n24484 ^ n24408 ;
  assign n24505 = n24504 ^ n24426 ;
  assign n24502 = n24457 ^ n24426 ;
  assign n24506 = n24505 ^ n24502 ;
  assign n24507 = n24502 ^ n24398 ;
  assign n24508 = n24507 ^ n24502 ;
  assign n24509 = n24506 & n24508 ;
  assign n24510 = n24509 ^ n24502 ;
  assign n24511 = ~n24399 & n24510 ;
  assign n24538 = n24537 ^ n24511 ;
  assign n24501 = n24422 & n24473 ;
  assign n24539 = n24538 ^ n24501 ;
  assign n24540 = n24539 ^ n22101 ;
  assign n24551 = n23376 ^ n23340 ;
  assign n24549 = n23368 ^ n23334 ;
  assign n24552 = n24551 ^ n24549 ;
  assign n24553 = ~n23206 & ~n24552 ;
  assign n24542 = n23376 ^ n23374 ;
  assign n24543 = n24542 ^ n23351 ;
  assign n24544 = ~n23206 & n24543 ;
  assign n24545 = n24544 ^ n23379 ;
  assign n24548 = n24545 ^ n23362 ;
  assign n24550 = n24549 ^ n24548 ;
  assign n24554 = n24553 ^ n24550 ;
  assign n24555 = ~n23447 & ~n24554 ;
  assign n24541 = n23445 ^ n23349 ;
  assign n24546 = n24545 ^ n24541 ;
  assign n24547 = n24546 ^ n23413 ;
  assign n24556 = n24555 ^ n24547 ;
  assign n24557 = ~n23475 & n24556 ;
  assign n24558 = n24557 ^ n21339 ;
  assign n24599 = n22466 ^ x112 ;
  assign n24559 = n22869 ^ x65 ;
  assign n24563 = n22743 ^ x72 ;
  assign n24561 = n21535 ^ x89 ;
  assign n24601 = n24563 ^ n24561 ;
  assign n24560 = n23515 ^ x98 ;
  assign n24568 = ~n24560 & ~n24563 ;
  assign n24575 = n24568 ^ n24560 ;
  assign n24573 = n24067 ^ x107 ;
  assign n24577 = n24573 ^ n24563 ;
  assign n24578 = n24575 & n24577 ;
  assign n24590 = n24561 & n24578 ;
  assign n24612 = n24590 ^ n24561 ;
  assign n24566 = n24560 & n24561 ;
  assign n24567 = n24563 & ~n24566 ;
  assign n24569 = n24568 ^ n24567 ;
  assign n24570 = n24569 ^ n24566 ;
  assign n24564 = n24563 ^ n24560 ;
  assign n24565 = ~n24561 & n24564 ;
  assign n24571 = n24570 ^ n24565 ;
  assign n24586 = n24575 ^ n24571 ;
  assign n24587 = ~n24573 & n24586 ;
  assign n24611 = n24587 ^ n24566 ;
  assign n24613 = n24612 ^ n24611 ;
  assign n24604 = ~n24573 & ~n24601 ;
  assign n24605 = n24604 ^ n24561 ;
  assign n24606 = n24560 & ~n24605 ;
  assign n24603 = n24577 ^ n24561 ;
  assign n24607 = n24606 ^ n24603 ;
  assign n24602 = n24573 ^ n24564 ;
  assign n24608 = n24607 ^ n24602 ;
  assign n24609 = n24608 ^ n24564 ;
  assign n24610 = n24609 ^ n24607 ;
  assign n24614 = n24613 ^ n24610 ;
  assign n24615 = ~n24601 & ~n24614 ;
  assign n24616 = n24615 ^ n24608 ;
  assign n24617 = ~n24559 & ~n24616 ;
  assign n24618 = n24617 ^ n24607 ;
  assign n24582 = n24570 ^ n24561 ;
  assign n24591 = n24590 ^ n24582 ;
  assign n24588 = n24587 ^ n24571 ;
  assign n24579 = n24578 ^ n24577 ;
  assign n24589 = n24588 ^ n24579 ;
  assign n24592 = n24591 ^ n24589 ;
  assign n24574 = n24563 & n24573 ;
  assign n24576 = n24575 ^ n24574 ;
  assign n24580 = n24579 ^ n24576 ;
  assign n24581 = n24580 ^ n24578 ;
  assign n24583 = n24582 ^ n24581 ;
  assign n24593 = n24592 ^ n24583 ;
  assign n24594 = n24593 ^ n24582 ;
  assign n24595 = n24594 ^ n24564 ;
  assign n24572 = n24571 ^ n24567 ;
  assign n24584 = n24583 ^ n24572 ;
  assign n24562 = n24561 ^ n24560 ;
  assign n24585 = n24584 ^ n24562 ;
  assign n24596 = n24595 ^ n24585 ;
  assign n24597 = n24559 & ~n24596 ;
  assign n24598 = n24597 ^ n24595 ;
  assign n24619 = n24618 ^ n24598 ;
  assign n24620 = n24599 & ~n24619 ;
  assign n24621 = n24620 ^ n24618 ;
  assign n24600 = n24599 ^ n24598 ;
  assign n24622 = n24621 ^ n24600 ;
  assign n24623 = n24622 ^ n24618 ;
  assign n24624 = n24623 ^ n20545 ;
  assign n24650 = n24293 ^ n24275 ;
  assign n24651 = n24650 ^ n24294 ;
  assign n24652 = n24651 ^ n24313 ;
  assign n24653 = ~n24254 & n24652 ;
  assign n24654 = n24653 ^ n24283 ;
  assign n24655 = n24255 & n24654 ;
  assign n24637 = n24303 ^ n24257 ;
  assign n24638 = n24294 ^ n24259 ;
  assign n24641 = ~n24303 & n24638 ;
  assign n24642 = n24641 ^ n24259 ;
  assign n24643 = n24637 & ~n24642 ;
  assign n24644 = n24643 ^ n24257 ;
  assign n24626 = n24310 ^ n24268 ;
  assign n24645 = n24644 ^ n24626 ;
  assign n24646 = n24645 ^ n24359 ;
  assign n24635 = n24256 & ~n24300 ;
  assign n24636 = n24635 ^ n24314 ;
  assign n24647 = n24646 ^ n24636 ;
  assign n24627 = n24626 ^ n24271 ;
  assign n24628 = n24627 ^ n24289 ;
  assign n24629 = n24628 ^ n24626 ;
  assign n24630 = n24626 ^ n24255 ;
  assign n24631 = n24630 ^ n24626 ;
  assign n24632 = n24629 & ~n24631 ;
  assign n24633 = n24632 ^ n24626 ;
  assign n24634 = n24338 & n24633 ;
  assign n24648 = n24647 ^ n24634 ;
  assign n24625 = ~n24259 & n24297 ;
  assign n24649 = n24648 ^ n24625 ;
  assign n24656 = n24655 ^ n24649 ;
  assign n24657 = n24656 ^ n24301 ;
  assign n24658 = n24657 ^ n21562 ;
  assign n24687 = n24080 ^ n22643 ;
  assign n24688 = ~n22652 & n24687 ;
  assign n24669 = n22621 ^ n22601 ;
  assign n24670 = n24669 ^ n22643 ;
  assign n24668 = n22676 ^ n22622 ;
  assign n24671 = n24670 ^ n24668 ;
  assign n24672 = n21536 & ~n24671 ;
  assign n24673 = n24672 ^ n24670 ;
  assign n24681 = n24673 ^ n22706 ;
  assign n24682 = n24681 ^ n22675 ;
  assign n24683 = n24682 ^ n22612 ;
  assign n24684 = n24683 ^ n22340 ;
  assign n24674 = n24673 ^ n22667 ;
  assign n24675 = n24674 ^ n22633 ;
  assign n24676 = n24675 ^ n22639 ;
  assign n24677 = n24676 ^ n24673 ;
  assign n24678 = ~n21536 & n24677 ;
  assign n24679 = n24678 ^ n24674 ;
  assign n24680 = n21824 & n24679 ;
  assign n24685 = n24684 ^ n24680 ;
  assign n24667 = ~n22651 & n22653 ;
  assign n24686 = n24685 ^ n24667 ;
  assign n24689 = n24688 ^ n24686 ;
  assign n24666 = ~n21824 & n22637 ;
  assign n24690 = n24689 ^ n24666 ;
  assign n24659 = n22638 ^ n22602 ;
  assign n24660 = n24659 ^ n22655 ;
  assign n24661 = n22655 ^ n21536 ;
  assign n24662 = n24661 ^ n22655 ;
  assign n24663 = n24660 & n24662 ;
  assign n24664 = n24663 ^ n22655 ;
  assign n24665 = ~n21823 & n24664 ;
  assign n24691 = n24690 ^ n24665 ;
  assign n24708 = n24514 ^ n24429 ;
  assign n24706 = n24432 ^ n24427 ;
  assign n24707 = n24471 & n24706 ;
  assign n24709 = n24708 ^ n24707 ;
  assign n24710 = n24709 ^ n24455 ;
  assign n24705 = n24473 & n24504 ;
  assign n24711 = n24710 ^ n24705 ;
  assign n24715 = n24711 ^ n24501 ;
  assign n24694 = n24439 ^ n24398 ;
  assign n24695 = n24694 ^ n24439 ;
  assign n24696 = n24440 & ~n24695 ;
  assign n24697 = n24696 ^ n24439 ;
  assign n24698 = n24399 & n24697 ;
  assign n24716 = n24715 ^ n24698 ;
  assign n24704 = n24454 ^ n24444 ;
  assign n24712 = n24711 ^ n24704 ;
  assign n24700 = n24428 ^ n24420 ;
  assign n24701 = n24700 ^ n24454 ;
  assign n24702 = n24701 ^ n24444 ;
  assign n24703 = n24398 & ~n24702 ;
  assign n24713 = n24712 ^ n24703 ;
  assign n24714 = ~n24399 & ~n24713 ;
  assign n24717 = n24716 ^ n24714 ;
  assign n24699 = n24397 & n24436 ;
  assign n24718 = n24717 ^ n24699 ;
  assign n24719 = n24718 ^ n24698 ;
  assign n24720 = n24473 ^ n24397 ;
  assign n24721 = n24427 & ~n24720 ;
  assign n24722 = ~n24719 & n24721 ;
  assign n24723 = n24722 ^ n24718 ;
  assign n24724 = n24441 ^ n24423 ;
  assign n24725 = n24398 & ~n24724 ;
  assign n24726 = n24725 ^ n24423 ;
  assign n24729 = n24726 ^ n24455 ;
  assign n24730 = n24729 ^ n24726 ;
  assign n24731 = n24398 & n24730 ;
  assign n24732 = n24731 ^ n24726 ;
  assign n24733 = n24397 & n24732 ;
  assign n24734 = n24733 ^ n24726 ;
  assign n24735 = ~n24723 & ~n24734 ;
  assign n24736 = ~n24474 & n24735 ;
  assign n24737 = n24736 ^ n21448 ;
  assign n24741 = n24456 ^ n24431 ;
  assign n24742 = n24741 ^ n24515 ;
  assign n24743 = ~n24398 & n24742 ;
  assign n24744 = n24743 ^ n24431 ;
  assign n24752 = n24744 ^ n24501 ;
  assign n24748 = n24514 ^ n24439 ;
  assign n24749 = ~n24398 & n24748 ;
  assign n24746 = n24427 & n24471 ;
  assign n24740 = n24527 ^ n24504 ;
  assign n24745 = n24744 ^ n24740 ;
  assign n24747 = n24746 ^ n24745 ;
  assign n24750 = n24749 ^ n24747 ;
  assign n24751 = n24399 & n24750 ;
  assign n24753 = n24752 ^ n24751 ;
  assign n24739 = ~n24445 & n24472 ;
  assign n24754 = n24753 ^ n24739 ;
  assign n24755 = ~n24397 & ~n24754 ;
  assign n24756 = n24432 ^ n24398 ;
  assign n24757 = n24756 ^ n24432 ;
  assign n24760 = n24484 & ~n24757 ;
  assign n24761 = n24760 ^ n24432 ;
  assign n24762 = n24755 & n24761 ;
  assign n24763 = n24762 ^ n24754 ;
  assign n24764 = ~n24734 & ~n24763 ;
  assign n24765 = n24764 ^ n19947 ;
  assign n24738 = n24399 & n24454 ;
  assign n24768 = n24765 ^ n24738 ;
  assign n24769 = n23667 ^ n23618 ;
  assign n24786 = n24769 ^ n23627 ;
  assign n24787 = n24786 ^ n24368 ;
  assign n24788 = n24787 ^ n24218 ;
  assign n24789 = n24788 ^ n24373 ;
  assign n24779 = n24368 ^ n24222 ;
  assign n24778 = n24375 ^ n24368 ;
  assign n24780 = n24779 ^ n24778 ;
  assign n24781 = n24779 ^ n23622 ;
  assign n24782 = n24781 ^ n24779 ;
  assign n24783 = n24780 & n24782 ;
  assign n24784 = n24783 ^ n24779 ;
  assign n24785 = ~n23528 & n24784 ;
  assign n24790 = n24789 ^ n24785 ;
  assign n24770 = n24769 ^ n23614 ;
  assign n24771 = n24770 ^ n23616 ;
  assign n24772 = n24771 ^ n24769 ;
  assign n24773 = n24769 ^ n23622 ;
  assign n24774 = n24773 ^ n24769 ;
  assign n24775 = ~n24772 & n24774 ;
  assign n24776 = n24775 ^ n24769 ;
  assign n24777 = ~n24212 & n24776 ;
  assign n24791 = n24790 ^ n24777 ;
  assign n24792 = n24791 ^ n24211 ;
  assign n24793 = n24792 ^ n23669 ;
  assign n24794 = n24793 ^ n22775 ;
  assign n24808 = n24361 ^ n24287 ;
  assign n24809 = n24808 ^ n24361 ;
  assign n24810 = n24809 ^ n24271 ;
  assign n24811 = n24810 ^ n24809 ;
  assign n24812 = n24809 ^ n24255 ;
  assign n24813 = n24812 ^ n24809 ;
  assign n24814 = n24811 & n24813 ;
  assign n24815 = n24814 ^ n24809 ;
  assign n24816 = n24338 & n24815 ;
  assign n24817 = n24816 ^ n24808 ;
  assign n24818 = n24817 ^ n24636 ;
  assign n24805 = n24293 ^ n24272 ;
  assign n24806 = n24805 ^ n24309 ;
  assign n24807 = n24257 & n24806 ;
  assign n24819 = n24818 ^ n24807 ;
  assign n24804 = ~n24299 & ~n24338 ;
  assign n24820 = n24819 ^ n24804 ;
  assign n24799 = n24306 ^ n24254 ;
  assign n24800 = n24799 ^ n24306 ;
  assign n24801 = n24312 & n24800 ;
  assign n24802 = n24801 ^ n24306 ;
  assign n24803 = ~n24255 & n24802 ;
  assign n24821 = n24820 ^ n24803 ;
  assign n24796 = n24258 & n24317 ;
  assign n24822 = n24821 ^ n24796 ;
  assign n24823 = ~n24344 & ~n24822 ;
  assign n24824 = ~n24351 & n24823 ;
  assign n24825 = n24824 ^ n22381 ;
  assign n24795 = ~n24259 & n24282 ;
  assign n24828 = n24825 ^ n24795 ;
  assign n24838 = n24566 & n24574 ;
  assign n24836 = n24580 ^ n24569 ;
  assign n24835 = n24605 ^ n24589 ;
  assign n24837 = n24836 ^ n24835 ;
  assign n24839 = n24838 ^ n24837 ;
  assign n24829 = n24566 ^ n24561 ;
  assign n24832 = n24577 & ~n24829 ;
  assign n24833 = n24832 ^ n24566 ;
  assign n24834 = n24588 & ~n24833 ;
  assign n24840 = n24839 ^ n24834 ;
  assign n24841 = ~n24559 & n24840 ;
  assign n24842 = n24841 ^ n24839 ;
  assign n24845 = n24842 ^ n24592 ;
  assign n24844 = n24842 ^ n24583 ;
  assign n24846 = n24845 ^ n24844 ;
  assign n24849 = ~n24559 & ~n24846 ;
  assign n24850 = n24849 ^ n24845 ;
  assign n24851 = n24599 & n24850 ;
  assign n24843 = n24842 ^ n21397 ;
  assign n24852 = n24851 ^ n24843 ;
  assign n24862 = n24309 ^ n24255 ;
  assign n24863 = n24338 & n24862 ;
  assign n24864 = n24863 ^ n24255 ;
  assign n24867 = n24309 ^ n24289 ;
  assign n24868 = ~n24864 & n24867 ;
  assign n24865 = n24289 ^ n24282 ;
  assign n24869 = n24868 ^ n24865 ;
  assign n24880 = n24869 ^ n24644 ;
  assign n24874 = n24265 ^ n24260 ;
  assign n24875 = n24261 & ~n24874 ;
  assign n24872 = n24869 ^ n24290 ;
  assign n24870 = n24265 ^ n24264 ;
  assign n24871 = n24870 ^ n24869 ;
  assign n24873 = n24872 ^ n24871 ;
  assign n24876 = n24875 ^ n24873 ;
  assign n24877 = ~n24255 & n24876 ;
  assign n24878 = n24877 ^ n24872 ;
  assign n24879 = n24338 & n24878 ;
  assign n24881 = n24880 ^ n24879 ;
  assign n24860 = n24313 ^ n24295 ;
  assign n24861 = ~n24259 & n24860 ;
  assign n24882 = n24881 ^ n24861 ;
  assign n24855 = n24272 ^ n24254 ;
  assign n24856 = n24855 ^ n24272 ;
  assign n24857 = n24279 & ~n24856 ;
  assign n24858 = n24857 ^ n24272 ;
  assign n24859 = n24255 & n24858 ;
  assign n24883 = n24882 ^ n24859 ;
  assign n24884 = ~n24301 & ~n24883 ;
  assign n24885 = n24884 ^ n20319 ;
  assign n24886 = n24621 ^ n22783 ;
  assign n24888 = n24592 ^ n24564 ;
  assign n24889 = n24888 ^ n24616 ;
  assign n24891 = ~n24559 & ~n24599 ;
  assign n24892 = n24889 & n24891 ;
  assign n24887 = n24589 ^ n24583 ;
  assign n24890 = n24889 ^ n24887 ;
  assign n24893 = n24892 ^ n24890 ;
  assign n24894 = n24834 ^ n24591 ;
  assign n24895 = ~n24559 & n24894 ;
  assign n24896 = n24895 ^ n24591 ;
  assign n24897 = n24896 ^ n24599 ;
  assign n24898 = n24897 ^ n24559 ;
  assign n24899 = n24898 ^ n24896 ;
  assign n24900 = n24559 & ~n24839 ;
  assign n24901 = n24900 ^ n24896 ;
  assign n24902 = ~n24899 & ~n24901 ;
  assign n24903 = n24902 ^ n24896 ;
  assign n24904 = ~n24893 & ~n24903 ;
  assign n24905 = n24904 ^ n24893 ;
  assign n24906 = n24589 & ~n24905 ;
  assign n24907 = n24906 ^ n21571 ;
  assign n24948 = n23756 & n23874 ;
  assign n24941 = n23913 ^ n23856 ;
  assign n24942 = n24941 ^ n23944 ;
  assign n24936 = n23895 ^ n23858 ;
  assign n24937 = n24936 ^ n23884 ;
  assign n24938 = n24937 ^ n23869 ;
  assign n24943 = n24942 ^ n24938 ;
  assign n24944 = n23756 & n24943 ;
  assign n24925 = n23869 ^ n23855 ;
  assign n24926 = n24925 ^ n23902 ;
  assign n24927 = n24926 ^ n23880 ;
  assign n24924 = n23868 ^ n23859 ;
  assign n24928 = n24927 ^ n24924 ;
  assign n24929 = n23756 & ~n24928 ;
  assign n24930 = n24929 ^ n24927 ;
  assign n24939 = n24938 ^ n24930 ;
  assign n24945 = n24944 ^ n24939 ;
  assign n24946 = ~n23757 & ~n24945 ;
  assign n24931 = n24930 ^ n23957 ;
  assign n24920 = n23884 ^ n23880 ;
  assign n24921 = n23952 & n24920 ;
  assign n24922 = n24921 ^ n23880 ;
  assign n24923 = ~n23758 & n24922 ;
  assign n24932 = n24931 ^ n24923 ;
  assign n24933 = n24932 ^ n23966 ;
  assign n24914 = n23913 ^ n23895 ;
  assign n24915 = n23895 ^ n23757 ;
  assign n24916 = n24915 ^ n23895 ;
  assign n24917 = n24914 & ~n24916 ;
  assign n24918 = n24917 ^ n23895 ;
  assign n24919 = ~n23758 & n24918 ;
  assign n24934 = n24933 ^ n24919 ;
  assign n24908 = n23944 ^ n23868 ;
  assign n24909 = n23868 ^ n23757 ;
  assign n24910 = n24909 ^ n23868 ;
  assign n24911 = n24908 & n24910 ;
  assign n24912 = n24911 ^ n23868 ;
  assign n24913 = n23758 & n24912 ;
  assign n24935 = n24934 ^ n24913 ;
  assign n24947 = n24946 ^ n24935 ;
  assign n24949 = n24948 ^ n24947 ;
  assign n24950 = ~n23899 & n24949 ;
  assign n24951 = n24950 ^ n21372 ;
  assign n24977 = ~n23899 & n23974 ;
  assign n24972 = n23897 ^ n23880 ;
  assign n24973 = n24972 ^ n23913 ;
  assign n24974 = n24973 ^ n24926 ;
  assign n24975 = n23756 & ~n24974 ;
  assign n24969 = n24926 ^ n23896 ;
  assign n24970 = n23887 & ~n24969 ;
  assign n24961 = n23899 ^ n23868 ;
  assign n24962 = n24961 ^ n24919 ;
  assign n24958 = n24923 ^ n23869 ;
  assign n24957 = n24913 ^ n23865 ;
  assign n24959 = n24958 ^ n24957 ;
  assign n24956 = n24926 ^ n23897 ;
  assign n24960 = n24959 ^ n24956 ;
  assign n24963 = n24962 ^ n24960 ;
  assign n24964 = n24963 ^ n23937 ;
  assign n24965 = n24964 ^ n23890 ;
  assign n24966 = n24965 ^ n20723 ;
  assign n24954 = n23907 ^ n23855 ;
  assign n24955 = ~n23757 & ~n24954 ;
  assign n24967 = n24966 ^ n24955 ;
  assign n24952 = n24926 ^ n23868 ;
  assign n24953 = ~n23869 & ~n24952 ;
  assign n24968 = n24967 ^ n24953 ;
  assign n24971 = n24970 ^ n24968 ;
  assign n24976 = n24975 ^ n24971 ;
  assign n24978 = n24977 ^ n24976 ;
  assign n24994 = n24080 ^ n22634 ;
  assign n24991 = n22641 ^ n22622 ;
  assign n24992 = ~n21536 & n24991 ;
  assign n24993 = n24992 ^ n22662 ;
  assign n24995 = n24994 ^ n24993 ;
  assign n24987 = n22659 ^ n22634 ;
  assign n24988 = n24987 ^ n22654 ;
  assign n24989 = n24988 ^ n24080 ;
  assign n24990 = ~n21536 & ~n24989 ;
  assign n24996 = n24995 ^ n24990 ;
  assign n24997 = n21824 & ~n24996 ;
  assign n24998 = n24997 ^ n24993 ;
  assign n24986 = n22640 & n22649 ;
  assign n24999 = n24998 ^ n24986 ;
  assign n24985 = ~n22650 & n24094 ;
  assign n25000 = n24999 ^ n24985 ;
  assign n24979 = n22656 ^ n22622 ;
  assign n24980 = n22622 ^ n21536 ;
  assign n24981 = n24980 ^ n22622 ;
  assign n24982 = n24979 & n24981 ;
  assign n24983 = n24982 ^ n22622 ;
  assign n24984 = n21823 & n24983 ;
  assign n25001 = n25000 ^ n24984 ;
  assign n25002 = ~n24104 & ~n25001 ;
  assign n25003 = ~n22697 & n25002 ;
  assign n25004 = n25003 ^ n21996 ;
  assign y0 = ~n20981 ;
  assign y1 = ~n22709 ;
  assign y2 = n21535 ;
  assign y3 = ~n23073 ;
  assign y4 = ~n23096 ;
  assign y5 = ~n23135 ;
  assign y6 = ~n23176 ;
  assign y7 = n23415 ;
  assign y8 = n23444 ;
  assign y9 = n23477 ;
  assign y10 = ~n23515 ;
  assign y11 = ~n23687 ;
  assign y12 = ~n23725 ;
  assign y13 = n23934 ;
  assign y14 = n23601 ;
  assign y15 = ~n23976 ;
  assign y16 = ~n24014 ;
  assign y17 = n24046 ;
  assign y18 = n24067 ;
  assign y19 = ~n24107 ;
  assign y20 = n24145 ;
  assign y21 = ~n24184 ;
  assign y22 = n23561 ;
  assign y23 = ~n24210 ;
  assign y24 = ~n23755 ;
  assign y25 = n24253 ;
  assign y26 = n22743 ;
  assign y27 = n24365 ;
  assign y28 = n21822 ;
  assign y29 = n24396 ;
  assign y30 = ~n23205 ;
  assign y31 = n24500 ;
  assign y32 = n23850 ;
  assign y33 = n24540 ;
  assign y34 = n22869 ;
  assign y35 = n24558 ;
  assign y36 = n22596 ;
  assign y37 = n24624 ;
  assign y38 = ~n23329 ;
  assign y39 = ~n24658 ;
  assign y40 = n23810 ;
  assign y41 = ~n24691 ;
  assign y42 = ~n22913 ;
  assign y43 = ~n24737 ;
  assign y44 = n22069 ;
  assign y45 = n24768 ;
  assign y46 = ~n23254 ;
  assign y47 = n24794 ;
  assign y48 = n23780 ;
  assign y49 = n24828 ;
  assign y50 = ~n22985 ;
  assign y51 = n24852 ;
  assign y52 = n22298 ;
  assign y53 = ~n24885 ;
  assign y54 = ~n23293 ;
  assign y55 = ~n24886 ;
  assign y56 = n23527 ;
  assign y57 = n24907 ;
  assign y58 = n22960 ;
  assign y59 = ~n24951 ;
  assign y60 = n22466 ;
  assign y61 = ~n24978 ;
  assign y62 = ~n23287 ;
  assign y63 = ~n25004 ;
endmodule
