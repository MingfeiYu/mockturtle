module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n800 , n801 , n802 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n821 , n822 , n823 , n824 , n825 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n987 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1366 , n1367 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2178 , n2179 , n2180 , n2181 ;
  assign n257 = ~x129 & ~x130 ;
  assign n258 = x1 & n257 ;
  assign n259 = x2 & ~x3 ;
  assign n260 = ~x130 & n259 ;
  assign n261 = n260 ^ x3 ;
  assign n262 = n258 & ~n261 ;
  assign n263 = n262 ^ n261 ;
  assign n264 = ~x131 & ~x132 ;
  assign n265 = x4 & ~x5 ;
  assign n266 = ~x132 & n265 ;
  assign n267 = n266 ^ x5 ;
  assign n268 = n264 & ~n267 ;
  assign n269 = n263 & n268 ;
  assign n270 = n269 ^ n267 ;
  assign n271 = ~x252 & ~x253 ;
  assign n272 = ~x254 & n271 ;
  assign n273 = ~x221 & ~x222 ;
  assign n274 = ~x248 & ~x250 ;
  assign n275 = ~x249 & n274 ;
  assign n276 = ~x247 & ~x251 ;
  assign n277 = n275 & n276 ;
  assign n278 = ~x246 & n277 ;
  assign n279 = ~x245 & n278 ;
  assign n280 = ~x241 & ~x242 ;
  assign n281 = ~x240 & n280 ;
  assign n282 = ~x243 & n281 ;
  assign n283 = ~x244 & n282 ;
  assign n284 = n279 & n283 ;
  assign n285 = ~x238 & ~x239 ;
  assign n286 = n284 & n285 ;
  assign n287 = ~x235 & ~x237 ;
  assign n288 = ~x236 & n287 ;
  assign n289 = ~x229 & ~x230 ;
  assign n290 = ~x228 & n289 ;
  assign n291 = ~x231 & n290 ;
  assign n292 = ~x227 & ~x232 ;
  assign n293 = n291 & n292 ;
  assign n294 = ~x226 & ~x233 ;
  assign n295 = n293 & n294 ;
  assign n296 = ~x234 & n295 ;
  assign n297 = n288 & n296 ;
  assign n298 = n286 & n297 ;
  assign n299 = ~x224 & ~x225 ;
  assign n300 = ~x223 & n299 ;
  assign n301 = n298 & n300 ;
  assign n302 = n273 & n301 ;
  assign n303 = ~x216 & ~x217 ;
  assign n304 = ~x218 & n303 ;
  assign n305 = ~x219 & n304 ;
  assign n306 = ~x212 & ~x213 ;
  assign n307 = ~x214 & n306 ;
  assign n308 = ~x215 & n307 ;
  assign n309 = ~x209 & ~x210 ;
  assign n310 = ~x208 & n309 ;
  assign n311 = ~x211 & n310 ;
  assign n312 = n308 & n311 ;
  assign n313 = n305 & n312 ;
  assign n314 = ~x205 & ~x206 ;
  assign n315 = ~x207 & n314 ;
  assign n316 = ~x203 & ~x204 ;
  assign n317 = n315 & n316 ;
  assign n318 = ~x200 & ~x202 ;
  assign n319 = ~x201 & n318 ;
  assign n320 = n317 & n319 ;
  assign n321 = n313 & n320 ;
  assign n322 = ~x220 & n321 ;
  assign n323 = n302 & n322 ;
  assign n324 = ~x197 & ~x198 ;
  assign n325 = ~x196 & n324 ;
  assign n326 = ~x199 & n325 ;
  assign n327 = ~x193 & ~x194 ;
  assign n328 = ~x192 & n327 ;
  assign n329 = ~x195 & n328 ;
  assign n330 = n326 & n329 ;
  assign n331 = ~x188 & ~x189 ;
  assign n332 = ~x190 & n331 ;
  assign n333 = ~x191 & n332 ;
  assign n334 = ~x184 & ~x185 ;
  assign n335 = ~x186 & n334 ;
  assign n336 = ~x187 & n335 ;
  assign n337 = n333 & n336 ;
  assign n338 = n330 & n337 ;
  assign n339 = n323 & n338 ;
  assign n340 = ~x180 & ~x181 ;
  assign n341 = ~x182 & n340 ;
  assign n342 = ~x183 & n341 ;
  assign n343 = ~x176 & ~x178 ;
  assign n344 = ~x177 & n343 ;
  assign n345 = ~x179 & n344 ;
  assign n346 = n342 & n345 ;
  assign n347 = n339 & n346 ;
  assign n348 = n272 & n347 ;
  assign n349 = ~x173 & ~x174 ;
  assign n350 = ~x172 & n349 ;
  assign n351 = ~x171 & ~x175 ;
  assign n352 = n350 & n351 ;
  assign n353 = ~x170 & n352 ;
  assign n354 = ~x168 & ~x169 ;
  assign n355 = n353 & n354 ;
  assign n356 = n348 & n355 ;
  assign n357 = ~x165 & ~x166 ;
  assign n358 = ~x164 & n357 ;
  assign n359 = ~x167 & n358 ;
  assign n360 = n356 & n359 ;
  assign n361 = ~x161 & ~x162 ;
  assign n362 = ~x160 & n361 ;
  assign n363 = ~x163 & n362 ;
  assign n364 = n360 & n363 ;
  assign n365 = ~x157 & ~x158 ;
  assign n366 = ~x156 & n365 ;
  assign n367 = ~x159 & n366 ;
  assign n368 = n364 & n367 ;
  assign n369 = ~x154 & ~x155 ;
  assign n370 = n368 & n369 ;
  assign n371 = ~x153 & n370 ;
  assign n372 = ~x150 & ~x151 ;
  assign n373 = ~x149 & n372 ;
  assign n374 = ~x147 & ~x148 ;
  assign n375 = n373 & n374 ;
  assign n376 = ~x146 & ~x152 ;
  assign n377 = n375 & n376 ;
  assign n378 = n371 & n377 ;
  assign n379 = ~x142 & ~x144 ;
  assign n380 = ~x143 & n379 ;
  assign n381 = ~x145 & n380 ;
  assign n382 = ~x141 & n381 ;
  assign n383 = n378 & n382 ;
  assign n384 = ~x139 & ~x140 ;
  assign n385 = ~x138 & n384 ;
  assign n386 = n383 & n385 ;
  assign n387 = ~x134 & ~x135 ;
  assign n388 = ~x136 & n387 ;
  assign n389 = ~x133 & ~x137 ;
  assign n390 = n388 & n389 ;
  assign n391 = ~x255 & n390 ;
  assign n392 = n386 & n391 ;
  assign n393 = x14 & n381 ;
  assign n394 = ~x18 & ~x145 ;
  assign n395 = ~x16 & ~x144 ;
  assign n403 = x15 & n395 ;
  assign n404 = ~x143 & n403 ;
  assign n405 = n404 ^ x143 ;
  assign n396 = n395 ^ x144 ;
  assign n397 = n396 ^ x143 ;
  assign n406 = n405 ^ n397 ;
  assign n407 = ~x17 & n406 ;
  assign n408 = n394 & ~n407 ;
  assign n409 = n408 ^ x18 ;
  assign n410 = n393 & ~n409 ;
  assign n411 = n410 ^ n409 ;
  assign n412 = x29 & n365 ;
  assign n413 = x30 & ~x31 ;
  assign n414 = ~x158 & n413 ;
  assign n415 = n414 ^ x31 ;
  assign n416 = n412 & ~n415 ;
  assign n417 = n416 ^ n415 ;
  assign n418 = ~x32 & ~x159 ;
  assign n419 = n417 & n418 ;
  assign n420 = n419 ^ x32 ;
  assign n421 = x37 & n357 ;
  assign n422 = x38 & ~x39 ;
  assign n423 = ~x166 & n422 ;
  assign n424 = n423 ^ x39 ;
  assign n425 = n421 & ~n424 ;
  assign n426 = n425 ^ n424 ;
  assign n427 = ~x40 & ~x167 ;
  assign n428 = n426 & n427 ;
  assign n429 = n428 ^ x40 ;
  assign n430 = x125 & ~x126 ;
  assign n431 = ~x253 & n430 ;
  assign n432 = n431 ^ x126 ;
  assign n433 = ~x127 & ~x254 ;
  assign n434 = n432 & n433 ;
  assign n435 = n434 ^ x127 ;
  assign n436 = n272 & ~n435 ;
  assign n437 = x65 & n327 ;
  assign n438 = x66 & ~x67 ;
  assign n439 = ~x194 & n438 ;
  assign n440 = n439 ^ x67 ;
  assign n441 = n437 & ~n440 ;
  assign n442 = n441 ^ n440 ;
  assign n443 = ~x68 & ~x195 ;
  assign n444 = n442 & n443 ;
  assign n445 = n444 ^ x68 ;
  assign n446 = x69 & n324 ;
  assign n447 = x70 & ~x71 ;
  assign n448 = ~x198 & n447 ;
  assign n449 = n448 ^ x71 ;
  assign n450 = n446 & ~n449 ;
  assign n451 = n450 ^ n449 ;
  assign n452 = ~x72 & ~x199 ;
  assign n453 = n451 & n452 ;
  assign n454 = n453 ^ x72 ;
  assign n455 = n326 & ~n454 ;
  assign n456 = n445 & n455 ;
  assign n457 = n456 ^ n454 ;
  assign n458 = n330 & ~n457 ;
  assign n459 = x57 & ~x58 ;
  assign n460 = ~x185 & n459 ;
  assign n461 = n460 ^ x58 ;
  assign n462 = ~x59 & ~x186 ;
  assign n463 = n461 & n462 ;
  assign n464 = n463 ^ x59 ;
  assign n465 = ~x60 & ~x187 ;
  assign n466 = n464 & n465 ;
  assign n467 = n466 ^ x60 ;
  assign n468 = x61 & ~x62 ;
  assign n469 = ~x189 & n468 ;
  assign n470 = n469 ^ x62 ;
  assign n471 = ~x63 & ~x190 ;
  assign n472 = n470 & n471 ;
  assign n473 = n472 ^ x63 ;
  assign n474 = ~x64 & ~x191 ;
  assign n475 = n473 & n474 ;
  assign n476 = n475 ^ x64 ;
  assign n477 = n333 & ~n476 ;
  assign n478 = n467 & n477 ;
  assign n479 = n478 ^ n476 ;
  assign n480 = n458 & n479 ;
  assign n481 = n480 ^ n457 ;
  assign n482 = x81 & n309 ;
  assign n483 = x82 & ~x83 ;
  assign n484 = ~x210 & n483 ;
  assign n485 = n484 ^ x83 ;
  assign n486 = n482 & ~n485 ;
  assign n487 = n486 ^ n485 ;
  assign n488 = ~x84 & ~x211 ;
  assign n489 = n487 & n488 ;
  assign n490 = n489 ^ x84 ;
  assign n491 = x85 & ~x86 ;
  assign n492 = ~x213 & n491 ;
  assign n493 = n492 ^ x86 ;
  assign n494 = ~x87 & ~x214 ;
  assign n495 = n493 & n494 ;
  assign n496 = n495 ^ x87 ;
  assign n497 = ~x88 & ~x215 ;
  assign n498 = n496 & n497 ;
  assign n499 = n498 ^ x88 ;
  assign n500 = n308 & ~n499 ;
  assign n501 = n490 & n500 ;
  assign n502 = n501 ^ n499 ;
  assign n503 = x89 & ~x90 ;
  assign n504 = ~x217 & n503 ;
  assign n505 = n504 ^ x90 ;
  assign n506 = ~x91 & ~x218 ;
  assign n507 = n505 & n506 ;
  assign n508 = n507 ^ x91 ;
  assign n509 = ~x92 & ~x219 ;
  assign n510 = n508 & n509 ;
  assign n511 = n510 ^ x92 ;
  assign n512 = n305 & ~n511 ;
  assign n513 = n502 & n512 ;
  assign n514 = n513 ^ n511 ;
  assign n515 = x76 & ~x77 ;
  assign n516 = ~x204 & n515 ;
  assign n517 = n516 ^ x77 ;
  assign n518 = x78 & ~x79 ;
  assign n519 = ~x206 & n518 ;
  assign n520 = n519 ^ x79 ;
  assign n521 = ~x80 & ~x207 ;
  assign n522 = n520 & n521 ;
  assign n523 = n522 ^ x80 ;
  assign n524 = n315 & ~n523 ;
  assign n525 = n517 & n524 ;
  assign n526 = n525 ^ n523 ;
  assign n527 = n317 & ~n526 ;
  assign n528 = ~x74 & ~x202 ;
  assign n536 = x73 & n528 ;
  assign n537 = ~x201 & n536 ;
  assign n538 = n537 ^ x201 ;
  assign n529 = n528 ^ x202 ;
  assign n530 = n529 ^ x201 ;
  assign n539 = n538 ^ n530 ;
  assign n540 = ~x75 & n539 ;
  assign n541 = n527 & ~n540 ;
  assign n542 = n541 ^ n526 ;
  assign n543 = n313 & n542 ;
  assign n544 = ~n514 & n543 ;
  assign n545 = n544 ^ n514 ;
  assign n546 = ~x220 & n545 ;
  assign n547 = n302 & n546 ;
  assign n650 = x94 & ~x222 ;
  assign n651 = ~x95 & ~n650 ;
  assign n652 = ~x97 & ~x98 ;
  assign n653 = n651 & n652 ;
  assign n654 = x93 & ~x96 ;
  assign n655 = n273 & n654 ;
  assign n656 = n655 ^ x96 ;
  assign n657 = n653 & ~n656 ;
  assign n658 = n298 & ~n657 ;
  assign n548 = ~x107 & ~x234 ;
  assign n549 = x101 & n289 ;
  assign n550 = x102 & ~x103 ;
  assign n551 = ~x230 & n550 ;
  assign n552 = n551 ^ x103 ;
  assign n553 = n549 & ~n552 ;
  assign n554 = n553 ^ n552 ;
  assign n555 = ~x104 & ~x231 ;
  assign n556 = n554 & n555 ;
  assign n557 = n556 ^ x104 ;
  assign n558 = ~x232 & ~n557 ;
  assign n566 = n291 & n558 ;
  assign n567 = x100 & n566 ;
  assign n568 = n567 ^ x100 ;
  assign n559 = n558 ^ x232 ;
  assign n560 = n559 ^ x100 ;
  assign n569 = n568 ^ n560 ;
  assign n570 = ~x105 & n569 ;
  assign n571 = ~x233 & n570 ;
  assign n579 = n293 & n571 ;
  assign n580 = x99 & n579 ;
  assign n581 = n580 ^ x99 ;
  assign n572 = n571 ^ x233 ;
  assign n573 = n572 ^ x99 ;
  assign n582 = n581 ^ n573 ;
  assign n583 = ~x106 & n582 ;
  assign n584 = n548 & ~n583 ;
  assign n585 = n584 ^ x107 ;
  assign n586 = n288 & n585 ;
  assign n587 = ~x109 & ~x237 ;
  assign n588 = ~x236 & n587 ;
  assign n589 = x108 & n588 ;
  assign n590 = n589 ^ n587 ;
  assign n591 = n590 ^ x237 ;
  assign n592 = ~x110 & n591 ;
  assign n593 = ~n586 & n592 ;
  assign n594 = x113 & n280 ;
  assign n595 = x114 & ~x115 ;
  assign n596 = ~x242 & n595 ;
  assign n597 = n596 ^ x115 ;
  assign n598 = n594 & ~n597 ;
  assign n599 = n598 ^ n597 ;
  assign n600 = ~x116 & ~x243 ;
  assign n601 = n599 & n600 ;
  assign n602 = n601 ^ x116 ;
  assign n603 = ~x117 & ~x244 ;
  assign n604 = n602 & n603 ;
  assign n605 = n604 ^ x117 ;
  assign n606 = x118 & n278 ;
  assign n607 = ~x122 & ~x250 ;
  assign n615 = x121 & n607 ;
  assign n616 = ~x249 & n615 ;
  assign n617 = n616 ^ x249 ;
  assign n608 = n607 ^ x250 ;
  assign n609 = n608 ^ x249 ;
  assign n618 = n617 ^ n609 ;
  assign n619 = ~x123 & n618 ;
  assign n620 = ~x251 & n619 ;
  assign n628 = n275 & n620 ;
  assign n629 = x120 & n628 ;
  assign n630 = n629 ^ x120 ;
  assign n621 = n620 ^ x251 ;
  assign n622 = n621 ^ x120 ;
  assign n631 = n630 ^ n622 ;
  assign n632 = ~x124 & n631 ;
  assign n633 = x119 & n277 ;
  assign n634 = n632 & n633 ;
  assign n635 = n634 ^ n632 ;
  assign n636 = n606 & n635 ;
  assign n637 = n636 ^ n635 ;
  assign n638 = n279 & n637 ;
  assign n639 = n605 & n638 ;
  assign n640 = n639 ^ n637 ;
  assign n641 = x111 & ~x112 ;
  assign n642 = ~x239 & n641 ;
  assign n643 = n642 ^ x112 ;
  assign n644 = n284 & n643 ;
  assign n645 = n640 & n644 ;
  assign n646 = n645 ^ n640 ;
  assign n647 = n286 & n646 ;
  assign n648 = ~n593 & n647 ;
  assign n649 = n648 ^ n646 ;
  assign n659 = x96 & n299 ;
  assign n660 = x97 & ~x98 ;
  assign n661 = ~x225 & n660 ;
  assign n662 = n661 ^ x98 ;
  assign n663 = n659 & ~n662 ;
  assign n664 = n663 ^ n662 ;
  assign n665 = ~n300 & ~n664 ;
  assign n666 = n649 & ~n665 ;
  assign n667 = n658 & n666 ;
  assign n668 = n667 ^ n649 ;
  assign n669 = n547 & n668 ;
  assign n670 = n669 ^ n668 ;
  assign n671 = n323 & n670 ;
  assign n672 = n481 & n671 ;
  assign n673 = n672 ^ n670 ;
  assign n674 = ~x52 & ~x179 ;
  assign n675 = ~x50 & ~x178 ;
  assign n683 = x49 & n675 ;
  assign n684 = ~x177 & n683 ;
  assign n685 = n684 ^ x177 ;
  assign n676 = n675 ^ x178 ;
  assign n677 = n676 ^ x177 ;
  assign n686 = n685 ^ n677 ;
  assign n687 = ~x51 & n686 ;
  assign n688 = n674 & ~n687 ;
  assign n689 = n688 ^ x52 ;
  assign n690 = x53 & ~x54 ;
  assign n691 = ~x181 & n690 ;
  assign n692 = n691 ^ x54 ;
  assign n693 = ~x55 & ~x182 ;
  assign n694 = n692 & n693 ;
  assign n695 = n694 ^ x55 ;
  assign n696 = ~x56 & ~x183 ;
  assign n697 = n695 & n696 ;
  assign n698 = n697 ^ x56 ;
  assign n699 = n342 & ~n698 ;
  assign n700 = n689 & n699 ;
  assign n701 = n700 ^ n698 ;
  assign n702 = n339 & n701 ;
  assign n703 = n673 & n702 ;
  assign n704 = n703 ^ n673 ;
  assign n705 = n436 & ~n704 ;
  assign n706 = n705 ^ n435 ;
  assign n707 = n348 & ~n706 ;
  assign n708 = x41 & ~x42 ;
  assign n709 = ~x169 & n708 ;
  assign n710 = n709 ^ x42 ;
  assign n711 = x45 & n349 ;
  assign n712 = x46 & ~x47 ;
  assign n713 = ~x174 & n712 ;
  assign n714 = n713 ^ x47 ;
  assign n715 = n711 & ~n714 ;
  assign n716 = n715 ^ n714 ;
  assign n717 = ~x175 & ~n716 ;
  assign n718 = n350 & n717 ;
  assign n719 = x44 & n718 ;
  assign n720 = n719 ^ n717 ;
  assign n721 = n720 ^ x175 ;
  assign n722 = ~x48 & n721 ;
  assign n723 = x43 & n352 ;
  assign n724 = n722 & n723 ;
  assign n725 = n724 ^ n722 ;
  assign n726 = n353 & n725 ;
  assign n727 = n710 & n726 ;
  assign n728 = n727 ^ n725 ;
  assign n729 = n707 & ~n728 ;
  assign n730 = n729 ^ n706 ;
  assign n731 = n356 & ~n730 ;
  assign n732 = n429 & n731 ;
  assign n733 = n732 ^ n730 ;
  assign n734 = x33 & n361 ;
  assign n735 = x34 & ~x35 ;
  assign n736 = ~x162 & n735 ;
  assign n737 = n736 ^ x35 ;
  assign n738 = n734 & ~n737 ;
  assign n739 = n738 ^ n737 ;
  assign n740 = ~x36 & ~x163 ;
  assign n741 = n739 & n740 ;
  assign n742 = n741 ^ x36 ;
  assign n743 = n360 & n742 ;
  assign n744 = ~n733 & n743 ;
  assign n745 = n744 ^ n733 ;
  assign n746 = n364 & ~n745 ;
  assign n747 = n420 & n746 ;
  assign n748 = n747 ^ n745 ;
  assign n749 = x27 & ~x28 ;
  assign n750 = ~x155 & n749 ;
  assign n751 = n750 ^ x28 ;
  assign n752 = n368 & n751 ;
  assign n753 = ~n748 & n752 ;
  assign n754 = n753 ^ n748 ;
  assign n755 = x26 & n370 ;
  assign n756 = ~n754 & n755 ;
  assign n757 = n756 ^ n754 ;
  assign n758 = n371 & ~n757 ;
  assign n759 = x20 & ~x148 ;
  assign n760 = n373 & n759 ;
  assign n761 = x21 & n373 ;
  assign n762 = x22 & n372 ;
  assign n763 = x23 & ~x24 ;
  assign n764 = ~x151 & n763 ;
  assign n765 = n764 ^ x24 ;
  assign n766 = n762 & ~n765 ;
  assign n767 = n766 ^ n765 ;
  assign n768 = n761 & ~n767 ;
  assign n769 = n768 ^ n767 ;
  assign n770 = ~n760 & ~n769 ;
  assign n771 = ~x152 & n770 ;
  assign n779 = n375 & n771 ;
  assign n780 = x19 & n779 ;
  assign n781 = n780 ^ x19 ;
  assign n772 = n771 ^ x152 ;
  assign n773 = n772 ^ x19 ;
  assign n782 = n781 ^ n773 ;
  assign n783 = ~x25 & n782 ;
  assign n784 = n758 & ~n783 ;
  assign n785 = n784 ^ n757 ;
  assign n786 = n378 & ~n785 ;
  assign n787 = n411 & n786 ;
  assign n788 = n787 ^ n785 ;
  assign n789 = x11 & n384 ;
  assign n790 = x12 & ~x140 ;
  assign n791 = ~x13 & ~n790 ;
  assign n792 = ~n789 & n791 ;
  assign n793 = n383 & ~n792 ;
  assign n794 = ~n788 & n793 ;
  assign n795 = n794 ^ n788 ;
  assign n796 = ~x255 & ~n795 ;
  assign n800 = ~x8 & ~x136 ;
  assign n808 = x7 & n800 ;
  assign n809 = ~x135 & n808 ;
  assign n810 = n809 ^ x135 ;
  assign n801 = n800 ^ x136 ;
  assign n802 = n801 ^ x135 ;
  assign n811 = n810 ^ n802 ;
  assign n812 = ~x9 & n811 ;
  assign n813 = ~x137 & n812 ;
  assign n821 = n388 & n813 ;
  assign n822 = x6 & n821 ;
  assign n823 = n822 ^ x6 ;
  assign n814 = n813 ^ x137 ;
  assign n815 = n814 ^ x6 ;
  assign n824 = n823 ^ n815 ;
  assign n825 = ~x10 & n824 ;
  assign n830 = n796 & ~n825 ;
  assign n831 = n386 & n830 ;
  assign n832 = n831 ^ n386 ;
  assign n797 = n796 ^ x255 ;
  assign n798 = n797 ^ n386 ;
  assign n833 = n832 ^ n798 ;
  assign n834 = ~x0 & n833 ;
  assign n835 = x128 & n834 ;
  assign n836 = n392 & n835 ;
  assign n837 = n270 & n836 ;
  assign n838 = n837 ^ n835 ;
  assign n839 = n838 ^ x128 ;
  assign n840 = ~x1 & ~x128 ;
  assign n841 = n392 & n834 ;
  assign n846 = n261 & n268 ;
  assign n847 = n846 ^ n267 ;
  assign n848 = n841 & n847 ;
  assign n849 = n848 ^ n834 ;
  assign n850 = n840 & ~n849 ;
  assign n851 = n850 ^ x1 ;
  assign n852 = x129 & n851 ;
  assign n853 = ~x128 & n834 ;
  assign n854 = ~n267 & n392 ;
  assign n855 = x3 & n854 ;
  assign n856 = n264 & n855 ;
  assign n857 = n856 ^ n854 ;
  assign n858 = n857 ^ n392 ;
  assign n859 = n853 & ~n858 ;
  assign n860 = n859 ^ x128 ;
  assign n861 = ~x1 & n860 ;
  assign n862 = ~x2 & x130 ;
  assign n863 = ~x129 & n862 ;
  assign n864 = ~n861 & n863 ;
  assign n865 = n864 ^ n862 ;
  assign n866 = n865 ^ x130 ;
  assign n867 = ~x128 & n257 ;
  assign n868 = x131 & ~n263 ;
  assign n869 = ~n861 & n868 ;
  assign n870 = n867 & n869 ;
  assign n871 = n870 ^ n868 ;
  assign n872 = n871 ^ x131 ;
  assign n873 = ~x131 & ~n263 ;
  assign n874 = n834 & n867 ;
  assign n875 = x5 & n874 ;
  assign n876 = n392 & n875 ;
  assign n877 = n876 ^ n874 ;
  assign n878 = n877 ^ n867 ;
  assign n879 = n873 & ~n878 ;
  assign n880 = n879 ^ x131 ;
  assign n881 = ~x4 & x132 ;
  assign n882 = n880 & n881 ;
  assign n883 = n882 ^ x132 ;
  assign n884 = n264 & n867 ;
  assign n885 = ~n270 & n884 ;
  assign n886 = ~n834 & n885 ;
  assign n887 = n886 ^ n270 ;
  assign n888 = ~x133 & n887 ;
  assign n889 = n888 ^ n887 ;
  assign n890 = ~x6 & ~n888 ;
  assign n891 = ~x134 & ~n890 ;
  assign n892 = n891 ^ n890 ;
  assign n893 = ~x7 & ~n891 ;
  assign n894 = ~x135 & ~n893 ;
  assign n895 = n894 ^ n893 ;
  assign n896 = ~x8 & x136 ;
  assign n897 = ~n894 & n896 ;
  assign n898 = n897 ^ x136 ;
  assign n899 = x137 & n812 ;
  assign n900 = ~n890 & n899 ;
  assign n901 = n388 & n900 ;
  assign n902 = n901 ^ n899 ;
  assign n903 = n902 ^ x137 ;
  assign n904 = n391 & n884 ;
  assign n905 = ~n270 & n390 ;
  assign n913 = x0 & n905 ;
  assign n914 = n884 & n913 ;
  assign n915 = n914 ^ n884 ;
  assign n906 = n905 ^ n390 ;
  assign n907 = n906 ^ n884 ;
  assign n916 = n915 ^ n907 ;
  assign n917 = n825 & ~n916 ;
  assign n918 = x138 & n917 ;
  assign n919 = n904 & n918 ;
  assign n920 = n795 & n919 ;
  assign n921 = n920 ^ n918 ;
  assign n922 = n921 ^ x138 ;
  assign n923 = ~x138 & n904 ;
  assign n924 = ~n788 & n923 ;
  assign n932 = x13 & n924 ;
  assign n933 = n383 & n932 ;
  assign n934 = n933 ^ n383 ;
  assign n925 = n924 ^ n923 ;
  assign n926 = n925 ^ n383 ;
  assign n935 = n934 ^ n926 ;
  assign n936 = ~x11 & ~n935 ;
  assign n937 = ~x138 & ~n917 ;
  assign n938 = n936 & n937 ;
  assign n939 = n938 ^ n936 ;
  assign n940 = n790 & n923 ;
  assign n941 = n383 & n940 ;
  assign n942 = n941 ^ x139 ;
  assign n943 = x139 & n942 ;
  assign n944 = n939 & n943 ;
  assign n945 = n944 ^ x139 ;
  assign n946 = ~x12 & x140 ;
  assign n947 = ~x139 & n946 ;
  assign n948 = ~n939 & n947 ;
  assign n949 = n948 ^ n946 ;
  assign n950 = n949 ^ x140 ;
  assign n951 = n385 & n904 ;
  assign n952 = n385 & n792 ;
  assign n953 = ~n917 & n952 ;
  assign n954 = n953 ^ n792 ;
  assign n955 = x141 & n954 ;
  assign n956 = n951 & n955 ;
  assign n957 = n788 & n956 ;
  assign n958 = n957 ^ n955 ;
  assign n959 = n958 ^ x141 ;
  assign n960 = ~x141 & n951 ;
  assign n961 = n378 & n960 ;
  assign n962 = n951 ^ x141 ;
  assign n963 = n962 ^ x14 ;
  assign n964 = n954 ^ n951 ;
  assign n965 = n964 ^ x14 ;
  assign n966 = n954 ^ n785 ;
  assign n967 = n966 ^ x141 ;
  assign n968 = ~n965 & ~n967 ;
  assign n969 = n963 & n968 ;
  assign n970 = n969 ^ n954 ;
  assign n971 = n970 ^ x141 ;
  assign n972 = ~x14 & ~n971 ;
  assign n973 = ~x141 & n972 ;
  assign n974 = n973 ^ x14 ;
  assign n975 = x142 & ~n974 ;
  assign n976 = n961 & n975 ;
  assign n977 = n409 & n976 ;
  assign n978 = n977 ^ n975 ;
  assign n979 = n978 ^ x142 ;
  assign n980 = x18 & n961 ;
  assign n981 = ~n974 & n980 ;
  assign n982 = n981 ^ n974 ;
  assign n983 = ~x142 & ~n982 ;
  assign n987 = ~x145 & n961 ;
  assign n992 = n983 & n987 ;
  assign n993 = x17 & n992 ;
  assign n994 = n993 ^ x17 ;
  assign n984 = n983 ^ x142 ;
  assign n985 = n984 ^ x17 ;
  assign n995 = n994 ^ n985 ;
  assign n996 = ~x15 & n995 ;
  assign n997 = n379 & n987 ;
  assign n998 = x16 & n997 ;
  assign n999 = n998 ^ x143 ;
  assign n1000 = x143 & n999 ;
  assign n1001 = n996 & n1000 ;
  assign n1002 = n1001 ^ x143 ;
  assign n1003 = ~x16 & x144 ;
  assign n1004 = ~x143 & n1003 ;
  assign n1005 = ~n996 & n1004 ;
  assign n1006 = n1005 ^ n1003 ;
  assign n1007 = n1006 ^ x144 ;
  assign n1008 = x145 & n407 ;
  assign n1009 = n982 & n1008 ;
  assign n1010 = n380 & n1009 ;
  assign n1011 = n1010 ^ n1008 ;
  assign n1012 = n1011 ^ x145 ;
  assign n1013 = x146 & ~n409 ;
  assign n1014 = n381 & n1013 ;
  assign n1015 = n974 & n1014 ;
  assign n1016 = n1015 ^ n1013 ;
  assign n1017 = n1016 ^ x146 ;
  assign n1018 = n382 & n951 ;
  assign n1019 = n376 & n1018 ;
  assign n1020 = n371 & n1019 ;
  assign n1021 = n382 & ~n411 ;
  assign n1022 = ~n954 & n1021 ;
  assign n1023 = n1022 ^ n411 ;
  assign n1024 = ~x146 & ~n1023 ;
  assign n1025 = ~n757 & n1018 ;
  assign n1026 = x25 & n1025 ;
  assign n1027 = n371 & n1026 ;
  assign n1028 = n1027 ^ n1025 ;
  assign n1029 = n1028 ^ n1018 ;
  assign n1030 = n1024 & ~n1029 ;
  assign n1031 = n1030 ^ x146 ;
  assign n1032 = ~x19 & n1031 ;
  assign n1033 = n769 & n1020 ;
  assign n1034 = n1032 & n1033 ;
  assign n1035 = n1034 ^ n1032 ;
  assign n1036 = x147 & n1035 ;
  assign n1037 = n1020 & n1036 ;
  assign n1038 = n760 & n1037 ;
  assign n1039 = n1038 ^ n1036 ;
  assign n1040 = n1039 ^ x147 ;
  assign n1041 = ~x20 & x148 ;
  assign n1042 = ~x147 & n1041 ;
  assign n1043 = ~n1035 & n1042 ;
  assign n1044 = n1043 ^ n1041 ;
  assign n1045 = n1044 ^ x148 ;
  assign n1046 = n374 & n1020 ;
  assign n1047 = n374 & ~n1032 ;
  assign n1048 = ~x21 & ~n759 ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1050 = x149 & n1049 ;
  assign n1051 = n1046 & n1050 ;
  assign n1052 = n767 & n1051 ;
  assign n1053 = n1052 ^ n1050 ;
  assign n1054 = n1053 ^ x149 ;
  assign n1055 = ~x22 & x150 ;
  assign n1056 = n765 & n1046 ;
  assign n1057 = ~x149 & n1049 ;
  assign n1060 = n1056 & n1057 ;
  assign n1058 = n1057 ^ x149 ;
  assign n1061 = n1060 ^ n1058 ;
  assign n1062 = n1055 & n1061 ;
  assign n1063 = n1062 ^ x150 ;
  assign n1064 = ~x22 & ~x150 ;
  assign n1065 = x24 & n1046 ;
  assign n1066 = n1057 & n1065 ;
  assign n1067 = n1066 ^ n1058 ;
  assign n1068 = n1064 & n1067 ;
  assign n1069 = n1068 ^ x150 ;
  assign n1070 = ~x23 & x151 ;
  assign n1071 = n1069 & n1070 ;
  assign n1072 = n1071 ^ x151 ;
  assign n1073 = x152 & ~n767 ;
  assign n1074 = n373 & n1073 ;
  assign n1075 = ~n1049 & n1074 ;
  assign n1076 = n1075 ^ n1073 ;
  assign n1077 = n1076 ^ x152 ;
  assign n1078 = n377 & n1018 ;
  assign n1079 = n377 & n1023 ;
  assign n1080 = n783 & n1079 ;
  assign n1081 = n1080 ^ n783 ;
  assign n1082 = x153 & n1081 ;
  assign n1083 = n1078 & n1082 ;
  assign n1084 = n757 & n1083 ;
  assign n1085 = n1084 ^ n1082 ;
  assign n1086 = n1085 ^ x153 ;
  assign n1087 = ~x153 & n1078 ;
  assign n1088 = ~x26 & ~x153 ;
  assign n1089 = ~n1081 & n1088 ;
  assign n1090 = n1089 ^ x26 ;
  assign n1091 = x154 & ~n1090 ;
  assign n1092 = n1087 & n1091 ;
  assign n1093 = n754 & n1092 ;
  assign n1094 = n1093 ^ n1091 ;
  assign n1095 = n1094 ^ x154 ;
  assign n1096 = ~x154 & ~n1090 ;
  assign n1097 = ~n748 & n1087 ;
  assign n1098 = x28 & n1097 ;
  assign n1099 = n368 & n1098 ;
  assign n1100 = n1099 ^ n1097 ;
  assign n1101 = n1100 ^ n1087 ;
  assign n1102 = n1096 & ~n1101 ;
  assign n1103 = n1102 ^ x154 ;
  assign n1104 = ~x27 & x155 ;
  assign n1105 = n1103 & n1104 ;
  assign n1106 = n1105 ^ x155 ;
  assign n1107 = n369 & n1087 ;
  assign n1108 = n369 & ~n751 ;
  assign n1109 = n1090 & n1108 ;
  assign n1110 = n1109 ^ n751 ;
  assign n1111 = x156 & ~n1110 ;
  assign n1112 = n1107 & n1111 ;
  assign n1113 = n748 & n1112 ;
  assign n1114 = n1113 ^ n1111 ;
  assign n1115 = n1114 ^ x156 ;
  assign n1116 = ~x29 & x157 ;
  assign n1117 = ~n745 & n1107 ;
  assign n1125 = x32 & n1117 ;
  assign n1126 = n364 & n1125 ;
  assign n1127 = n1126 ^ n364 ;
  assign n1118 = n1117 ^ n1107 ;
  assign n1119 = n1118 ^ n364 ;
  assign n1128 = n1127 ^ n1119 ;
  assign n1129 = ~n1110 & ~n1128 ;
  assign n1130 = ~x156 & n1129 ;
  assign n1135 = n1130 ^ x156 ;
  assign n1131 = ~x159 & n364 ;
  assign n1132 = n1107 & n1131 ;
  assign n1133 = n415 & n1132 ;
  assign n1134 = n1130 & n1133 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1137 = n1116 & n1136 ;
  assign n1138 = n1137 ^ x157 ;
  assign n1139 = ~x29 & ~x157 ;
  assign n1140 = x31 & n1132 ;
  assign n1142 = n1130 & n1140 ;
  assign n1143 = n1142 ^ n1135 ;
  assign n1144 = n1139 & n1143 ;
  assign n1145 = n1144 ^ x157 ;
  assign n1146 = ~x30 & x158 ;
  assign n1147 = n1145 & n1146 ;
  assign n1148 = n1147 ^ x158 ;
  assign n1149 = x159 & ~n417 ;
  assign n1150 = n366 & n1149 ;
  assign n1151 = ~n1129 & n1150 ;
  assign n1152 = n1151 ^ n1149 ;
  assign n1153 = n1152 ^ x159 ;
  assign n1154 = n367 & n1107 ;
  assign n1155 = n367 & ~n420 ;
  assign n1156 = n1110 & n1155 ;
  assign n1157 = n1156 ^ n420 ;
  assign n1158 = x160 & ~n1157 ;
  assign n1159 = n1154 & n1158 ;
  assign n1160 = n745 & n1159 ;
  assign n1161 = n1160 ^ n1158 ;
  assign n1162 = n1161 ^ x160 ;
  assign n1163 = ~x33 & x161 ;
  assign n1164 = ~n733 & n1154 ;
  assign n1172 = x36 & n1164 ;
  assign n1173 = n360 & n1172 ;
  assign n1174 = n1173 ^ n360 ;
  assign n1165 = n1164 ^ n1154 ;
  assign n1166 = n1165 ^ n360 ;
  assign n1175 = n1174 ^ n1166 ;
  assign n1176 = ~n1157 & ~n1175 ;
  assign n1177 = ~x160 & n1176 ;
  assign n1182 = n1177 ^ x160 ;
  assign n1178 = ~x163 & n360 ;
  assign n1179 = n1154 & n1178 ;
  assign n1180 = n737 & n1179 ;
  assign n1181 = n1177 & n1180 ;
  assign n1183 = n1182 ^ n1181 ;
  assign n1184 = n1163 & n1183 ;
  assign n1185 = n1184 ^ x161 ;
  assign n1186 = ~x33 & ~x161 ;
  assign n1187 = x35 & n1179 ;
  assign n1189 = n1177 & n1187 ;
  assign n1190 = n1189 ^ n1182 ;
  assign n1191 = n1186 & n1190 ;
  assign n1192 = n1191 ^ x161 ;
  assign n1193 = ~x34 & x162 ;
  assign n1194 = n1192 & n1193 ;
  assign n1195 = n1194 ^ x162 ;
  assign n1196 = x163 & ~n739 ;
  assign n1197 = n362 & n1196 ;
  assign n1198 = ~n1176 & n1197 ;
  assign n1199 = n1198 ^ n1196 ;
  assign n1200 = n1199 ^ x163 ;
  assign n1201 = n363 & n1154 ;
  assign n1202 = n363 & ~n742 ;
  assign n1203 = n1157 & n1202 ;
  assign n1204 = n1203 ^ n742 ;
  assign n1205 = x164 & ~n1204 ;
  assign n1206 = n1201 & n1205 ;
  assign n1207 = n733 & n1206 ;
  assign n1208 = n1207 ^ n1205 ;
  assign n1209 = n1208 ^ x164 ;
  assign n1210 = ~x37 & x165 ;
  assign n1211 = ~n730 & n1201 ;
  assign n1219 = x40 & n1211 ;
  assign n1220 = n356 & n1219 ;
  assign n1221 = n1220 ^ n356 ;
  assign n1212 = n1211 ^ n1201 ;
  assign n1213 = n1212 ^ n356 ;
  assign n1222 = n1221 ^ n1213 ;
  assign n1223 = ~n1204 & ~n1222 ;
  assign n1224 = ~x164 & n1223 ;
  assign n1229 = n1224 ^ x164 ;
  assign n1225 = ~x167 & n356 ;
  assign n1226 = n1201 & n1225 ;
  assign n1227 = n424 & n1226 ;
  assign n1228 = n1224 & n1227 ;
  assign n1230 = n1229 ^ n1228 ;
  assign n1231 = n1210 & n1230 ;
  assign n1232 = n1231 ^ x165 ;
  assign n1233 = ~x37 & ~x165 ;
  assign n1234 = x39 & n1226 ;
  assign n1236 = n1224 & n1234 ;
  assign n1237 = n1236 ^ n1229 ;
  assign n1238 = n1233 & n1237 ;
  assign n1239 = n1238 ^ x165 ;
  assign n1240 = ~x38 & x166 ;
  assign n1241 = n1239 & n1240 ;
  assign n1242 = n1241 ^ x166 ;
  assign n1243 = x167 & ~n426 ;
  assign n1244 = n358 & n1243 ;
  assign n1245 = ~n1223 & n1244 ;
  assign n1246 = n1245 ^ n1243 ;
  assign n1247 = n1246 ^ x167 ;
  assign n1248 = n359 & n1201 ;
  assign n1249 = n359 & ~n429 ;
  assign n1250 = n1204 & n1249 ;
  assign n1251 = n1250 ^ n429 ;
  assign n1252 = x168 & ~n1251 ;
  assign n1253 = n1248 & n1252 ;
  assign n1254 = n730 & n1253 ;
  assign n1255 = n1254 ^ n1252 ;
  assign n1256 = n1255 ^ x168 ;
  assign n1257 = n706 & n1248 ;
  assign n1258 = ~n1251 & n1257 ;
  assign n1259 = n1258 ^ n1251 ;
  assign n1260 = ~x168 & ~n1259 ;
  assign n1261 = n348 & n1248 ;
  assign n1262 = n725 & n1261 ;
  assign n1263 = x42 & n1262 ;
  assign n1264 = n353 & n1263 ;
  assign n1265 = n1264 ^ n1262 ;
  assign n1266 = n1265 ^ n1261 ;
  assign n1267 = n1260 & ~n1266 ;
  assign n1268 = n1267 ^ x168 ;
  assign n1269 = ~x41 & x169 ;
  assign n1270 = n1268 & n1269 ;
  assign n1271 = n1270 ^ x169 ;
  assign n1272 = n354 & n1261 ;
  assign n1273 = n354 & ~n710 ;
  assign n1274 = n1259 & n1273 ;
  assign n1275 = n1274 ^ n710 ;
  assign n1276 = x170 & ~n1275 ;
  assign n1277 = n1272 & n1276 ;
  assign n1278 = ~n725 & n1277 ;
  assign n1279 = n1278 ^ n1276 ;
  assign n1280 = n1279 ^ x170 ;
  assign n1281 = ~x170 & n1272 ;
  assign n1282 = n1272 ^ x170 ;
  assign n1283 = n1282 ^ x43 ;
  assign n1284 = n1275 ^ n1272 ;
  assign n1285 = n1284 ^ x43 ;
  assign n1286 = n1275 ^ x48 ;
  assign n1287 = n1286 ^ x170 ;
  assign n1288 = n1285 & n1287 ;
  assign n1289 = n1283 & n1288 ;
  assign n1290 = n1289 ^ n1275 ;
  assign n1291 = n1290 ^ x170 ;
  assign n1292 = ~x43 & n1291 ;
  assign n1293 = ~x170 & n1292 ;
  assign n1294 = n1293 ^ x43 ;
  assign n1295 = x171 & ~n1294 ;
  assign n1296 = n1281 & n1295 ;
  assign n1297 = ~n721 & n1296 ;
  assign n1298 = n1297 ^ n1295 ;
  assign n1299 = n1298 ^ x171 ;
  assign n1300 = n351 & n1281 ;
  assign n1301 = ~x44 & ~x171 ;
  assign n1302 = n1294 & n1301 ;
  assign n1303 = n1302 ^ x44 ;
  assign n1304 = x172 & ~n1303 ;
  assign n1305 = n1300 & n1304 ;
  assign n1306 = n716 & n1305 ;
  assign n1307 = n1306 ^ n1304 ;
  assign n1308 = n1307 ^ x172 ;
  assign n1309 = ~x45 & x173 ;
  assign n1310 = n714 & n1300 ;
  assign n1311 = ~x172 & ~n1303 ;
  assign n1314 = n1310 & n1311 ;
  assign n1312 = n1311 ^ x172 ;
  assign n1315 = n1314 ^ n1312 ;
  assign n1316 = n1309 & n1315 ;
  assign n1317 = n1316 ^ x173 ;
  assign n1318 = ~x45 & ~x173 ;
  assign n1319 = x47 & n1300 ;
  assign n1320 = n1311 & n1319 ;
  assign n1321 = n1320 ^ n1312 ;
  assign n1322 = n1318 & n1321 ;
  assign n1323 = n1322 ^ x173 ;
  assign n1324 = ~x46 & x174 ;
  assign n1325 = n1323 & n1324 ;
  assign n1326 = n1325 ^ x174 ;
  assign n1327 = x175 & ~n716 ;
  assign n1328 = n350 & n1327 ;
  assign n1329 = n1303 & n1328 ;
  assign n1330 = n1329 ^ n1327 ;
  assign n1331 = n1330 ^ x175 ;
  assign n1332 = x176 & n728 ;
  assign n1333 = n1259 & n1332 ;
  assign n1334 = n355 & n1333 ;
  assign n1335 = n1334 ^ n1332 ;
  assign n1336 = n1335 ^ x176 ;
  assign n1337 = n355 & n1248 ;
  assign n1338 = n272 & n1337 ;
  assign n1339 = n355 & n1251 ;
  assign n1340 = n728 & n1339 ;
  assign n1341 = n1340 ^ n728 ;
  assign n1342 = n435 & n1337 ;
  assign n1343 = n1341 & n1342 ;
  assign n1344 = n1343 ^ n1341 ;
  assign n1345 = n1338 & n1344 ;
  assign n1346 = ~n673 & n1345 ;
  assign n1347 = n1346 ^ n1344 ;
  assign n1348 = n339 & n1338 ;
  assign n1349 = ~n698 & n1348 ;
  assign n1357 = n342 & n1349 ;
  assign n1358 = x52 & n1357 ;
  assign n1359 = n1358 ^ x52 ;
  assign n1350 = n1349 ^ n1348 ;
  assign n1351 = n1350 ^ x52 ;
  assign n1360 = n1359 ^ n1351 ;
  assign n1361 = n1347 & ~n1360 ;
  assign n1362 = ~x176 & n1361 ;
  assign n1366 = ~x179 & n342 ;
  assign n1367 = n1348 & n1366 ;
  assign n1372 = n1362 & n1367 ;
  assign n1373 = x51 & n1372 ;
  assign n1374 = n1373 ^ x51 ;
  assign n1363 = n1362 ^ x176 ;
  assign n1364 = n1363 ^ x51 ;
  assign n1375 = n1374 ^ n1364 ;
  assign n1376 = ~x49 & n1375 ;
  assign n1377 = n343 & n1367 ;
  assign n1378 = x50 & n1377 ;
  assign n1379 = n1378 ^ x177 ;
  assign n1380 = x177 & n1379 ;
  assign n1381 = n1376 & n1380 ;
  assign n1382 = n1381 ^ x177 ;
  assign n1383 = ~x50 & x178 ;
  assign n1384 = ~x177 & n1383 ;
  assign n1385 = ~n1376 & n1384 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1387 = n1386 ^ x178 ;
  assign n1388 = x179 & n687 ;
  assign n1389 = n344 & n1388 ;
  assign n1390 = ~n1361 & n1389 ;
  assign n1391 = n1390 ^ n1388 ;
  assign n1392 = n1391 ^ x179 ;
  assign n1393 = n345 & n1348 ;
  assign n1394 = n345 & ~n689 ;
  assign n1395 = ~n1347 & n1394 ;
  assign n1396 = n1395 ^ n689 ;
  assign n1397 = x180 & ~n1396 ;
  assign n1398 = n1393 & n1397 ;
  assign n1399 = n698 & n1398 ;
  assign n1400 = n1399 ^ n1397 ;
  assign n1401 = n1400 ^ x180 ;
  assign n1402 = ~x183 & n1393 ;
  assign n1403 = x55 & n1402 ;
  assign n1404 = x56 & n1393 ;
  assign n1405 = ~n1396 & n1404 ;
  assign n1406 = n1405 ^ n1396 ;
  assign n1407 = n1403 & ~n1406 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1409 = ~x182 & n1402 ;
  assign n1410 = x54 & n1409 ;
  assign n1411 = n1410 ^ x180 ;
  assign n1412 = ~x180 & ~n1411 ;
  assign n1413 = ~n1408 & n1412 ;
  assign n1414 = n1413 ^ x180 ;
  assign n1415 = ~x53 & x181 ;
  assign n1416 = n1414 & n1415 ;
  assign n1417 = n1416 ^ x181 ;
  assign n1418 = x182 & ~n692 ;
  assign n1419 = n340 & n1418 ;
  assign n1420 = n1408 & n1419 ;
  assign n1421 = n1420 ^ n1418 ;
  assign n1422 = n1421 ^ x182 ;
  assign n1423 = x183 & ~n695 ;
  assign n1424 = n341 & n1423 ;
  assign n1425 = n1406 & n1424 ;
  assign n1426 = n1425 ^ n1423 ;
  assign n1427 = n1426 ^ x183 ;
  assign n1432 = n699 & n1396 ;
  assign n1433 = n1432 ^ n698 ;
  assign n1434 = x184 & n1433 ;
  assign n1435 = n346 & n1338 ;
  assign n1436 = n323 & n1435 ;
  assign n1437 = n330 & n1436 ;
  assign n1438 = n333 & n1437 ;
  assign n1439 = ~x187 & n1438 ;
  assign n1440 = x59 & n1439 ;
  assign n1441 = x60 & n1438 ;
  assign n1442 = ~n670 & n1435 ;
  assign n1443 = n346 & ~n701 ;
  assign n1444 = ~n1344 & n1443 ;
  assign n1445 = n1444 ^ n701 ;
  assign n1446 = n1442 & ~n1445 ;
  assign n1447 = n1446 ^ n1445 ;
  assign n1448 = n1436 & ~n1447 ;
  assign n1449 = n457 & n1448 ;
  assign n1450 = n1449 ^ n1447 ;
  assign n1451 = n476 & n1437 ;
  assign n1452 = ~n1450 & n1451 ;
  assign n1453 = n1452 ^ n1450 ;
  assign n1454 = n1441 & ~n1453 ;
  assign n1455 = n1454 ^ n1453 ;
  assign n1456 = n1440 & ~n1455 ;
  assign n1457 = n1456 ^ n1455 ;
  assign n1458 = ~x186 & n1439 ;
  assign n1459 = x58 & n1458 ;
  assign n1460 = n1459 ^ x184 ;
  assign n1461 = ~x184 & ~n1460 ;
  assign n1462 = ~n1457 & n1461 ;
  assign n1463 = n1462 ^ x184 ;
  assign n1464 = ~x57 & x185 ;
  assign n1465 = n1463 & n1464 ;
  assign n1466 = n1465 ^ x185 ;
  assign n1467 = x186 & ~n461 ;
  assign n1468 = n334 & n1467 ;
  assign n1469 = n1457 & n1468 ;
  assign n1470 = n1469 ^ n1467 ;
  assign n1471 = n1470 ^ x186 ;
  assign n1472 = x187 & ~n464 ;
  assign n1473 = n335 & n1472 ;
  assign n1474 = n1455 & n1473 ;
  assign n1475 = n1474 ^ n1472 ;
  assign n1476 = n1475 ^ x187 ;
  assign n1477 = x188 & ~n467 ;
  assign n1478 = n336 & n1477 ;
  assign n1479 = n1453 & n1478 ;
  assign n1480 = n1479 ^ n1477 ;
  assign n1481 = n1480 ^ x188 ;
  assign n1482 = n336 & ~n1450 ;
  assign n1490 = n1437 & n1482 ;
  assign n1491 = x64 & n1490 ;
  assign n1492 = n1491 ^ x64 ;
  assign n1483 = n1482 ^ n336 ;
  assign n1484 = n1483 ^ x64 ;
  assign n1493 = n1492 ^ n1484 ;
  assign n1494 = ~n467 & ~n1493 ;
  assign n1495 = ~x191 & n336 ;
  assign n1496 = n1437 & n1495 ;
  assign n1497 = x63 & n1496 ;
  assign n1498 = n1494 & n1497 ;
  assign n1499 = n1498 ^ n1494 ;
  assign n1500 = ~x190 & n1496 ;
  assign n1501 = x62 & n1500 ;
  assign n1502 = n1501 ^ x188 ;
  assign n1503 = ~x188 & ~n1502 ;
  assign n1504 = n1499 & n1503 ;
  assign n1505 = n1504 ^ x188 ;
  assign n1506 = ~x61 & x189 ;
  assign n1507 = n1505 & n1506 ;
  assign n1508 = n1507 ^ x189 ;
  assign n1509 = x190 & ~n470 ;
  assign n1510 = n331 & n1509 ;
  assign n1511 = ~n1499 & n1510 ;
  assign n1512 = n1511 ^ n1509 ;
  assign n1513 = n1512 ^ x190 ;
  assign n1514 = x191 & ~n473 ;
  assign n1515 = n332 & n1514 ;
  assign n1516 = ~n1494 & n1515 ;
  assign n1517 = n1516 ^ n1514 ;
  assign n1518 = n1517 ^ x191 ;
  assign n1519 = x192 & ~n479 ;
  assign n1520 = n1450 & n1519 ;
  assign n1521 = n337 & n1520 ;
  assign n1522 = n1521 ^ n1519 ;
  assign n1523 = n1522 ^ x192 ;
  assign n1524 = ~x65 & x193 ;
  assign n1525 = n337 & n1436 ;
  assign n1526 = n326 & n1525 ;
  assign n1527 = x68 & n1526 ;
  assign n1528 = n337 & n1447 ;
  assign n1529 = ~n479 & n1528 ;
  assign n1530 = n1529 ^ n479 ;
  assign n1531 = n454 & n1525 ;
  assign n1532 = ~n1530 & n1531 ;
  assign n1533 = n1532 ^ n1530 ;
  assign n1534 = n1527 & ~n1533 ;
  assign n1535 = n1534 ^ n1533 ;
  assign n1536 = ~x192 & ~n1535 ;
  assign n1540 = n1536 ^ x192 ;
  assign n1537 = ~x195 & n1526 ;
  assign n1538 = n440 & n1537 ;
  assign n1539 = n1536 & n1538 ;
  assign n1541 = n1540 ^ n1539 ;
  assign n1542 = n1524 & n1541 ;
  assign n1543 = n1542 ^ x193 ;
  assign n1544 = ~x65 & ~x193 ;
  assign n1545 = x67 & n1537 ;
  assign n1547 = n1536 & n1545 ;
  assign n1548 = n1547 ^ n1540 ;
  assign n1549 = n1544 & n1548 ;
  assign n1550 = n1549 ^ x193 ;
  assign n1551 = ~x66 & x194 ;
  assign n1552 = n1550 & n1551 ;
  assign n1553 = n1552 ^ x194 ;
  assign n1554 = x195 & ~n442 ;
  assign n1555 = n328 & n1554 ;
  assign n1556 = n1535 & n1555 ;
  assign n1557 = n1556 ^ n1554 ;
  assign n1558 = n1557 ^ x195 ;
  assign n1559 = x196 & ~n445 ;
  assign n1560 = n329 & n1559 ;
  assign n1561 = n1533 & n1560 ;
  assign n1562 = n1561 ^ n1559 ;
  assign n1563 = n1562 ^ x196 ;
  assign n1564 = ~x69 & x197 ;
  assign n1565 = n329 & ~n1530 ;
  assign n1573 = n1525 & n1565 ;
  assign n1574 = x72 & n1573 ;
  assign n1575 = n1574 ^ x72 ;
  assign n1566 = n1565 ^ n329 ;
  assign n1567 = n1566 ^ x72 ;
  assign n1576 = n1575 ^ n1567 ;
  assign n1577 = ~n445 & ~n1576 ;
  assign n1578 = ~x196 & n1577 ;
  assign n1583 = n1578 ^ x196 ;
  assign n1579 = ~x199 & n329 ;
  assign n1580 = n1525 & n1579 ;
  assign n1581 = n449 & n1580 ;
  assign n1582 = n1578 & n1581 ;
  assign n1584 = n1583 ^ n1582 ;
  assign n1585 = n1564 & n1584 ;
  assign n1586 = n1585 ^ x197 ;
  assign n1587 = ~x69 & ~x197 ;
  assign n1588 = x71 & n1580 ;
  assign n1590 = n1578 & n1588 ;
  assign n1591 = n1590 ^ n1583 ;
  assign n1592 = n1587 & n1591 ;
  assign n1593 = n1592 ^ x197 ;
  assign n1594 = ~x70 & x198 ;
  assign n1595 = n1593 & n1594 ;
  assign n1596 = n1595 ^ x198 ;
  assign n1597 = x199 & ~n451 ;
  assign n1598 = n325 & n1597 ;
  assign n1599 = ~n1577 & n1598 ;
  assign n1600 = n1599 ^ n1597 ;
  assign n1601 = n1600 ^ x199 ;
  assign n1606 = n458 & n1530 ;
  assign n1607 = n1606 ^ n457 ;
  assign n1608 = x200 & n1607 ;
  assign n1609 = n338 & n1435 ;
  assign n1610 = ~x220 & n302 ;
  assign n1611 = n1609 & n1610 ;
  assign n1612 = n313 & n1611 ;
  assign n1613 = ~n526 & n1612 ;
  assign n1621 = x75 & n1613 ;
  assign n1622 = n317 & n1621 ;
  assign n1623 = n1622 ^ n317 ;
  assign n1614 = n1613 ^ n1612 ;
  assign n1615 = n1614 ^ n317 ;
  assign n1624 = n1623 ^ n1615 ;
  assign n1625 = ~n668 & n1609 ;
  assign n1626 = n338 & ~n481 ;
  assign n1627 = n1445 & n1626 ;
  assign n1628 = n1627 ^ n481 ;
  assign n1629 = n1625 & ~n1628 ;
  assign n1630 = n1629 ^ n1628 ;
  assign n1631 = n1611 & ~n1630 ;
  assign n1632 = n514 & n1631 ;
  assign n1633 = n1632 ^ n1630 ;
  assign n1634 = ~x200 & ~n1633 ;
  assign n1635 = ~n1624 & n1634 ;
  assign n1636 = n1635 ^ x200 ;
  assign n1637 = ~x73 & n1636 ;
  assign n1638 = x74 & n318 ;
  assign n1639 = n317 & n1638 ;
  assign n1640 = n1612 & n1639 ;
  assign n1641 = n1637 & ~n1640 ;
  assign n1642 = x201 & ~n1641 ;
  assign n1643 = ~x74 & x202 ;
  assign n1644 = ~x201 & n1643 ;
  assign n1645 = ~n1637 & n1644 ;
  assign n1646 = n1645 ^ n1643 ;
  assign n1647 = n1646 ^ x202 ;
  assign n1648 = n319 & n1612 ;
  assign n1649 = n319 & n1633 ;
  assign n1650 = n540 & n1649 ;
  assign n1651 = n1650 ^ n540 ;
  assign n1652 = x203 & n1651 ;
  assign n1653 = n1648 & n1652 ;
  assign n1654 = n526 & n1653 ;
  assign n1655 = n1654 ^ n1652 ;
  assign n1656 = n1655 ^ x203 ;
  assign n1657 = ~x203 & n1651 ;
  assign n1658 = ~n523 & n1648 ;
  assign n1659 = x77 & n1658 ;
  assign n1660 = n315 & n1659 ;
  assign n1661 = n1660 ^ n1658 ;
  assign n1662 = n1661 ^ n1648 ;
  assign n1663 = n1657 & ~n1662 ;
  assign n1664 = n1663 ^ x203 ;
  assign n1665 = ~x76 & x204 ;
  assign n1666 = n1664 & n1665 ;
  assign n1667 = n1666 ^ x204 ;
  assign n1668 = n316 & n1648 ;
  assign n1669 = n316 & ~n517 ;
  assign n1670 = ~n1651 & n1669 ;
  assign n1671 = n1670 ^ n517 ;
  assign n1672 = x205 & ~n1671 ;
  assign n1673 = n1668 & n1672 ;
  assign n1674 = n523 & n1673 ;
  assign n1675 = n1674 ^ n1672 ;
  assign n1676 = n1675 ^ x205 ;
  assign n1677 = x80 & n1668 ;
  assign n1678 = ~n1671 & n1677 ;
  assign n1679 = n1678 ^ n1671 ;
  assign n1680 = ~x207 & n1668 ;
  assign n1681 = x79 & n1680 ;
  assign n1682 = n1681 ^ x205 ;
  assign n1683 = ~x205 & ~n1682 ;
  assign n1684 = ~n1679 & n1683 ;
  assign n1685 = n1684 ^ x205 ;
  assign n1686 = ~x78 & x206 ;
  assign n1687 = n1685 & n1686 ;
  assign n1688 = n1687 ^ x206 ;
  assign n1689 = x207 & ~n520 ;
  assign n1690 = n314 & n1689 ;
  assign n1691 = n1679 & n1690 ;
  assign n1692 = n1691 ^ n1689 ;
  assign n1693 = n1692 ^ x207 ;
  assign n1698 = n524 & n1671 ;
  assign n1699 = n1698 ^ n523 ;
  assign n1700 = x208 & n1699 ;
  assign n1701 = ~x81 & x209 ;
  assign n1702 = n320 & n1611 ;
  assign n1703 = n511 & n1702 ;
  assign n1704 = n320 & ~n542 ;
  assign n1705 = n1630 & n1704 ;
  assign n1706 = n1705 ^ n542 ;
  assign n1707 = n1703 & ~n1706 ;
  assign n1708 = n1707 ^ n1706 ;
  assign n1709 = n305 & n1702 ;
  assign n1710 = ~n499 & n1709 ;
  assign n1718 = x84 & n1710 ;
  assign n1719 = n308 & n1718 ;
  assign n1720 = n1719 ^ n308 ;
  assign n1711 = n1710 ^ n1709 ;
  assign n1712 = n1711 ^ n308 ;
  assign n1721 = n1720 ^ n1712 ;
  assign n1722 = ~n1708 & ~n1721 ;
  assign n1723 = ~x208 & n1722 ;
  assign n1728 = n1723 ^ x208 ;
  assign n1724 = ~x211 & n308 ;
  assign n1725 = n1709 & n1724 ;
  assign n1726 = n485 & n1725 ;
  assign n1727 = n1723 & n1726 ;
  assign n1729 = n1728 ^ n1727 ;
  assign n1730 = n1701 & n1729 ;
  assign n1731 = n1730 ^ x209 ;
  assign n1732 = ~x81 & ~x209 ;
  assign n1733 = x83 & n1725 ;
  assign n1735 = n1723 & n1733 ;
  assign n1736 = n1735 ^ n1728 ;
  assign n1737 = n1732 & n1736 ;
  assign n1738 = n1737 ^ x209 ;
  assign n1739 = ~x82 & x210 ;
  assign n1740 = n1738 & n1739 ;
  assign n1741 = n1740 ^ x210 ;
  assign n1742 = x211 & ~n487 ;
  assign n1743 = n310 & n1742 ;
  assign n1744 = ~n1722 & n1743 ;
  assign n1745 = n1744 ^ n1742 ;
  assign n1746 = n1745 ^ x211 ;
  assign n1747 = n311 & n1709 ;
  assign n1748 = n311 & ~n490 ;
  assign n1749 = n1708 & n1748 ;
  assign n1750 = n1749 ^ n490 ;
  assign n1751 = x212 & ~n1750 ;
  assign n1752 = n1747 & n1751 ;
  assign n1753 = n499 & n1752 ;
  assign n1754 = n1753 ^ n1751 ;
  assign n1755 = n1754 ^ x212 ;
  assign n1756 = ~x215 & n1747 ;
  assign n1757 = x87 & n1756 ;
  assign n1758 = x88 & n1747 ;
  assign n1759 = ~n1750 & n1758 ;
  assign n1760 = n1759 ^ n1750 ;
  assign n1761 = n1757 & ~n1760 ;
  assign n1762 = n1761 ^ n1760 ;
  assign n1763 = ~x214 & n1756 ;
  assign n1764 = x86 & n1763 ;
  assign n1765 = n1764 ^ x212 ;
  assign n1766 = ~x212 & ~n1765 ;
  assign n1767 = ~n1762 & n1766 ;
  assign n1768 = n1767 ^ x212 ;
  assign n1769 = ~x85 & x213 ;
  assign n1770 = n1768 & n1769 ;
  assign n1771 = n1770 ^ x213 ;
  assign n1772 = x214 & ~n493 ;
  assign n1773 = n306 & n1772 ;
  assign n1774 = n1762 & n1773 ;
  assign n1775 = n1774 ^ n1772 ;
  assign n1776 = n1775 ^ x214 ;
  assign n1777 = x215 & ~n496 ;
  assign n1778 = n307 & n1777 ;
  assign n1779 = n1760 & n1778 ;
  assign n1780 = n1779 ^ n1777 ;
  assign n1781 = n1780 ^ x215 ;
  assign n1786 = n500 & n1750 ;
  assign n1787 = n1786 ^ n499 ;
  assign n1788 = x216 & n1787 ;
  assign n1789 = n312 & ~n1706 ;
  assign n1797 = n1702 & n1789 ;
  assign n1798 = x92 & n1797 ;
  assign n1799 = n1798 ^ x92 ;
  assign n1790 = n1789 ^ n312 ;
  assign n1791 = n1790 ^ x92 ;
  assign n1800 = n1799 ^ n1791 ;
  assign n1801 = ~n502 & ~n1800 ;
  assign n1802 = ~x219 & n312 ;
  assign n1803 = n1702 & n1802 ;
  assign n1804 = x91 & n1803 ;
  assign n1805 = n1801 & n1804 ;
  assign n1806 = n1805 ^ n1801 ;
  assign n1807 = ~x218 & n1803 ;
  assign n1808 = x90 & n1807 ;
  assign n1809 = n1808 ^ x216 ;
  assign n1810 = ~x216 & ~n1809 ;
  assign n1811 = n1806 & n1810 ;
  assign n1812 = n1811 ^ x216 ;
  assign n1813 = ~x89 & x217 ;
  assign n1814 = n1812 & n1813 ;
  assign n1815 = n1814 ^ x217 ;
  assign n1816 = x218 & ~n505 ;
  assign n1817 = n303 & n1816 ;
  assign n1818 = ~n1806 & n1817 ;
  assign n1819 = n1818 ^ n1816 ;
  assign n1820 = n1819 ^ x218 ;
  assign n1821 = x219 & ~n508 ;
  assign n1822 = n304 & n1821 ;
  assign n1823 = ~n1801 & n1822 ;
  assign n1824 = n1823 ^ n1821 ;
  assign n1825 = n1824 ^ x219 ;
  assign n1826 = x220 & ~n545 ;
  assign n1827 = n321 & n1826 ;
  assign n1828 = n1630 & n1827 ;
  assign n1829 = n1828 ^ n1826 ;
  assign n1830 = n1829 ^ x220 ;
  assign n1831 = n322 & n1628 ;
  assign n1832 = ~x93 & ~n546 ;
  assign n1833 = ~n1831 & n1832 ;
  assign n1834 = n322 & n1609 ;
  assign n1835 = n298 & n664 ;
  assign n1836 = n649 & n1835 ;
  assign n1837 = n1836 ^ n649 ;
  assign n1838 = n1834 & n1837 ;
  assign n1846 = n301 & n1838 ;
  assign n1847 = x95 & n1846 ;
  assign n1848 = n1847 ^ x95 ;
  assign n1839 = n1838 ^ n1834 ;
  assign n1840 = n1839 ^ x95 ;
  assign n1849 = n1848 ^ n1840 ;
  assign n1850 = n1833 & ~n1849 ;
  assign n1851 = n650 & n1834 ;
  assign n1852 = n301 & n1851 ;
  assign n1853 = n1852 ^ x221 ;
  assign n1854 = x221 & n1853 ;
  assign n1855 = n1850 & n1854 ;
  assign n1856 = n1855 ^ x221 ;
  assign n1857 = ~x94 & x222 ;
  assign n1858 = ~x221 & n1857 ;
  assign n1859 = ~n1850 & n1858 ;
  assign n1860 = n1859 ^ n1857 ;
  assign n1861 = n1860 ^ x222 ;
  assign n1862 = n273 & n1834 ;
  assign n1863 = n273 & ~n1833 ;
  assign n1864 = n651 & ~n1863 ;
  assign n1865 = x223 & n1864 ;
  assign n1866 = n1862 & n1865 ;
  assign n1867 = ~n1837 & n1866 ;
  assign n1868 = n1867 ^ n1865 ;
  assign n1869 = n1868 ^ x223 ;
  assign n1870 = ~x96 & x224 ;
  assign n1871 = ~n649 & n1862 ;
  assign n1872 = n1864 & ~n1871 ;
  assign n1873 = ~x223 & n1872 ;
  assign n1877 = n1873 ^ x223 ;
  assign n1874 = n298 & n1862 ;
  assign n1875 = n662 & n1874 ;
  assign n1876 = n1873 & n1875 ;
  assign n1878 = n1877 ^ n1876 ;
  assign n1879 = n1870 & n1878 ;
  assign n1880 = n1879 ^ x224 ;
  assign n1881 = ~x96 & ~x224 ;
  assign n1882 = x98 & n1874 ;
  assign n1884 = n1873 & n1882 ;
  assign n1885 = n1884 ^ n1877 ;
  assign n1886 = n1881 & n1885 ;
  assign n1887 = n1886 ^ x224 ;
  assign n1888 = ~x97 & x225 ;
  assign n1889 = n1887 & n1888 ;
  assign n1890 = n1889 ^ x225 ;
  assign n1891 = n657 & ~n1863 ;
  assign n1892 = ~n1871 & n1891 ;
  assign n1893 = x226 & ~n665 ;
  assign n1894 = ~n1892 & n1893 ;
  assign n1895 = n300 & n1862 ;
  assign n1896 = n286 & n1895 ;
  assign n1897 = n288 & n1896 ;
  assign n1898 = ~x234 & n1897 ;
  assign n1899 = n294 & n1898 ;
  assign n1900 = ~n591 & n1896 ;
  assign n1901 = ~n665 & ~n1891 ;
  assign n1902 = n646 & n1895 ;
  assign n1910 = x110 & n1902 ;
  assign n1911 = n286 & n1910 ;
  assign n1912 = n1911 ^ n286 ;
  assign n1903 = n1902 ^ n1895 ;
  assign n1904 = n1903 ^ n286 ;
  assign n1913 = n1912 ^ n1904 ;
  assign n1914 = ~n1901 & ~n1913 ;
  assign n1915 = ~n1900 & n1914 ;
  assign n1916 = x107 & n1897 ;
  assign n1917 = n1915 & n1916 ;
  assign n1918 = n1917 ^ n1915 ;
  assign n1919 = ~x226 & n1918 ;
  assign n1927 = n1898 & n1919 ;
  assign n1928 = x106 & n1927 ;
  assign n1929 = n1928 ^ x106 ;
  assign n1920 = n1919 ^ x226 ;
  assign n1921 = n1920 ^ x106 ;
  assign n1930 = n1929 ^ n1921 ;
  assign n1931 = ~x99 & n1930 ;
  assign n1932 = x227 & n1931 ;
  assign n1933 = ~n570 & n1932 ;
  assign n1934 = n1899 & n1933 ;
  assign n1935 = n1934 ^ n1932 ;
  assign n1936 = n1935 ^ x227 ;
  assign n1937 = n1899 & n1931 ;
  assign n1938 = ~x105 & ~x232 ;
  assign n1943 = n552 & n555 ;
  assign n1944 = n1943 ^ x104 ;
  assign n1945 = n1938 & n1944 ;
  assign n1946 = n1945 ^ x105 ;
  assign n1947 = n1937 & n1946 ;
  assign n1948 = n1947 ^ n1931 ;
  assign n1949 = ~x100 & ~x227 ;
  assign n1950 = ~n1948 & n1949 ;
  assign n1951 = n1950 ^ x100 ;
  assign n1952 = n557 & n1899 ;
  assign n1953 = n292 & n1952 ;
  assign n1954 = n1953 ^ x228 ;
  assign n1955 = x228 & n1954 ;
  assign n1956 = ~n1951 & n1955 ;
  assign n1957 = n1956 ^ x228 ;
  assign n1958 = ~x101 & ~x228 ;
  assign n1959 = n1951 & n1958 ;
  assign n1960 = n1959 ^ x101 ;
  assign n1961 = ~x229 & n1960 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1963 = ~x102 & x230 ;
  assign n1964 = ~n1961 & n1963 ;
  assign n1965 = n1964 ^ x230 ;
  assign n1966 = n290 & ~n554 ;
  assign n1967 = n1951 & n1966 ;
  assign n1968 = n1967 ^ n554 ;
  assign n1969 = ~x231 & n1968 ;
  assign n1970 = n1969 ^ n1968 ;
  assign n1971 = ~x104 & x232 ;
  assign n1972 = ~n1969 & n1971 ;
  assign n1973 = n1972 ^ x232 ;
  assign n1974 = x233 & n570 ;
  assign n1975 = n293 & n1974 ;
  assign n1976 = ~n1931 & n1975 ;
  assign n1977 = n1976 ^ n1974 ;
  assign n1978 = n1977 ^ x233 ;
  assign n1979 = x234 & n583 ;
  assign n1980 = ~n1918 & n1979 ;
  assign n1981 = n295 & n1980 ;
  assign n1982 = n1981 ^ n1979 ;
  assign n1983 = n1982 ^ x234 ;
  assign n1984 = n296 & ~n585 ;
  assign n1985 = ~n1914 & n1984 ;
  assign n1986 = n1985 ^ n585 ;
  assign n1987 = x235 & ~n1986 ;
  assign n1988 = n1900 & n1987 ;
  assign n1989 = n296 & n1988 ;
  assign n1990 = n1989 ^ n1987 ;
  assign n1991 = n1990 ^ x235 ;
  assign n1992 = x109 & n287 ;
  assign n1993 = n296 & n1992 ;
  assign n1994 = n1896 & n1993 ;
  assign n1995 = ~x108 & ~x235 ;
  assign n1996 = n1986 & n1995 ;
  assign n1997 = n1996 ^ x108 ;
  assign n1998 = ~n1994 & ~n1997 ;
  assign n1999 = x236 & ~n1998 ;
  assign n2000 = ~x109 & x237 ;
  assign n2001 = ~x236 & n2000 ;
  assign n2002 = n1997 & n2001 ;
  assign n2003 = n2002 ^ n2000 ;
  assign n2004 = n2003 ^ x237 ;
  assign n2005 = n297 & n593 ;
  assign n2006 = ~n1914 & n2005 ;
  assign n2007 = n2006 ^ n593 ;
  assign n2008 = ~x238 & ~n2007 ;
  assign n2009 = n2008 ^ n2007 ;
  assign n2010 = ~x111 & x239 ;
  assign n2011 = ~n2008 & n2010 ;
  assign n2012 = n2011 ^ x239 ;
  assign n2013 = n285 & n297 ;
  assign n2014 = n1895 & n2013 ;
  assign n2015 = n643 ^ n297 ;
  assign n2016 = n2015 ^ n285 ;
  assign n2017 = n593 ^ n297 ;
  assign n2018 = n2017 ^ n285 ;
  assign n2019 = n1901 ^ n593 ;
  assign n2020 = n2019 ^ n643 ;
  assign n2021 = n2018 & ~n2020 ;
  assign n2022 = ~n2016 & n2021 ;
  assign n2023 = n2022 ^ n593 ;
  assign n2024 = n2023 ^ n643 ;
  assign n2025 = n285 & ~n2024 ;
  assign n2026 = ~n643 & n2025 ;
  assign n2027 = n2026 ^ n643 ;
  assign n2028 = x240 & ~n2027 ;
  assign n2029 = ~n640 & n2028 ;
  assign n2030 = n2014 & n2029 ;
  assign n2031 = n2030 ^ n2028 ;
  assign n2032 = n2031 ^ x240 ;
  assign n2033 = ~x113 & x241 ;
  assign n2034 = ~n637 & n2014 ;
  assign n2035 = ~n2027 & n2034 ;
  assign n2036 = n2035 ^ n2027 ;
  assign n2037 = n279 & n2014 ;
  assign n2038 = x117 & n2037 ;
  assign n2039 = ~n2036 & n2038 ;
  assign n2040 = n2039 ^ n2036 ;
  assign n2041 = ~x244 & n2037 ;
  assign n2042 = x116 & n2041 ;
  assign n2043 = ~n2040 & n2042 ;
  assign n2044 = n2043 ^ n2040 ;
  assign n2045 = ~x240 & ~n2044 ;
  assign n2049 = n2045 ^ x240 ;
  assign n2046 = ~x243 & n2041 ;
  assign n2047 = n597 & n2046 ;
  assign n2048 = n2045 & n2047 ;
  assign n2050 = n2049 ^ n2048 ;
  assign n2051 = n2033 & n2050 ;
  assign n2052 = n2051 ^ x241 ;
  assign n2053 = ~x113 & ~x241 ;
  assign n2054 = x115 & n2046 ;
  assign n2056 = n2045 & n2054 ;
  assign n2057 = n2056 ^ n2049 ;
  assign n2058 = n2053 & n2057 ;
  assign n2059 = n2058 ^ x241 ;
  assign n2060 = ~x114 & x242 ;
  assign n2061 = n2059 & n2060 ;
  assign n2062 = n2061 ^ x242 ;
  assign n2063 = x243 & ~n599 ;
  assign n2064 = n281 & n2063 ;
  assign n2065 = n2044 & n2064 ;
  assign n2066 = n2065 ^ n2063 ;
  assign n2067 = n2066 ^ x243 ;
  assign n2068 = x244 & ~n602 ;
  assign n2069 = n282 & n2068 ;
  assign n2070 = n2040 & n2069 ;
  assign n2071 = n2070 ^ n2068 ;
  assign n2072 = n2071 ^ x244 ;
  assign n2073 = x245 & ~n605 ;
  assign n2074 = n283 & n2073 ;
  assign n2075 = n2036 & n2074 ;
  assign n2076 = n2075 ^ n2073 ;
  assign n2077 = n2076 ^ x245 ;
  assign n2078 = ~x245 & n283 ;
  assign n2079 = n2014 & n2078 ;
  assign n2080 = n283 ^ x245 ;
  assign n2081 = n2080 ^ x118 ;
  assign n2082 = n605 ^ n283 ;
  assign n2083 = n2082 ^ x118 ;
  assign n2084 = n2027 ^ n605 ;
  assign n2085 = n2084 ^ x245 ;
  assign n2086 = n2083 & n2085 ;
  assign n2087 = n2081 & n2086 ;
  assign n2088 = n2087 ^ n605 ;
  assign n2089 = n2088 ^ x245 ;
  assign n2090 = ~x118 & n2089 ;
  assign n2091 = ~x245 & n2090 ;
  assign n2092 = n2091 ^ x118 ;
  assign n2093 = x246 & ~n2092 ;
  assign n2094 = n2079 & n2093 ;
  assign n2095 = ~n635 & n2094 ;
  assign n2096 = n2095 ^ n2093 ;
  assign n2097 = n2096 ^ x246 ;
  assign n2098 = ~x246 & n2079 ;
  assign n2099 = ~x119 & ~x246 ;
  assign n2100 = n2092 & n2099 ;
  assign n2101 = n2100 ^ x119 ;
  assign n2102 = x247 & ~n2101 ;
  assign n2103 = n2098 & n2102 ;
  assign n2104 = ~n632 & n2103 ;
  assign n2105 = n2104 ^ n2102 ;
  assign n2106 = n2105 ^ x247 ;
  assign n2107 = n276 & n2098 ;
  assign n2108 = ~x247 & ~n2101 ;
  assign n2116 = n2098 & n2108 ;
  assign n2117 = x124 & n2116 ;
  assign n2118 = n2117 ^ x124 ;
  assign n2109 = n2108 ^ x247 ;
  assign n2110 = n2109 ^ x124 ;
  assign n2119 = n2118 ^ n2110 ;
  assign n2120 = ~x120 & n2119 ;
  assign n2121 = x248 & n2120 ;
  assign n2122 = ~n619 & n2121 ;
  assign n2123 = n2107 & n2122 ;
  assign n2124 = n2123 ^ n2121 ;
  assign n2125 = n2124 ^ x248 ;
  assign n2126 = ~x248 & n2120 ;
  assign n2134 = n2107 & n2126 ;
  assign n2135 = x123 & n2134 ;
  assign n2136 = n2135 ^ x123 ;
  assign n2127 = n2126 ^ x248 ;
  assign n2128 = n2127 ^ x123 ;
  assign n2137 = n2136 ^ n2128 ;
  assign n2138 = ~x121 & n2137 ;
  assign n2139 = n274 & n2107 ;
  assign n2140 = x122 & n2139 ;
  assign n2141 = n2140 ^ x249 ;
  assign n2142 = x249 & n2141 ;
  assign n2143 = n2138 & n2142 ;
  assign n2144 = n2143 ^ x249 ;
  assign n2145 = ~x122 & x250 ;
  assign n2146 = ~x249 & n2145 ;
  assign n2147 = ~n2138 & n2146 ;
  assign n2148 = n2147 ^ n2145 ;
  assign n2149 = n2148 ^ x250 ;
  assign n2150 = x251 & n619 ;
  assign n2151 = n275 & n2150 ;
  assign n2152 = ~n2120 & n2151 ;
  assign n2153 = n2152 ^ n2150 ;
  assign n2154 = n2153 ^ x251 ;
  assign n2155 = n347 & n704 ;
  assign n2156 = n1445 & n2155 ;
  assign n2157 = n2156 ^ n704 ;
  assign n2158 = ~x252 & ~n2157 ;
  assign n2159 = n2158 ^ n2157 ;
  assign n2160 = ~x125 & x253 ;
  assign n2161 = ~n2158 & n2160 ;
  assign n2162 = n2161 ^ x253 ;
  assign n2163 = n271 & n704 ;
  assign n2164 = n347 & n1341 ;
  assign n2165 = n1337 & n2164 ;
  assign n2166 = x127 & n2165 ;
  assign n2167 = n2166 ^ n2164 ;
  assign n2168 = n2167 ^ n347 ;
  assign n2169 = n2163 & ~n2168 ;
  assign n2170 = n2169 ^ n271 ;
  assign n2171 = x254 & ~n432 ;
  assign n2172 = ~n2170 & n2171 ;
  assign n2173 = n2172 ^ x254 ;
  assign n2178 = n707 & ~n1341 ;
  assign n2179 = n2178 ^ n706 ;
  assign n2180 = x255 & n2179 ;
  assign n2181 = n348 & n1337 ;
  assign y0 = n839 ;
  assign y1 = n852 ;
  assign y2 = n866 ;
  assign y3 = n872 ;
  assign y4 = n883 ;
  assign y5 = n889 ;
  assign y6 = ~n892 ;
  assign y7 = ~n895 ;
  assign y8 = n898 ;
  assign y9 = n903 ;
  assign y10 = n922 ;
  assign y11 = n945 ;
  assign y12 = n950 ;
  assign y13 = n959 ;
  assign y14 = n979 ;
  assign y15 = n1002 ;
  assign y16 = n1007 ;
  assign y17 = n1012 ;
  assign y18 = n1017 ;
  assign y19 = n1040 ;
  assign y20 = n1045 ;
  assign y21 = n1054 ;
  assign y22 = n1063 ;
  assign y23 = n1072 ;
  assign y24 = n1077 ;
  assign y25 = n1086 ;
  assign y26 = n1095 ;
  assign y27 = n1106 ;
  assign y28 = n1115 ;
  assign y29 = n1138 ;
  assign y30 = n1148 ;
  assign y31 = n1153 ;
  assign y32 = n1162 ;
  assign y33 = n1185 ;
  assign y34 = n1195 ;
  assign y35 = n1200 ;
  assign y36 = n1209 ;
  assign y37 = n1232 ;
  assign y38 = n1242 ;
  assign y39 = n1247 ;
  assign y40 = n1256 ;
  assign y41 = n1271 ;
  assign y42 = n1280 ;
  assign y43 = n1299 ;
  assign y44 = n1308 ;
  assign y45 = n1317 ;
  assign y46 = n1326 ;
  assign y47 = n1331 ;
  assign y48 = n1336 ;
  assign y49 = n1382 ;
  assign y50 = n1387 ;
  assign y51 = n1392 ;
  assign y52 = n1401 ;
  assign y53 = n1417 ;
  assign y54 = n1422 ;
  assign y55 = n1427 ;
  assign y56 = n1434 ;
  assign y57 = n1466 ;
  assign y58 = n1471 ;
  assign y59 = n1476 ;
  assign y60 = n1481 ;
  assign y61 = n1508 ;
  assign y62 = n1513 ;
  assign y63 = n1518 ;
  assign y64 = n1523 ;
  assign y65 = n1543 ;
  assign y66 = n1553 ;
  assign y67 = n1558 ;
  assign y68 = n1563 ;
  assign y69 = n1586 ;
  assign y70 = n1596 ;
  assign y71 = n1601 ;
  assign y72 = n1608 ;
  assign y73 = n1642 ;
  assign y74 = n1647 ;
  assign y75 = n1656 ;
  assign y76 = n1667 ;
  assign y77 = n1676 ;
  assign y78 = n1688 ;
  assign y79 = n1693 ;
  assign y80 = n1700 ;
  assign y81 = n1731 ;
  assign y82 = n1741 ;
  assign y83 = n1746 ;
  assign y84 = n1755 ;
  assign y85 = n1771 ;
  assign y86 = n1776 ;
  assign y87 = n1781 ;
  assign y88 = n1788 ;
  assign y89 = n1815 ;
  assign y90 = n1820 ;
  assign y91 = n1825 ;
  assign y92 = n1830 ;
  assign y93 = n1856 ;
  assign y94 = n1861 ;
  assign y95 = n1869 ;
  assign y96 = n1880 ;
  assign y97 = n1890 ;
  assign y98 = n1894 ;
  assign y99 = n1936 ;
  assign y100 = n1957 ;
  assign y101 = n1962 ;
  assign y102 = n1965 ;
  assign y103 = n1970 ;
  assign y104 = n1973 ;
  assign y105 = n1978 ;
  assign y106 = n1983 ;
  assign y107 = n1991 ;
  assign y108 = n1999 ;
  assign y109 = n2004 ;
  assign y110 = ~n2009 ;
  assign y111 = n2012 ;
  assign y112 = n2032 ;
  assign y113 = n2052 ;
  assign y114 = n2062 ;
  assign y115 = n2067 ;
  assign y116 = n2072 ;
  assign y117 = n2077 ;
  assign y118 = n2097 ;
  assign y119 = n2106 ;
  assign y120 = n2125 ;
  assign y121 = n2144 ;
  assign y122 = n2149 ;
  assign y123 = n2154 ;
  assign y124 = ~n2159 ;
  assign y125 = n2162 ;
  assign y126 = n2173 ;
  assign y127 = n2180 ;
  assign y128 = ~n2181 ;
endmodule
