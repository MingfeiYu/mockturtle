module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, y0, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, y1, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528, n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552, n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677, n_5678, n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705, n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713, n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743, n_5744, n_5745, n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772, n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789, n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907, n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983, n_5984, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208, n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263, n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311, n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319, n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359, n_6360, n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408, n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416, n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424, n_6425, n_6426, n_6427, n_6428, n_6429, n_6430, n_6431, n_6432, n_6433, n_6434, n_6435, n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443, n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457, n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, n_6465, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472, n_6473, n_6474, n_6475, n_6476, n_6477, n_6478, n_6479, n_6480, n_6481, n_6482, n_6483, n_6484, n_6485, n_6486, n_6487, n_6488, n_6489, n_6490, n_6491, n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504, n_6505, n_6506, n_6507, n_6508, n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524, n_6525, n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540, n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556, n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564, n_6565, n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572, n_6573, n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592, n_6593, n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608, n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617, n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704, n_6705, n_6706, n_6707, n_6708, n_6709, n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723, n_6724, n_6725, y2, n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740, n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748, n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764, n_6765, n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772, n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788, n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796, n_6797, n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804, n_6805, n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812, n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820, n_6821, n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828, n_6829, n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6839, n_6840, n_6841, n_6842, n_6843, n_6844, n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853, n_6854, n_6855, n_6856, n_6857, n_6858, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864, n_6865, n_6866, n_6867, n_6868, n_6869, n_6870, n_6871, n_6872, n_6873, n_6874, n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881, n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888, n_6889, n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6898, n_6899, n_6900, n_6901, n_6902, n_6903, n_6904, n_6905, n_6906, n_6907, n_6908, n_6909, n_6910, n_6911, n_6912, n_6913, n_6914, n_6915, n_6916, n_6917, n_6918, n_6919, n_6920, n_6921, n_6922, n_6923, n_6924, n_6925, n_6926, n_6927, n_6928, n_6929, n_6930, n_6931, n_6932, n_6933, n_6934, n_6935, n_6936, n_6937, n_6938, n_6939, n_6940, n_6941, n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948, n_6949, n_6950, n_6951, n_6952, n_6953, n_6954, n_6955, n_6956, n_6957, n_6958, n_6959, n_6960, n_6961, n_6962, n_6963, n_6964, n_6965, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971, n_6972, n_6973, n_6974, n_6975, n_6976, n_6977, n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, n_7003, n_7004, n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012, n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020, n_7021, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030, n_7031, n_7032, n_7033, n_7034, n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041, n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7056, n_7057, n_7058, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065, n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073, n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081, n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089, n_7090, n_7091, n_7092, n_7093, n_7094, n_7095, n_7096, n_7097, n_7098, n_7099, n_7100, n_7101, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108, n_7109, n_7110, n_7111, n_7112, n_7113, n_7114, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129, n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136, n_7137, n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145, n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153, n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7160, n_7161, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172, n_7173, n_7174, y3, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181, n_7182, n_7183, n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198, n_7199, n_7200, n_7201, n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212, n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220, n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228, n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236, n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7256, n_7257, n_7258, n_7259, n_7260, n_7261, n_7262, n_7263, n_7264, n_7265, n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273, n_7274, n_7275, n_7276, n_7277, n_7278, n_7279, n_7280, n_7281, n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288, n_7289, n_7290, n_7291, n_7292, n_7293, n_7294, n_7295, n_7296, n_7297, n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304, n_7305, n_7306, n_7307, n_7308, n_7309, n_7310, n_7311, n_7312, n_7313, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332, n_7333, n_7334, n_7335, n_7336, n_7337, n_7338, n_7339, n_7340, n_7341, n_7342, n_7343, n_7344, n_7345, n_7346, n_7347, n_7348, n_7349, n_7350, n_7351, n_7352, n_7353, n_7354, n_7355, n_7356, n_7357, n_7358, n_7359, n_7360, n_7361, n_7362, n_7363, n_7364, n_7365, n_7366, n_7367, n_7368, n_7369, n_7370, n_7371, n_7372, n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, n_7380, n_7381, n_7382, n_7383, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389, n_7390, n_7391, n_7392, n_7393, n_7394, n_7395, n_7396, n_7397, n_7398, n_7399, n_7400, n_7401, n_7402, n_7403, n_7404, n_7405, n_7406, n_7407, n_7408, n_7409, n_7410, n_7411, n_7412, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7421, n_7422, n_7423, n_7424, n_7425, n_7426, n_7427, n_7428, n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7435, n_7436, n_7437, n_7438, n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7446, n_7447, n_7448, y4, n_7449, n_7450, n_7451, n_7452, n_7453, n_7454, n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461, n_7462, n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469, n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502, n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518, n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541, n_7542, n_7543, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552, n_7553, n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565, n_7566, n_7567, n_7568, n_7569, n_7570, n_7571, n_7572, n_7573, n_7574, n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7584, n_7585, n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596, n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603, n_7604, n_7605, n_7606, n_7607, n_7608, n_7609, n_7610, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625, n_7626, n_7627, n_7628, n_7629, n_7630, n_7631, n_7632, n_7633, n_7634, n_7635, n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643, n_7644, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650, n_7651, n_7652, n_7653, n_7654, n_7655, n_7656, n_7657, n_7658, n_7659, n_7660, n_7661, n_7662, n_7663, n_7664, n_7665, n_7666, n_7667, n_7668, n_7669, n_7670, n_7671, n_7672, n_7673, n_7674, n_7675, n_7676, n_7677, n_7678, n_7679, n_7680, n_7681, n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688, n_7689, n_7690, n_7691, n_7692, n_7693, n_7694, n_7695, n_7696, n_7697, n_7698, n_7699, n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, y5, n_7706, n_7707, n_7708, n_7709, n_7710, n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717, n_7718, n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726, n_7727, n_7728, n_7729, n_7730, n_7731, n_7732, n_7733, n_7734, n_7735, n_7736, n_7737, n_7738, n_7739, n_7740, n_7741, n_7742, n_7743, n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750, n_7751, n_7752, n_7753, n_7754, n_7755, n_7756, n_7757, n_7758, n_7759, n_7760, n_7761, n_7762, n_7763, n_7764, n_7765, n_7766, n_7767, n_7768, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781, n_7782, n_7783, n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7806, n_7807, n_7808, n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816, n_7817, n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824, n_7825, n_7826, n_7827, n_7828, n_7829, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835, n_7836, n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7843, n_7844, n_7845, n_7846, n_7847, n_7848, n_7849, n_7850, n_7851, n_7852, n_7853, n_7854, n_7855, n_7856, n_7857, n_7858, n_7859, n_7860, n_7861, n_7862, n_7863, n_7864, n_7865, n_7866, n_7867, n_7868, n_7869, n_7870, n_7871, n_7872, n_7873, n_7874, n_7875, n_7876, n_7877, n_7878, n_7879, n_7880, n_7881, n_7882, n_7883, n_7884, n_7885, n_7886, n_7887, n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, n_7895, n_7896, n_7897, n_7898, n_7899, n_7900, n_7901, n_7902, n_7903, n_7904, n_7905, n_7906, n_7907, n_7908, n_7909, n_7910, n_7911, n_7912, n_7913, n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920, n_7921, n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928, n_7929, n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937, n_7938, n_7939, n_7940, n_7941, n_7942, n_7943, n_7944, n_7945, n_7946, n_7947, n_7948, n_7949, n_7950, n_7951, n_7952, n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960, n_7961, n_7962, n_7963, n_7964, n_7965, n_7966, n_7967, n_7968, n_7969, n_7970, n_7971, n_7972, n_7973, n_7974, n_7975, n_7976, n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991, n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999, n_8000, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007, n_8008, n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016, n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025, n_8026, n_8027, n_8028, n_8029, n_8030, n_8031, n_8032, n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, n_8039, n_8040, n_8041, n_8042, n_8043, n_8044, n_8045, n_8046, n_8047, n_8048, n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055, n_8056, n_8057, n_8058, n_8059, n_8060, n_8061, n_8062, n_8063, n_8064, n_8065, n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072, n_8073, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080, n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088, n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096, n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104, n_8105, n_8106, y6, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112, n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120, n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128, n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136, n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144, n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152, n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160, n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168, n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176, n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184, n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192, n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200, n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208, n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216, n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224, n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232, n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240, n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248, n_8249, n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256, n_8257, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272, n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280, n_8281, n_8282, n_8283, n_8284, n_8285, n_8286, n_8287, n_8288, n_8289, n_8290, n_8291, n_8292, n_8293, n_8294, n_8295, n_8296, n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304, n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320, n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328, n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354, n_8355, n_8356, n_8357, n_8358, n_8359, n_8360, n_8361, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367, n_8368, n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376, n_8377, n_8378, n_8379, n_8380, n_8381, n_8382, n_8383, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389, n_8390, n_8391, n_8392, n_8393, n_8394, n_8395, n_8396, n_8397, n_8398, n_8399, n_8400, n_8401, n_8402, n_8403, n_8404, n_8405, n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416, n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424, n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432, n_8433, n_8434, n_8435, n_8436, n_8437, y7, n_8438, n_8439, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448, n_8449, n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456, n_8457, n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464, n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472, n_8473, n_8474, n_8475, n_8476, n_8477, n_8478, n_8479, n_8480, n_8481, n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488, n_8489, n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496, n_8497, n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, n_8504, n_8505, n_8506, n_8507, n_8508, n_8509, n_8510, n_8511, n_8512, n_8513, n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528, n_8529, n_8530, n_8531, n_8532, n_8533, n_8534, n_8535, n_8536, n_8537, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544, n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552, n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560, n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568, n_8569, n_8570, n_8571, n_8572, n_8573, n_8574, n_8575, n_8576, n_8577, n_8578, n_8579, n_8580, n_8581, n_8582, n_8583, n_8584, n_8585, n_8586, n_8587, n_8588, n_8589, n_8590, n_8591, n_8592, n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600, n_8601, n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613, n_8614, n_8615, n_8616, n_8617, n_8618, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8625, n_8626, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632, n_8633, n_8634, n_8635, n_8636, n_8637, n_8638, n_8639, n_8640, n_8641, n_8642, n_8643, n_8644, n_8645, n_8646, n_8647, n_8648, n_8649, n_8650, n_8651, n_8652, n_8653, n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8660, n_8661, n_8662, n_8663, n_8664, n_8665, n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, n_8672, n_8673, n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681, n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689, n_8690, n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697, n_8698, n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705, n_8706, n_8707, n_8708, n_8709, n_8710, n_8711, n_8712, n_8713, n_8714, n_8715, n_8716, n_8717, n_8718, n_8719, n_8720, n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727, n_8728, n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735, n_8736, n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743, n_8744, n_8745, n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8752, n_8753, n_8754, n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761, n_8762, n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769, n_8770, n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777, n_8778, n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786, n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793, n_8794, n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802, n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8809, n_8810, n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817, n_8818, y8, n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, n_8825, n_8826, n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833, n_8834, n_8835, n_8836, n_8837, n_8838, n_8839, n_8840, n_8841, n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8848, n_8849, n_8850, n_8851, n_8852, n_8853, n_8854, n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861, n_8862, n_8863, n_8864, n_8865, n_8866, n_8867, n_8868, n_8869, n_8870, n_8871, n_8872, n_8873, n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881, n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889, n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897, n_8898, n_8899, n_8900, n_8901, n_8902, n_8903, n_8904, n_8905, n_8906, n_8907, n_8908, n_8909, n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916, n_8917, n_8918, n_8919, n_8920, n_8921, n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928, n_8929, n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936, n_8937, n_8938, n_8939, n_8940, n_8941, n_8942, n_8943, n_8944, n_8945, n_8946, n_8947, n_8948, n_8949, n_8950, n_8951, n_8952, n_8953, n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960, n_8961, n_8962, n_8963, n_8964, n_8965, n_8966, n_8967, n_8968, n_8969, n_8970, n_8971, n_8972, n_8973, n_8974, n_8975, n_8976, n_8977, n_8978, n_8979, n_8980, n_8981, n_8982, n_8983, n_8984, n_8985, n_8986, n_8987, n_8988, n_8989, n_8990, n_8991, n_8992, n_8993, n_8994, n_8995, n_8996, n_8997, n_8998, n_8999, n_9000, n_9001, n_9002, n_9003, n_9004, n_9005, n_9006, n_9007, n_9008, n_9009, n_9010, n_9011, n_9012, n_9013, n_9014, n_9015, n_9016, n_9017, n_9018, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024, n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032, n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040, n_9041, n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048, n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056, n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9064, n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071, n_9072, n_9073, n_9074, n_9075, n_9076, n_9077, n_9078, n_9079, n_9080, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087, n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095, n_9096, n_9097, n_9098, n_9099, n_9100, n_9101, n_9102, n_9103, n_9104, n_9105, n_9106, n_9107, n_9108, n_9109, n_9110, n_9111, n_9112, n_9113, n_9114, n_9115, n_9116, n_9117, n_9118, n_9119, n_9120, n_9121, n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128, n_9129, n_9130, n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137, n_9138, n_9139, n_9140, n_9141, n_9142, n_9143, n_9144, n_9145, n_9146, n_9147, n_9148, n_9149, n_9150, n_9151, n_9152, n_9153, n_9154, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160, n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9168, n_9169, n_9170, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176, n_9177, n_9178, n_9179, n_9180, n_9181, n_9182, n_9183, n_9184, n_9185, n_9186, n_9187, n_9188, n_9189, n_9190, n_9191, n_9192, n_9193, n_9194, n_9195, n_9196, n_9197, n_9198, n_9199, n_9200, n_9201, n_9202, n_9203, n_9204, n_9205, n_9206, n_9207, n_9208, n_9209, n_9210, n_9211, n_9212, n_9213, n_9214, n_9215, n_9216, n_9217, n_9218, n_9219, n_9220, n_9221, n_9222, n_9223, n_9224, n_9225, n_9226, n_9227, n_9228, n_9229, n_9230, n_9231, n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9239, y9, n_9240, n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9247, n_9248, n_9249, n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256, n_9257, n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265, n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, n_9273, n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281, n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288, n_9289, n_9290, n_9291, n_9292, n_9293, n_9294, n_9295, n_9296, n_9297, n_9298, n_9299, n_9300, n_9301, n_9302, n_9303, n_9304, n_9305, n_9306, n_9307, n_9308, n_9309, n_9310, n_9311, n_9312, n_9313, n_9314, n_9315, n_9316, n_9317, n_9318, n_9319, n_9320, n_9321, n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9328, n_9329, n_9330, n_9331, n_9332, n_9333, n_9334, n_9335, n_9336, n_9337, n_9338, n_9339, n_9340, n_9341, n_9342, n_9343, n_9344, n_9345, n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353, n_9354, n_9355, n_9356, n_9357, n_9358, n_9359, n_9360, n_9361, n_9362, n_9363, n_9364, n_9365, n_9366, n_9367, n_9368, n_9369, n_9370, n_9371, n_9372, n_9373, n_9374, n_9375, n_9376, n_9377, n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9384, n_9385, n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396, n_9397, n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405, n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413, n_9414, n_9415, n_9416, n_9417, n_9418, n_9419, n_9420, n_9421, n_9422, n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430, n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438, n_9439, n_9440, n_9441, n_9442, n_9443, n_9444, n_9445, n_9446, n_9447, n_9448, n_9449, n_9450, n_9451, n_9452, n_9453, n_9454, n_9455, n_9456, n_9457, n_9458, n_9459, n_9460, n_9461, n_9462, n_9463, n_9464, n_9465, n_9466, n_9467, n_9468, n_9469, n_9470, n_9471, n_9472, n_9473, n_9474, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480, n_9481, n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489, n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496, n_9497, n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504, n_9505, n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512, n_9513, n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520, n_9521, n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, n_9528, n_9529, n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536, n_9537, n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545, n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552, n_9553, n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561, n_9562, n_9563, n_9564, n_9565, n_9566, n_9567, n_9568, n_9569, n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576, n_9577, n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584, n_9585, n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, n_9596, n_9597, n_9598, n_9599, n_9600, n_9601, n_9602, n_9603, n_9604, n_9605, n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612, n_9613, n_9614, n_9615, n_9616, n_9617, n_9618, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624, n_9625, n_9626, n_9627, n_9628, n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635, n_9636, n_9637, n_9638, n_9639, n_9640, n_9641, n_9642, n_9643, n_9644, n_9645, n_9646, n_9647, n_9648, n_9649, n_9650, n_9651, n_9652, n_9653, n_9654, n_9655, n_9656, n_9657, n_9658, n_9659, n_9660, n_9661, n_9662, n_9663, n_9664, n_9665, n_9666, n_9667, y10, n_9668, n_9669, n_9670, n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677, n_9678, n_9679, n_9680, n_9681, n_9682, n_9683, n_9684, n_9685, n_9686, n_9687, n_9688, n_9689, n_9690, n_9691, n_9692, n_9693, n_9694, n_9695, n_9696, n_9697, n_9698, n_9699, n_9700, n_9701, n_9702, n_9703, n_9704, n_9705, n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712, n_9713, n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720, n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728, n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736, n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744, n_9745, n_9746, n_9747, n_9748, n_9749, n_9750, n_9751, n_9752, n_9753, n_9754, n_9755, n_9756, n_9757, n_9758, n_9759, n_9760, n_9761, n_9762, n_9763, n_9764, n_9765, n_9766, n_9767, n_9768, n_9769, n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776, n_9777, n_9778, n_9779, n_9780, n_9781, n_9782, n_9783, n_9784, n_9785, n_9786, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792, n_9793, n_9794, n_9795, n_9796, n_9797, n_9798, n_9799, n_9800, n_9801, n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808, n_9809, n_9810, n_9811, n_9812, n_9813, n_9814, n_9815, n_9816, n_9817, n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_9825, n_9826, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832, n_9833, n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848, n_9849, n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856, n_9857, n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864, n_9865, n_9866, n_9867, n_9868, n_9869, n_9870, n_9871, n_9872, n_9873, n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880, n_9881, n_9882, n_9883, n_9884, n_9885, n_9886, n_9887, n_9888, n_9889, n_9890, n_9891, n_9892, n_9893, n_9894, n_9895, n_9896, n_9897, n_9898, n_9899, n_9900, n_9901, n_9902, n_9903, n_9904, n_9905, n_9906, n_9907, n_9908, n_9909, n_9910, n_9911, n_9912, n_9913, n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920, n_9921, n_9922, n_9923, n_9924, n_9925, n_9926, n_9927, n_9928, n_9929, n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937, n_9938, n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945, n_9946, n_9947, n_9948, n_9949, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955, n_9956, n_9957, n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964, n_9965, n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972, n_9973, n_9974, n_9975, n_9976, n_9977, n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984, n_9985, n_9986, n_9987, n_9988, n_9989, n_9990, n_9991, n_9992, n_9993, n_9994, n_9995, n_9996, n_9997, n_9998, n_9999, n_10000, n_10001, n_10002, n_10003, n_10004, n_10005, n_10006, n_10007, n_10008, n_10009, n_10010, n_10011, n_10012, n_10013, n_10014, n_10015, n_10016, n_10017, n_10018, n_10019, n_10020, n_10021, n_10022, n_10023, n_10024, n_10025, n_10026, n_10027, n_10028, n_10029, n_10030, n_10031, n_10032, n_10033, n_10034, n_10035, n_10036, n_10037, n_10038, n_10039, n_10040, n_10041, n_10042, n_10043, n_10044, n_10045, n_10046, n_10047, n_10048, n_10049, n_10050, n_10051, n_10052, n_10053, n_10054, n_10055, n_10056, n_10057, n_10058, n_10059, n_10060, n_10061, n_10062, n_10063, n_10064, n_10065, n_10066, n_10067, n_10068, n_10069, n_10070, n_10071, n_10072, n_10073, n_10074, n_10075, n_10076, n_10077, n_10078, n_10079, n_10080, n_10081, n_10082, n_10083, n_10084, n_10085, n_10086, n_10087, n_10088, n_10089, n_10090, n_10091, n_10092, n_10093, y11, n_10094, n_10095, n_10096, n_10097, n_10098, n_10099, n_10100, n_10101, n_10102, n_10103, n_10104, n_10105, n_10106, n_10107, n_10108, n_10109, n_10110, n_10111, n_10112, n_10113, n_10114, n_10115, n_10116, n_10117, n_10118, n_10119, n_10120, n_10121, n_10122, n_10123, n_10124, n_10125, n_10126, n_10127, n_10128, n_10129, n_10130, n_10131, n_10132, n_10133, n_10134, n_10135, n_10136, n_10137, n_10138, n_10139, n_10140, n_10141, n_10142, n_10143, n_10144, n_10145, n_10146, n_10147, n_10148, n_10149, n_10150, n_10151, n_10152, n_10153, n_10154, n_10155, n_10156, n_10157, n_10158, n_10159, n_10160, n_10161, n_10162, n_10163, n_10164, n_10165, n_10166, n_10167, n_10168, n_10169, n_10170, n_10171, n_10172, n_10173, n_10174, n_10175, n_10176, n_10177, n_10178, n_10179, n_10180, n_10181, n_10182, n_10183, n_10184, n_10185, n_10186, n_10187, n_10188, n_10189, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195, n_10196, n_10197, n_10198, n_10199, n_10200, n_10201, n_10202, n_10203, n_10204, n_10205, n_10206, n_10207, n_10208, n_10209, n_10210, n_10211, n_10212, n_10213, n_10214, n_10215, n_10216, n_10217, n_10218, n_10219, n_10220, n_10221, n_10222, n_10223, n_10224, n_10225, n_10226, n_10227, n_10228, n_10229, n_10230, n_10231, n_10232, n_10233, n_10234, n_10235, n_10236, n_10237, n_10238, n_10239, n_10240, n_10241, n_10242, n_10243, n_10244, n_10245, n_10246, n_10247, n_10248, n_10249, n_10250, n_10251, n_10252, n_10253, n_10254, n_10255, n_10256, n_10257, n_10258, n_10259, n_10260, n_10261, n_10262, n_10263, n_10264, n_10265, n_10266, n_10267, n_10268, n_10269, n_10270, n_10271, n_10272, n_10273, n_10274, n_10275, n_10276, n_10277, n_10278, n_10279, n_10280, n_10281, n_10282, n_10283, n_10284, n_10285, n_10286, n_10287, n_10288, n_10289, n_10290, n_10291, n_10292, n_10293, n_10294, n_10295, n_10296, n_10297, n_10298, n_10299, n_10300, n_10301, n_10302, n_10303, n_10304, n_10305, n_10306, n_10307, n_10308, n_10309, n_10310, n_10311, n_10312, n_10313, n_10314, n_10315, n_10316, n_10317, n_10318, n_10319, n_10320, n_10321, n_10322, n_10323, n_10324, n_10325, n_10326, n_10327, n_10328, n_10329, n_10330, n_10331, n_10332, n_10333, n_10334, n_10335, n_10336, n_10337, n_10338, n_10339, n_10340, n_10341, n_10342, n_10343, n_10344, n_10345, n_10346, n_10347, n_10348, n_10349, n_10350, n_10351, n_10352, n_10353, n_10354, n_10355, n_10356, n_10357, n_10358, n_10359, n_10360, n_10361, n_10362, n_10363, n_10364, n_10365, n_10366, n_10367, n_10368, n_10369, n_10370, n_10371, n_10372, n_10373, n_10374, n_10375, n_10376, n_10377, n_10378, n_10379, n_10380, n_10381, n_10382, n_10383, n_10384, n_10385, n_10386, n_10387, n_10388, n_10389, n_10390, n_10391, n_10392, n_10393, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399, n_10400, n_10401, n_10402, n_10403, n_10404, n_10405, n_10406, n_10407, n_10408, n_10409, n_10410, n_10411, n_10412, n_10413, n_10414, n_10415, n_10416, n_10417, n_10418, n_10419, n_10420, n_10421, n_10422, n_10423, n_10424, n_10425, n_10426, n_10427, n_10428, n_10429, n_10430, n_10431, n_10432, n_10433, n_10434, n_10435, n_10436, n_10437, n_10438, n_10439, n_10440, n_10441, n_10442, n_10443, n_10444, n_10445, n_10446, n_10447, n_10448, n_10449, n_10450, n_10451, n_10452, n_10453, n_10454, n_10455, n_10456, n_10457, n_10458, n_10459, n_10460, n_10461, n_10462, n_10463, n_10464, n_10465, n_10466, n_10467, n_10468, n_10469, n_10470, n_10471, n_10472, n_10473, n_10474, n_10475, n_10476, n_10477, n_10478, n_10479, n_10480, n_10481, y12, n_10482, n_10483, n_10484, n_10485, n_10486, n_10487, n_10488, n_10489, n_10490, n_10491, n_10492, n_10493, n_10494, n_10495, n_10496, n_10497, n_10498, n_10499, n_10500, n_10501, n_10502, n_10503, n_10504, n_10505, n_10506, n_10507, n_10508, n_10509, n_10510, n_10511, n_10512, n_10513, n_10514, n_10515, n_10516, n_10517, n_10518, n_10519, n_10520, n_10521, n_10522, n_10523, n_10524, n_10525, n_10526, n_10527, n_10528, n_10529, n_10530, n_10531, n_10532, n_10533, n_10534, n_10535, n_10536, n_10537, n_10538, n_10539, n_10540, n_10541, n_10542, n_10543, n_10544, n_10545, n_10546, n_10547, n_10548, n_10549, n_10550, n_10551, n_10552, n_10553, n_10554, n_10555, n_10556, n_10557, n_10558, n_10559, n_10560, n_10561, n_10562, n_10563, n_10564, n_10565, n_10566, n_10567, n_10568, n_10569, n_10570, n_10571, n_10572, n_10573, n_10574, n_10575, n_10576, n_10577, n_10578, n_10579, n_10580, n_10581, n_10582, n_10583, n_10584, n_10585, n_10586, n_10587, n_10588, n_10589, n_10590, n_10591, n_10592, n_10593, n_10594, n_10595, n_10596, n_10597, n_10598, n_10599, n_10600, n_10601, n_10602, n_10603, n_10604, n_10605, n_10606, n_10607, n_10608, n_10609, n_10610, n_10611, n_10612, n_10613, n_10614, n_10615, n_10616, n_10617, n_10618, n_10619, n_10620, n_10621, n_10622, n_10623, n_10624, n_10625, n_10626, n_10627, n_10628, n_10629, n_10630, n_10631, n_10632, n_10633, n_10634, n_10635, n_10636, n_10637, n_10638, n_10639, n_10640, n_10641, n_10642, n_10643, n_10644, n_10645, n_10646, n_10647, n_10648, n_10649, n_10650, n_10651, n_10652, n_10653, n_10654, n_10655, n_10656, n_10657, n_10658, n_10659, n_10660, n_10661, n_10662, n_10663, n_10664, n_10665, n_10666, n_10667, n_10668, n_10669, n_10670, n_10671, n_10672, n_10673, n_10674, n_10675, n_10676, n_10677, n_10678, n_10679, n_10680, n_10681, n_10682, n_10683, n_10684, n_10685, n_10686, n_10687, n_10688, n_10689, n_10690, n_10691, n_10692, n_10693, n_10694, n_10695, n_10696, n_10697, n_10698, n_10699, n_10700, n_10701, n_10702, n_10703, n_10704, n_10705, n_10706, n_10707, n_10708, n_10709, n_10710, n_10711, n_10712, n_10713, n_10714, n_10715, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721, n_10722, n_10723, n_10724, n_10725, n_10726, n_10727, n_10728, n_10729, n_10730, n_10731, n_10732, n_10733, n_10734, n_10735, n_10736, n_10737, n_10738, n_10739, n_10740, n_10741, n_10742, n_10743, n_10744, n_10745, n_10746, n_10747, n_10748, n_10749, n_10750, n_10751, n_10752, n_10753, n_10754, n_10755, n_10756, n_10757, n_10758, n_10759, n_10760, n_10761, n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768, n_10769, n_10770, n_10771, n_10772, n_10773, n_10774, n_10775, n_10776, n_10777, n_10778, n_10779, n_10780, n_10781, n_10782, n_10783, n_10784, n_10785, n_10786, n_10787, n_10788, n_10789, n_10790, n_10791, n_10792, n_10793, n_10794, n_10795, n_10796, n_10797, n_10798, n_10799, n_10800, n_10801, n_10802, n_10803, n_10804, n_10805, n_10806, n_10807, n_10808, n_10809, n_10810, n_10811, n_10812, n_10813, n_10814, n_10815, n_10816, n_10817, n_10818, n_10819, n_10820, n_10821, n_10822, n_10823, n_10824, n_10825, n_10826, n_10827, n_10828, n_10829, n_10830, n_10831, n_10832, n_10833, n_10834, n_10835, n_10836, y13, n_10837, n_10838, n_10839, n_10840, n_10841, n_10842, n_10843, n_10844, n_10845, n_10846, n_10847, n_10848, n_10849, n_10850, n_10851, n_10852, n_10853, n_10854, n_10855, n_10856, n_10857, n_10858, n_10859, n_10860, n_10861, n_10862, n_10863, n_10864, n_10865, n_10866, n_10867, n_10868, n_10869, n_10870, n_10871, n_10872, n_10873, n_10874, n_10875, n_10876, n_10877, n_10878, n_10879, n_10880, n_10881, n_10882, n_10883, n_10884, n_10885, n_10886, n_10887, n_10888, n_10889, n_10890, n_10891, n_10892, n_10893, n_10894, n_10895, n_10896, n_10897, n_10898, n_10899, n_10900, n_10901, n_10902, n_10903, n_10904, n_10905, n_10906, n_10907, n_10908, n_10909, n_10910, n_10911, n_10912, n_10913, n_10914, n_10915, n_10916, n_10917, n_10918, n_10919, n_10920, n_10921, n_10922, n_10923, n_10924, n_10925, n_10926, n_10927, n_10928, n_10929, n_10930, n_10931, n_10932, n_10933, n_10934, n_10935, n_10936, n_10937, n_10938, n_10939, n_10940, n_10941, n_10942, n_10943, n_10944, n_10945, n_10946, n_10947, n_10948, n_10949, n_10950, n_10951, n_10952, n_10953, n_10954, n_10955, n_10956, n_10957, n_10958, n_10959, n_10960, n_10961, n_10962, n_10963, n_10964, n_10965, n_10966, n_10967, n_10968, n_10969, n_10970, n_10971, n_10972, n_10973, n_10974, n_10975, n_10976, n_10977, n_10978, n_10979, n_10980, n_10981, n_10982, n_10983, n_10984, n_10985, n_10986, n_10987, n_10988, n_10989, n_10990, n_10991, n_10992, n_10993, n_10994, n_10995, n_10996, n_10997, n_10998, n_10999, n_11000, n_11001, n_11002, n_11003, n_11004, n_11005, n_11006, n_11007, n_11008, n_11009, n_11010, n_11011, n_11012, n_11013, n_11014, n_11015, n_11016, n_11017, n_11018, n_11019, n_11020, n_11021, n_11022, n_11023, n_11024, n_11025, n_11026, n_11027, n_11028, n_11029, n_11030, n_11031, n_11032, n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, n_11039, n_11040, n_11041, n_11042, n_11043, n_11044, n_11045, n_11046, n_11047, n_11048, n_11049, n_11050, n_11051, n_11052, n_11053, n_11054, n_11055, n_11056, n_11057, n_11058, n_11059, n_11060, n_11061, n_11062, n_11063, n_11064, n_11065, n_11066, n_11067, n_11068, n_11069, n_11070, n_11071, n_11072, n_11073, n_11074, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080, n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087, n_11088, n_11089, n_11090, n_11091, n_11092, n_11093, n_11094, n_11095, n_11096, n_11097, n_11098, n_11099, n_11100, n_11101, n_11102, n_11103, n_11104, n_11105, y14, n_11106, n_11107, n_11108, n_11109, n_11110, n_11111, n_11112, n_11113, n_11114, n_11115, n_11116, n_11117, n_11118, n_11119, n_11120, n_11121, n_11122, n_11123, n_11124, n_11125, n_11126, n_11127, n_11128, n_11129, n_11130, n_11131, n_11132, n_11133, n_11134, n_11135, n_11136, n_11137, n_11138, n_11139, n_11140, n_11141, n_11142, n_11143, n_11144, n_11145, n_11146, n_11147, n_11148, n_11149, n_11150, n_11151, n_11152, n_11153, n_11154, n_11155, n_11156, n_11157, n_11158, n_11159, n_11160, n_11161, n_11162, n_11163, n_11164, n_11165, n_11166, n_11167, n_11168, n_11169, n_11170, n_11171, n_11172, n_11173, n_11174, n_11175, n_11176, n_11177, n_11178, n_11179, n_11180, n_11181, n_11182, n_11183, n_11184, n_11185, n_11186, n_11187, n_11188, n_11189, n_11190, n_11191, n_11192, n_11193, n_11194, n_11195, n_11196, n_11197, n_11198, n_11199, n_11200, n_11201, n_11202, n_11203, n_11204, n_11205, n_11206, n_11207, n_11208, n_11209, n_11210, n_11211, n_11212, n_11213, n_11214, n_11215, n_11216, n_11217, n_11218, n_11219, n_11220, n_11221, n_11222, n_11223, n_11224, n_11225, n_11226, n_11227, n_11228, n_11229, n_11230, n_11231, n_11232, n_11233, n_11234, n_11235, n_11236, n_11237, n_11238, n_11239, n_11240, n_11241, n_11242, n_11243, n_11244, n_11245, n_11246, n_11247, n_11248, n_11249, n_11250, n_11251, n_11252, n_11253, n_11254, n_11255, n_11256, n_11257, n_11258, n_11259, n_11260, n_11261, n_11262, n_11263, n_11264, n_11265, n_11266, n_11267, n_11268, n_11269, n_11270, n_11271, n_11272, n_11273, n_11274, n_11275, n_11276, n_11277, n_11278, n_11279, n_11280, n_11281, n_11282, n_11283, n_11284, n_11285, n_11286, n_11287, n_11288, n_11289, n_11290, n_11291, n_11292, n_11293, n_11294, n_11295, n_11296, n_11297, n_11298, n_11299, n_11300, n_11301, n_11302, n_11303, n_11304, n_11305, n_11306, n_11307, n_11308, n_11309, n_11310, n_11311, n_11312, n_11313, n_11314, n_11315, n_11316, n_11317, n_11318, n_11319, n_11320, n_11321, n_11322, n_11323, n_11324, n_11325, n_11326, n_11327, n_11328, n_11329, n_11330, n_11331, n_11332, n_11333, n_11334, n_11335, n_11336, n_11337, n_11338, n_11339, n_11340, n_11341, n_11342, n_11343, n_11344, n_11345, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351, n_11352, n_11353, n_11354, n_11355, n_11356, n_11357, n_11358, n_11359, n_11360, n_11361, n_11362, n_11363, n_11364, n_11365, n_11366, n_11367, n_11368, n_11369, n_11370, n_11371, n_11372, n_11373, n_11374, n_11375, n_11376, y15, n_11377, n_11378, n_11379, n_11380, n_11381, n_11382, n_11383, n_11384, n_11385, n_11386, n_11387, n_11388, n_11389, n_11390, n_11391, n_11392, n_11393, n_11394, n_11395, n_11396, n_11397, n_11398, n_11399, n_11400, n_11401, n_11402, n_11403, n_11404, n_11405, n_11406, n_11407, n_11408, n_11409, n_11410, n_11411, n_11412, n_11413, n_11414, n_11415, n_11416, n_11417, n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424, n_11425, n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432, n_11433, n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440, n_11441, n_11442, n_11443, n_11444, n_11445, n_11446, n_11447, n_11448, n_11449, n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11456, n_11457, n_11458, n_11459, n_11460, n_11461, n_11462, n_11463, n_11464, n_11465, n_11466, n_11467, n_11468, n_11469, n_11470, n_11471, n_11472, n_11473, n_11474, n_11475, n_11476, n_11477, n_11478, n_11479, n_11480, n_11481, n_11482, n_11483, n_11484, n_11485, n_11486, n_11487, n_11488, n_11489, n_11490, n_11491, n_11492, n_11493, n_11494, n_11495, n_11496, n_11497, n_11498, n_11499, n_11500, n_11501, n_11502, n_11503, n_11504, n_11505, n_11506, n_11507, n_11508, n_11509, n_11510, n_11511, n_11512, n_11513, n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520, n_11521, n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528, n_11529, n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536, n_11537, n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544, n_11545, n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552, n_11553, n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560, n_11561, n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568, n_11569, n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576, n_11577, n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584, n_11585, n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592, n_11593, n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600, n_11601, n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11608, n_11609, n_11610, n_11611, n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618, n_11619, n_11620, n_11621, n_11622, n_11623, n_11624, n_11625, n_11626, n_11627, n_11628, n_11629, n_11630, n_11631, n_11632, n_11633, n_11634, n_11635, n_11636, n_11637, n_11638, n_11639, n_11640, n_11641, n_11642, n_11643, n_11644, n_11645, n_11646, n_11647, n_11648, n_11649, n_11650, n_11651, n_11652, n_11653, n_11654, n_11655, n_11656, n_11657, n_11658, n_11659, n_11660, n_11661, n_11662, n_11663, n_11664, n_11665, n_11666, n_11667, n_11668, n_11669, n_11670, n_11671, n_11672, n_11673, n_11674, n_11675, n_11676, n_11677, n_11678, n_11679, n_11680, n_11681, n_11682, n_11683, n_11684, n_11685, n_11686, n_11687, y16, n_11688, n_11689, n_11690, n_11691, n_11692, n_11693, n_11694, n_11695, n_11696, n_11697, n_11698, n_11699, n_11700, n_11701, n_11702, n_11703, n_11704, n_11705, n_11706, n_11707, n_11708, n_11709, n_11710, n_11711, n_11712, n_11713, n_11714, n_11715, n_11716, n_11717, n_11718, n_11719, n_11720, n_11721, n_11722, n_11723, n_11724, n_11725, n_11726, n_11727, n_11728, n_11729, n_11730, n_11731, n_11732, n_11733, n_11734, n_11735, n_11736, n_11737, n_11738, n_11739, n_11740, n_11741, n_11742, n_11743, n_11744, n_11745, n_11746, n_11747, n_11748, n_11749, n_11750, n_11751, n_11752, n_11753, n_11754, n_11755, n_11756, n_11757, n_11758, n_11759, n_11760, n_11761, n_11762, n_11763, n_11764, n_11765, n_11766, n_11767, n_11768, n_11769, n_11770, n_11771, n_11772, n_11773, n_11774, n_11775, n_11776, n_11777, n_11778, n_11779, n_11780, n_11781, n_11782, n_11783, n_11784, n_11785, n_11786, n_11787, n_11788, n_11789, n_11790, n_11791, n_11792, n_11793, n_11794, n_11795, n_11796, n_11797, n_11798, n_11799, n_11800, n_11801, n_11802, n_11803, n_11804, n_11805, n_11806, n_11807, n_11808, n_11809, n_11810, n_11811, n_11812, n_11813, n_11814, n_11815, n_11816, n_11817, n_11818, n_11819, n_11820, n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827, n_11828, n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835, n_11836, n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843, n_11844, n_11845, n_11846, n_11847, n_11848, n_11849, n_11850, n_11851, n_11852, n_11853, n_11854, n_11855, n_11856, n_11857, n_11858, n_11859, n_11860, n_11861, n_11862, n_11863, n_11864, n_11865, n_11866, n_11867, n_11868, n_11869, n_11870, n_11871, n_11872, n_11873, n_11874, n_11875, n_11876, n_11877, n_11878, n_11879, n_11880, n_11881, n_11882, n_11883, n_11884, n_11885, n_11886, n_11887, n_11888, n_11889, n_11890, n_11891, n_11892, n_11893, n_11894, n_11895, n_11896, n_11897, n_11898, n_11899, n_11900, n_11901, n_11902, n_11903, n_11904, n_11905, n_11906, n_11907, n_11908, n_11909, n_11910, n_11911, n_11912, n_11913, n_11914, n_11915, n_11916, n_11917, n_11918, n_11919, n_11920, n_11921, n_11922, n_11923, n_11924, n_11925, n_11926, n_11927, n_11928, n_11929, n_11930, n_11931, n_11932, y17, n_11933, n_11934, n_11935, n_11936, n_11937, n_11938, n_11939, n_11940, n_11941, n_11942, n_11943, n_11944, n_11945, n_11946, n_11947, n_11948, n_11949, n_11950, n_11951, n_11952, n_11953, n_11954, n_11955, n_11956, n_11957, n_11958, n_11959, n_11960, n_11961, n_11962, n_11963, n_11964, n_11965, n_11966, n_11967, n_11968, n_11969, n_11970, n_11971, n_11972, n_11973, n_11974, n_11975, n_11976, n_11977, n_11978, n_11979, n_11980, n_11981, n_11982, n_11983, n_11984, n_11985, n_11986, n_11987, n_11988, n_11989, n_11990, n_11991, n_11992, n_11993, n_11994, n_11995, n_11996, n_11997, n_11998, n_11999, n_12000, n_12001, n_12002, n_12003, n_12004, n_12005, n_12006, n_12007, n_12008, n_12009, n_12010, n_12011, n_12012, n_12013, n_12014, n_12015, n_12016, n_12017, n_12018, n_12019, n_12020, n_12021, n_12022, n_12023, n_12024, n_12025, n_12026, n_12027, n_12028, n_12029, n_12030, n_12031, n_12032, n_12033, n_12034, n_12035, n_12036, n_12037, n_12038, n_12039, n_12040, n_12041, n_12042, n_12043, n_12044, n_12045, n_12046, n_12047, n_12048, n_12049, n_12050, n_12051, n_12052, n_12053, n_12054, n_12055, n_12056, n_12057, n_12058, n_12059, n_12060, n_12061, n_12062, n_12063, n_12064, n_12065, n_12066, n_12067, n_12068, n_12069, n_12070, n_12071, n_12072, n_12073, n_12074, n_12075, n_12076, n_12077, n_12078, n_12079, n_12080, n_12081, n_12082, n_12083, n_12084, n_12085, n_12086, n_12087, n_12088, n_12089, n_12090, n_12091, n_12092, n_12093, n_12094, n_12095, n_12096, n_12097, n_12098, n_12099, n_12100, n_12101, n_12102, n_12103, n_12104, n_12105, n_12106, n_12107, n_12108, n_12109, n_12110, n_12111, n_12112, n_12113, n_12114, n_12115, n_12116, n_12117, n_12118, n_12119, n_12120, n_12121, n_12122, n_12123, n_12124, n_12125, n_12126, n_12127, n_12128, n_12129, n_12130, n_12131, n_12132, n_12133, n_12134, n_12135, n_12136, n_12137, n_12138, n_12139, n_12140, n_12141, n_12142, n_12143, y18, n_12144, n_12145, n_12146, n_12147, n_12148, n_12149, n_12150, n_12151, n_12152, n_12153, n_12154, n_12155, n_12156, n_12157, n_12158, n_12159, n_12160, n_12161, n_12162, n_12163, n_12164, n_12165, n_12166, n_12167, n_12168, n_12169, n_12170, n_12171, n_12172, n_12173, n_12174, n_12175, n_12176, n_12177, n_12178, n_12179, n_12180, n_12181, n_12182, n_12183, n_12184, n_12185, n_12186, n_12187, n_12188, n_12189, n_12190, n_12191, n_12192, n_12193, n_12194, n_12195, n_12196, n_12197, n_12198, n_12199, n_12200, n_12201, n_12202, n_12203, n_12204, n_12205, n_12206, n_12207, n_12208, n_12209, n_12210, n_12211, n_12212, n_12213, n_12214, n_12215, n_12216, n_12217, n_12218, n_12219, n_12220, n_12221, n_12222, n_12223, n_12224, n_12225, n_12226, n_12227, n_12228, n_12229, n_12230, n_12231, n_12232, n_12233, n_12234, n_12235, n_12236, n_12237, n_12238, n_12239, n_12240, n_12241, n_12242, n_12243, n_12244, n_12245, n_12246, n_12247, n_12248, n_12249, n_12250, n_12251, n_12252, n_12253, n_12254, n_12255, n_12256, n_12257, n_12258, n_12259, n_12260, n_12261, n_12262, n_12263, n_12264, n_12265, n_12266, n_12267, n_12268, n_12269, n_12270, n_12271, n_12272, n_12273, n_12274, n_12275, n_12276, n_12277, n_12278, n_12279, n_12280, n_12281, n_12282, n_12283, n_12284, n_12285, n_12286, n_12287, n_12288, n_12289, n_12290, n_12291, n_12292, n_12293, n_12294, n_12295, n_12296, n_12297, n_12298, n_12299, n_12300, n_12301, n_12302, n_12303, n_12304, n_12305, n_12306, n_12307, n_12308, n_12309, n_12310, n_12311, n_12312, n_12313, n_12314, n_12315, n_12316, n_12317, n_12318, n_12319, n_12320, n_12321, n_12322, n_12323, n_12324, n_12325, n_12326, n_12327, n_12328, n_12329, n_12330, n_12331, n_12332, n_12333, n_12334, n_12335, n_12336, n_12337, n_12338, n_12339, n_12340, n_12341, n_12342, n_12343, n_12344, n_12345, n_12346, n_12347, n_12348, n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355, n_12356, n_12357, n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364, n_12365, n_12366, n_12367, n_12368, n_12369, n_12370, n_12371, n_12372, n_12373, n_12374, n_12375, n_12376, n_12377, n_12378, n_12379, n_12380, y19, n_12381, n_12382, n_12383, n_12384, n_12385, n_12386, n_12387, n_12388, n_12389, n_12390, n_12391, n_12392, n_12393, n_12394, n_12395, n_12396, n_12397, n_12398, n_12399, n_12400, n_12401, n_12402, n_12403, n_12404, n_12405, n_12406, n_12407, n_12408, n_12409, n_12410, n_12411, n_12412, n_12413, n_12414, n_12415, n_12416, n_12417, n_12418, n_12419, n_12420, n_12421, n_12422, n_12423, n_12424, n_12425, n_12426, n_12427, n_12428, n_12429, n_12430, n_12431, n_12432, n_12433, n_12434, n_12435, n_12436, n_12437, n_12438, n_12439, n_12440, n_12441, n_12442, n_12443, n_12444, n_12445, n_12446, n_12447, n_12448, n_12449, n_12450, n_12451, n_12452, n_12453, n_12454, n_12455, n_12456, n_12457, n_12458, n_12459, n_12460, n_12461, n_12462, n_12463, n_12464, n_12465, n_12466, n_12467, n_12468, n_12469, n_12470, n_12471, n_12472, n_12473, n_12474, n_12475, n_12476, n_12477, n_12478, n_12479, n_12480, n_12481, n_12482, n_12483, n_12484, n_12485, n_12486, n_12487, n_12488, n_12489, n_12490, n_12491, n_12492, n_12493, n_12494, n_12495, n_12496, n_12497, n_12498, n_12499, n_12500, n_12501, n_12502, n_12503, n_12504, n_12505, n_12506, n_12507, n_12508, n_12509, n_12510, n_12511, n_12512, n_12513, n_12514, n_12515, n_12516, n_12517, n_12518, n_12519, n_12520, n_12521, n_12522, n_12523, n_12524, n_12525, n_12526, n_12527, n_12528, n_12529, n_12530, n_12531, n_12532, n_12533, n_12534, n_12535, n_12536, n_12537, n_12538, n_12539, n_12540, n_12541, n_12542, n_12543, n_12544, n_12545, n_12546, n_12547, n_12548, n_12549, n_12550, n_12551, n_12552, n_12553, n_12554, n_12555, n_12556, n_12557, n_12558, n_12559, n_12560, n_12561, n_12562, n_12563, n_12564, n_12565, n_12566, n_12567, n_12568, n_12569, n_12570, n_12571, n_12572, n_12573, n_12574, n_12575, n_12576, n_12577, n_12578, n_12579, n_12580, n_12581, n_12582, n_12583, n_12584, n_12585, n_12586, n_12587, n_12588, n_12589, n_12590, n_12591, n_12592, n_12593, n_12594, n_12595, n_12596, n_12597, n_12598, n_12599, n_12600, n_12601, n_12602, n_12603, n_12604, n_12605, n_12606, n_12607, n_12608, n_12609, n_12610, n_12611, n_12612, n_12613, n_12614, n_12615, n_12616, n_12617, n_12618, n_12619, n_12620, n_12621, n_12622, n_12623, n_12624, n_12625, n_12626, n_12627, n_12628, n_12629, n_12630, n_12631, n_12632, n_12633, n_12634, n_12635, n_12636, n_12637, n_12638, n_12639, n_12640, n_12641, n_12642, n_12643, n_12644, n_12645, n_12646, n_12647, n_12648, n_12649, n_12650, n_12651, n_12652, n_12653, n_12654, n_12655, n_12656, n_12657, n_12658, n_12659, n_12660, n_12661, n_12662, n_12663, n_12664, n_12665, n_12666, n_12667, n_12668, n_12669, n_12670, n_12671, n_12672, n_12673, n_12674, n_12675, n_12676, n_12677, n_12678, n_12679, n_12680, n_12681, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687, n_12688, n_12689, n_12690, n_12691, n_12692, n_12693, n_12694, n_12695, n_12696, n_12697, n_12698, n_12699, n_12700, n_12701, n_12702, n_12703, n_12704, n_12705, n_12706, n_12707, n_12708, n_12709, n_12710, n_12711, n_12712, n_12713, n_12714, n_12715, n_12716, n_12717, n_12718, n_12719, n_12720, n_12721, n_12722, n_12723, n_12724, n_12725, n_12726, n_12727, n_12728, n_12729, n_12730, n_12731, n_12732, n_12733, n_12734, n_12735, n_12736, n_12737, n_12738, n_12739, n_12740, n_12741, n_12742, n_12743, n_12744, n_12745, n_12746, n_12747, n_12748, n_12749, n_12750, n_12751, n_12752, n_12753, n_12754, n_12755, n_12756, n_12757, y20, n_12758, n_12759, n_12760, n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767, n_12768, n_12769, n_12770, n_12771, n_12772, n_12773, n_12774, n_12775, n_12776, n_12777, n_12778, n_12779, n_12780, n_12781, n_12782, n_12783, n_12784, n_12785, n_12786, n_12787, n_12788, n_12789, n_12790, n_12791, n_12792, n_12793, n_12794, n_12795, n_12796, n_12797, n_12798, n_12799, n_12800, n_12801, n_12802, n_12803, n_12804, n_12805, n_12806, n_12807, n_12808, n_12809, n_12810, n_12811, n_12812, n_12813, n_12814, n_12815, n_12816, n_12817, n_12818, n_12819, n_12820, n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827, n_12828, n_12829, n_12830, n_12831, n_12832, n_12833, n_12834, n_12835, n_12836, n_12837, n_12838, n_12839, n_12840, n_12841, n_12842, n_12843, n_12844, n_12845, n_12846, n_12847, n_12848, n_12849, n_12850, n_12851, n_12852, n_12853, n_12854, n_12855, n_12856, n_12857, n_12858, n_12859, n_12860, n_12861, n_12862, n_12863, n_12864, n_12865, n_12866, n_12867, n_12868, n_12869, n_12870, n_12871, n_12872, n_12873, n_12874, n_12875, n_12876, n_12877, n_12878, n_12879, n_12880, n_12881, n_12882, n_12883, n_12884, n_12885, n_12886, n_12887, n_12888, n_12889, n_12890, n_12891, n_12892, n_12893, n_12894, n_12895, n_12896, n_12897, n_12898, n_12899, n_12900, n_12901, n_12902, n_12903, n_12904, n_12905, n_12906, n_12907, n_12908, n_12909, n_12910, n_12911, n_12912, n_12913, n_12914, n_12915, n_12916, n_12917, n_12918, n_12919, n_12920, n_12921, n_12922, n_12923, n_12924, n_12925, n_12926, n_12927, n_12928, n_12929, n_12930, n_12931, n_12932, n_12933, n_12934, n_12935, n_12936, n_12937, n_12938, n_12939, n_12940, n_12941, n_12942, n_12943, n_12944, n_12945, n_12946, n_12947, n_12948, n_12949, n_12950, n_12951, n_12952, n_12953, n_12954, n_12955, n_12956, n_12957, n_12958, n_12959, n_12960, n_12961, n_12962, n_12963, n_12964, n_12965, n_12966, n_12967, n_12968, n_12969, n_12970, n_12971, n_12972, n_12973, n_12974, n_12975, n_12976, n_12977, n_12978, n_12979, n_12980, n_12981, n_12982, n_12983, n_12984, n_12985, n_12986, n_12987, n_12988, n_12989, n_12990, n_12991, n_12992, n_12993, n_12994, n_12995, n_12996, n_12997, n_12998, n_12999, n_13000, n_13001, n_13002, n_13003, n_13004, n_13005, n_13006, n_13007, n_13008, n_13009, n_13010, n_13011, n_13012, n_13013, n_13014, n_13015, n_13016, n_13017, n_13018, n_13019, n_13020, n_13021, n_13022, n_13023, n_13024, n_13025, n_13026, n_13027, n_13028, n_13029, n_13030, n_13031, n_13032, n_13033, n_13034, n_13035, n_13036, n_13037, n_13038, n_13039, n_13040, n_13041, n_13042, n_13043, n_13044, n_13045, n_13046, n_13047, n_13048, n_13049, n_13050, n_13051, n_13052, n_13053, n_13054, n_13055, n_13056, n_13057, n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064, n_13065, n_13066, n_13067, n_13068, n_13069, n_13070, n_13071, n_13072, n_13073, n_13074, n_13075, n_13076, n_13077, n_13078, n_13079, n_13080, n_13081, n_13082, n_13083, n_13084, n_13085, n_13086, n_13087, n_13088, n_13089, n_13090, n_13091, n_13092, n_13093, n_13094, n_13095, n_13096, n_13097, n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104, n_13105, n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13112, n_13113, n_13114, n_13115, n_13116, n_13117, n_13118, n_13119, n_13120, n_13121, n_13122, n_13123, n_13124, n_13125, n_13126, n_13127, n_13128, n_13129, n_13130, n_13131, n_13132, n_13133, n_13134, n_13135, n_13136, n_13137, n_13138, n_13139, n_13140, n_13141, n_13142, n_13143, n_13144, n_13145, n_13146, n_13147, n_13148, n_13149, n_13150, n_13151, n_13152, n_13153, n_13154, y21, n_13155, n_13156, n_13157, n_13158, n_13159, n_13160, n_13161, n_13162, n_13163, n_13164, n_13165, n_13166, n_13167, n_13168, n_13169, n_13170, n_13171, n_13172, n_13173, n_13174, n_13175, n_13176, n_13177, n_13178, n_13179, n_13180, n_13181, n_13182, n_13183, n_13184, n_13185, n_13186, n_13187, n_13188, n_13189, n_13190, n_13191, n_13192, n_13193, n_13194, n_13195, n_13196, n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203, n_13204, n_13205, n_13206, n_13207, n_13208, n_13209, n_13210, n_13211, n_13212, n_13213, n_13214, n_13215, n_13216, n_13217, n_13218, n_13219, n_13220, n_13221, n_13222, n_13223, n_13224, n_13225, n_13226, n_13227, n_13228, n_13229, n_13230, n_13231, n_13232, n_13233, n_13234, n_13235, n_13236, n_13237, n_13238, n_13239, n_13240, n_13241, n_13242, n_13243, n_13244, n_13245, n_13246, n_13247, n_13248, n_13249, n_13250, n_13251, n_13252, n_13253, n_13254, n_13255, n_13256, n_13257, n_13258, n_13259, n_13260, n_13261, n_13262, n_13263, n_13264, n_13265, n_13266, n_13267, n_13268, n_13269, n_13270, n_13271, n_13272, n_13273, n_13274, n_13275, n_13276, n_13277, n_13278, n_13279, n_13280, n_13281, n_13282, n_13283, n_13284, n_13285, n_13286, n_13287, n_13288, n_13289, n_13290, n_13291, n_13292, n_13293, n_13294, n_13295, n_13296, n_13297, n_13298, n_13299, n_13300, n_13301, n_13302, n_13303, n_13304, n_13305, n_13306, n_13307, n_13308, n_13309, n_13310, n_13311, n_13312, n_13313, n_13314, n_13315, n_13316, n_13317, n_13318, n_13319, n_13320, n_13321, n_13322, n_13323, n_13324, n_13325, n_13326, n_13327, n_13328, n_13329, n_13330, n_13331, n_13332, n_13333, n_13334, n_13335, n_13336, n_13337, n_13338, n_13339, n_13340, n_13341, n_13342, n_13343, n_13344, n_13345, n_13346, n_13347, n_13348, n_13349, n_13350, n_13351, n_13352, n_13353, n_13354, n_13355, n_13356, n_13357, n_13358, n_13359, n_13360, n_13361, n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368, n_13369, n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376, n_13377, n_13378, n_13379, n_13380, n_13381, n_13382, n_13383, n_13384, n_13385, n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392, n_13393, n_13394, n_13395, n_13396, n_13397, n_13398, n_13399, n_13400, n_13401, n_13402, n_13403, n_13404, n_13405, n_13406, n_13407, n_13408, n_13409, n_13410, n_13411, n_13412, n_13413, n_13414, n_13415, n_13416, n_13417, n_13418, n_13419, n_13420, n_13421, n_13422, n_13423, n_13424, n_13425, n_13426, n_13427, n_13428, n_13429, n_13430, n_13431, n_13432, n_13433, n_13434, n_13435, n_13436, n_13437, n_13438, n_13439, n_13440, n_13441, n_13442, n_13443, n_13444, n_13445, n_13446, n_13447, n_13448, n_13449, n_13450, n_13451, n_13452, n_13453, n_13454, n_13455, n_13456, n_13457, n_13458, n_13459, n_13460, n_13461, n_13462, n_13463, n_13464, n_13465, n_13466, n_13467, n_13468, n_13469, n_13470, n_13471, n_13472, n_13473, n_13474, n_13475, n_13476, n_13477, n_13478, n_13479, n_13480, n_13481, n_13482, n_13483, n_13484, n_13485, n_13486, n_13487, n_13488, n_13489, n_13490, n_13491, n_13492, n_13493, n_13494, n_13495, n_13496, n_13497, n_13498, n_13499, n_13500, n_13501, n_13502, n_13503, n_13504, n_13505, n_13506, y22, n_13507, n_13508, n_13509, n_13510, n_13511, n_13512, n_13513, n_13514, n_13515, n_13516, n_13517, n_13518, n_13519, n_13520, n_13521, n_13522, n_13523, n_13524, n_13525, n_13526, n_13527, n_13528, n_13529, n_13530, n_13531, n_13532, n_13533, n_13534, n_13535, n_13536, n_13537, n_13538, n_13539, n_13540, n_13541, n_13542, n_13543, n_13544, n_13545, n_13546, n_13547, n_13548, n_13549, n_13550, n_13551, n_13552, n_13553, n_13554, n_13555, n_13556, n_13557, n_13558, n_13559, n_13560, n_13561, n_13562, n_13563, n_13564, n_13565, n_13566, n_13567, n_13568, n_13569, n_13570, n_13571, n_13572, n_13573, n_13574, n_13575, n_13576, n_13577, n_13578, n_13579, n_13580, n_13581, n_13582, n_13583, n_13584, n_13585, n_13586, n_13587, n_13588, n_13589, n_13590, n_13591, n_13592, n_13593, n_13594, n_13595, n_13596, n_13597, n_13598, n_13599, n_13600, n_13601, n_13602, n_13603, n_13604, n_13605, n_13606, n_13607, n_13608, n_13609, n_13610, n_13611, n_13612, n_13613, n_13614, n_13615, n_13616, n_13617, n_13618, n_13619, n_13620, n_13621, n_13622, n_13623, n_13624, n_13625, n_13626, n_13627, n_13628, n_13629, n_13630, n_13631, n_13632, n_13633, n_13634, n_13635, n_13636, n_13637, n_13638, n_13639, n_13640, n_13641, n_13642, n_13643, n_13644, n_13645, n_13646, n_13647, n_13648, n_13649, n_13650, n_13651, n_13652, n_13653, n_13654, n_13655, n_13656, n_13657, n_13658, n_13659, n_13660, n_13661, n_13662, n_13663, n_13664, n_13665, n_13666, n_13667, n_13668, n_13669, n_13670, n_13671, n_13672, n_13673, n_13674, n_13675, n_13676, n_13677, n_13678, n_13679, n_13680, n_13681, n_13682, n_13683, n_13684, n_13685, n_13686, n_13687, n_13688, n_13689, n_13690, n_13691, n_13692, n_13693, n_13694, n_13695, n_13696, n_13697, n_13698, n_13699, n_13700, n_13701, n_13702, n_13703, n_13704, n_13705, n_13706, n_13707, n_13708, n_13709, n_13710, n_13711, n_13712, n_13713, n_13714, n_13715, n_13716, n_13717, n_13718, n_13719, n_13720, n_13721, n_13722, n_13723, n_13724, n_13725, n_13726, n_13727, n_13728, n_13729, n_13730, n_13731, n_13732, n_13733, n_13734, n_13735, n_13736, n_13737, n_13738, n_13739, n_13740, n_13741, n_13742, n_13743, n_13744, n_13745, n_13746, n_13747, n_13748, n_13749, n_13750, n_13751, n_13752, n_13753, n_13754, n_13755, n_13756, n_13757, n_13758, n_13759, n_13760, n_13761, n_13762, n_13763, n_13764, n_13765, n_13766, n_13767, n_13768, n_13769, y23, n_13770, n_13771, n_13772, n_13773, n_13774, n_13775, n_13776, n_13777, n_13778, n_13779, n_13780, n_13781, n_13782, n_13783, n_13784, n_13785, n_13786, n_13787, n_13788, n_13789, n_13790, n_13791, n_13792, n_13793, n_13794, n_13795, n_13796, n_13797, n_13798, n_13799, n_13800, n_13801, n_13802, n_13803, n_13804, n_13805, n_13806, n_13807, n_13808, n_13809, n_13810, n_13811, n_13812, n_13813, n_13814, n_13815, n_13816, n_13817, n_13818, n_13819, n_13820, n_13821, n_13822, n_13823, n_13824, n_13825, n_13826, n_13827, n_13828, n_13829, n_13830, n_13831, n_13832, n_13833, n_13834, n_13835, n_13836, n_13837, n_13838, n_13839, n_13840, n_13841, n_13842, n_13843, n_13844, n_13845, n_13846, n_13847, n_13848, n_13849, n_13850, n_13851, n_13852, n_13853, n_13854, n_13855, n_13856, n_13857, n_13858, n_13859, n_13860, n_13861, n_13862, n_13863, n_13864, n_13865, n_13866, n_13867, n_13868, n_13869, n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13876, n_13877, n_13878, n_13879, n_13880, n_13881, n_13882, n_13883, n_13884, n_13885, n_13886, n_13887, n_13888, n_13889, n_13890, n_13891, n_13892, n_13893, n_13894, n_13895, n_13896, n_13897, n_13898, n_13899, n_13900, n_13901, n_13902, n_13903, n_13904, n_13905, n_13906, n_13907, n_13908, n_13909, n_13910, n_13911, n_13912, n_13913, n_13914, n_13915, n_13916, n_13917, n_13918, n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925, n_13926, n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933, n_13934, n_13935, n_13936, n_13937, n_13938, n_13939, n_13940, n_13941, n_13942, n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949, n_13950, n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957, n_13958, n_13959, n_13960, n_13961, n_13962, n_13963, n_13964, n_13965, n_13966, n_13967, n_13968, n_13969, n_13970, n_13971, n_13972, n_13973, n_13974, n_13975, n_13976, n_13977, n_13978, n_13979, n_13980, n_13981, n_13982, n_13983, n_13984, n_13985, n_13986, n_13987, n_13988, n_13989, n_13990, n_13991, n_13992, n_13993, n_13994, n_13995, n_13996, n_13997, n_13998, n_13999, n_14000, n_14001, n_14002, n_14003, n_14004, n_14005, n_14006, n_14007, n_14008, n_14009, n_14010, n_14011, n_14012, n_14013, n_14014, n_14015, n_14016, n_14017, n_14018, n_14019, n_14020, n_14021, n_14022, n_14023, n_14024, n_14025, n_14026, n_14027, n_14028, n_14029, n_14030, n_14031, n_14032, n_14033, n_14034, n_14035, n_14036, n_14037, n_14038, n_14039, n_14040, n_14041, n_14042, n_14043, n_14044, n_14045, n_14046, n_14047, n_14048, n_14049, n_14050, n_14051, n_14052, n_14053, n_14054, n_14055, n_14056, n_14057, n_14058, n_14059, n_14060, n_14061, n_14062, n_14063, n_14064, n_14065, n_14066, n_14067, n_14068, n_14069, n_14070, n_14071, n_14072, n_14073, n_14074, n_14075, n_14076, n_14077, n_14078, n_14079, n_14080, n_14081, n_14082, n_14083, n_14084, n_14085, n_14086, n_14087, n_14088, n_14089, n_14090, n_14091, n_14092, n_14093, n_14094, n_14095, n_14096, n_14097, n_14098, n_14099, n_14100, n_14101, n_14102, n_14103, n_14104, n_14105, n_14106, n_14107, n_14108, n_14109, n_14110, n_14111, n_14112, n_14113, n_14114, n_14115, n_14116, n_14117, n_14118, n_14119, n_14120, n_14121, n_14122, n_14123, n_14124, n_14125, n_14126, n_14127, y24, n_14128, n_14129, n_14130, n_14131, n_14132, n_14133, n_14134, n_14135, n_14136, n_14137, n_14138, n_14139, n_14140, n_14141, n_14142, n_14143, n_14144, n_14145, n_14146, n_14147, n_14148, n_14149, n_14150, n_14151, n_14152, n_14153, n_14154, n_14155, n_14156, n_14157, n_14158, n_14159, n_14160, n_14161, n_14162, n_14163, n_14164, n_14165, n_14166, n_14167, n_14168, n_14169, n_14170, n_14171, n_14172, n_14173, n_14174, n_14175, n_14176, n_14177, n_14178, n_14179, n_14180, n_14181, n_14182, n_14183, n_14184, n_14185, n_14186, n_14187, n_14188, n_14189, n_14190, n_14191, n_14192, n_14193, n_14194, n_14195, n_14196, n_14197, n_14198, n_14199, n_14200, n_14201, n_14202, n_14203, n_14204, n_14205, n_14206, n_14207, n_14208, n_14209, n_14210, n_14211, n_14212, n_14213, n_14214, n_14215, n_14216, n_14217, n_14218, n_14219, n_14220, n_14221, n_14222, n_14223, n_14224, n_14225, n_14226, n_14227, n_14228, n_14229, n_14230, n_14231, n_14232, n_14233, n_14234, n_14235, n_14236, n_14237, n_14238, n_14239, n_14240, n_14241, n_14242, n_14243, n_14244, n_14245, n_14246, n_14247, n_14248, n_14249, n_14250, n_14251, n_14252, n_14253, n_14254, n_14255, n_14256, n_14257, n_14258, n_14259, n_14260, n_14261, n_14262, n_14263, n_14264, n_14265, n_14266, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272, n_14273, n_14274, n_14275, n_14276, n_14277, n_14278, n_14279, n_14280, n_14281, n_14282, n_14283, n_14284, n_14285, n_14286, n_14287, n_14288, n_14289, n_14290, n_14291, n_14292, n_14293, n_14294, n_14295, n_14296, n_14297, n_14298, n_14299, n_14300, n_14301, n_14302, n_14303, n_14304, n_14305, n_14306, n_14307, n_14308, n_14309, n_14310, n_14311, n_14312, n_14313, n_14314, n_14315, n_14316, n_14317, n_14318, n_14319, n_14320, n_14321, n_14322, n_14323, n_14324, n_14325, n_14326, n_14327, n_14328, n_14329, n_14330, n_14331, n_14332, n_14333, n_14334, n_14335, n_14336, n_14337, n_14338, n_14339, n_14340, n_14341, n_14342, n_14343, n_14344, n_14345, n_14346, n_14347, n_14348, n_14349, n_14350, n_14351, n_14352, n_14353, n_14354, n_14355, n_14356, n_14357, n_14358, n_14359, n_14360, n_14361, n_14362, n_14363, n_14364, n_14365, n_14366, n_14367, n_14368, n_14369, n_14370, n_14371, n_14372, n_14373, n_14374, n_14375, n_14376, n_14377, n_14378, n_14379, n_14380, n_14381, n_14382, n_14383, n_14384, n_14385, n_14386, n_14387, n_14388, n_14389, n_14390, n_14391, n_14392, n_14393, n_14394, n_14395, n_14396, n_14397, n_14398, n_14399, n_14400, n_14401, n_14402, n_14403, n_14404, n_14405, n_14406, n_14407, n_14408, n_14409, n_14410, n_14411, n_14412, n_14413, n_14414, n_14415, n_14416, n_14417, n_14418, n_14419, n_14420, n_14421, n_14422, n_14423, n_14424, n_14425, n_14426, n_14427, n_14428, n_14429, n_14430, n_14431, n_14432, n_14433, n_14434, n_14435, n_14436, n_14437, n_14438, n_14439, n_14440, n_14441, n_14442, n_14443, n_14444, n_14445, n_14446, n_14447, n_14448, n_14449, n_14450, n_14451, n_14452, n_14453, n_14454, n_14455, n_14456, n_14457, n_14458, n_14459, n_14460, n_14461, n_14462, n_14463, n_14464, n_14465, n_14466, n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, n_14473, n_14474, n_14475, n_14476, n_14477, n_14478, n_14479, n_14480, n_14481, n_14482, n_14483, n_14484, n_14485, n_14486, n_14487, n_14488, n_14489, n_14490, n_14491, n_14492, n_14493, n_14494, n_14495, n_14496, n_14497, n_14498, n_14499, n_14500, n_14501, n_14502, n_14503, n_14504, n_14505, n_14506, n_14507, n_14508, n_14509, n_14510, n_14511, n_14512, n_14513, n_14514, n_14515, n_14516, n_14517, n_14518, n_14519, n_14520, n_14521, n_14522, n_14523, n_14524, n_14525, n_14526, n_14527, n_14528, n_14529, n_14530, n_14531, n_14532, n_14533, n_14534, n_14535, n_14536, n_14537, n_14538, n_14539, n_14540, n_14541, n_14542, n_14543, n_14544, n_14545, n_14546, n_14547, n_14548, n_14549, n_14550, n_14551, n_14552, n_14553, n_14554, n_14555, n_14556, n_14557, n_14558, n_14559, n_14560, n_14561, n_14562, n_14563, n_14564, n_14565, n_14566, n_14567, n_14568, y25, n_14569, n_14570, n_14571, n_14572, n_14573, n_14574, n_14575, n_14576, n_14577, n_14578, n_14579, n_14580, n_14581, n_14582, n_14583, n_14584, n_14585, n_14586, n_14587, n_14588, n_14589, n_14590, n_14591, n_14592, n_14593, n_14594, n_14595, n_14596, n_14597, n_14598, n_14599, n_14600, n_14601, n_14602, n_14603, n_14604, n_14605, n_14606, n_14607, n_14608, n_14609, n_14610, n_14611, n_14612, n_14613, n_14614, n_14615, n_14616, n_14617, n_14618, n_14619, n_14620, n_14621, n_14622, n_14623, n_14624, n_14625, n_14626, n_14627, n_14628, n_14629, n_14630, n_14631, n_14632, n_14633, n_14634, n_14635, n_14636, n_14637, n_14638, n_14639, n_14640, n_14641, n_14642, n_14643, n_14644, n_14645, n_14646, n_14647, n_14648, n_14649, n_14650, n_14651, n_14652, n_14653, n_14654, n_14655, n_14656, n_14657, n_14658, n_14659, n_14660, n_14661, n_14662, n_14663, n_14664, n_14665, n_14666, n_14667, n_14668, n_14669, n_14670, n_14671, n_14672, n_14673, n_14674, n_14675, n_14676, n_14677, n_14678, n_14679, n_14680, n_14681, n_14682, n_14683, n_14684, n_14685, n_14686, n_14687, n_14688, n_14689, n_14690, n_14691, n_14692, n_14693, n_14694, n_14695, n_14696, n_14697, n_14698, n_14699, n_14700, n_14701, n_14702, n_14703, n_14704, n_14705, n_14706, n_14707, n_14708, n_14709, n_14710, n_14711, n_14712, n_14713, n_14714, n_14715, n_14716, n_14717, n_14718, n_14719, n_14720, n_14721, n_14722, n_14723, n_14724, n_14725, n_14726, n_14727, n_14728, n_14729, n_14730, n_14731, n_14732, n_14733, n_14734, n_14735, n_14736, n_14737, n_14738, n_14739, n_14740, n_14741, n_14742, n_14743, n_14744, n_14745, n_14746, n_14747, n_14748, n_14749, n_14750, n_14751, n_14752, n_14753, n_14754, n_14755, n_14756, n_14757, n_14758, n_14759, n_14760, n_14761, n_14762, n_14763, n_14764, n_14765, n_14766, n_14767, n_14768, n_14769, n_14770, n_14771, n_14772, n_14773, n_14774, n_14775, n_14776, n_14777, n_14778, n_14779, n_14780, n_14781, n_14782, n_14783, n_14784, n_14785, n_14786, n_14787, n_14788, n_14789, n_14790, n_14791, n_14792, n_14793, n_14794, n_14795, n_14796, n_14797, n_14798, n_14799, n_14800, n_14801, n_14802, n_14803, n_14804, n_14805, n_14806, n_14807, n_14808, n_14809, n_14810, n_14811, n_14812, n_14813, n_14814, n_14815, n_14816, n_14817, n_14818, n_14819, n_14820, n_14821, n_14822, n_14823, n_14824, n_14825, n_14826, n_14827, n_14828, n_14829, n_14830, n_14831, n_14832, n_14833, n_14834, n_14835, n_14836, n_14837, n_14838, n_14839, n_14840, n_14841, n_14842, n_14843, n_14844, n_14845, n_14846, n_14847, n_14848, n_14849, n_14850, n_14851, n_14852, n_14853, n_14854, n_14855, n_14856, n_14857, n_14858, n_14859, n_14860, n_14861, n_14862, n_14863, n_14864, n_14865, n_14866, n_14867, n_14868, n_14869, n_14870, n_14871, n_14872, n_14873, n_14874, n_14875, n_14876, n_14877, n_14878, n_14879, n_14880, n_14881, n_14882, n_14883, n_14884, n_14885, n_14886, n_14887, n_14888, n_14889, n_14890, n_14891, n_14892, n_14893, n_14894, n_14895, n_14896, n_14897, n_14898, n_14899, n_14900, n_14901, n_14902, n_14903, n_14904, n_14905, n_14906, n_14907, n_14908, n_14909, n_14910, n_14911, n_14912, n_14913, n_14914, n_14915, n_14916, n_14917, n_14918, n_14919, n_14920, n_14921, n_14922, n_14923, n_14924, n_14925, n_14926, n_14927, n_14928, n_14929, n_14930, n_14931, n_14932, n_14933, n_14934, n_14935, n_14936, n_14937, n_14938, n_14939, n_14940, n_14941, n_14942, n_14943, n_14944, n_14945, n_14946, n_14947, n_14948, n_14949, n_14950, n_14951, n_14952, n_14953, n_14954, n_14955, n_14956, n_14957, n_14958, n_14959, n_14960, n_14961, n_14962, n_14963, n_14964, n_14965, n_14966, n_14967, n_14968, n_14969, n_14970, n_14971, n_14972, n_14973, n_14974, n_14975, n_14976, n_14977, n_14978, n_14979, n_14980, n_14981, n_14982, n_14983, n_14984, n_14985, n_14986, n_14987, n_14988, n_14989, n_14990, n_14991, n_14992, n_14993, n_14994, n_14995, n_14996, n_14997, n_14998, n_14999, n_15000, n_15001, n_15002, n_15003, n_15004, n_15005, n_15006, n_15007, n_15008, n_15009, n_15010, n_15011, n_15012, n_15013, n_15014, n_15015, n_15016, n_15017, n_15018, n_15019, n_15020, n_15021, n_15022, n_15023, n_15024, n_15025, n_15026, n_15027, n_15028, n_15029, y26, n_15030, n_15031, n_15032, n_15033, n_15034, n_15035, n_15036, n_15037, n_15038, n_15039, n_15040, n_15041, n_15042, n_15043, n_15044, n_15045, n_15046, n_15047, n_15048, n_15049, n_15050, n_15051, n_15052, n_15053, n_15054, n_15055, n_15056, n_15057, n_15058, n_15059, n_15060, n_15061, n_15062, n_15063, n_15064, n_15065, n_15066, n_15067, n_15068, n_15069, n_15070, n_15071, n_15072, n_15073, n_15074, n_15075, n_15076, n_15077, n_15078, n_15079, n_15080, n_15081, n_15082, n_15083, n_15084, n_15085, n_15086, n_15087, n_15088, n_15089, n_15090, n_15091, n_15092, n_15093, n_15094, n_15095, n_15096, n_15097, n_15098, n_15099, n_15100, n_15101, n_15102, n_15103, n_15104, n_15105, n_15106, n_15107, n_15108, n_15109, n_15110, n_15111, n_15112, n_15113, n_15114, n_15115, n_15116, n_15117, n_15118, n_15119, n_15120, n_15121, n_15122, n_15123, n_15124, n_15125, n_15126, n_15127, n_15128, n_15129, n_15130, n_15131, n_15132, n_15133, n_15134, n_15135, n_15136, n_15137, n_15138, n_15139, n_15140, n_15141, n_15142, n_15143, n_15144, n_15145, n_15146, n_15147, n_15148, n_15149, n_15150, n_15151, n_15152, n_15153, n_15154, n_15155, n_15156, n_15157, n_15158, n_15159, n_15160, n_15161, n_15162, n_15163, n_15164, n_15165, n_15166, n_15167, n_15168, n_15169, n_15170, n_15171, n_15172, n_15173, n_15174, n_15175, n_15176, n_15177, n_15178, n_15179, n_15180, n_15181, n_15182, n_15183, n_15184, n_15185, n_15186, n_15187, n_15188, n_15189, n_15190, n_15191, n_15192, n_15193, n_15194, n_15195, n_15196, n_15197, n_15198, n_15199, n_15200, n_15201, n_15202, n_15203, n_15204, n_15205, n_15206, n_15207, n_15208, n_15209, n_15210, n_15211, n_15212, n_15213, n_15214, n_15215, n_15216, n_15217, n_15218, n_15219, n_15220, n_15221, n_15222, n_15223, n_15224, n_15225, n_15226, n_15227, n_15228, n_15229, n_15230, n_15231, n_15232, n_15233, n_15234, n_15235, n_15236, n_15237, n_15238, n_15239, n_15240, n_15241, n_15242, n_15243, n_15244, n_15245, n_15246, n_15247, n_15248, n_15249, n_15250, n_15251, n_15252, n_15253, n_15254, n_15255, n_15256, n_15257, n_15258, n_15259, n_15260, n_15261, n_15262, n_15263, n_15264, n_15265, n_15266, n_15267, n_15268, n_15269, n_15270, n_15271, n_15272, n_15273, n_15274, n_15275, n_15276, n_15277, n_15278, n_15279, n_15280, n_15281, n_15282, n_15283, n_15284, n_15285, n_15286, n_15287, n_15288, n_15289, n_15290, n_15291, n_15292, n_15293, n_15294, n_15295, n_15296, n_15297, n_15298, n_15299, n_15300, n_15301, n_15302, n_15303, n_15304, n_15305, n_15306, n_15307, n_15308, n_15309, n_15310, n_15311, n_15312, n_15313, n_15314, n_15315, n_15316, n_15317, n_15318, n_15319, n_15320, n_15321, n_15322, n_15323, n_15324, n_15325, n_15326, n_15327, n_15328, n_15329, n_15330, n_15331, n_15332, n_15333, n_15334, n_15335, n_15336, n_15337, n_15338, n_15339, n_15340, n_15341, n_15342, n_15343, n_15344, n_15345, n_15346, n_15347, n_15348, n_15349, n_15350, n_15351, n_15352, n_15353, n_15354, n_15355, n_15356, n_15357, n_15358, n_15359, n_15360, n_15361, n_15362, n_15363, n_15364, n_15365, n_15366, n_15367, n_15368, n_15369, n_15370, n_15371, n_15372, n_15373, n_15374, n_15375, n_15376, n_15377, n_15378, n_15379, n_15380, n_15381, n_15382, n_15383, n_15384, n_15385, n_15386, n_15387, n_15388, n_15389, n_15390, n_15391, n_15392, n_15393, n_15394, n_15395, n_15396, n_15397, n_15398, n_15399, n_15400, n_15401, n_15402, n_15403, n_15404, n_15405, n_15406, n_15407, n_15408, n_15409, n_15410, n_15411, n_15412, n_15413, n_15414, n_15415, n_15416, n_15417, n_15418, n_15419, n_15420, n_15421, n_15422, n_15423, n_15424, n_15425, n_15426, n_15427, n_15428, n_15429, n_15430, n_15431, n_15432, n_15433, n_15434, n_15435, n_15436, n_15437, n_15438, n_15439, n_15440, n_15441, n_15442, n_15443, n_15444, n_15445, n_15446, n_15447, n_15448, n_15449, n_15450, n_15451, n_15452, n_15453, n_15454, n_15455, n_15456, n_15457, n_15458, n_15459, n_15460, n_15461, n_15462, n_15463, n_15464, n_15465, n_15466, n_15467, n_15468, n_15469, n_15470, n_15471, n_15472, n_15473, n_15474, n_15475, n_15476, n_15477, n_15478, n_15479, n_15480, n_15481, n_15482, n_15483, n_15484, n_15485, n_15486, n_15487, n_15488, n_15489, n_15490, y27, n_15491, n_15492, n_15493, n_15494, n_15495, n_15496, n_15497, n_15498, n_15499, n_15500, n_15501, n_15502, n_15503, n_15504, n_15505, n_15506, n_15507, n_15508, n_15509, n_15510, n_15511, n_15512, n_15513, n_15514, n_15515, n_15516, n_15517, n_15518, n_15519, n_15520, n_15521, n_15522, n_15523, n_15524, n_15525, n_15526, n_15527, n_15528, n_15529, n_15530, n_15531, n_15532, n_15533, n_15534, n_15535, n_15536, n_15537, n_15538, n_15539, n_15540, n_15541, n_15542, n_15543, n_15544, n_15545, n_15546, n_15547, n_15548, n_15549, n_15550, n_15551, n_15552, n_15553, n_15554, n_15555, n_15556, n_15557, n_15558, n_15559, n_15560, n_15561, n_15562, n_15563, n_15564, n_15565, n_15566, n_15567, n_15568, n_15569, n_15570, n_15571, n_15572, n_15573, n_15574, n_15575, n_15576, n_15577, n_15578, n_15579, n_15580, n_15581, n_15582, n_15583, n_15584, n_15585, n_15586, n_15587, n_15588, n_15589, n_15590, n_15591, n_15592, n_15593, n_15594, n_15595, n_15596, n_15597, n_15598, n_15599, n_15600, n_15601, n_15602, n_15603, n_15604, n_15605, n_15606, n_15607, n_15608, n_15609, n_15610, n_15611, n_15612, n_15613, n_15614, n_15615, n_15616, n_15617, n_15618, n_15619, n_15620, n_15621, n_15622, n_15623, n_15624, n_15625, n_15626, n_15627, n_15628, n_15629, n_15630, n_15631, n_15632, n_15633, n_15634, n_15635, n_15636, n_15637, n_15638, n_15639, n_15640, n_15641, n_15642, n_15643, n_15644, n_15645, n_15646, n_15647, n_15648, n_15649, n_15650, n_15651, n_15652, n_15653, n_15654, n_15655, n_15656, n_15657, n_15658, n_15659, n_15660, n_15661, n_15662, n_15663, n_15664, n_15665, n_15666, n_15667, n_15668, n_15669, n_15670, n_15671, n_15672, n_15673, n_15674, n_15675, n_15676, n_15677, n_15678, n_15679, n_15680, n_15681, n_15682, n_15683, n_15684, n_15685, n_15686, n_15687, n_15688, n_15689, n_15690, n_15691, n_15692, n_15693, n_15694, n_15695, n_15696, n_15697, n_15698, n_15699, n_15700, n_15701, n_15702, n_15703, n_15704, n_15705, n_15706, n_15707, n_15708, n_15709, n_15710, n_15711, n_15712, n_15713, n_15714, n_15715, n_15716, n_15717, n_15718, n_15719, n_15720, n_15721, n_15722, n_15723, n_15724, n_15725, n_15726, n_15727, n_15728, n_15729, n_15730, n_15731, n_15732, n_15733, n_15734, n_15735, n_15736, n_15737, n_15738, n_15739, n_15740, n_15741, n_15742, n_15743, n_15744, n_15745, n_15746, n_15747, n_15748, n_15749, n_15750, n_15751, n_15752, n_15753, n_15754, n_15755, n_15756, n_15757, n_15758, n_15759, n_15760, n_15761, n_15762, n_15763, n_15764, n_15765, n_15766, n_15767, n_15768, n_15769, n_15770, n_15771, n_15772, n_15773, n_15774, n_15775, n_15776, n_15777, n_15778, n_15779, n_15780, n_15781, n_15782, n_15783, n_15784, n_15785, n_15786, n_15787, n_15788, n_15789, n_15790, n_15791, n_15792, n_15793, n_15794, n_15795, n_15796, n_15797, n_15798, n_15799, n_15800, n_15801, n_15802, n_15803, n_15804, n_15805, n_15806, n_15807, n_15808, n_15809, n_15810, n_15811, n_15812, n_15813, n_15814, n_15815, n_15816, n_15817, n_15818, n_15819, n_15820, n_15821, n_15822, n_15823, n_15824, n_15825, n_15826, n_15827, n_15828, n_15829, n_15830, n_15831, n_15832, n_15833, n_15834, n_15835, n_15836, n_15837, n_15838, n_15839, n_15840, n_15841, n_15842, n_15843, n_15844, n_15845, n_15846, n_15847, n_15848, n_15849, n_15850, n_15851, n_15852, n_15853, n_15854, n_15855, n_15856, n_15857, n_15858, n_15859, n_15860, n_15861, n_15862, n_15863, n_15864, n_15865, n_15866, n_15867, n_15868, n_15869, n_15870, n_15871, n_15872, n_15873, n_15874, n_15875, n_15876, n_15877, n_15878, y28, n_15879, n_15880, n_15881, n_15882, n_15883, n_15884, n_15885, n_15886, n_15887, n_15888, n_15889, n_15890, n_15891, n_15892, n_15893, n_15894, n_15895, n_15896, n_15897, n_15898, n_15899, n_15900, n_15901, n_15902, n_15903, n_15904, n_15905, n_15906, n_15907, n_15908, n_15909, n_15910, n_15911, n_15912, n_15913, n_15914, n_15915, n_15916, n_15917, n_15918, n_15919, n_15920, n_15921, n_15922, n_15923, n_15924, n_15925, n_15926, n_15927, n_15928, n_15929, n_15930, n_15931, n_15932, n_15933, n_15934, n_15935, n_15936, n_15937, n_15938, n_15939, n_15940, n_15941, n_15942, n_15943, n_15944, n_15945, n_15946, n_15947, n_15948, n_15949, n_15950, n_15951, n_15952, n_15953, n_15954, n_15955, n_15956, n_15957, n_15958, n_15959, n_15960, n_15961, n_15962, n_15963, n_15964, n_15965, n_15966, n_15967, n_15968, n_15969, n_15970, n_15971, n_15972, n_15973, n_15974, n_15975, n_15976, n_15977, n_15978, n_15979, n_15980, n_15981, n_15982, n_15983, n_15984, n_15985, n_15986, n_15987, n_15988, n_15989, n_15990, n_15991, n_15992, n_15993, n_15994, n_15995, n_15996, n_15997, n_15998, n_15999, n_16000, n_16001, n_16002, n_16003, n_16004, n_16005, n_16006, n_16007, n_16008, n_16009, n_16010, n_16011, n_16012, n_16013, n_16014, n_16015, n_16016, n_16017, n_16018, n_16019, n_16020, n_16021, n_16022, n_16023, n_16024, n_16025, n_16026, n_16027, n_16028, n_16029, n_16030, n_16031, n_16032, n_16033, n_16034, n_16035, n_16036, n_16037, n_16038, n_16039, n_16040, n_16041, n_16042, n_16043, n_16044, n_16045, n_16046, n_16047, n_16048, n_16049, n_16050, n_16051, n_16052, n_16053, n_16054, n_16055, n_16056, n_16057, n_16058, n_16059, n_16060, n_16061, n_16062, n_16063, n_16064, n_16065, n_16066, n_16067, n_16068, n_16069, n_16070, n_16071, n_16072, n_16073, n_16074, n_16075, n_16076, n_16077, n_16078, n_16079, n_16080, n_16081, n_16082, n_16083, n_16084, n_16085, n_16086, n_16087, n_16088, n_16089, n_16090, n_16091, n_16092, n_16093, n_16094, n_16095, n_16096, n_16097, n_16098, n_16099, n_16100, n_16101, n_16102, n_16103, n_16104, n_16105, n_16106, n_16107, n_16108, n_16109, n_16110, n_16111, n_16112, n_16113, n_16114, n_16115, n_16116, n_16117, n_16118, n_16119, n_16120, n_16121, n_16122, n_16123, n_16124, n_16125, n_16126, n_16127, n_16128, n_16129, n_16130, n_16131, n_16132, n_16133, n_16134, n_16135, n_16136, n_16137, n_16138, n_16139, n_16140, n_16141, n_16142, n_16143, n_16144, n_16145, n_16146, n_16147, n_16148, n_16149, n_16150, n_16151, n_16152, n_16153, n_16154, n_16155, n_16156, n_16157, n_16158, n_16159, n_16160, n_16161, n_16162, n_16163, n_16164, n_16165, n_16166, n_16167, n_16168, n_16169, n_16170, n_16171, n_16172, n_16173, n_16174, n_16175, n_16176, n_16177, n_16178, n_16179, n_16180, n_16181, n_16182, n_16183, n_16184, n_16185, n_16186, n_16187, n_16188, n_16189, n_16190, n_16191, n_16192, n_16193, n_16194, n_16195, n_16196, n_16197, n_16198, n_16199, n_16200, n_16201, n_16202, n_16203, n_16204, n_16205, n_16206, n_16207, n_16208, n_16209, n_16210, n_16211, n_16212, n_16213, n_16214, n_16215, n_16216, n_16217, n_16218, n_16219, n_16220, n_16221, n_16222, n_16223, n_16224, n_16225, n_16226, n_16227, n_16228, n_16229, n_16230, n_16231, n_16232, n_16233, n_16234, n_16235, n_16236, n_16237, n_16238, n_16239, n_16240, n_16241, n_16242, n_16243, n_16244, n_16245, n_16246, n_16247, n_16248, n_16249, n_16250, n_16251, n_16252, n_16253, n_16254, n_16255, n_16256, n_16257, n_16258, n_16259, n_16260, n_16261, n_16262, n_16263, n_16264, n_16265, n_16266, n_16267, n_16268, n_16269, n_16270, n_16271, n_16272, n_16273, n_16274, n_16275, n_16276, n_16277, n_16278, n_16279, n_16280, n_16281, n_16282, n_16283, n_16284, n_16285, n_16286, n_16287, n_16288, n_16289, n_16290, n_16291, n_16292, n_16293, n_16294, n_16295, n_16296, n_16297, y29, n_16298, n_16299, n_16300, n_16301, n_16302, n_16303, n_16304, n_16305, n_16306, n_16307, n_16308, n_16309, n_16310, n_16311, n_16312, n_16313, n_16314, n_16315, n_16316, n_16317, n_16318, n_16319, n_16320, n_16321, n_16322, n_16323, n_16324, n_16325, n_16326, n_16327, n_16328, n_16329, n_16330, n_16331, n_16332, n_16333, n_16334, n_16335, n_16336, n_16337, n_16338, n_16339, n_16340, n_16341, n_16342, n_16343, n_16344, n_16345, n_16346, n_16347, n_16348, n_16349, n_16350, n_16351, n_16352, n_16353, n_16354, n_16355, n_16356, n_16357, n_16358, n_16359, n_16360, n_16361, n_16362, n_16363, n_16364, n_16365, n_16366, n_16367, n_16368, n_16369, n_16370, n_16371, n_16372, n_16373, n_16374, n_16375, n_16376, n_16377, n_16378, n_16379, n_16380, n_16381, n_16382, n_16383, n_16384, n_16385, n_16386, n_16387, n_16388, n_16389, n_16390, n_16391, n_16392, n_16393, n_16394, n_16395, n_16396, n_16397, n_16398, n_16399, n_16400, n_16401, n_16402, n_16403, n_16404, n_16405, n_16406, n_16407, n_16408, n_16409, n_16410, n_16411, n_16412, n_16413, n_16414, n_16415, n_16416, n_16417, n_16418, n_16419, n_16420, n_16421, n_16422, n_16423, n_16424, n_16425, n_16426, n_16427, n_16428, n_16429, n_16430, n_16431, n_16432, n_16433, n_16434, n_16435, n_16436, n_16437, n_16438, n_16439, n_16440, n_16441, n_16442, n_16443, n_16444, n_16445, n_16446, n_16447, n_16448, n_16449, n_16450, n_16451, n_16452, n_16453, n_16454, n_16455, n_16456, n_16457, n_16458, n_16459, n_16460, n_16461, n_16462, n_16463, n_16464, n_16465, n_16466, n_16467, n_16468, n_16469, n_16470, n_16471, n_16472, n_16473, n_16474, n_16475, n_16476, n_16477, n_16478, n_16479, n_16480, n_16481, n_16482, n_16483, n_16484, n_16485, n_16486, n_16487, n_16488, n_16489, n_16490, n_16491, n_16492, n_16493, n_16494, n_16495, n_16496, n_16497, n_16498, n_16499, n_16500, n_16501, n_16502, n_16503, n_16504, n_16505, n_16506, n_16507, n_16508, n_16509, n_16510, n_16511, n_16512, n_16513, n_16514, n_16515, n_16516, n_16517, n_16518, n_16519, n_16520, n_16521, n_16522, n_16523, n_16524, n_16525, n_16526, n_16527, n_16528, n_16529, n_16530, n_16531, n_16532, n_16533, n_16534, n_16535, n_16536, n_16537, n_16538, n_16539, n_16540, n_16541, n_16542, n_16543, n_16544, n_16545, n_16546, n_16547, n_16548, n_16549, n_16550, n_16551, n_16552, n_16553, n_16554, n_16555, n_16556, n_16557, n_16558, n_16559, n_16560, n_16561, n_16562, n_16563, n_16564, n_16565, n_16566, n_16567, n_16568, n_16569, n_16570, n_16571, n_16572, n_16573, n_16574, n_16575, n_16576, n_16577, n_16578, n_16579, n_16580, n_16581, n_16582, n_16583, n_16584, n_16585, n_16586, n_16587, n_16588, n_16589, n_16590, n_16591, n_16592, n_16593, n_16594, n_16595, n_16596, n_16597, n_16598, n_16599, n_16600, n_16601, n_16602, n_16603, n_16604, n_16605, n_16606, n_16607, n_16608, n_16609, n_16610, n_16611, n_16612, n_16613, n_16614, n_16615, n_16616, n_16617, n_16618, n_16619, n_16620, n_16621, n_16622, n_16623, n_16624, n_16625, n_16626, n_16627, n_16628, n_16629, n_16630, n_16631, n_16632, n_16633, n_16634, n_16635, n_16636, n_16637, n_16638, n_16639, n_16640, n_16641, n_16642, n_16643, n_16644, n_16645, n_16646, n_16647, n_16648, n_16649, n_16650, n_16651, n_16652, n_16653, n_16654, n_16655, n_16656, n_16657, n_16658, n_16659, n_16660, n_16661, n_16662, n_16663, n_16664, n_16665, n_16666, n_16667, n_16668, n_16669, n_16670, n_16671, n_16672, n_16673, n_16674, n_16675, n_16676, n_16677, n_16678, n_16679, n_16680, n_16681, n_16682, n_16683, n_16684, n_16685, n_16686, n_16687, n_16688, n_16689, n_16690, n_16691, n_16692, n_16693, n_16694, n_16695, n_16696, n_16697, n_16698, n_16699, n_16700, n_16701, n_16702, n_16703, n_16704, n_16705, n_16706, n_16707, n_16708, n_16709, n_16710, n_16711, n_16712, n_16713, n_16714, n_16715, n_16716, n_16717, n_16718, n_16719, n_16720, n_16721, n_16722, n_16723, n_16724, n_16725, n_16726, n_16727, n_16728, n_16729, n_16730, n_16731, n_16732, n_16733, n_16734, n_16735, n_16736, n_16737, n_16738, n_16739, n_16740, n_16741, n_16742, n_16743, n_16744, n_16745, n_16746, n_16747, n_16748, n_16749, n_16750, n_16751, n_16752, n_16753, n_16754, n_16755, n_16756, n_16757, n_16758, n_16759, n_16760, n_16761, n_16762, n_16763, n_16764, n_16765, n_16766, n_16767, n_16768, n_16769, n_16770, n_16771, n_16772, n_16773, n_16774, n_16775, n_16776, n_16777, n_16778, n_16779, n_16780, n_16781, n_16782, n_16783, n_16784, n_16785, n_16786, n_16787, n_16788, n_16789, n_16790, n_16791, n_16792, n_16793, n_16794, n_16795, n_16796, n_16797, n_16798, n_16799, n_16800, n_16801, n_16802, n_16803, n_16804, n_16805, n_16806, n_16807, n_16808, n_16809, n_16810, n_16811, n_16812, n_16813, n_16814, n_16815, n_16816, n_16817, n_16818, n_16819, n_16820, y30, n_16821, n_16822, n_16823, n_16824, n_16825, n_16826, n_16827, n_16828, n_16829, n_16830, n_16831, n_16832, n_16833, n_16834, n_16835, n_16836, n_16837, n_16838, n_16839, n_16840, n_16841, n_16842, n_16843, n_16844, n_16845, n_16846, n_16847, n_16848, n_16849, n_16850, n_16851, n_16852, n_16853, n_16854, n_16855, n_16856, n_16857, n_16858, n_16859, n_16860, n_16861, n_16862, n_16863, n_16864, n_16865, n_16866, n_16867, n_16868, n_16869, n_16870, n_16871, n_16872, n_16873, n_16874, n_16875, n_16876, n_16877, n_16878, n_16879, n_16880, n_16881, n_16882, n_16883, n_16884, n_16885, n_16886, n_16887, n_16888, n_16889, n_16890, n_16891, n_16892, n_16893, n_16894, n_16895, n_16896, n_16897, n_16898, n_16899, n_16900, n_16901, n_16902, n_16903, n_16904, n_16905, n_16906, n_16907, n_16908, n_16909, n_16910, n_16911, n_16912, n_16913, n_16914, n_16915, n_16916, n_16917, n_16918, n_16919, n_16920, n_16921, n_16922, n_16923, n_16924, n_16925, n_16926, n_16927, n_16928, n_16929, n_16930, n_16931, n_16932, n_16933, n_16934, n_16935, n_16936, n_16937, n_16938, n_16939, n_16940, n_16941, n_16942, n_16943, n_16944, n_16945, n_16946, n_16947, n_16948, n_16949, n_16950, n_16951, n_16952, n_16953, n_16954, n_16955, n_16956, n_16957, n_16958, n_16959, n_16960, n_16961, n_16962, n_16963, n_16964, n_16965, n_16966, n_16967, n_16968, n_16969, n_16970, n_16971, n_16972, n_16973, n_16974, n_16975, n_16976, n_16977, n_16978, n_16979, n_16980, n_16981, n_16982, n_16983, n_16984, n_16985, n_16986, n_16987, n_16988, n_16989, n_16990, n_16991, n_16992, n_16993, n_16994, n_16995, n_16996, n_16997, n_16998, n_16999, n_17000, n_17001, n_17002, n_17003, n_17004, n_17005, n_17006, n_17007, n_17008, n_17009, n_17010, n_17011, n_17012, n_17013, n_17014, n_17015, n_17016, n_17017, n_17018, n_17019, n_17020, n_17021, n_17022, n_17023, n_17024, n_17025, n_17026, n_17027, n_17028, n_17029, n_17030, n_17031, n_17032, n_17033, n_17034, n_17035, n_17036, n_17037, n_17038, n_17039, n_17040, n_17041, n_17042, n_17043, n_17044, n_17045, n_17046, n_17047, n_17048, n_17049, n_17050, n_17051, n_17052, n_17053, n_17054, n_17055, n_17056, n_17057, n_17058, n_17059, n_17060, n_17061, n_17062, n_17063, n_17064, n_17065, n_17066, n_17067, n_17068, n_17069, n_17070, n_17071, n_17072, n_17073, n_17074, n_17075, n_17076, n_17077, n_17078, n_17079, n_17080, n_17081, n_17082, n_17083, n_17084, n_17085, n_17086, n_17087, n_17088, n_17089, n_17090, n_17091, n_17092, n_17093, n_17094, n_17095, n_17096, n_17097, n_17098, n_17099, n_17100, n_17101, n_17102, n_17103, n_17104, n_17105, n_17106, n_17107, n_17108, n_17109, n_17110, n_17111, n_17112, n_17113, n_17114, n_17115, n_17116, n_17117, n_17118, n_17119, n_17120, n_17121, n_17122, n_17123, n_17124, n_17125, n_17126, n_17127, n_17128, n_17129, n_17130, n_17131, n_17132, n_17133, n_17134, n_17135, n_17136, n_17137, n_17138, n_17139, n_17140, n_17141, n_17142, n_17143, n_17144, n_17145, n_17146, n_17147, n_17148, n_17149, n_17150, n_17151, n_17152, n_17153, n_17154, n_17155, n_17156, n_17157, n_17158, n_17159, n_17160, n_17161, n_17162, n_17163, n_17164, n_17165, n_17166, n_17167, n_17168, n_17169, n_17170, n_17171, n_17172, n_17173, n_17174, n_17175, n_17176, n_17177, n_17178, n_17179, n_17180, n_17181, n_17182, n_17183, n_17184, n_17185, n_17186, n_17187, n_17188, n_17189, n_17190, n_17191, n_17192, n_17193, n_17194, n_17195, n_17196, n_17197, n_17198, n_17199, n_17200, n_17201, n_17202, n_17203, n_17204, n_17205, n_17206, n_17207, n_17208, n_17209, n_17210, n_17211, n_17212, n_17213, n_17214, n_17215, n_17216, n_17217, n_17218, n_17219, n_17220, n_17221, n_17222, n_17223, n_17224, n_17225, n_17226, n_17227, n_17228, n_17229, n_17230, n_17231, n_17232, n_17233, n_17234, n_17235, n_17236, n_17237, n_17238, n_17239, n_17240, n_17241, n_17242, n_17243, n_17244, n_17245, n_17246, n_17247, n_17248, n_17249, n_17250, n_17251, y31, n_17252, n_17253, n_17254, n_17255, n_17256, n_17257, n_17258, n_17259, n_17260, n_17261, n_17262, n_17263, n_17264, n_17265, n_17266, n_17267, n_17268, n_17269, n_17270, n_17271, n_17272, n_17273, n_17274, n_17275, n_17276, n_17277, n_17278, n_17279, n_17280, n_17281, n_17282, n_17283, n_17284, n_17285, n_17286, n_17287, n_17288, n_17289, n_17290, n_17291, n_17292, n_17293, n_17294, n_17295, n_17296, n_17297, n_17298, n_17299, n_17300, n_17301, n_17302, n_17303, n_17304, n_17305, n_17306, n_17307, n_17308, n_17309, n_17310, n_17311, n_17312, n_17313, n_17314, n_17315, n_17316, n_17317, n_17318, n_17319, n_17320, n_17321, n_17322, n_17323, n_17324, n_17325, n_17326, n_17327, n_17328, n_17329, n_17330, n_17331, n_17332, n_17333, n_17334, n_17335, n_17336, n_17337, n_17338, n_17339, n_17340, n_17341, n_17342, n_17343, n_17344, n_17345, n_17346, n_17347, n_17348, n_17349, n_17350, n_17351, n_17352, n_17353, n_17354, n_17355, n_17356, n_17357, n_17358, n_17359, n_17360, n_17361, n_17362, n_17363, n_17364, n_17365, n_17366, n_17367, n_17368, n_17369, n_17370, n_17371, n_17372, n_17373, n_17374, n_17375, n_17376, n_17377, n_17378, n_17379, n_17380, n_17381, n_17382, n_17383, n_17384, n_17385, n_17386, n_17387, n_17388, n_17389, n_17390, n_17391, n_17392, n_17393, n_17394, n_17395, n_17396, n_17397, n_17398, n_17399, n_17400, n_17401, n_17402, n_17403, n_17404, n_17405, n_17406, n_17407, n_17408, n_17409, n_17410, n_17411, n_17412, n_17413, n_17414, n_17415, n_17416, n_17417, n_17418, n_17419, n_17420, n_17421, n_17422, n_17423, n_17424, n_17425, n_17426, n_17427, n_17428, n_17429, n_17430, n_17431, n_17432, n_17433, n_17434, n_17435, n_17436, n_17437, n_17438, n_17439, n_17440, n_17441, n_17442, n_17443, n_17444, n_17445, n_17446, n_17447, n_17448, n_17449, n_17450, n_17451, n_17452, n_17453, n_17454, n_17455, n_17456, n_17457, n_17458, n_17459, n_17460, n_17461, n_17462, n_17463, n_17464, n_17465, n_17466, n_17467, n_17468, n_17469, n_17470, n_17471, n_17472, n_17473, n_17474, n_17475, n_17476, n_17477, n_17478, n_17479, n_17480, n_17481, n_17482, n_17483, n_17484, n_17485, n_17486, n_17487, n_17488, n_17489, n_17490, n_17491, n_17492, n_17493, n_17494, n_17495, n_17496, n_17497, n_17498, n_17499, n_17500, n_17501, n_17502, n_17503, n_17504, n_17505, n_17506, n_17507, n_17508, n_17509, n_17510, n_17511, n_17512, n_17513, n_17514, n_17515, n_17516, n_17517, n_17518, n_17519, n_17520, n_17521, n_17522, n_17523, n_17524, n_17525, n_17526, n_17527, n_17528, n_17529, y32, n_17530, n_17531, n_17532, n_17533, n_17534, n_17535, n_17536, n_17537, n_17538, n_17539, n_17540, n_17541, n_17542, n_17543, n_17544, n_17545, n_17546, n_17547, n_17548, n_17549, n_17550, n_17551, n_17552, n_17553, n_17554, n_17555, n_17556, n_17557, n_17558, n_17559, n_17560, n_17561, n_17562, n_17563, n_17564, n_17565, n_17566, n_17567, n_17568, n_17569, n_17570, n_17571, n_17572, n_17573, n_17574, n_17575, n_17576, n_17577, n_17578, n_17579, n_17580, n_17581, n_17582, n_17583, n_17584, n_17585, n_17586, n_17587, n_17588, n_17589, n_17590, n_17591, n_17592, n_17593, n_17594, n_17595, n_17596, n_17597, n_17598, n_17599, n_17600, n_17601, n_17602, n_17603, n_17604, n_17605, n_17606, n_17607, n_17608, n_17609, n_17610, n_17611, n_17612, n_17613, n_17614, n_17615, n_17616, n_17617, n_17618, n_17619, n_17620, n_17621, n_17622, n_17623, n_17624, n_17625, n_17626, n_17627, n_17628, n_17629, n_17630, n_17631, n_17632, n_17633, n_17634, n_17635, n_17636, n_17637, n_17638, n_17639, n_17640, n_17641, n_17642, n_17643, n_17644, n_17645, n_17646, n_17647, n_17648, n_17649, n_17650, n_17651, n_17652, n_17653, n_17654, n_17655, n_17656, n_17657, n_17658, n_17659, n_17660, n_17661, n_17662, n_17663, n_17664, n_17665, n_17666, n_17667, n_17668, n_17669, n_17670, n_17671, n_17672, n_17673, n_17674, n_17675, n_17676, n_17677, n_17678, n_17679, n_17680, n_17681, n_17682, n_17683, n_17684, n_17685, n_17686, n_17687, n_17688, n_17689, n_17690, n_17691, n_17692, n_17693, n_17694, n_17695, n_17696, n_17697, n_17698, n_17699, n_17700, n_17701, n_17702, n_17703, n_17704, n_17705, n_17706, n_17707, n_17708, n_17709, n_17710, n_17711, n_17712, n_17713, n_17714, n_17715, n_17716, n_17717, n_17718, n_17719, n_17720, n_17721, n_17722, n_17723, n_17724, n_17725, n_17726, n_17727, n_17728, n_17729, n_17730, n_17731, n_17732, n_17733, n_17734, n_17735, n_17736, n_17737, n_17738, n_17739, n_17740, n_17741, n_17742, n_17743, n_17744, n_17745, n_17746, n_17747, n_17748, n_17749, n_17750, n_17751, n_17752, n_17753, n_17754, n_17755, n_17756, n_17757, n_17758, n_17759, n_17760, n_17761, n_17762, n_17763, n_17764, n_17765, n_17766, n_17767, n_17768, n_17769, n_17770, n_17771, y33, n_17772, n_17773, n_17774, n_17775, n_17776, n_17777, n_17778, n_17779, n_17780, n_17781, n_17782, n_17783, n_17784, n_17785, n_17786, n_17787, n_17788, n_17789, n_17790, n_17791, n_17792, n_17793, n_17794, n_17795, n_17796, n_17797, n_17798, n_17799, n_17800, n_17801, n_17802, n_17803, n_17804, n_17805, n_17806, n_17807, n_17808, n_17809, n_17810, n_17811, n_17812, n_17813, n_17814, n_17815, n_17816, n_17817, n_17818, n_17819, n_17820, n_17821, n_17822, n_17823, n_17824, n_17825, n_17826, n_17827, n_17828, n_17829, n_17830, n_17831, n_17832, n_17833, n_17834, n_17835, n_17836, n_17837, n_17838, n_17839, n_17840, n_17841, n_17842, n_17843, n_17844, n_17845, n_17846, n_17847, n_17848, n_17849, n_17850, n_17851, n_17852, n_17853, n_17854, n_17855, n_17856, n_17857, n_17858, n_17859, n_17860, n_17861, n_17862, n_17863, n_17864, n_17865, n_17866, n_17867, n_17868, n_17869, n_17870, n_17871, n_17872, n_17873, n_17874, n_17875, n_17876, n_17877, n_17878, n_17879, n_17880, n_17881, n_17882, n_17883, n_17884, n_17885, n_17886, n_17887, n_17888, n_17889, n_17890, n_17891, n_17892, n_17893, n_17894, n_17895, n_17896, n_17897, n_17898, n_17899, n_17900, n_17901, n_17902, n_17903, n_17904, n_17905, n_17906, n_17907, n_17908, n_17909, n_17910, n_17911, n_17912, n_17913, n_17914, n_17915, y34, n_17916, n_17917, n_17918, n_17919, n_17920, n_17921, n_17922, n_17923, n_17924, n_17925, n_17926, n_17927, n_17928, n_17929, n_17930, n_17931, n_17932, n_17933, n_17934, n_17935, n_17936, n_17937, n_17938, n_17939, n_17940, n_17941, n_17942, n_17943, n_17944, n_17945, n_17946, n_17947, n_17948, n_17949, n_17950, n_17951, n_17952, n_17953, n_17954, n_17955, n_17956, n_17957, n_17958, n_17959, n_17960, n_17961, n_17962, n_17963, n_17964, n_17965, n_17966, n_17967, n_17968, n_17969, n_17970, n_17971, n_17972, n_17973, n_17974, n_17975, n_17976, n_17977, n_17978, n_17979, n_17980, n_17981, n_17982, n_17983, n_17984, n_17985, n_17986, n_17987, n_17988, n_17989, n_17990, n_17991, n_17992, n_17993, n_17994, n_17995, n_17996, n_17997, n_17998, n_17999, y35, n_18000, n_18001, n_18002, n_18003, n_18004, n_18005, n_18006, n_18007, n_18008, n_18009, n_18010, n_18011, n_18012, n_18013, n_18014, n_18015, n_18016, n_18017, n_18018, n_18019, n_18020, n_18021, n_18022, n_18023, n_18024, n_18025, n_18026, n_18027, n_18028, n_18029, n_18030, n_18031, n_18032, n_18033, n_18034, n_18035, n_18036, n_18037, n_18038, n_18039, n_18040, n_18041, n_18042, n_18043, n_18044, n_18045, n_18046, n_18047, n_18048, n_18049, n_18050, n_18051, n_18052, n_18053, n_18054, n_18055, n_18056, n_18057, n_18058, n_18059, n_18060, n_18061, n_18062, n_18063, n_18064, n_18065, n_18066, n_18067, n_18068, n_18069, n_18070, n_18071, n_18072, n_18073, n_18074, y36, n_18075, n_18076, n_18077, n_18078, n_18079, n_18080, n_18081, n_18082, n_18083, n_18084, n_18085, n_18086, n_18087, n_18088, n_18089, n_18090, n_18091, n_18092, n_18093, n_18094, n_18095, n_18096, n_18097, n_18098, n_18099, n_18100, n_18101, n_18102, n_18103, n_18104, n_18105, n_18106, n_18107, n_18108, n_18109, n_18110, n_18111, n_18112, n_18113, n_18114, n_18115, n_18116, n_18117, n_18118, n_18119, n_18120, n_18121, n_18122, n_18123, n_18124, n_18125, n_18126, n_18127, n_18128, n_18129, n_18130, n_18131, n_18132, n_18133, n_18134, n_18135, n_18136, n_18137, n_18138, n_18139, n_18140, n_18141, n_18142, n_18143, n_18144, n_18145, n_18146, n_18147, n_18148, n_18149, y37, n_18150, n_18151, n_18152, n_18153, n_18154, n_18155, n_18156, n_18157, n_18158, n_18159, n_18160, n_18161, n_18162, n_18163, n_18164, n_18165, n_18166, n_18167, n_18168, n_18169, n_18170, n_18171, n_18172, n_18173, n_18174, n_18175, n_18176, n_18177, n_18178, n_18179, n_18180, n_18181, n_18182, n_18183, n_18184, n_18185, n_18186, n_18187, n_18188, n_18189, n_18190, n_18191, n_18192, n_18193, n_18194, n_18195, n_18196, n_18197, n_18198, n_18199, n_18200, n_18201, n_18202, n_18203, n_18204, n_18205, n_18206, n_18207, n_18208, n_18209, n_18210, n_18211, n_18212, n_18213, n_18214, n_18215, n_18216, n_18217, n_18218, n_18219, n_18220, n_18221, n_18222, n_18223, n_18224, n_18225, n_18226, n_18227, n_18228, y38, n_18229, n_18230, n_18231, n_18232, n_18233, n_18234, n_18235, n_18236, n_18237, n_18238, n_18239, n_18240, n_18241, n_18242, n_18243, n_18244, n_18245, n_18246, n_18247, n_18248, n_18249, n_18250, n_18251, n_18252, n_18253, n_18254, n_18255, n_18256, n_18257, n_18258, n_18259, n_18260, n_18261, n_18262, n_18263, n_18264, n_18265, n_18266, n_18267, n_18268, n_18269, n_18270, n_18271, n_18272, n_18273, n_18274, n_18275, n_18276, n_18277, n_18278, n_18279, n_18280, n_18281, n_18282, n_18283, n_18284, n_18285, n_18286, n_18287, n_18288, n_18289, n_18290, n_18291, n_18292, n_18293, y39, n_18294, n_18295, n_18296, n_18297, n_18298, n_18299, n_18300, n_18301, n_18302, n_18303, n_18304, n_18305, n_18306, n_18307, n_18308, n_18309, n_18310, n_18311, n_18312, n_18313, n_18314, n_18315, n_18316, n_18317, n_18318, n_18319, n_18320, n_18321, n_18322, n_18323, n_18324, n_18325, n_18326, n_18327, n_18328, n_18329, n_18330, n_18331, n_18332, n_18333, n_18334, n_18335, n_18336, n_18337, n_18338, n_18339, n_18340, n_18341, n_18342, n_18343, n_18344, n_18345, n_18346, n_18347, n_18348, n_18349, n_18350, n_18351, n_18352, n_18353, n_18354, n_18355, n_18356, n_18357, y40, n_18358, n_18359, n_18360, n_18361, n_18362, n_18363, n_18364, n_18365, n_18366, n_18367, n_18368, n_18369, n_18370, n_18371, n_18372, n_18373, n_18374, n_18375, n_18376, n_18377, n_18378, n_18379, n_18380, n_18381, n_18382, n_18383, n_18384, n_18385, n_18386, n_18387, n_18388, n_18389, n_18390, n_18391, n_18392, n_18393, n_18394, n_18395, n_18396, n_18397, n_18398, n_18399, n_18400, n_18401, n_18402, n_18403, n_18404, n_18405, n_18406, n_18407, n_18408, n_18409, n_18410, n_18411, n_18412, n_18413, n_18414, n_18415, n_18416, n_18417, n_18418, n_18419, n_18420, y41, n_18421, n_18422, n_18423, n_18424, n_18425, n_18426, n_18427, n_18428, n_18429, n_18430, n_18431, n_18432, n_18433, n_18434, n_18435, n_18436, n_18437, n_18438, n_18439, n_18440, n_18441, n_18442, n_18443, n_18444, n_18445, n_18446, n_18447, n_18448, n_18449, n_18450, n_18451, n_18452, n_18453, n_18454, n_18455, n_18456, n_18457, n_18458, n_18459, n_18460, n_18461, n_18462, n_18463, n_18464, n_18465, n_18466, n_18467, n_18468, n_18469, n_18470, n_18471, n_18472, n_18473, n_18474, n_18475, n_18476, n_18477, n_18478, n_18479, n_18480, n_18481, n_18482, n_18483, n_18484, n_18485, n_18486, n_18487, n_18488, y42, n_18489, n_18490, n_18491, n_18492, n_18493, n_18494, n_18495, n_18496, n_18497, n_18498, n_18499, n_18500, n_18501, n_18502, n_18503, n_18504, n_18505, n_18506, n_18507, n_18508, n_18509, n_18510, n_18511, n_18512, n_18513, n_18514, n_18515, n_18516, n_18517, n_18518, n_18519, n_18520, n_18521, n_18522, n_18523, n_18524, n_18525, n_18526, n_18527, n_18528, n_18529, n_18530, n_18531, n_18532, n_18533, n_18534, n_18535, n_18536, n_18537, n_18538, n_18539, n_18540, n_18541, n_18542, n_18543, n_18544, n_18545, n_18546, n_18547, y43, n_18548, n_18549, n_18550, n_18551, n_18552, n_18553, n_18554, n_18555, n_18556, n_18557, n_18558, n_18559, n_18560, n_18561, n_18562, n_18563, n_18564, n_18565, n_18566, n_18567, n_18568, n_18569, n_18570, n_18571, n_18572, n_18573, n_18574, n_18575, n_18576, n_18577, n_18578, n_18579, n_18580, n_18581, n_18582, n_18583, n_18584, n_18585, n_18586, n_18587, n_18588, n_18589, n_18590, n_18591, n_18592, n_18593, n_18594, n_18595, n_18596, n_18597, n_18598, n_18599, n_18600, n_18601, n_18602, y44, n_18603, n_18604, n_18605, n_18606, n_18607, n_18608, n_18609, n_18610, n_18611, n_18612, n_18613, n_18614, n_18615, n_18616, n_18617, n_18618, n_18619, n_18620, n_18621, n_18622, n_18623, n_18624, n_18625, n_18626, n_18627, n_18628, n_18629, n_18630, n_18631, n_18632, n_18633, n_18634, n_18635, n_18636, n_18637, n_18638, n_18639, n_18640, n_18641, n_18642, n_18643, n_18644, n_18645, n_18646, n_18647, n_18648, n_18649, n_18650, n_18651, n_18652, n_18653, n_18654, n_18655, y45, n_18656, n_18657, n_18658, n_18659, n_18660, n_18661, n_18662, n_18663, n_18664, n_18665, n_18666, n_18667, n_18668, n_18669, n_18670, n_18671, n_18672, n_18673, n_18674, n_18675, n_18676, n_18677, n_18678, n_18679, n_18680, n_18681, n_18682, n_18683, n_18684, n_18685, n_18686, n_18687, n_18688, n_18689, n_18690, n_18691, n_18692, n_18693, n_18694, n_18695, n_18696, n_18697, n_18698, n_18699, n_18700, n_18701, n_18702, n_18703, n_18704, y46, n_18705, n_18706, n_18707, n_18708, n_18709, n_18710, n_18711, n_18712, n_18713, n_18714, n_18715, n_18716, n_18717, n_18718, n_18719, n_18720, n_18721, n_18722, n_18723, n_18724, n_18725, n_18726, n_18727, n_18728, n_18729, n_18730, n_18731, n_18732, n_18733, n_18734, n_18735, n_18736, n_18737, n_18738, n_18739, n_18740, n_18741, n_18742, n_18743, n_18744, n_18745, n_18746, n_18747, n_18748, n_18749, n_18750, n_18751, y47, n_18752, n_18753, n_18754, n_18755, n_18756, n_18757, n_18758, n_18759, n_18760, n_18761, n_18762, n_18763, n_18764, n_18765, n_18766, n_18767, n_18768, n_18769, n_18770, n_18771, n_18772, n_18773, n_18774, n_18775, n_18776, n_18777, n_18778, n_18779, n_18780, n_18781, n_18782, n_18783, n_18784, n_18785, n_18786, n_18787, n_18788, n_18789, n_18790, n_18791, n_18792, n_18793, n_18794, n_18795, y48, n_18796, n_18797, n_18798, n_18799, n_18800, n_18801, n_18802, n_18803, n_18804, n_18805, n_18806, n_18807, n_18808, n_18809, n_18810, n_18811, n_18812, n_18813, n_18814, n_18815, n_18816, n_18817, n_18818, n_18819, n_18820, n_18821, n_18822, n_18823, n_18824, n_18825, n_18826, n_18827, n_18828, n_18829, n_18830, n_18831, n_18832, n_18833, n_18834, n_18835, n_18836, y49, n_18837, n_18838, n_18839, n_18840, n_18841, n_18842, n_18843, n_18844, n_18845, n_18846, n_18847, n_18848, n_18849, n_18850, n_18851, n_18852, n_18853, n_18854, n_18855, n_18856, n_18857, n_18858, n_18859, n_18860, n_18861, n_18862, n_18863, n_18864, n_18865, n_18866, n_18867, n_18868, n_18869, n_18870, n_18871, n_18872, n_18873, n_18874, n_18875, y50, n_18876, n_18877, n_18878, n_18879, n_18880, n_18881, n_18882, n_18883, n_18884, n_18885, n_18886, n_18887, n_18888, n_18889, n_18890, n_18891, n_18892, n_18893, n_18894, n_18895, n_18896, n_18897, n_18898, n_18899, n_18900, n_18901, n_18902, n_18903, n_18904, n_18905, n_18906, n_18907, n_18908, n_18909, n_18910, n_18911, n_18912, n_18913, n_18914, n_18915, n_18916, y51, n_18917, n_18918, n_18919, n_18920, n_18921, n_18922, n_18923, n_18924, n_18925, n_18926, n_18927, n_18928, n_18929, n_18930, n_18931, n_18932, n_18933, n_18934, n_18935, n_18936, n_18937, n_18938, n_18939, n_18940, n_18941, n_18942, n_18943, n_18944, n_18945, n_18946, n_18947, n_18948, n_18949, n_18950, n_18951, n_18952, n_18953, n_18954, n_18955, n_18956, n_18957, y52, n_18958, n_18959, n_18960, n_18961, n_18962, n_18963, n_18964, n_18965, n_18966, n_18967, n_18968, n_18969, n_18970, n_18971, n_18972, n_18973, n_18974, n_18975, n_18976, n_18977, n_18978, n_18979, n_18980, n_18981, n_18982, n_18983, n_18984, n_18985, n_18986, n_18987, n_18988, n_18989, n_18990, n_18991, n_18992, n_18993, n_18994, n_18995, n_18996, y53, n_18997, n_18998, n_18999, n_19000, n_19001, n_19002, n_19003, n_19004, n_19005, n_19006, n_19007, n_19008, n_19009, n_19010, n_19011, n_19012, n_19013, n_19014, n_19015, n_19016, n_19017, n_19018, n_19019, n_19020, n_19021, n_19022, n_19023, n_19024, n_19025, n_19026, n_19027, n_19028, n_19029, n_19030, n_19031, n_19032, n_19033, n_19034, n_19035, n_19036, n_19037, n_19038, n_19039, n_19040, n_19041, n_19042, n_19043, n_19044, n_19045, n_19046, n_19047, n_19048, n_19049, y54, n_19050, n_19051, n_19052, n_19053, n_19054, n_19055, n_19056, n_19057, n_19058, n_19059, n_19060, n_19061, n_19062, n_19063, n_19064, n_19065, n_19066, n_19067, n_19068, n_19069, n_19070, n_19071, n_19072, n_19073, n_19074, n_19075, n_19076, n_19077, n_19078, n_19079, n_19080, n_19081, n_19082, n_19083, n_19084, n_19085, n_19086, n_19087, n_19088, n_19089, n_19090, n_19091, n_19092, n_19093, n_19094, n_19095, n_19096, n_19097, n_19098, n_19099, n_19100, n_19101, n_19102, n_19103, n_19104, n_19105, n_19106, n_19107, n_19108, n_19109, n_19110, y55, n_19111, n_19112, n_19113, n_19114, n_19115, n_19116, n_19117, n_19118, n_19119, n_19120, n_19121, n_19122, n_19123, n_19124, n_19125, n_19126, n_19127, n_19128, n_19129, n_19130, n_19131, n_19132, n_19133, n_19134, n_19135, n_19136, n_19137, n_19138, n_19139, n_19140, n_19141, n_19142, n_19143, n_19144, n_19145, n_19146, n_19147, n_19148, n_19149, n_19150, n_19151, n_19152, n_19153, n_19154, n_19155, n_19156, n_19157, n_19158, y56, n_19159, n_19160, n_19161, n_19162, n_19163, n_19164, n_19165, n_19166, n_19167, n_19168, n_19169, n_19170, n_19171, n_19172, n_19173, n_19174, n_19175, n_19176, n_19177, n_19178, n_19179, n_19180, y57, n_19181, n_19182, n_19183, n_19184, n_19185, n_19186, n_19187, n_19188, y58, n_19189, n_19190, n_19191, n_19192, n_19193, n_19194, n_19195, y60, n_19196, n_19197, y59, n_19198, n_19199, n_19200, n_19201, n_19202, y61, y62, n_19203, n_19204, n_19205, n_19206, y63, n_19207, n_19208, n_19209, n_19210, y64, n_19211, n_19212, n_19213, n_19214, y65, n_19215, n_19216, n_19217, n_19218, y66, n_19219, n_19220, n_19221, n_19222, y67, n_19223, n_19224, n_19225, n_19226, n_19227, n_19228, y68, n_19229, n_19230, n_19231, n_19232, n_19233, n_19234, n_19235, n_19236, n_19237, n_19238, n_19239, y69, y70, n_19240, n_19241, n_19242, n_19243, n_19244, y71, n_19245, n_19246, n_19247, n_19248, n_19249, n_19250, y73, n_19251, y72, n_19252, n_19253, n_19254, y74, n_19255, n_19256, n_19257, n_19258, y75, n_19259, n_19260, n_19261, n_19262, y76, n_19263, n_19264, n_19265, n_19266, n_19267, n_19268, y77, n_19269, n_19270, n_19271, n_19272, n_19273, n_19274, n_19275, y78, n_19276, n_19277, n_19278, n_19279, n_19280, n_19281, y79, n_19282, n_19283, n_19284, n_19285, n_19286, n_19287, n_19288, n_19289, n_19290, n_19291, n_19292, y80, n_19293, n_19294, n_19295, n_19296, y81, n_19297, n_19298, n_19299, n_19300, n_19301, n_19302, n_19303, y82, n_19304, n_19305, n_19306, n_19307, y83, n_19308, n_19309, n_19310, n_19311, n_19312, n_19313, y85, n_19314, y84, n_19315, n_19316, n_19317, y86, n_19318, n_19319, n_19320, n_19321, n_19322, n_19323, y87, n_19324, n_19325, n_19326, n_19327, n_19328, n_19329, n_19330, y88, n_19331, n_19332, n_19333, n_19334, n_19335, y89, n_19336, n_19337, n_19338, n_19339, n_19340, n_19341, n_19342, n_19343, n_19344, y91, n_19345, n_19346, n_19347, n_19348, n_19349, n_19350, y90, y92, n_19351, n_19352, n_19353, n_19354, n_19355, n_19356, y93, n_19357, n_19358, n_19359, n_19360, n_19361, n_19362, n_19363, y95, n_19364, n_19365, n_19366, y94, n_19367, n_19368, y96, n_19369, n_19370, n_19371, n_19372, n_19373, y97, n_19374, n_19375, n_19376, n_19377, n_19378, n_19379, n_19380, y99, n_19381, n_19382, n_19383, y98, n_19384, n_19385, y100, n_19386, n_19387, n_19388, n_19389, y101, n_19390, n_19391, n_19392, n_19393, n_19394, n_19395, n_19396, y102, n_19397, n_19398, n_19399, n_19400, n_19401, n_19402, n_19403, n_19404, n_19405, n_19406, y103, n_19407, n_19408, n_19409, y104, n_19410, n_19411, n_19412, n_19413, n_19414, n_19415, y106, n_19416, y105, n_19417, n_19418, n_19419, n_19420, n_19421, n_19422, y107, n_19423, n_19424, n_19425, n_19426, n_19427, n_19428, n_19429, n_19430, n_19431, n_19432, y108, n_19433, n_19434, n_19435, n_19436, n_19437, y109, n_19438, n_19439, n_19440, n_19441, n_19442, n_19443, n_19444, n_19445, n_19446, n_19447, y110, n_19448, n_19449, n_19450, n_19451, n_19452, y111, n_19453, n_19454, n_19455, n_19456, n_19457, n_19458, n_19459, n_19460, n_19461, n_19462, n_19463, n_19464, n_19465, n_19466, y113, n_19467, n_19468, n_19469, n_19470, n_19471, n_19472, n_19473, n_19474, n_19475, n_19476, n_19477, n_19478, y112, n_19479, y115, n_19480, n_19481, n_19482, n_19483, n_19484, n_19485, y114, y116, n_19486, n_19487, n_19488, n_19489, n_19490, n_19491, n_19492, y117, n_19493, n_19494, n_19495, n_19496, n_19497, n_19498, n_19499, n_19500, n_19501, n_19502, n_19503, n_19504, y118, y119, n_19505, n_19506, n_19507, n_19508, n_19509, n_19510, n_19511, n_19512, n_19513, n_19514, y121, n_19515, n_19516, n_19517, y120, n_19518, n_19519, n_19520, n_19521, y122, n_19522, n_19523, n_19524, n_19525, n_19526, n_19527, n_19528, n_19529, y124, n_19530, n_19531, n_19532, y123, n_19533, n_19534, y125, n_19535, n_19536, n_19537, n_19538, y126, n_19539, n_19540, n_19541, y127;
assign n_0 = x1 ^ x0;
assign n_1 = x2 ^ x1;
assign n_2 = ~x1 & x2;
assign n_3 = x3 ^ x2;
assign n_4 = x2 & x3;
assign n_5 = x4 ^ x2;
assign n_6 = x5 ^ x4;
assign n_7 = x5 ^ x2;
assign n_8 = x6 ^ x5;
assign n_9 = ~x5 & ~x6;
assign n_10 = x7 ^ x6;
assign n_11 = x8 ^ x7;
assign n_12 = x9 ^ x8;
assign n_13 = ~x8 & ~x9;
assign n_14 = x11 ^ x10;
assign n_15 = x12 ^ x11;
assign n_16 = x11 & x12;
assign n_17 = x14 ^ x13;
assign n_18 = x15 ^ x14;
assign n_19 = ~x14 & ~x15;
assign n_20 = x17 ^ x16;
assign n_21 = x18 ^ x17;
assign n_22 = ~x17 & ~x18;
assign n_23 = x20 ^ x19;
assign n_24 = x21 ^ x20;
assign n_25 = ~x20 & ~x21;
assign n_26 = x23 ^ x22;
assign n_27 = x24 ^ x23;
assign n_28 = x23 & x24;
assign n_29 = x26 ^ x25;
assign n_30 = x27 ^ x26;
assign n_31 = x26 & x27;
assign n_32 = x29 ^ x28;
assign n_33 = x30 ^ x29;
assign n_34 = ~x29 & ~x30;
assign n_35 = x32 ^ x31;
assign n_36 = x33 ^ x32;
assign n_37 = ~x32 & ~x33;
assign n_38 = x35 ^ x34;
assign n_39 = x36 ^ x35;
assign n_40 = ~x35 & ~x36;
assign n_41 = x38 ^ x37;
assign n_42 = x39 ^ x38;
assign n_43 = ~x38 & ~x39;
assign n_44 = x41 ^ x40;
assign n_45 = x42 ^ x41;
assign n_46 = ~x41 & ~x42;
assign n_47 = x44 ^ x43;
assign n_48 = x45 ^ x44;
assign n_49 = ~x44 & ~x45;
assign n_50 = x47 ^ x46;
assign n_51 = x48 ^ x47;
assign n_52 = ~x47 & ~x48;
assign n_53 = x50 ^ x49;
assign n_54 = x51 ^ x50;
assign n_55 = ~x50 & ~x51;
assign n_56 = x53 ^ x52;
assign n_57 = x54 ^ x53;
assign n_58 = x53 & x54;
assign n_59 = x56 ^ x55;
assign n_60 = x57 ^ x56;
assign n_61 = x56 & x57;
assign n_62 = x59 ^ x58;
assign n_63 = x60 ^ x59;
assign n_64 = x59 & x60;
assign n_65 = x62 ^ x61;
assign n_66 = x63 ^ x62;
assign n_67 = x62 & ~x63;
assign n_68 = x0 & x64;
assign n_69 = x1 & x64;
assign n_70 = x2 & x64;
assign n_71 = x3 & x64;
assign n_72 = ~x7 & x64;
assign n_73 = ~x10 & x64;
assign n_74 = x13 & x64;
assign n_75 = x28 & x64;
assign n_76 = ~x49 & x64;
assign n_77 = ~x52 & x64;
assign n_78 = x63 & x64;
assign n_79 = x0 & x65;
assign n_80 = x1 & x65;
assign n_81 = x2 & ~x65;
assign n_82 = ~x64 & ~x65;
assign n_83 = x65 ^ x3;
assign n_84 = x65 ^ x9;
assign n_85 = x65 ^ x12;
assign n_86 = x65 ^ x15;
assign n_87 = x65 ^ x18;
assign n_88 = x65 ^ x21;
assign n_89 = x65 ^ x24;
assign n_90 = x65 ^ x27;
assign n_91 = x65 ^ x30;
assign n_92 = x65 ^ x33;
assign n_93 = x65 ^ x36;
assign n_94 = x65 ^ x39;
assign n_95 = x65 ^ x42;
assign n_96 = x65 ^ x45;
assign n_97 = x65 ^ x48;
assign n_98 = x65 ^ x51;
assign n_99 = x65 ^ x54;
assign n_100 = x65 ^ x57;
assign n_101 = x65 ^ x60;
assign n_102 = x63 & x65;
assign n_103 = x66 ^ x2;
assign n_104 = ~x64 & x66;
assign n_105 = x65 & x66;
assign n_106 = x66 ^ x65;
assign n_107 = x1 & x67;
assign n_108 = x67 ^ x2;
assign n_109 = x67 ^ x66;
assign n_110 = x63 & x67;
assign n_111 = x68 ^ x2;
assign n_112 = x63 & x68;
assign n_113 = x1 & x69;
assign n_114 = x2 & ~x69;
assign n_115 = x63 & x69;
assign n_116 = x70 ^ x2;
assign n_117 = x71 ^ x70;
assign n_118 = x1 & x71;
assign n_119 = x2 & ~x71;
assign n_120 = x71 & ~x72;
assign n_121 = x72 ^ x71;
assign n_122 = x72 ^ x2;
assign n_123 = x2 & ~x72;
assign n_124 = x72 ^ x8;
assign n_125 = x72 & ~x73;
assign n_126 = x73 ^ x2;
assign n_127 = x73 ^ x71;
assign n_128 = x1 & x74;
assign n_129 = x2 & ~x74;
assign n_130 = x74 ^ x73;
assign n_131 = x75 ^ x2;
assign n_132 = ~x74 & x75;
assign n_133 = x63 & x75;
assign n_134 = x1 & x76;
assign n_135 = x63 & x76;
assign n_136 = x1 & x77;
assign n_137 = x2 & ~x77;
assign n_138 = x77 ^ x76;
assign n_139 = x78 ^ x77;
assign n_140 = x78 ^ x2;
assign n_141 = x63 & x78;
assign n_142 = x79 ^ x78;
assign n_143 = x1 & x79;
assign n_144 = x79 ^ x2;
assign n_145 = x80 ^ x79;
assign n_146 = x80 ^ x2;
assign n_147 = x2 & ~x80;
assign n_148 = x63 & x80;
assign n_149 = x81 ^ x80;
assign n_150 = x81 ^ x2;
assign n_151 = ~x80 & x81;
assign n_152 = x81 ^ x17;
assign n_153 = x82 ^ x81;
assign n_154 = x1 & x82;
assign n_155 = x82 ^ x2;
assign n_156 = x82 ^ x80;
assign n_157 = x83 ^ x82;
assign n_158 = x83 ^ x2;
assign n_159 = x2 & ~x83;
assign n_160 = x84 ^ x83;
assign n_161 = x84 ^ x2;
assign n_162 = x2 & ~x84;
assign n_163 = x84 ^ x20;
assign n_164 = x85 ^ x84;
assign n_165 = x85 ^ x2;
assign n_166 = x2 & ~x85;
assign n_167 = x85 ^ x83;
assign n_168 = x86 ^ x85;
assign n_169 = x86 ^ x2;
assign n_170 = x2 & ~x86;
assign n_171 = x87 ^ x86;
assign n_172 = x87 ^ x2;
assign n_173 = x2 & ~x87;
assign n_174 = x87 ^ x23;
assign n_175 = x88 ^ x87;
assign n_176 = x88 ^ x2;
assign n_177 = x2 & ~x88;
assign n_178 = x88 ^ x86;
assign n_179 = x89 ^ x88;
assign n_180 = x89 ^ x2;
assign n_181 = x2 & ~x89;
assign n_182 = x90 ^ x89;
assign n_183 = x90 ^ x2;
assign n_184 = x90 ^ x26;
assign n_185 = x91 ^ x90;
assign n_186 = x91 ^ x2;
assign n_187 = x91 ^ x89;
assign n_188 = x63 & x91;
assign n_189 = x92 ^ x91;
assign n_190 = x92 ^ x2;
assign n_191 = x2 & ~x92;
assign n_192 = ~x91 & x92;
assign n_193 = x93 ^ x92;
assign n_194 = x93 ^ x91;
assign n_195 = x93 ^ x2;
assign n_196 = ~x92 & x93;
assign n_197 = x93 ^ x29;
assign n_198 = x94 ^ x93;
assign n_199 = x94 ^ x2;
assign n_200 = x2 & ~x94;
assign n_201 = x94 ^ x92;
assign n_202 = x95 ^ x94;
assign n_203 = x95 ^ x2;
assign n_204 = x2 & ~x95;
assign n_205 = x96 ^ x95;
assign n_206 = x96 ^ x94;
assign n_207 = x96 ^ x2;
assign n_208 = x96 ^ x32;
assign n_209 = x97 ^ x96;
assign n_210 = x97 ^ x94;
assign n_211 = x1 & x97;
assign n_212 = x2 & ~x97;
assign n_213 = x97 ^ x95;
assign n_214 = x98 ^ x97;
assign n_215 = x98 ^ x2;
assign n_216 = x99 ^ x98;
assign n_217 = x1 & x99;
assign n_218 = x99 ^ x2;
assign n_219 = x99 ^ x35;
assign n_220 = x100 ^ x99;
assign n_221 = x100 ^ x2;
assign n_222 = x2 & x100;
assign n_223 = x100 ^ x98;
assign n_224 = x101 ^ x100;
assign n_225 = x101 ^ x98;
assign n_226 = x2 & ~x101;
assign n_227 = ~x100 ^ x101;
assign n_228 = x102 ^ x2;
assign n_229 = x2 & ~x102;
assign n_230 = ~x101 ^ x102;
assign n_231 = x63 & x102;
assign n_232 = x103 ^ x2;
assign n_233 = x63 & x103;
assign n_234 = x1 & x104;
assign n_235 = x2 & ~x104;
assign n_236 = x63 & x104;
assign n_237 = x105 ^ x2;
assign n_238 = x63 & x105;
assign n_239 = x1 & x106;
assign n_240 = x2 & ~x106;
assign n_241 = x63 & x106;
assign n_242 = x107 ^ x106;
assign n_243 = x107 ^ x2;
assign n_244 = x108 ^ x107;
assign n_245 = x108 ^ x2;
assign n_246 = ~x107 & x108;
assign n_247 = x63 & x108;
assign n_248 = x109 ^ x108;
assign n_249 = x109 ^ x2;
assign n_250 = x2 & ~x109;
assign n_251 = x110 ^ x2;
assign n_252 = x2 & ~x110;
assign n_253 = x110 ^ x109;
assign n_254 = x111 ^ x2;
assign n_255 = x111 ^ x110;
assign n_256 = x111 ^ x47;
assign n_257 = x1 & x112;
assign n_258 = x2 & ~x112;
assign n_259 = x112 ^ x110;
assign n_260 = x63 & x112;
assign n_261 = x113 ^ x2;
assign n_262 = x2 & ~x113;
assign n_263 = x113 ^ x112;
assign n_264 = x114 ^ x2;
assign n_265 = x114 ^ x113;
assign n_266 = x113 & ~x114;
assign n_267 = x63 & x114;
assign n_268 = x115 ^ x2;
assign n_269 = x116 ^ x2;
assign n_270 = x1 & x117;
assign n_271 = x117 ^ x53;
assign n_272 = x118 ^ x117;
assign n_273 = x1 & x118;
assign n_274 = x118 ^ x116;
assign n_275 = x118 ^ x63;
assign n_276 = x119 ^ x118;
assign n_277 = x1 & x119;
assign n_278 = ~x117 & ~x119;
assign n_279 = ~x118 & x119;
assign n_280 = ~x118 & ~x120;
assign n_281 = ~x119 & x120;
assign n_282 = x1 & x120;
assign n_283 = x63 & x120;
assign n_284 = x1 & x121;
assign n_285 = x1 & x122;
assign n_286 = x123 ^ x122;
assign n_287 = x1 & x123;
assign n_288 = x123 ^ x59;
assign n_289 = x1 & x124;
assign n_290 = x124 ^ x2;
assign n_291 = x124 ^ x122;
assign n_292 = ~x124 & x125;
assign n_293 = x125 ^ x124;
assign n_294 = x125 ^ x2;
assign n_295 = x2 & ~x125;
assign n_296 = x125 & ~x126;
assign n_297 = x126 ^ x125;
assign n_298 = x126 ^ x2;
assign n_299 = ~x1 & x126;
assign n_300 = x126 ^ x124;
assign n_301 = x124 & x126;
assign n_302 = x2 & ~x127;
assign n_303 = ~x126 & x127;
assign n_304 = x127 ^ x126;
assign n_305 = ~x7 & x127;
assign n_306 = ~x10 & x127;
assign n_307 = ~x31 & x127;
assign n_308 = x127 ^ x125;
assign n_309 = x127 ^ x62;
assign n_310 = x125 & x127;
assign n_311 = n_1 ^ x127;
assign n_312 = x66 & n_2;
assign n_313 = x68 & n_2;
assign n_314 = x70 & n_2;
assign n_315 = x73 & n_2;
assign n_316 = x75 & n_2;
assign n_317 = x76 & n_2;
assign n_318 = x78 & n_2;
assign n_319 = x81 & n_2;
assign n_320 = x96 & n_2;
assign n_321 = x98 & n_2;
assign n_322 = x103 & n_2;
assign n_323 = x105 & n_2;
assign n_324 = x111 & n_2;
assign n_325 = x116 & n_2;
assign n_326 = x117 & n_2;
assign n_327 = x118 & n_2;
assign n_328 = x119 & n_2;
assign n_329 = x120 & n_2;
assign n_330 = x121 & n_2;
assign n_331 = x122 & n_2;
assign n_332 = x123 & n_2;
assign n_333 = x4 & ~n_3;
assign n_334 = x66 & n_3;
assign n_335 = x5 & ~n_3;
assign n_336 = n_4 ^ x4;
assign n_337 = x64 & n_5;
assign n_338 = n_3 & ~n_6;
assign n_339 = x64 & n_8;
assign n_340 = x66 & n_8;
assign n_341 = ~x8 & ~n_8;
assign n_342 = n_9 ^ n_8;
assign n_343 = x65 & ~n_9;
assign n_344 = n_9 ^ x7;
assign n_345 = ~n_8 & n_10;
assign n_346 = n_8 & ~n_11;
assign n_347 = x64 & n_12;
assign n_348 = ~x10 & ~n_12;
assign n_349 = x66 & n_12;
assign n_350 = x11 & ~n_12;
assign n_351 = n_13 ^ n_12;
assign n_352 = n_13 ^ x10;
assign n_353 = x64 & n_15;
assign n_354 = x13 & ~n_15;
assign n_355 = x66 & n_15;
assign n_356 = x14 & ~n_15;
assign n_357 = n_15 & ~n_17;
assign n_358 = x64 & n_18;
assign n_359 = x16 & ~n_18;
assign n_360 = x66 & n_18;
assign n_361 = x17 & ~n_18;
assign n_362 = n_19 ^ n_18;
assign n_363 = n_18 & ~n_20;
assign n_364 = x64 & n_21;
assign n_365 = x19 & ~n_21;
assign n_366 = x66 & n_21;
assign n_367 = x20 & ~n_21;
assign n_368 = n_22 ^ n_21;
assign n_369 = n_21 & ~n_23;
assign n_370 = x64 & n_24;
assign n_371 = x22 & ~n_24;
assign n_372 = x66 & n_24;
assign n_373 = x23 & ~n_24;
assign n_374 = n_25 ^ n_24;
assign n_375 = n_24 & ~n_26;
assign n_376 = x64 & n_27;
assign n_377 = x25 & ~n_27;
assign n_378 = x66 & n_27;
assign n_379 = x26 & ~n_27;
assign n_380 = n_28 ^ x25;
assign n_381 = n_27 & ~n_29;
assign n_382 = x64 & n_30;
assign n_383 = x28 & ~n_30;
assign n_384 = x66 & n_30;
assign n_385 = x29 & ~n_30;
assign n_386 = n_31 ^ x28;
assign n_387 = n_30 & ~n_32;
assign n_388 = x64 & n_33;
assign n_389 = x31 & ~n_33;
assign n_390 = x66 & n_33;
assign n_391 = x32 & ~n_33;
assign n_392 = n_34 ^ n_33;
assign n_393 = n_34 ^ x31;
assign n_394 = n_33 & ~n_35;
assign n_395 = x64 & n_36;
assign n_396 = x34 & ~n_36;
assign n_397 = x66 & n_36;
assign n_398 = x35 & ~n_36;
assign n_399 = n_37 ^ n_36;
assign n_400 = n_36 & ~n_38;
assign n_401 = x64 & n_39;
assign n_402 = x37 & ~n_39;
assign n_403 = x66 & n_39;
assign n_404 = x38 & ~n_39;
assign n_405 = n_40 ^ n_39;
assign n_406 = n_39 & ~n_41;
assign n_407 = x64 & n_42;
assign n_408 = x40 & ~n_42;
assign n_409 = x66 & n_42;
assign n_410 = x41 & ~n_42;
assign n_411 = n_43 ^ x40;
assign n_412 = n_43 ^ n_42;
assign n_413 = n_42 & ~n_44;
assign n_414 = x64 & n_45;
assign n_415 = x43 & ~n_45;
assign n_416 = x66 & n_45;
assign n_417 = x44 & ~n_45;
assign n_418 = n_46 ^ n_45;
assign n_419 = n_45 & ~n_47;
assign n_420 = x64 & n_48;
assign n_421 = x47 & ~n_48;
assign n_422 = x46 & ~n_48;
assign n_423 = x66 & n_48;
assign n_424 = n_49 ^ n_48;
assign n_425 = n_48 & ~n_50;
assign n_426 = x64 & n_51;
assign n_427 = x49 & ~n_51;
assign n_428 = x66 & n_51;
assign n_429 = x50 & ~n_51;
assign n_430 = n_52 ^ n_51;
assign n_431 = n_51 & ~n_53;
assign n_432 = x64 & n_54;
assign n_433 = x53 & ~n_54;
assign n_434 = x52 & ~n_54;
assign n_435 = x66 & n_54;
assign n_436 = n_55 ^ n_54;
assign n_437 = n_54 & ~n_56;
assign n_438 = x64 & n_57;
assign n_439 = x55 & ~n_57;
assign n_440 = x66 & n_57;
assign n_441 = x56 & ~n_57;
assign n_442 = n_58 ^ x55;
assign n_443 = n_57 & ~n_59;
assign n_444 = x64 & n_60;
assign n_445 = x58 & ~n_60;
assign n_446 = x66 & n_60;
assign n_447 = x59 & ~n_60;
assign n_448 = n_61 ^ x58;
assign n_449 = n_60 & ~n_62;
assign n_450 = x64 & n_63;
assign n_451 = x61 & ~n_63;
assign n_452 = x66 & n_63;
assign n_453 = x62 & ~n_63;
assign n_454 = n_64 ^ x61;
assign n_455 = n_63 & ~n_65;
assign n_456 = x64 & n_66;
assign n_457 = x71 & n_66;
assign n_458 = n_66 ^ x71;
assign n_459 = ~x72 & n_66;
assign n_460 = x74 & n_66;
assign n_461 = x83 & n_66;
assign n_462 = ~x84 & n_66;
assign n_463 = n_66 ^ x83;
assign n_464 = x86 & n_66;
assign n_465 = x89 & n_66;
assign n_466 = ~x90 & n_66;
assign n_467 = n_66 ^ x89;
assign n_468 = x95 & n_66;
assign n_469 = n_66 ^ x95;
assign n_470 = ~x96 & n_66;
assign n_471 = x98 & n_66;
assign n_472 = n_66 ^ x98;
assign n_473 = ~x99 & n_66;
assign n_474 = x101 & n_66;
assign n_475 = ~x102 & n_66;
assign n_476 = x110 & n_66;
assign n_477 = n_66 ^ x110;
assign n_478 = ~x111 & n_66;
assign n_479 = x116 & n_66;
assign n_480 = ~x117 & n_66;
assign n_481 = n_66 ^ x116;
assign n_482 = n_66 ^ x119;
assign n_483 = x122 & n_66;
assign n_484 = ~x123 & n_66;
assign n_485 = n_66 ^ x122;
assign n_486 = x125 & n_66;
assign n_487 = n_67 ^ x62;
assign n_488 = n_67 ^ x63;
assign y0 = n_68;
assign n_489 = ~x0 & ~n_70;
assign n_490 = n_71 ^ x2;
assign n_491 = n_72 ^ x64;
assign n_492 = n_9 & n_72;
assign n_493 = n_13 & n_73;
assign n_494 = n_16 & n_74;
assign n_495 = n_31 & n_75;
assign n_496 = n_75 ^ x64;
assign n_497 = n_52 & n_76;
assign n_498 = n_55 & n_77;
assign n_499 = n_78 ^ x65;
assign n_500 = n_79 ^ n_69;
assign n_501 = ~x0 & ~n_80;
assign n_502 = n_82 ^ x64;
assign n_503 = x41 & ~n_82;
assign n_504 = n_3 & ~n_83;
assign n_505 = n_12 & ~n_84;
assign n_506 = n_15 & ~n_85;
assign n_507 = n_18 & ~n_86;
assign n_508 = n_21 & ~n_87;
assign n_509 = n_24 & ~n_88;
assign n_510 = n_27 & ~n_89;
assign n_511 = n_30 & ~n_90;
assign n_512 = n_33 & ~n_91;
assign n_513 = n_36 & ~n_92;
assign n_514 = n_39 & ~n_93;
assign n_515 = n_42 & ~n_94;
assign n_516 = n_45 & ~n_95;
assign n_517 = n_48 & ~n_96;
assign n_518 = n_51 & ~n_97;
assign n_519 = n_54 & ~n_98;
assign n_520 = n_57 & ~n_99;
assign n_521 = n_60 & ~n_100;
assign n_522 = n_63 & ~n_101;
assign n_523 = n_102 ^ x66;
assign n_524 = n_68 & ~n_103;
assign n_525 = n_81 ^ n_103;
assign n_526 = n_104 ^ x64;
assign n_527 = n_104 ^ x0;
assign n_528 = ~x67 & ~n_105;
assign n_529 = n_106 ^ n_104;
assign n_530 = ~x67 & ~n_108;
assign n_531 = ~x63 & n_109;
assign n_532 = n_110 ^ x2;
assign n_533 = n_112 ^ x68;
assign n_534 = n_112 ^ x2;
assign n_535 = n_115 ^ x69;
assign n_536 = n_115 ^ x2;
assign n_537 = n_115 ^ x70;
assign n_538 = n_116 ^ n_114;
assign n_539 = n_120 ^ n_121;
assign n_540 = n_119 ^ n_122;
assign n_541 = n_123 ^ n_126;
assign n_542 = n_129 ^ n_131;
assign n_543 = n_132 ^ n_130;
assign n_544 = n_133 ^ x76;
assign n_545 = n_135 ^ x77;
assign n_546 = x63 & n_138;
assign n_547 = n_139 ^ x62;
assign n_548 = x63 & n_139;
assign n_549 = n_137 ^ n_140;
assign n_550 = n_141 ^ x79;
assign n_551 = ~x79 & ~n_144;
assign n_552 = ~x63 & n_145;
assign n_553 = n_149 ^ x62;
assign n_554 = n_147 ^ n_150;
assign n_555 = n_151 ^ n_149;
assign n_556 = ~x82 & ~n_155;
assign n_557 = n_161 ^ n_159;
assign n_558 = n_162 ^ n_165;
assign n_559 = x63 & n_168;
assign n_560 = n_166 ^ n_169;
assign n_561 = n_170 ^ n_172;
assign n_562 = n_173 ^ n_176;
assign n_563 = n_180 ^ n_177;
assign n_564 = n_183 ^ n_181;
assign n_565 = ~x90 & ~n_183;
assign n_566 = ~x91 & ~n_186;
assign n_567 = n_188 ^ x92;
assign n_568 = n_192 ^ n_189;
assign n_569 = x63 & n_192;
assign n_570 = n_191 ^ n_195;
assign n_571 = ~x93 & ~n_195;
assign n_572 = n_196 ^ n_193;
assign n_573 = n_200 ^ n_203;
assign n_574 = n_204 ^ n_207;
assign n_575 = n_210 ^ n_205;
assign n_576 = n_215 ^ n_212;
assign n_577 = ~x99 & ~n_218;
assign n_578 = n_222 ^ x101;
assign n_579 = n_225 ^ n_220;
assign n_580 = n_226 ^ n_228;
assign n_581 = ~n_230 ^ ~n_227;
assign n_582 = n_231 ^ x103;
assign n_583 = n_232 ^ n_229;
assign n_584 = n_233 ^ x104;
assign n_585 = n_236 ^ x105;
assign n_586 = n_235 ^ n_237;
assign n_587 = n_238 ^ x106;
assign n_588 = n_241 ^ x107;
assign n_589 = x63 & n_242;
assign n_590 = n_240 ^ n_243;
assign n_591 = ~x107 & ~n_243;
assign n_592 = n_244 ^ x62;
assign n_593 = ~x108 & ~n_245;
assign n_594 = n_246 ^ n_244;
assign n_595 = x63 & n_246;
assign n_596 = n_67 & ~n_246;
assign n_597 = n_247 ^ x109;
assign n_598 = n_250 ^ n_251;
assign n_599 = n_252 ^ n_254;
assign n_600 = n_260 ^ x113;
assign n_601 = n_258 ^ n_261;
assign n_602 = x63 & n_263;
assign n_603 = n_262 ^ n_264;
assign n_604 = ~x114 & ~n_264;
assign n_605 = n_265 ^ x62;
assign n_606 = n_266 ^ n_265;
assign n_607 = n_267 ^ x115;
assign n_608 = ~x115 & ~n_268;
assign n_609 = x118 & n_275;
assign n_610 = ~x117 & n_280;
assign n_611 = n_278 ^ n_280;
assign n_612 = x118 & n_281;
assign n_613 = n_279 ^ n_281;
assign n_614 = n_283 ^ x121;
assign n_615 = ~x124 & ~n_290;
assign n_616 = n_292 ^ n_293;
assign n_617 = n_296 ^ n_297;
assign n_618 = ~n_297 & n_66;
assign n_619 = n_295 ^ n_298;
assign n_620 = n_301 ^ x125;
assign n_621 = ~n_299 & n_302;
assign n_622 = n_303 ^ n_304;
assign n_623 = ~x2 & ~n_304;
assign n_624 = n_305 ^ x8;
assign n_625 = n_306 ^ x11;
assign n_626 = n_307 ^ x32;
assign n_627 = n_300 ^ n_308;
assign n_628 = n_308 ^ x62;
assign n_629 = n_67 & n_310;
assign n_630 = n_107 ^ n_312;
assign n_631 = n_113 ^ n_313;
assign n_632 = n_118 ^ n_314;
assign n_633 = n_128 ^ n_315;
assign n_634 = n_134 ^ n_316;
assign n_635 = n_136 ^ n_317;
assign n_636 = n_143 ^ n_318;
assign n_637 = n_154 ^ n_319;
assign n_638 = n_211 ^ n_320;
assign n_639 = n_217 ^ n_321;
assign n_640 = n_234 ^ n_322;
assign n_641 = n_239 ^ n_323;
assign n_642 = n_257 ^ n_324;
assign n_643 = n_270 ^ n_325;
assign n_644 = n_273 ^ n_326;
assign n_645 = n_277 ^ n_327;
assign n_646 = n_282 ^ n_328;
assign n_647 = n_284 ^ n_329;
assign n_648 = n_285 ^ n_330;
assign n_649 = n_287 ^ n_331;
assign n_650 = n_289 ^ n_332;
assign n_651 = n_333 ^ n_4;
assign n_652 = n_335 ^ n_4;
assign n_653 = ~x64 & n_336;
assign n_654 = n_337 ^ n_82;
assign n_655 = n_338 ^ n_3;
assign n_656 = x67 & n_338;
assign n_657 = x68 & n_338;
assign n_658 = x69 & n_338;
assign n_659 = x70 & n_338;
assign n_660 = x71 & n_338;
assign n_661 = x72 & n_338;
assign n_662 = x73 & n_338;
assign n_663 = x74 & n_338;
assign n_664 = x75 & n_338;
assign n_665 = x76 & n_338;
assign n_666 = x77 & n_338;
assign n_667 = x78 & n_338;
assign n_668 = x79 & n_338;
assign n_669 = x80 & n_338;
assign n_670 = x81 & n_338;
assign n_671 = x82 & n_338;
assign n_672 = x83 & n_338;
assign n_673 = x84 & n_338;
assign n_674 = x85 & n_338;
assign n_675 = x86 & n_338;
assign n_676 = x87 & n_338;
assign n_677 = x88 & n_338;
assign n_678 = x89 & n_338;
assign n_679 = x90 & n_338;
assign n_680 = x91 & n_338;
assign n_681 = x92 & n_338;
assign n_682 = x93 & n_338;
assign n_683 = x94 & n_338;
assign n_684 = x95 & n_338;
assign n_685 = x96 & n_338;
assign n_686 = x97 & n_338;
assign n_687 = x98 & n_338;
assign n_688 = x99 & n_338;
assign n_689 = x100 & n_338;
assign n_690 = x101 & n_338;
assign n_691 = x102 & n_338;
assign n_692 = x103 & n_338;
assign n_693 = x104 & n_338;
assign n_694 = x105 & n_338;
assign n_695 = x106 & n_338;
assign n_696 = x107 & n_338;
assign n_697 = x108 & n_338;
assign n_698 = x109 & n_338;
assign n_699 = x110 & n_338;
assign n_700 = x111 & n_338;
assign n_701 = x112 & n_338;
assign n_702 = x113 & n_338;
assign n_703 = x114 & n_338;
assign n_704 = x115 & n_338;
assign n_705 = x116 & n_338;
assign n_706 = x117 & n_338;
assign n_707 = x118 & n_338;
assign n_708 = x119 & n_338;
assign n_709 = x120 & n_338;
assign n_710 = x121 & n_338;
assign n_711 = x122 & n_338;
assign n_712 = x123 & n_338;
assign n_713 = x124 & n_338;
assign n_714 = x125 & n_338;
assign n_715 = x126 & n_338;
assign n_716 = x127 & n_338;
assign n_717 = n_341 ^ n_9;
assign n_718 = ~n_342 & ~n_72;
assign n_719 = x64 & ~n_342;
assign n_720 = n_11 & n_344;
assign n_721 = x65 & n_345;
assign n_722 = x66 & n_345;
assign n_723 = x67 & n_345;
assign n_724 = x68 & n_345;
assign n_725 = x69 & n_345;
assign n_726 = x70 & n_345;
assign n_727 = x71 & n_345;
assign n_728 = x72 & n_345;
assign n_729 = x73 & n_345;
assign n_730 = x74 & n_345;
assign n_731 = x75 & n_345;
assign n_732 = x76 & n_345;
assign n_733 = x77 & n_345;
assign n_734 = x78 & n_345;
assign n_735 = x79 & n_345;
assign n_736 = x80 & n_345;
assign n_737 = x81 & n_345;
assign n_738 = x82 & n_345;
assign n_739 = x83 & n_345;
assign n_740 = x84 & n_345;
assign n_741 = x85 & n_345;
assign n_742 = x86 & n_345;
assign n_743 = x87 & n_345;
assign n_744 = x88 & n_345;
assign n_745 = x89 & n_345;
assign n_746 = x90 & n_345;
assign n_747 = x91 & n_345;
assign n_748 = x92 & n_345;
assign n_749 = x93 & n_345;
assign n_750 = x94 & n_345;
assign n_751 = x95 & n_345;
assign n_752 = x96 & n_345;
assign n_753 = x97 & n_345;
assign n_754 = x98 & n_345;
assign n_755 = x99 & n_345;
assign n_756 = x100 & n_345;
assign n_757 = x101 & n_345;
assign n_758 = x102 & n_345;
assign n_759 = x103 & n_345;
assign n_760 = x104 & n_345;
assign n_761 = x105 & n_345;
assign n_762 = x106 & n_345;
assign n_763 = x107 & n_345;
assign n_764 = x108 & n_345;
assign n_765 = x109 & n_345;
assign n_766 = x110 & n_345;
assign n_767 = x111 & n_345;
assign n_768 = x112 & n_345;
assign n_769 = x113 & n_345;
assign n_770 = x114 & n_345;
assign n_771 = x115 & n_345;
assign n_772 = x116 & n_345;
assign n_773 = x117 & n_345;
assign n_774 = x118 & n_345;
assign n_775 = x119 & n_345;
assign n_776 = x120 & n_345;
assign n_777 = x121 & n_345;
assign n_778 = x122 & n_345;
assign n_779 = x123 & n_345;
assign n_780 = x124 & n_345;
assign n_781 = x125 & n_345;
assign n_782 = x126 & n_345;
assign n_783 = x127 & n_345;
assign n_784 = n_346 ^ n_8;
assign n_785 = x67 & n_346;
assign n_786 = x68 & n_346;
assign n_787 = x69 & n_346;
assign n_788 = x70 & n_346;
assign n_789 = x71 & n_346;
assign n_790 = x72 & n_346;
assign n_791 = x73 & n_346;
assign n_792 = x74 & n_346;
assign n_793 = x75 & n_346;
assign n_794 = x76 & n_346;
assign n_795 = x77 & n_346;
assign n_796 = x78 & n_346;
assign n_797 = x79 & n_346;
assign n_798 = x80 & n_346;
assign n_799 = x81 & n_346;
assign n_800 = x82 & n_346;
assign n_801 = x83 & n_346;
assign n_802 = x84 & n_346;
assign n_803 = x85 & n_346;
assign n_804 = x86 & n_346;
assign n_805 = x87 & n_346;
assign n_806 = x88 & n_346;
assign n_807 = x89 & n_346;
assign n_808 = x90 & n_346;
assign n_809 = x91 & n_346;
assign n_810 = x92 & n_346;
assign n_811 = x93 & n_346;
assign n_812 = x94 & n_346;
assign n_813 = x95 & n_346;
assign n_814 = x96 & n_346;
assign n_815 = x97 & n_346;
assign n_816 = x98 & n_346;
assign n_817 = x99 & n_346;
assign n_818 = x100 & n_346;
assign n_819 = x101 & n_346;
assign n_820 = x102 & n_346;
assign n_821 = x103 & n_346;
assign n_822 = x104 & n_346;
assign n_823 = x105 & n_346;
assign n_824 = x106 & n_346;
assign n_825 = x107 & n_346;
assign n_826 = x108 & n_346;
assign n_827 = x109 & n_346;
assign n_828 = x110 & n_346;
assign n_829 = x111 & n_346;
assign n_830 = x112 & n_346;
assign n_831 = x113 & n_346;
assign n_832 = x114 & n_346;
assign n_833 = x115 & n_346;
assign n_834 = x116 & n_346;
assign n_835 = x117 & n_346;
assign n_836 = x118 & n_346;
assign n_837 = x119 & n_346;
assign n_838 = x120 & n_346;
assign n_839 = x121 & n_346;
assign n_840 = x122 & n_346;
assign n_841 = x123 & n_346;
assign n_842 = x124 & n_346;
assign n_843 = x125 & n_346;
assign n_844 = x126 & n_346;
assign n_845 = x127 & n_346;
assign n_846 = n_348 ^ n_13;
assign n_847 = n_348 ^ n_14;
assign n_848 = n_351 ^ x10;
assign n_849 = x10 & ~n_351;
assign n_850 = n_350 ^ n_351;
assign n_851 = n_14 & n_352;
assign n_852 = n_16 ^ n_354;
assign n_853 = n_356 ^ n_16;
assign n_854 = n_357 ^ n_15;
assign n_855 = x67 & n_357;
assign n_856 = x68 & n_357;
assign n_857 = x69 & n_357;
assign n_858 = x70 & n_357;
assign n_859 = x71 & n_357;
assign n_860 = x72 & n_357;
assign n_861 = x73 & n_357;
assign n_862 = x74 & n_357;
assign n_863 = x75 & n_357;
assign n_864 = x76 & n_357;
assign n_865 = x77 & n_357;
assign n_866 = x78 & n_357;
assign n_867 = x79 & n_357;
assign n_868 = x80 & n_357;
assign n_869 = x81 & n_357;
assign n_870 = x82 & n_357;
assign n_871 = x83 & n_357;
assign n_872 = x84 & n_357;
assign n_873 = x85 & n_357;
assign n_874 = x86 & n_357;
assign n_875 = x87 & n_357;
assign n_876 = x88 & n_357;
assign n_877 = x89 & n_357;
assign n_878 = x90 & n_357;
assign n_879 = x91 & n_357;
assign n_880 = x92 & n_357;
assign n_881 = x93 & n_357;
assign n_882 = x94 & n_357;
assign n_883 = x95 & n_357;
assign n_884 = x96 & n_357;
assign n_885 = x97 & n_357;
assign n_886 = x98 & n_357;
assign n_887 = x99 & n_357;
assign n_888 = x100 & n_357;
assign n_889 = x101 & n_357;
assign n_890 = x102 & n_357;
assign n_891 = x103 & n_357;
assign n_892 = x104 & n_357;
assign n_893 = x105 & n_357;
assign n_894 = x106 & n_357;
assign n_895 = x107 & n_357;
assign n_896 = x108 & n_357;
assign n_897 = x109 & n_357;
assign n_898 = x110 & n_357;
assign n_899 = x111 & n_357;
assign n_900 = x112 & n_357;
assign n_901 = x113 & n_357;
assign n_902 = x114 & n_357;
assign n_903 = x115 & n_357;
assign n_904 = x116 & n_357;
assign n_905 = x117 & n_357;
assign n_906 = x118 & n_357;
assign n_907 = x119 & n_357;
assign n_908 = x120 & n_357;
assign n_909 = x121 & n_357;
assign n_910 = x122 & n_357;
assign n_911 = x123 & n_357;
assign n_912 = x124 & n_357;
assign n_913 = x125 & n_357;
assign n_914 = x126 & n_357;
assign n_915 = x127 & n_357;
assign n_916 = n_362 ^ x16;
assign n_917 = x16 & ~n_362;
assign n_918 = n_359 ^ n_362;
assign n_919 = n_361 ^ n_362;
assign n_920 = n_363 ^ n_18;
assign n_921 = x67 & n_363;
assign n_922 = x68 & n_363;
assign n_923 = x69 & n_363;
assign n_924 = x70 & n_363;
assign n_925 = x71 & n_363;
assign n_926 = x72 & n_363;
assign n_927 = x73 & n_363;
assign n_928 = x74 & n_363;
assign n_929 = x75 & n_363;
assign n_930 = x76 & n_363;
assign n_931 = x77 & n_363;
assign n_932 = x78 & n_363;
assign n_933 = x79 & n_363;
assign n_934 = x80 & n_363;
assign n_935 = x81 & n_363;
assign n_936 = x82 & n_363;
assign n_937 = x83 & n_363;
assign n_938 = x84 & n_363;
assign n_939 = x85 & n_363;
assign n_940 = x86 & n_363;
assign n_941 = x87 & n_363;
assign n_942 = x88 & n_363;
assign n_943 = x89 & n_363;
assign n_944 = x90 & n_363;
assign n_945 = x91 & n_363;
assign n_946 = x92 & n_363;
assign n_947 = x93 & n_363;
assign n_948 = x94 & n_363;
assign n_949 = x95 & n_363;
assign n_950 = x96 & n_363;
assign n_951 = x97 & n_363;
assign n_952 = x98 & n_363;
assign n_953 = x99 & n_363;
assign n_954 = x100 & n_363;
assign n_955 = x101 & n_363;
assign n_956 = x102 & n_363;
assign n_957 = x103 & n_363;
assign n_958 = x104 & n_363;
assign n_959 = x105 & n_363;
assign n_960 = x106 & n_363;
assign n_961 = x107 & n_363;
assign n_962 = x108 & n_363;
assign n_963 = x109 & n_363;
assign n_964 = x110 & n_363;
assign n_965 = x111 & n_363;
assign n_966 = x112 & n_363;
assign n_967 = x113 & n_363;
assign n_968 = x114 & n_363;
assign n_969 = x115 & n_363;
assign n_970 = x116 & n_363;
assign n_971 = x117 & n_363;
assign n_972 = x118 & n_363;
assign n_973 = x119 & n_363;
assign n_974 = x120 & n_363;
assign n_975 = x121 & n_363;
assign n_976 = x122 & n_363;
assign n_977 = x123 & n_363;
assign n_978 = x124 & n_363;
assign n_979 = x125 & n_363;
assign n_980 = x126 & n_363;
assign n_981 = x127 & n_363;
assign n_982 = n_368 ^ x19;
assign n_983 = x19 & ~n_368;
assign n_984 = n_365 ^ n_368;
assign n_985 = n_367 ^ n_368;
assign n_986 = n_369 ^ n_21;
assign n_987 = x67 & n_369;
assign n_988 = x68 & n_369;
assign n_989 = x69 & n_369;
assign n_990 = x70 & n_369;
assign n_991 = x71 & n_369;
assign n_992 = x72 & n_369;
assign n_993 = x73 & n_369;
assign n_994 = x74 & n_369;
assign n_995 = x75 & n_369;
assign n_996 = x76 & n_369;
assign n_997 = x77 & n_369;
assign n_998 = x78 & n_369;
assign n_999 = x79 & n_369;
assign n_1000 = x80 & n_369;
assign n_1001 = x81 & n_369;
assign n_1002 = x82 & n_369;
assign n_1003 = x83 & n_369;
assign n_1004 = x84 & n_369;
assign n_1005 = x85 & n_369;
assign n_1006 = x86 & n_369;
assign n_1007 = x87 & n_369;
assign n_1008 = x88 & n_369;
assign n_1009 = x89 & n_369;
assign n_1010 = x90 & n_369;
assign n_1011 = x91 & n_369;
assign n_1012 = x92 & n_369;
assign n_1013 = x93 & n_369;
assign n_1014 = x94 & n_369;
assign n_1015 = x95 & n_369;
assign n_1016 = x96 & n_369;
assign n_1017 = x97 & n_369;
assign n_1018 = x98 & n_369;
assign n_1019 = x99 & n_369;
assign n_1020 = x100 & n_369;
assign n_1021 = x101 & n_369;
assign n_1022 = x102 & n_369;
assign n_1023 = x103 & n_369;
assign n_1024 = x104 & n_369;
assign n_1025 = x105 & n_369;
assign n_1026 = x106 & n_369;
assign n_1027 = x107 & n_369;
assign n_1028 = x108 & n_369;
assign n_1029 = x109 & n_369;
assign n_1030 = x110 & n_369;
assign n_1031 = x111 & n_369;
assign n_1032 = x112 & n_369;
assign n_1033 = x113 & n_369;
assign n_1034 = x114 & n_369;
assign n_1035 = x115 & n_369;
assign n_1036 = x116 & n_369;
assign n_1037 = x117 & n_369;
assign n_1038 = x118 & n_369;
assign n_1039 = x119 & n_369;
assign n_1040 = x120 & n_369;
assign n_1041 = x121 & n_369;
assign n_1042 = x122 & n_369;
assign n_1043 = x123 & n_369;
assign n_1044 = x124 & n_369;
assign n_1045 = x125 & n_369;
assign n_1046 = x126 & n_369;
assign n_1047 = x127 & n_369;
assign n_1048 = n_374 ^ x22;
assign n_1049 = x22 & ~n_374;
assign n_1050 = n_371 ^ n_374;
assign n_1051 = n_373 ^ n_374;
assign n_1052 = n_375 ^ n_24;
assign n_1053 = x67 & n_375;
assign n_1054 = x68 & n_375;
assign n_1055 = x69 & n_375;
assign n_1056 = x70 & n_375;
assign n_1057 = x71 & n_375;
assign n_1058 = x72 & n_375;
assign n_1059 = x73 & n_375;
assign n_1060 = x74 & n_375;
assign n_1061 = x75 & n_375;
assign n_1062 = x76 & n_375;
assign n_1063 = x77 & n_375;
assign n_1064 = x78 & n_375;
assign n_1065 = x79 & n_375;
assign n_1066 = x80 & n_375;
assign n_1067 = x81 & n_375;
assign n_1068 = x82 & n_375;
assign n_1069 = x83 & n_375;
assign n_1070 = x84 & n_375;
assign n_1071 = x85 & n_375;
assign n_1072 = x86 & n_375;
assign n_1073 = x87 & n_375;
assign n_1074 = x88 & n_375;
assign n_1075 = x89 & n_375;
assign n_1076 = x90 & n_375;
assign n_1077 = x91 & n_375;
assign n_1078 = x92 & n_375;
assign n_1079 = x93 & n_375;
assign n_1080 = x94 & n_375;
assign n_1081 = x95 & n_375;
assign n_1082 = x96 & n_375;
assign n_1083 = x97 & n_375;
assign n_1084 = x98 & n_375;
assign n_1085 = x99 & n_375;
assign n_1086 = x100 & n_375;
assign n_1087 = x101 & n_375;
assign n_1088 = x102 & n_375;
assign n_1089 = x103 & n_375;
assign n_1090 = x104 & n_375;
assign n_1091 = x105 & n_375;
assign n_1092 = x106 & n_375;
assign n_1093 = x107 & n_375;
assign n_1094 = x108 & n_375;
assign n_1095 = x109 & n_375;
assign n_1096 = x110 & n_375;
assign n_1097 = x111 & n_375;
assign n_1098 = x112 & n_375;
assign n_1099 = x113 & n_375;
assign n_1100 = x114 & n_375;
assign n_1101 = x115 & n_375;
assign n_1102 = x116 & n_375;
assign n_1103 = x117 & n_375;
assign n_1104 = x118 & n_375;
assign n_1105 = x119 & n_375;
assign n_1106 = x120 & n_375;
assign n_1107 = x121 & n_375;
assign n_1108 = x122 & n_375;
assign n_1109 = x123 & n_375;
assign n_1110 = x124 & n_375;
assign n_1111 = x125 & n_375;
assign n_1112 = x126 & n_375;
assign n_1113 = x127 & n_375;
assign n_1114 = n_377 ^ n_28;
assign n_1115 = n_379 ^ n_28;
assign n_1116 = ~x64 & n_380;
assign n_1117 = n_381 ^ n_27;
assign n_1118 = x68 & n_381;
assign n_1119 = x69 & n_381;
assign n_1120 = x70 & n_381;
assign n_1121 = x71 & n_381;
assign n_1122 = x72 & n_381;
assign n_1123 = x73 & n_381;
assign n_1124 = x74 & n_381;
assign n_1125 = x75 & n_381;
assign n_1126 = x76 & n_381;
assign n_1127 = x77 & n_381;
assign n_1128 = x78 & n_381;
assign n_1129 = x79 & n_381;
assign n_1130 = x80 & n_381;
assign n_1131 = x81 & n_381;
assign n_1132 = x82 & n_381;
assign n_1133 = x83 & n_381;
assign n_1134 = x84 & n_381;
assign n_1135 = x85 & n_381;
assign n_1136 = x86 & n_381;
assign n_1137 = x87 & n_381;
assign n_1138 = x88 & n_381;
assign n_1139 = x89 & n_381;
assign n_1140 = x90 & n_381;
assign n_1141 = x91 & n_381;
assign n_1142 = x92 & n_381;
assign n_1143 = x93 & n_381;
assign n_1144 = x94 & n_381;
assign n_1145 = x95 & n_381;
assign n_1146 = x96 & n_381;
assign n_1147 = x97 & n_381;
assign n_1148 = x98 & n_381;
assign n_1149 = x99 & n_381;
assign n_1150 = x100 & n_381;
assign n_1151 = x101 & n_381;
assign n_1152 = x102 & n_381;
assign n_1153 = x103 & n_381;
assign n_1154 = x104 & n_381;
assign n_1155 = x105 & n_381;
assign n_1156 = x106 & n_381;
assign n_1157 = x107 & n_381;
assign n_1158 = x108 & n_381;
assign n_1159 = x109 & n_381;
assign n_1160 = x110 & n_381;
assign n_1161 = x111 & n_381;
assign n_1162 = x112 & n_381;
assign n_1163 = x113 & n_381;
assign n_1164 = x114 & n_381;
assign n_1165 = x115 & n_381;
assign n_1166 = x116 & n_381;
assign n_1167 = x117 & n_381;
assign n_1168 = x118 & n_381;
assign n_1169 = x119 & n_381;
assign n_1170 = x120 & n_381;
assign n_1171 = x121 & n_381;
assign n_1172 = x122 & n_381;
assign n_1173 = x123 & n_381;
assign n_1174 = x124 & n_381;
assign n_1175 = x125 & n_381;
assign n_1176 = x126 & n_381;
assign n_1177 = x127 & n_381;
assign n_1178 = n_383 ^ n_31;
assign n_1179 = n_385 ^ n_31;
assign n_1180 = ~x64 & n_386;
assign n_1181 = n_387 ^ n_30;
assign n_1182 = x67 & n_387;
assign n_1183 = x68 & n_387;
assign n_1184 = x69 & n_387;
assign n_1185 = x70 & n_387;
assign n_1186 = x71 & n_387;
assign n_1187 = x72 & n_387;
assign n_1188 = x73 & n_387;
assign n_1189 = x74 & n_387;
assign n_1190 = x75 & n_387;
assign n_1191 = x76 & n_387;
assign n_1192 = x77 & n_387;
assign n_1193 = x78 & n_387;
assign n_1194 = x79 & n_387;
assign n_1195 = x80 & n_387;
assign n_1196 = x81 & n_387;
assign n_1197 = x82 & n_387;
assign n_1198 = x83 & n_387;
assign n_1199 = x84 & n_387;
assign n_1200 = x85 & n_387;
assign n_1201 = x86 & n_387;
assign n_1202 = x87 & n_387;
assign n_1203 = x88 & n_387;
assign n_1204 = x89 & n_387;
assign n_1205 = x90 & n_387;
assign n_1206 = x91 & n_387;
assign n_1207 = x92 & n_387;
assign n_1208 = x93 & n_387;
assign n_1209 = x94 & n_387;
assign n_1210 = x95 & n_387;
assign n_1211 = x96 & n_387;
assign n_1212 = x97 & n_387;
assign n_1213 = x98 & n_387;
assign n_1214 = x99 & n_387;
assign n_1215 = x100 & n_387;
assign n_1216 = x101 & n_387;
assign n_1217 = x102 & n_387;
assign n_1218 = x103 & n_387;
assign n_1219 = x104 & n_387;
assign n_1220 = x105 & n_387;
assign n_1221 = x106 & n_387;
assign n_1222 = x107 & n_387;
assign n_1223 = x108 & n_387;
assign n_1224 = x109 & n_387;
assign n_1225 = x110 & n_387;
assign n_1226 = x111 & n_387;
assign n_1227 = x112 & n_387;
assign n_1228 = x113 & n_387;
assign n_1229 = x114 & n_387;
assign n_1230 = x115 & n_387;
assign n_1231 = x116 & n_387;
assign n_1232 = x117 & n_387;
assign n_1233 = x118 & n_387;
assign n_1234 = x119 & n_387;
assign n_1235 = x120 & n_387;
assign n_1236 = x121 & n_387;
assign n_1237 = x122 & n_387;
assign n_1238 = x123 & n_387;
assign n_1239 = x124 & n_387;
assign n_1240 = x125 & n_387;
assign n_1241 = x126 & n_387;
assign n_1242 = x127 & n_387;
assign n_1243 = n_392 ^ x31;
assign n_1244 = x31 & ~n_392;
assign n_1245 = n_389 ^ n_392;
assign n_1246 = n_391 ^ n_392;
assign n_1247 = n_35 & n_393;
assign n_1248 = n_394 ^ n_33;
assign n_1249 = x67 & n_394;
assign n_1250 = x68 & n_394;
assign n_1251 = x69 & n_394;
assign n_1252 = x70 & n_394;
assign n_1253 = x71 & n_394;
assign n_1254 = x72 & n_394;
assign n_1255 = x73 & n_394;
assign n_1256 = x74 & n_394;
assign n_1257 = x75 & n_394;
assign n_1258 = x76 & n_394;
assign n_1259 = x77 & n_394;
assign n_1260 = x78 & n_394;
assign n_1261 = x79 & n_394;
assign n_1262 = x80 & n_394;
assign n_1263 = x81 & n_394;
assign n_1264 = x82 & n_394;
assign n_1265 = x83 & n_394;
assign n_1266 = x84 & n_394;
assign n_1267 = x85 & n_394;
assign n_1268 = x86 & n_394;
assign n_1269 = x87 & n_394;
assign n_1270 = x88 & n_394;
assign n_1271 = x89 & n_394;
assign n_1272 = x90 & n_394;
assign n_1273 = x91 & n_394;
assign n_1274 = x92 & n_394;
assign n_1275 = x93 & n_394;
assign n_1276 = x94 & n_394;
assign n_1277 = x95 & n_394;
assign n_1278 = x96 & n_394;
assign n_1279 = x97 & n_394;
assign n_1280 = x98 & n_394;
assign n_1281 = x99 & n_394;
assign n_1282 = x100 & n_394;
assign n_1283 = x101 & n_394;
assign n_1284 = x102 & n_394;
assign n_1285 = x103 & n_394;
assign n_1286 = x104 & n_394;
assign n_1287 = x105 & n_394;
assign n_1288 = x106 & n_394;
assign n_1289 = x107 & n_394;
assign n_1290 = x108 & n_394;
assign n_1291 = x109 & n_394;
assign n_1292 = x110 & n_394;
assign n_1293 = x111 & n_394;
assign n_1294 = x112 & n_394;
assign n_1295 = x113 & n_394;
assign n_1296 = x114 & n_394;
assign n_1297 = x115 & n_394;
assign n_1298 = x116 & n_394;
assign n_1299 = x117 & n_394;
assign n_1300 = x118 & n_394;
assign n_1301 = x119 & n_394;
assign n_1302 = x120 & n_394;
assign n_1303 = x121 & n_394;
assign n_1304 = x122 & n_394;
assign n_1305 = x123 & n_394;
assign n_1306 = x124 & n_394;
assign n_1307 = x125 & n_394;
assign n_1308 = x126 & n_394;
assign n_1309 = x127 & n_394;
assign n_1310 = n_399 ^ x34;
assign n_1311 = x34 & ~n_399;
assign n_1312 = n_396 ^ n_399;
assign n_1313 = n_398 ^ n_399;
assign n_1314 = n_400 ^ n_36;
assign n_1315 = x67 & n_400;
assign n_1316 = x68 & n_400;
assign n_1317 = x69 & n_400;
assign n_1318 = x70 & n_400;
assign n_1319 = x71 & n_400;
assign n_1320 = x72 & n_400;
assign n_1321 = x73 & n_400;
assign n_1322 = x74 & n_400;
assign n_1323 = x75 & n_400;
assign n_1324 = x76 & n_400;
assign n_1325 = x77 & n_400;
assign n_1326 = x78 & n_400;
assign n_1327 = x79 & n_400;
assign n_1328 = x80 & n_400;
assign n_1329 = x81 & n_400;
assign n_1330 = x82 & n_400;
assign n_1331 = x83 & n_400;
assign n_1332 = x84 & n_400;
assign n_1333 = x85 & n_400;
assign n_1334 = x86 & n_400;
assign n_1335 = x87 & n_400;
assign n_1336 = x88 & n_400;
assign n_1337 = x89 & n_400;
assign n_1338 = x90 & n_400;
assign n_1339 = x91 & n_400;
assign n_1340 = x92 & n_400;
assign n_1341 = x93 & n_400;
assign n_1342 = x94 & n_400;
assign n_1343 = x95 & n_400;
assign n_1344 = x96 & n_400;
assign n_1345 = x97 & n_400;
assign n_1346 = x98 & n_400;
assign n_1347 = x99 & n_400;
assign n_1348 = x100 & n_400;
assign n_1349 = x101 & n_400;
assign n_1350 = x102 & n_400;
assign n_1351 = x103 & n_400;
assign n_1352 = x104 & n_400;
assign n_1353 = x105 & n_400;
assign n_1354 = x106 & n_400;
assign n_1355 = x107 & n_400;
assign n_1356 = x108 & n_400;
assign n_1357 = x109 & n_400;
assign n_1358 = x110 & n_400;
assign n_1359 = x111 & n_400;
assign n_1360 = x112 & n_400;
assign n_1361 = x113 & n_400;
assign n_1362 = x114 & n_400;
assign n_1363 = x115 & n_400;
assign n_1364 = x116 & n_400;
assign n_1365 = x117 & n_400;
assign n_1366 = x118 & n_400;
assign n_1367 = x119 & n_400;
assign n_1368 = x120 & n_400;
assign n_1369 = x121 & n_400;
assign n_1370 = x122 & n_400;
assign n_1371 = x123 & n_400;
assign n_1372 = x124 & n_400;
assign n_1373 = x125 & n_400;
assign n_1374 = x126 & n_400;
assign n_1375 = x127 & n_400;
assign n_1376 = n_405 ^ x37;
assign n_1377 = x37 & ~n_405;
assign n_1378 = n_402 ^ n_405;
assign n_1379 = n_404 ^ n_405;
assign n_1380 = n_406 ^ n_39;
assign n_1381 = x67 & n_406;
assign n_1382 = x68 & n_406;
assign n_1383 = x69 & n_406;
assign n_1384 = x70 & n_406;
assign n_1385 = x71 & n_406;
assign n_1386 = x72 & n_406;
assign n_1387 = x73 & n_406;
assign n_1388 = x74 & n_406;
assign n_1389 = x75 & n_406;
assign n_1390 = x76 & n_406;
assign n_1391 = x77 & n_406;
assign n_1392 = x78 & n_406;
assign n_1393 = x79 & n_406;
assign n_1394 = x80 & n_406;
assign n_1395 = x81 & n_406;
assign n_1396 = x82 & n_406;
assign n_1397 = x83 & n_406;
assign n_1398 = x84 & n_406;
assign n_1399 = x85 & n_406;
assign n_1400 = x86 & n_406;
assign n_1401 = x87 & n_406;
assign n_1402 = x88 & n_406;
assign n_1403 = x89 & n_406;
assign n_1404 = x90 & n_406;
assign n_1405 = x91 & n_406;
assign n_1406 = x92 & n_406;
assign n_1407 = x93 & n_406;
assign n_1408 = x94 & n_406;
assign n_1409 = x95 & n_406;
assign n_1410 = x96 & n_406;
assign n_1411 = x97 & n_406;
assign n_1412 = x98 & n_406;
assign n_1413 = x99 & n_406;
assign n_1414 = x100 & n_406;
assign n_1415 = x101 & n_406;
assign n_1416 = x102 & n_406;
assign n_1417 = x103 & n_406;
assign n_1418 = x104 & n_406;
assign n_1419 = x105 & n_406;
assign n_1420 = x106 & n_406;
assign n_1421 = x107 & n_406;
assign n_1422 = x108 & n_406;
assign n_1423 = x109 & n_406;
assign n_1424 = x110 & n_406;
assign n_1425 = x111 & n_406;
assign n_1426 = x112 & n_406;
assign n_1427 = x113 & n_406;
assign n_1428 = x114 & n_406;
assign n_1429 = x115 & n_406;
assign n_1430 = x116 & n_406;
assign n_1431 = x117 & n_406;
assign n_1432 = x118 & n_406;
assign n_1433 = x119 & n_406;
assign n_1434 = x120 & n_406;
assign n_1435 = x121 & n_406;
assign n_1436 = x122 & n_406;
assign n_1437 = x123 & n_406;
assign n_1438 = x124 & n_406;
assign n_1439 = x125 & n_406;
assign n_1440 = x126 & n_406;
assign n_1441 = x127 & n_406;
assign n_1442 = ~x64 & ~n_411;
assign n_1443 = n_408 ^ n_412;
assign n_1444 = n_412 ^ n_410;
assign n_1445 = n_413 ^ n_42;
assign n_1446 = x68 & n_413;
assign n_1447 = x69 & n_413;
assign n_1448 = x70 & n_413;
assign n_1449 = x71 & n_413;
assign n_1450 = x72 & n_413;
assign n_1451 = x73 & n_413;
assign n_1452 = x74 & n_413;
assign n_1453 = x75 & n_413;
assign n_1454 = x76 & n_413;
assign n_1455 = x77 & n_413;
assign n_1456 = x78 & n_413;
assign n_1457 = x79 & n_413;
assign n_1458 = x80 & n_413;
assign n_1459 = x81 & n_413;
assign n_1460 = x82 & n_413;
assign n_1461 = x83 & n_413;
assign n_1462 = x84 & n_413;
assign n_1463 = x85 & n_413;
assign n_1464 = x86 & n_413;
assign n_1465 = x87 & n_413;
assign n_1466 = x88 & n_413;
assign n_1467 = x89 & n_413;
assign n_1468 = x90 & n_413;
assign n_1469 = x91 & n_413;
assign n_1470 = x92 & n_413;
assign n_1471 = x93 & n_413;
assign n_1472 = x94 & n_413;
assign n_1473 = x95 & n_413;
assign n_1474 = x96 & n_413;
assign n_1475 = x97 & n_413;
assign n_1476 = x98 & n_413;
assign n_1477 = x99 & n_413;
assign n_1478 = x100 & n_413;
assign n_1479 = x101 & n_413;
assign n_1480 = x102 & n_413;
assign n_1481 = x103 & n_413;
assign n_1482 = x104 & n_413;
assign n_1483 = x105 & n_413;
assign n_1484 = x106 & n_413;
assign n_1485 = x107 & n_413;
assign n_1486 = x108 & n_413;
assign n_1487 = x109 & n_413;
assign n_1488 = x110 & n_413;
assign n_1489 = x111 & n_413;
assign n_1490 = x112 & n_413;
assign n_1491 = x113 & n_413;
assign n_1492 = x114 & n_413;
assign n_1493 = x115 & n_413;
assign n_1494 = x116 & n_413;
assign n_1495 = x117 & n_413;
assign n_1496 = x118 & n_413;
assign n_1497 = x119 & n_413;
assign n_1498 = x120 & n_413;
assign n_1499 = x121 & n_413;
assign n_1500 = x122 & n_413;
assign n_1501 = x123 & n_413;
assign n_1502 = x124 & n_413;
assign n_1503 = x125 & n_413;
assign n_1504 = x126 & n_413;
assign n_1505 = x127 & n_413;
assign n_1506 = n_418 ^ x43;
assign n_1507 = x43 & ~n_418;
assign n_1508 = n_415 ^ n_418;
assign n_1509 = n_417 ^ n_418;
assign n_1510 = n_419 ^ n_45;
assign n_1511 = x67 & n_419;
assign n_1512 = x68 & n_419;
assign n_1513 = x69 & n_419;
assign n_1514 = x70 & n_419;
assign n_1515 = x71 & n_419;
assign n_1516 = x72 & n_419;
assign n_1517 = x73 & n_419;
assign n_1518 = x74 & n_419;
assign n_1519 = x75 & n_419;
assign n_1520 = x76 & n_419;
assign n_1521 = x77 & n_419;
assign n_1522 = x78 & n_419;
assign n_1523 = x79 & n_419;
assign n_1524 = x80 & n_419;
assign n_1525 = x81 & n_419;
assign n_1526 = x82 & n_419;
assign n_1527 = x83 & n_419;
assign n_1528 = x84 & n_419;
assign n_1529 = x85 & n_419;
assign n_1530 = x86 & n_419;
assign n_1531 = x87 & n_419;
assign n_1532 = x88 & n_419;
assign n_1533 = x89 & n_419;
assign n_1534 = x90 & n_419;
assign n_1535 = x91 & n_419;
assign n_1536 = x92 & n_419;
assign n_1537 = x93 & n_419;
assign n_1538 = x94 & n_419;
assign n_1539 = x95 & n_419;
assign n_1540 = x96 & n_419;
assign n_1541 = x97 & n_419;
assign n_1542 = x98 & n_419;
assign n_1543 = x99 & n_419;
assign n_1544 = x100 & n_419;
assign n_1545 = x101 & n_419;
assign n_1546 = x102 & n_419;
assign n_1547 = x103 & n_419;
assign n_1548 = x104 & n_419;
assign n_1549 = x105 & n_419;
assign n_1550 = x106 & n_419;
assign n_1551 = x107 & n_419;
assign n_1552 = x108 & n_419;
assign n_1553 = x109 & n_419;
assign n_1554 = x110 & n_419;
assign n_1555 = x111 & n_419;
assign n_1556 = x112 & n_419;
assign n_1557 = x113 & n_419;
assign n_1558 = x114 & n_419;
assign n_1559 = x115 & n_419;
assign n_1560 = x116 & n_419;
assign n_1561 = x117 & n_419;
assign n_1562 = x118 & n_419;
assign n_1563 = x119 & n_419;
assign n_1564 = x120 & n_419;
assign n_1565 = x121 & n_419;
assign n_1566 = x122 & n_419;
assign n_1567 = x123 & n_419;
assign n_1568 = x124 & n_419;
assign n_1569 = x125 & n_419;
assign n_1570 = x126 & n_419;
assign n_1571 = x127 & n_419;
assign n_1572 = n_424 ^ x46;
assign n_1573 = n_421 ^ n_424;
assign n_1574 = n_422 ^ n_424;
assign n_1575 = x46 & ~n_424;
assign n_1576 = n_425 ^ n_48;
assign n_1577 = x68 & n_425;
assign n_1578 = x69 & n_425;
assign n_1579 = x70 & n_425;
assign n_1580 = x71 & n_425;
assign n_1581 = x72 & n_425;
assign n_1582 = x73 & n_425;
assign n_1583 = x74 & n_425;
assign n_1584 = x75 & n_425;
assign n_1585 = x76 & n_425;
assign n_1586 = x77 & n_425;
assign n_1587 = x78 & n_425;
assign n_1588 = x79 & n_425;
assign n_1589 = x80 & n_425;
assign n_1590 = x81 & n_425;
assign n_1591 = x82 & n_425;
assign n_1592 = x83 & n_425;
assign n_1593 = x84 & n_425;
assign n_1594 = x85 & n_425;
assign n_1595 = x86 & n_425;
assign n_1596 = x87 & n_425;
assign n_1597 = x88 & n_425;
assign n_1598 = x89 & n_425;
assign n_1599 = x90 & n_425;
assign n_1600 = x91 & n_425;
assign n_1601 = x92 & n_425;
assign n_1602 = x93 & n_425;
assign n_1603 = x94 & n_425;
assign n_1604 = x95 & n_425;
assign n_1605 = x96 & n_425;
assign n_1606 = x97 & n_425;
assign n_1607 = x98 & n_425;
assign n_1608 = x99 & n_425;
assign n_1609 = x100 & n_425;
assign n_1610 = x101 & n_425;
assign n_1611 = x102 & n_425;
assign n_1612 = x103 & n_425;
assign n_1613 = x104 & n_425;
assign n_1614 = x105 & n_425;
assign n_1615 = x106 & n_425;
assign n_1616 = x107 & n_425;
assign n_1617 = x108 & n_425;
assign n_1618 = x109 & n_425;
assign n_1619 = x110 & n_425;
assign n_1620 = x111 & n_425;
assign n_1621 = x112 & n_425;
assign n_1622 = x113 & n_425;
assign n_1623 = x114 & n_425;
assign n_1624 = x115 & n_425;
assign n_1625 = x116 & n_425;
assign n_1626 = x117 & n_425;
assign n_1627 = x118 & n_425;
assign n_1628 = x119 & n_425;
assign n_1629 = x120 & n_425;
assign n_1630 = x121 & n_425;
assign n_1631 = x122 & n_425;
assign n_1632 = x123 & n_425;
assign n_1633 = x124 & n_425;
assign n_1634 = x125 & n_425;
assign n_1635 = x126 & n_425;
assign n_1636 = x127 & n_425;
assign n_1637 = n_430 ^ x49;
assign n_1638 = x49 & ~n_430;
assign n_1639 = n_427 ^ n_430;
assign n_1640 = n_429 ^ n_430;
assign n_1641 = n_431 ^ n_51;
assign n_1642 = x67 & n_431;
assign n_1643 = x68 & n_431;
assign n_1644 = x69 & n_431;
assign n_1645 = x70 & n_431;
assign n_1646 = x71 & n_431;
assign n_1647 = x72 & n_431;
assign n_1648 = x73 & n_431;
assign n_1649 = x74 & n_431;
assign n_1650 = x75 & n_431;
assign n_1651 = x76 & n_431;
assign n_1652 = x77 & n_431;
assign n_1653 = x78 & n_431;
assign n_1654 = x79 & n_431;
assign n_1655 = x80 & n_431;
assign n_1656 = x81 & n_431;
assign n_1657 = x82 & n_431;
assign n_1658 = x83 & n_431;
assign n_1659 = x84 & n_431;
assign n_1660 = x85 & n_431;
assign n_1661 = x86 & n_431;
assign n_1662 = x87 & n_431;
assign n_1663 = x88 & n_431;
assign n_1664 = x89 & n_431;
assign n_1665 = x90 & n_431;
assign n_1666 = x91 & n_431;
assign n_1667 = x92 & n_431;
assign n_1668 = x93 & n_431;
assign n_1669 = x94 & n_431;
assign n_1670 = x95 & n_431;
assign n_1671 = x96 & n_431;
assign n_1672 = x97 & n_431;
assign n_1673 = x98 & n_431;
assign n_1674 = x99 & n_431;
assign n_1675 = x100 & n_431;
assign n_1676 = x101 & n_431;
assign n_1677 = x102 & n_431;
assign n_1678 = x103 & n_431;
assign n_1679 = x104 & n_431;
assign n_1680 = x105 & n_431;
assign n_1681 = x106 & n_431;
assign n_1682 = x107 & n_431;
assign n_1683 = x108 & n_431;
assign n_1684 = x109 & n_431;
assign n_1685 = x110 & n_431;
assign n_1686 = x111 & n_431;
assign n_1687 = x112 & n_431;
assign n_1688 = x113 & n_431;
assign n_1689 = x114 & n_431;
assign n_1690 = x115 & n_431;
assign n_1691 = x116 & n_431;
assign n_1692 = x117 & n_431;
assign n_1693 = x118 & n_431;
assign n_1694 = x119 & n_431;
assign n_1695 = x120 & n_431;
assign n_1696 = x121 & n_431;
assign n_1697 = x122 & n_431;
assign n_1698 = x123 & n_431;
assign n_1699 = x124 & n_431;
assign n_1700 = x125 & n_431;
assign n_1701 = x126 & n_431;
assign n_1702 = x127 & n_431;
assign n_1703 = n_436 ^ x52;
assign n_1704 = n_433 ^ n_436;
assign n_1705 = n_434 ^ n_436;
assign n_1706 = n_437 ^ n_54;
assign n_1707 = x67 & n_437;
assign n_1708 = x68 & n_437;
assign n_1709 = x69 & n_437;
assign n_1710 = x70 & n_437;
assign n_1711 = x71 & n_437;
assign n_1712 = x72 & n_437;
assign n_1713 = x73 & n_437;
assign n_1714 = x74 & n_437;
assign n_1715 = x75 & n_437;
assign n_1716 = x76 & n_437;
assign n_1717 = x77 & n_437;
assign n_1718 = x78 & n_437;
assign n_1719 = x79 & n_437;
assign n_1720 = x80 & n_437;
assign n_1721 = x81 & n_437;
assign n_1722 = x82 & n_437;
assign n_1723 = x83 & n_437;
assign n_1724 = x84 & n_437;
assign n_1725 = x85 & n_437;
assign n_1726 = x86 & n_437;
assign n_1727 = x87 & n_437;
assign n_1728 = x88 & n_437;
assign n_1729 = x89 & n_437;
assign n_1730 = x90 & n_437;
assign n_1731 = x91 & n_437;
assign n_1732 = x92 & n_437;
assign n_1733 = x93 & n_437;
assign n_1734 = x94 & n_437;
assign n_1735 = x95 & n_437;
assign n_1736 = x96 & n_437;
assign n_1737 = x97 & n_437;
assign n_1738 = x98 & n_437;
assign n_1739 = x99 & n_437;
assign n_1740 = x100 & n_437;
assign n_1741 = x101 & n_437;
assign n_1742 = x102 & n_437;
assign n_1743 = x103 & n_437;
assign n_1744 = x104 & n_437;
assign n_1745 = x105 & n_437;
assign n_1746 = x106 & n_437;
assign n_1747 = x107 & n_437;
assign n_1748 = x108 & n_437;
assign n_1749 = x109 & n_437;
assign n_1750 = x110 & n_437;
assign n_1751 = x111 & n_437;
assign n_1752 = x112 & n_437;
assign n_1753 = x113 & n_437;
assign n_1754 = x114 & n_437;
assign n_1755 = x115 & n_437;
assign n_1756 = x116 & n_437;
assign n_1757 = x117 & n_437;
assign n_1758 = x118 & n_437;
assign n_1759 = x119 & n_437;
assign n_1760 = x120 & n_437;
assign n_1761 = x121 & n_437;
assign n_1762 = x122 & n_437;
assign n_1763 = x123 & n_437;
assign n_1764 = x124 & n_437;
assign n_1765 = x125 & n_437;
assign n_1766 = x126 & n_437;
assign n_1767 = x127 & n_437;
assign n_1768 = n_439 ^ n_58;
assign n_1769 = n_441 ^ n_58;
assign n_1770 = ~x64 & n_442;
assign n_1771 = n_443 ^ n_57;
assign n_1772 = x68 & n_443;
assign n_1773 = x69 & n_443;
assign n_1774 = x70 & n_443;
assign n_1775 = x71 & n_443;
assign n_1776 = x72 & n_443;
assign n_1777 = x73 & n_443;
assign n_1778 = x74 & n_443;
assign n_1779 = x75 & n_443;
assign n_1780 = x76 & n_443;
assign n_1781 = x77 & n_443;
assign n_1782 = x78 & n_443;
assign n_1783 = x79 & n_443;
assign n_1784 = x80 & n_443;
assign n_1785 = x81 & n_443;
assign n_1786 = x82 & n_443;
assign n_1787 = x83 & n_443;
assign n_1788 = x84 & n_443;
assign n_1789 = x85 & n_443;
assign n_1790 = x86 & n_443;
assign n_1791 = x87 & n_443;
assign n_1792 = x88 & n_443;
assign n_1793 = x89 & n_443;
assign n_1794 = x90 & n_443;
assign n_1795 = x91 & n_443;
assign n_1796 = x92 & n_443;
assign n_1797 = x93 & n_443;
assign n_1798 = x94 & n_443;
assign n_1799 = x95 & n_443;
assign n_1800 = x96 & n_443;
assign n_1801 = x97 & n_443;
assign n_1802 = x98 & n_443;
assign n_1803 = x99 & n_443;
assign n_1804 = x100 & n_443;
assign n_1805 = x101 & n_443;
assign n_1806 = x102 & n_443;
assign n_1807 = x103 & n_443;
assign n_1808 = x104 & n_443;
assign n_1809 = x105 & n_443;
assign n_1810 = x106 & n_443;
assign n_1811 = x107 & n_443;
assign n_1812 = x108 & n_443;
assign n_1813 = x109 & n_443;
assign n_1814 = x110 & n_443;
assign n_1815 = x111 & n_443;
assign n_1816 = x112 & n_443;
assign n_1817 = x113 & n_443;
assign n_1818 = x114 & n_443;
assign n_1819 = x115 & n_443;
assign n_1820 = x116 & n_443;
assign n_1821 = x117 & n_443;
assign n_1822 = x118 & n_443;
assign n_1823 = x119 & n_443;
assign n_1824 = x120 & n_443;
assign n_1825 = x121 & n_443;
assign n_1826 = x122 & n_443;
assign n_1827 = x123 & n_443;
assign n_1828 = x124 & n_443;
assign n_1829 = x125 & n_443;
assign n_1830 = x126 & n_443;
assign n_1831 = x127 & n_443;
assign n_1832 = n_445 ^ n_61;
assign n_1833 = n_447 ^ n_61;
assign n_1834 = ~x64 & n_448;
assign n_1835 = n_449 ^ n_60;
assign n_1836 = x68 & n_449;
assign n_1837 = x69 & n_449;
assign n_1838 = x70 & n_449;
assign n_1839 = x71 & n_449;
assign n_1840 = x72 & n_449;
assign n_1841 = x73 & n_449;
assign n_1842 = x74 & n_449;
assign n_1843 = x75 & n_449;
assign n_1844 = x76 & n_449;
assign n_1845 = x77 & n_449;
assign n_1846 = x78 & n_449;
assign n_1847 = x79 & n_449;
assign n_1848 = x80 & n_449;
assign n_1849 = x81 & n_449;
assign n_1850 = x82 & n_449;
assign n_1851 = x83 & n_449;
assign n_1852 = x84 & n_449;
assign n_1853 = x85 & n_449;
assign n_1854 = x86 & n_449;
assign n_1855 = x87 & n_449;
assign n_1856 = x88 & n_449;
assign n_1857 = x89 & n_449;
assign n_1858 = x90 & n_449;
assign n_1859 = x91 & n_449;
assign n_1860 = x92 & n_449;
assign n_1861 = x93 & n_449;
assign n_1862 = x94 & n_449;
assign n_1863 = x95 & n_449;
assign n_1864 = x96 & n_449;
assign n_1865 = x97 & n_449;
assign n_1866 = x98 & n_449;
assign n_1867 = x99 & n_449;
assign n_1868 = x100 & n_449;
assign n_1869 = x101 & n_449;
assign n_1870 = x102 & n_449;
assign n_1871 = x103 & n_449;
assign n_1872 = x104 & n_449;
assign n_1873 = x105 & n_449;
assign n_1874 = x106 & n_449;
assign n_1875 = x107 & n_449;
assign n_1876 = x108 & n_449;
assign n_1877 = x109 & n_449;
assign n_1878 = x110 & n_449;
assign n_1879 = x111 & n_449;
assign n_1880 = x112 & n_449;
assign n_1881 = x113 & n_449;
assign n_1882 = x114 & n_449;
assign n_1883 = x115 & n_449;
assign n_1884 = x116 & n_449;
assign n_1885 = x117 & n_449;
assign n_1886 = x118 & n_449;
assign n_1887 = x119 & n_449;
assign n_1888 = x120 & n_449;
assign n_1889 = x121 & n_449;
assign n_1890 = x122 & n_449;
assign n_1891 = x123 & n_449;
assign n_1892 = x124 & n_449;
assign n_1893 = x125 & n_449;
assign n_1894 = x126 & n_449;
assign n_1895 = x127 & n_449;
assign n_1896 = n_451 ^ n_64;
assign n_1897 = n_453 ^ n_64;
assign n_1898 = ~x64 & n_454;
assign n_1899 = n_455 ^ n_63;
assign n_1900 = x68 & n_455;
assign n_1901 = x69 & n_455;
assign n_1902 = x70 & n_455;
assign n_1903 = x71 & n_455;
assign n_1904 = x72 & n_455;
assign n_1905 = x73 & n_455;
assign n_1906 = x74 & n_455;
assign n_1907 = x75 & n_455;
assign n_1908 = x76 & n_455;
assign n_1909 = x77 & n_455;
assign n_1910 = x78 & n_455;
assign n_1911 = x79 & n_455;
assign n_1912 = x80 & n_455;
assign n_1913 = x81 & n_455;
assign n_1914 = x82 & n_455;
assign n_1915 = x83 & n_455;
assign n_1916 = x84 & n_455;
assign n_1917 = x85 & n_455;
assign n_1918 = x86 & n_455;
assign n_1919 = x87 & n_455;
assign n_1920 = x88 & n_455;
assign n_1921 = x89 & n_455;
assign n_1922 = x90 & n_455;
assign n_1923 = x91 & n_455;
assign n_1924 = x92 & n_455;
assign n_1925 = x93 & n_455;
assign n_1926 = x94 & n_455;
assign n_1927 = x95 & n_455;
assign n_1928 = x96 & n_455;
assign n_1929 = x97 & n_455;
assign n_1930 = x98 & n_455;
assign n_1931 = x99 & n_455;
assign n_1932 = x100 & n_455;
assign n_1933 = x101 & n_455;
assign n_1934 = x102 & n_455;
assign n_1935 = x103 & n_455;
assign n_1936 = x104 & n_455;
assign n_1937 = x105 & n_455;
assign n_1938 = x106 & n_455;
assign n_1939 = x107 & n_455;
assign n_1940 = x108 & n_455;
assign n_1941 = x109 & n_455;
assign n_1942 = x110 & n_455;
assign n_1943 = x111 & n_455;
assign n_1944 = x112 & n_455;
assign n_1945 = x113 & n_455;
assign n_1946 = x114 & n_455;
assign n_1947 = x115 & n_455;
assign n_1948 = x116 & n_455;
assign n_1949 = x117 & n_455;
assign n_1950 = x118 & n_455;
assign n_1951 = x119 & n_455;
assign n_1952 = x120 & n_455;
assign n_1953 = x121 & n_455;
assign n_1954 = x122 & n_455;
assign n_1955 = x123 & n_455;
assign n_1956 = x124 & n_455;
assign n_1957 = x125 & n_455;
assign n_1958 = x126 & n_455;
assign n_1959 = x127 & n_455;
assign n_1960 = ~x75 & n_460;
assign n_1961 = x70 & n_487;
assign n_1962 = ~n_487 & n_127;
assign n_1963 = x73 & n_487;
assign n_1964 = n_487 & n_156;
assign n_1965 = x82 & n_487;
assign n_1966 = n_487 & n_167;
assign n_1967 = x85 & n_487;
assign n_1968 = n_487 & n_178;
assign n_1969 = x88 & n_487;
assign n_1970 = ~n_487 & n_187;
assign n_1971 = n_487 & n_201;
assign n_1972 = x94 & n_487;
assign n_1973 = ~n_487 & n_213;
assign n_1974 = x97 & n_487;
assign n_1975 = ~n_487 & n_223;
assign n_1976 = x100 & n_487;
assign n_1977 = x109 & n_487;
assign n_1978 = ~n_487 & n_259;
assign n_1979 = x115 & n_487;
assign n_1980 = ~n_487 & n_274;
assign n_1981 = x121 & n_487;
assign n_1982 = ~n_487 & n_291;
assign n_1983 = x124 & n_487;
assign n_1984 = n_293 & n_487;
assign n_1985 = n_488 ^ x70;
assign n_1986 = n_488 ^ x82;
assign n_1987 = n_488 ^ x88;
assign n_1988 = n_488 ^ x94;
assign n_1989 = n_488 ^ x97;
assign n_1990 = n_488 ^ x109;
assign n_1991 = n_488 ^ x115;
assign n_1992 = n_488 ^ x121;
assign n_1993 = n_491 ^ n_343;
assign n_1994 = x29 & ~n_496;
assign n_1995 = ~n_66 & n_499;
assign y1 = n_500;
assign n_1996 = n_502 ^ x65;
assign n_1997 = ~n_502 & n_15;
assign n_1998 = n_504 ^ x2;
assign n_1999 = n_505 ^ x8;
assign n_2000 = n_506 ^ x11;
assign n_2001 = n_507 ^ x14;
assign n_2002 = n_508 ^ x17;
assign n_2003 = n_509 ^ x20;
assign n_2004 = n_510 ^ x23;
assign n_2005 = n_511 ^ x26;
assign n_2006 = n_512 ^ x29;
assign n_2007 = n_513 ^ x32;
assign n_2008 = n_514 ^ x35;
assign n_2009 = n_515 ^ x38;
assign n_2010 = n_516 ^ x41;
assign n_2011 = n_517 ^ x44;
assign n_2012 = n_518 ^ x47;
assign n_2013 = n_519 ^ x50;
assign n_2014 = n_520 ^ x53;
assign n_2015 = n_521 ^ x56;
assign n_2016 = n_522 ^ x59;
assign n_2017 = ~n_66 & n_523;
assign n_2018 = ~x1 & n_525;
assign n_2019 = n_526 ^ n_527;
assign n_2020 = x68 & ~n_528;
assign n_2021 = n_530 ^ n_111;
assign n_2022 = n_531 ^ x66;
assign n_2023 = n_533 ^ n_110;
assign n_2024 = n_535 ^ n_533;
assign n_2025 = ~n_66 & n_537;
assign n_2026 = x1 & n_538;
assign n_2027 = ~x1 & n_540;
assign n_2028 = ~x1 & n_541;
assign n_2029 = ~x1 & n_542;
assign n_2030 = n_543 ^ n_132;
assign n_2031 = ~n_66 & n_544;
assign n_2032 = ~n_66 & n_545;
assign n_2033 = n_546 ^ n_139;
assign n_2034 = x78 & n_548;
assign n_2035 = ~x1 & n_549;
assign n_2036 = ~n_66 & n_550;
assign n_2037 = n_551 ^ n_146;
assign n_2038 = n_552 ^ x79;
assign n_2039 = ~x1 & n_554;
assign n_2040 = x63 & n_555;
assign n_2041 = n_556 ^ n_158;
assign n_2042 = x1 & n_557;
assign n_2043 = ~x1 & n_558;
assign n_2044 = n_559 ^ n_171;
assign n_2045 = ~x1 & n_560;
assign n_2046 = ~x1 & n_561;
assign n_2047 = ~x1 & n_562;
assign n_2048 = x1 & n_563;
assign n_2049 = x1 & n_564;
assign n_2050 = n_565 ^ n_186;
assign n_2051 = n_566 ^ n_190;
assign n_2052 = ~n_66 & n_567;
assign n_2053 = n_569 ^ n_196;
assign n_2054 = ~x1 & n_570;
assign n_2055 = n_571 ^ n_199;
assign n_2056 = n_572 ^ n_568;
assign n_2057 = ~x1 & n_573;
assign n_2058 = ~x1 & n_574;
assign n_2059 = n_210 & n_575;
assign n_2060 = x1 & n_576;
assign n_2061 = n_577 ^ n_221;
assign n_2062 = ~x1 & n_578;
assign n_2063 = n_225 & n_579;
assign n_2064 = ~x1 & n_580;
assign n_2065 = n_581 ^ ~n_230;
assign n_2066 = ~n_66 & n_582;
assign n_2067 = ~x1 & n_583;
assign n_2068 = ~n_66 & n_584;
assign n_2069 = ~n_66 & n_585;
assign n_2070 = ~x1 & n_586;
assign n_2071 = ~n_66 & n_587;
assign n_2072 = ~n_66 & n_588;
assign n_2073 = n_589 ^ n_244;
assign n_2074 = ~x1 & n_590;
assign n_2075 = n_591 ^ n_245;
assign n_2076 = n_593 ^ n_249;
assign n_2077 = ~x62 & ~n_595;
assign n_2078 = ~n_66 & n_597;
assign n_2079 = ~x1 & n_598;
assign n_2080 = ~x1 & n_599;
assign n_2081 = ~n_66 & n_600;
assign n_2082 = ~x1 & n_601;
assign n_2083 = n_602 ^ n_265;
assign n_2084 = ~x1 & n_603;
assign n_2085 = n_604 ^ n_268;
assign n_2086 = x63 & n_606;
assign n_2087 = ~n_66 & n_607;
assign n_2088 = n_608 ^ n_269;
assign n_2089 = n_609 ^ x118;
assign n_2090 = n_609 ^ x120;
assign n_2091 = n_612 ^ x119;
assign n_2092 = n_613 ^ n_281;
assign n_2093 = ~n_66 & n_614;
assign n_2094 = n_615 ^ n_294;
assign n_2095 = n_618 ^ x63;
assign n_2096 = ~x1 & n_619;
assign n_2097 = x127 & n_620;
assign n_2098 = n_623 ^ x126;
assign n_2099 = n_627 ^ n_308;
assign n_2100 = n_630 ^ x2;
assign n_2101 = n_631 ^ x2;
assign n_2102 = n_632 ^ x2;
assign n_2103 = n_633 ^ x2;
assign n_2104 = n_634 ^ x2;
assign n_2105 = n_635 ^ x2;
assign n_2106 = n_636 ^ x2;
assign n_2107 = n_637 ^ x2;
assign n_2108 = n_638 ^ x2;
assign n_2109 = n_639 ^ x2;
assign n_2110 = n_640 ^ x2;
assign n_2111 = n_641 ^ x2;
assign n_2112 = n_642 ^ x2;
assign n_2113 = n_643 ^ x2;
assign n_2114 = n_644 ^ x2;
assign n_2115 = n_645 ^ x2;
assign n_2116 = n_646 ^ x2;
assign n_2117 = n_647 ^ x2;
assign n_2118 = n_648 ^ x2;
assign n_2119 = n_649 ^ x2;
assign n_2120 = n_650 ^ x2;
assign n_2121 = x65 & n_651;
assign n_2122 = x66 & n_651;
assign n_2123 = x67 & n_651;
assign n_2124 = x68 & n_651;
assign n_2125 = x69 & n_651;
assign n_2126 = x70 & n_651;
assign n_2127 = x71 & n_651;
assign n_2128 = x72 & n_651;
assign n_2129 = x73 & n_651;
assign n_2130 = x74 & n_651;
assign n_2131 = x75 & n_651;
assign n_2132 = x76 & n_651;
assign n_2133 = x77 & n_651;
assign n_2134 = x78 & n_651;
assign n_2135 = x79 & n_651;
assign n_2136 = x80 & n_651;
assign n_2137 = x81 & n_651;
assign n_2138 = x82 & n_651;
assign n_2139 = x83 & n_651;
assign n_2140 = x84 & n_651;
assign n_2141 = x85 & n_651;
assign n_2142 = x86 & n_651;
assign n_2143 = x87 & n_651;
assign n_2144 = x88 & n_651;
assign n_2145 = x89 & n_651;
assign n_2146 = x90 & n_651;
assign n_2147 = x91 & n_651;
assign n_2148 = x92 & n_651;
assign n_2149 = x93 & n_651;
assign n_2150 = x94 & n_651;
assign n_2151 = x95 & n_651;
assign n_2152 = x96 & n_651;
assign n_2153 = x97 & n_651;
assign n_2154 = x98 & n_651;
assign n_2155 = x99 & n_651;
assign n_2156 = x100 & n_651;
assign n_2157 = x101 & n_651;
assign n_2158 = x102 & n_651;
assign n_2159 = x103 & n_651;
assign n_2160 = x104 & n_651;
assign n_2161 = x105 & n_651;
assign n_2162 = x106 & n_651;
assign n_2163 = x107 & n_651;
assign n_2164 = x108 & n_651;
assign n_2165 = x109 & n_651;
assign n_2166 = x110 & n_651;
assign n_2167 = x111 & n_651;
assign n_2168 = x112 & n_651;
assign n_2169 = x113 & n_651;
assign n_2170 = x114 & n_651;
assign n_2171 = x115 & n_651;
assign n_2172 = x116 & n_651;
assign n_2173 = x117 & n_651;
assign n_2174 = x118 & n_651;
assign n_2175 = x119 & n_651;
assign n_2176 = x120 & n_651;
assign n_2177 = x121 & n_651;
assign n_2178 = x122 & n_651;
assign n_2179 = x123 & n_651;
assign n_2180 = x124 & n_651;
assign n_2181 = x125 & n_651;
assign n_2182 = x126 & n_651;
assign n_2183 = x127 & n_651;
assign n_2184 = n_6 & n_652;
assign n_2185 = x127 & n_652;
assign n_2186 = ~n_3 & ~n_654;
assign n_2187 = ~n_502 & n_655;
assign n_2188 = n_11 & n_717;
assign n_2189 = n_718 ^ n_342;
assign n_2190 = x127 & n_720;
assign n_2191 = ~n_502 & n_784;
assign n_2192 = x65 & n_846;
assign n_2193 = x66 & n_846;
assign n_2194 = x67 & n_846;
assign n_2195 = x68 & n_846;
assign n_2196 = x69 & n_846;
assign n_2197 = x70 & n_846;
assign n_2198 = x71 & n_846;
assign n_2199 = x72 & n_846;
assign n_2200 = x73 & n_846;
assign n_2201 = x74 & n_846;
assign n_2202 = x75 & n_846;
assign n_2203 = x76 & n_846;
assign n_2204 = x77 & n_846;
assign n_2205 = x78 & n_846;
assign n_2206 = x79 & n_846;
assign n_2207 = x80 & n_846;
assign n_2208 = x81 & n_846;
assign n_2209 = x82 & n_846;
assign n_2210 = x83 & n_846;
assign n_2211 = x84 & n_846;
assign n_2212 = x85 & n_846;
assign n_2213 = x86 & n_846;
assign n_2214 = x87 & n_846;
assign n_2215 = x88 & n_846;
assign n_2216 = x89 & n_846;
assign n_2217 = x90 & n_846;
assign n_2218 = x91 & n_846;
assign n_2219 = x92 & n_846;
assign n_2220 = x93 & n_846;
assign n_2221 = x94 & n_846;
assign n_2222 = x95 & n_846;
assign n_2223 = x96 & n_846;
assign n_2224 = x97 & n_846;
assign n_2225 = x98 & n_846;
assign n_2226 = x99 & n_846;
assign n_2227 = x100 & n_846;
assign n_2228 = x101 & n_846;
assign n_2229 = x102 & n_846;
assign n_2230 = x103 & n_846;
assign n_2231 = x104 & n_846;
assign n_2232 = x105 & n_846;
assign n_2233 = x106 & n_846;
assign n_2234 = x107 & n_846;
assign n_2235 = x108 & n_846;
assign n_2236 = x109 & n_846;
assign n_2237 = x110 & n_846;
assign n_2238 = x111 & n_846;
assign n_2239 = x112 & n_846;
assign n_2240 = x113 & n_846;
assign n_2241 = x114 & n_846;
assign n_2242 = x115 & n_846;
assign n_2243 = x116 & n_846;
assign n_2244 = x117 & n_846;
assign n_2245 = x118 & n_846;
assign n_2246 = x119 & n_846;
assign n_2247 = x120 & n_846;
assign n_2248 = x121 & n_846;
assign n_2249 = x122 & n_846;
assign n_2250 = x123 & n_846;
assign n_2251 = x124 & n_846;
assign n_2252 = x125 & n_846;
assign n_2253 = x126 & n_846;
assign n_2254 = x127 & n_846;
assign n_2255 = n_847 ^ n_350;
assign n_2256 = ~x64 & ~n_848;
assign n_2257 = x64 & n_849;
assign n_2258 = n_14 & ~n_850;
assign n_2259 = x127 & n_851;
assign n_2260 = x65 & n_852;
assign n_2261 = x66 & n_852;
assign n_2262 = x67 & n_852;
assign n_2263 = x68 & n_852;
assign n_2264 = x69 & n_852;
assign n_2265 = x70 & n_852;
assign n_2266 = x71 & n_852;
assign n_2267 = x72 & n_852;
assign n_2268 = x73 & n_852;
assign n_2269 = x74 & n_852;
assign n_2270 = x75 & n_852;
assign n_2271 = x76 & n_852;
assign n_2272 = x77 & n_852;
assign n_2273 = x78 & n_852;
assign n_2274 = x79 & n_852;
assign n_2275 = x80 & n_852;
assign n_2276 = x81 & n_852;
assign n_2277 = x82 & n_852;
assign n_2278 = x83 & n_852;
assign n_2279 = x84 & n_852;
assign n_2280 = x85 & n_852;
assign n_2281 = x86 & n_852;
assign n_2282 = x87 & n_852;
assign n_2283 = x88 & n_852;
assign n_2284 = x89 & n_852;
assign n_2285 = x90 & n_852;
assign n_2286 = x91 & n_852;
assign n_2287 = x92 & n_852;
assign n_2288 = x93 & n_852;
assign n_2289 = x94 & n_852;
assign n_2290 = x95 & n_852;
assign n_2291 = x96 & n_852;
assign n_2292 = x97 & n_852;
assign n_2293 = x98 & n_852;
assign n_2294 = x99 & n_852;
assign n_2295 = x100 & n_852;
assign n_2296 = x101 & n_852;
assign n_2297 = x102 & n_852;
assign n_2298 = x103 & n_852;
assign n_2299 = x104 & n_852;
assign n_2300 = x105 & n_852;
assign n_2301 = x106 & n_852;
assign n_2302 = x107 & n_852;
assign n_2303 = x108 & n_852;
assign n_2304 = x109 & n_852;
assign n_2305 = x110 & n_852;
assign n_2306 = x111 & n_852;
assign n_2307 = x112 & n_852;
assign n_2308 = x113 & n_852;
assign n_2309 = x114 & n_852;
assign n_2310 = x115 & n_852;
assign n_2311 = x116 & n_852;
assign n_2312 = x117 & n_852;
assign n_2313 = x118 & n_852;
assign n_2314 = x119 & n_852;
assign n_2315 = x120 & n_852;
assign n_2316 = x121 & n_852;
assign n_2317 = x122 & n_852;
assign n_2318 = x123 & n_852;
assign n_2319 = x124 & n_852;
assign n_2320 = x125 & n_852;
assign n_2321 = x126 & n_852;
assign n_2322 = x127 & n_852;
assign n_2323 = n_17 & n_853;
assign n_2324 = x127 & n_853;
assign n_2325 = ~n_502 & n_854;
assign n_2326 = ~x64 & ~n_916;
assign n_2327 = x65 & ~n_918;
assign n_2328 = x66 & ~n_918;
assign n_2329 = x67 & ~n_918;
assign n_2330 = x68 & ~n_918;
assign n_2331 = x69 & ~n_918;
assign n_2332 = x70 & ~n_918;
assign n_2333 = x71 & ~n_918;
assign n_2334 = x72 & ~n_918;
assign n_2335 = x73 & ~n_918;
assign n_2336 = x74 & ~n_918;
assign n_2337 = x75 & ~n_918;
assign n_2338 = x76 & ~n_918;
assign n_2339 = x77 & ~n_918;
assign n_2340 = x78 & ~n_918;
assign n_2341 = x79 & ~n_918;
assign n_2342 = x80 & ~n_918;
assign n_2343 = x81 & ~n_918;
assign n_2344 = x82 & ~n_918;
assign n_2345 = x83 & ~n_918;
assign n_2346 = x84 & ~n_918;
assign n_2347 = x85 & ~n_918;
assign n_2348 = x86 & ~n_918;
assign n_2349 = x87 & ~n_918;
assign n_2350 = x88 & ~n_918;
assign n_2351 = x89 & ~n_918;
assign n_2352 = x90 & ~n_918;
assign n_2353 = x91 & ~n_918;
assign n_2354 = x92 & ~n_918;
assign n_2355 = x93 & ~n_918;
assign n_2356 = x94 & ~n_918;
assign n_2357 = x95 & ~n_918;
assign n_2358 = x96 & ~n_918;
assign n_2359 = x97 & ~n_918;
assign n_2360 = x98 & ~n_918;
assign n_2361 = x99 & ~n_918;
assign n_2362 = x100 & ~n_918;
assign n_2363 = x101 & ~n_918;
assign n_2364 = x102 & ~n_918;
assign n_2365 = x103 & ~n_918;
assign n_2366 = x104 & ~n_918;
assign n_2367 = x105 & ~n_918;
assign n_2368 = x106 & ~n_918;
assign n_2369 = x107 & ~n_918;
assign n_2370 = x108 & ~n_918;
assign n_2371 = x109 & ~n_918;
assign n_2372 = x110 & ~n_918;
assign n_2373 = x111 & ~n_918;
assign n_2374 = x112 & ~n_918;
assign n_2375 = x113 & ~n_918;
assign n_2376 = x114 & ~n_918;
assign n_2377 = x115 & ~n_918;
assign n_2378 = x116 & ~n_918;
assign n_2379 = x117 & ~n_918;
assign n_2380 = x118 & ~n_918;
assign n_2381 = x119 & ~n_918;
assign n_2382 = x120 & ~n_918;
assign n_2383 = x121 & ~n_918;
assign n_2384 = x122 & ~n_918;
assign n_2385 = x123 & ~n_918;
assign n_2386 = x124 & ~n_918;
assign n_2387 = x125 & ~n_918;
assign n_2388 = x126 & ~n_918;
assign n_2389 = x127 & ~n_918;
assign n_2390 = n_20 & ~n_919;
assign n_2391 = x127 & ~n_919;
assign n_2392 = ~n_502 & n_920;
assign n_2393 = ~x64 & ~n_982;
assign n_2394 = x65 & ~n_984;
assign n_2395 = x66 & ~n_984;
assign n_2396 = x67 & ~n_984;
assign n_2397 = x68 & ~n_984;
assign n_2398 = x69 & ~n_984;
assign n_2399 = x70 & ~n_984;
assign n_2400 = x71 & ~n_984;
assign n_2401 = x72 & ~n_984;
assign n_2402 = x73 & ~n_984;
assign n_2403 = x74 & ~n_984;
assign n_2404 = x75 & ~n_984;
assign n_2405 = x76 & ~n_984;
assign n_2406 = x77 & ~n_984;
assign n_2407 = x78 & ~n_984;
assign n_2408 = x79 & ~n_984;
assign n_2409 = x80 & ~n_984;
assign n_2410 = x81 & ~n_984;
assign n_2411 = x82 & ~n_984;
assign n_2412 = x83 & ~n_984;
assign n_2413 = x84 & ~n_984;
assign n_2414 = x85 & ~n_984;
assign n_2415 = x86 & ~n_984;
assign n_2416 = x87 & ~n_984;
assign n_2417 = x88 & ~n_984;
assign n_2418 = x89 & ~n_984;
assign n_2419 = x90 & ~n_984;
assign n_2420 = x91 & ~n_984;
assign n_2421 = x92 & ~n_984;
assign n_2422 = x93 & ~n_984;
assign n_2423 = x94 & ~n_984;
assign n_2424 = x95 & ~n_984;
assign n_2425 = x96 & ~n_984;
assign n_2426 = x97 & ~n_984;
assign n_2427 = x98 & ~n_984;
assign n_2428 = x99 & ~n_984;
assign n_2429 = x100 & ~n_984;
assign n_2430 = x101 & ~n_984;
assign n_2431 = x102 & ~n_984;
assign n_2432 = x103 & ~n_984;
assign n_2433 = x104 & ~n_984;
assign n_2434 = x105 & ~n_984;
assign n_2435 = x106 & ~n_984;
assign n_2436 = x107 & ~n_984;
assign n_2437 = x108 & ~n_984;
assign n_2438 = x109 & ~n_984;
assign n_2439 = x110 & ~n_984;
assign n_2440 = x111 & ~n_984;
assign n_2441 = x112 & ~n_984;
assign n_2442 = x113 & ~n_984;
assign n_2443 = x114 & ~n_984;
assign n_2444 = x115 & ~n_984;
assign n_2445 = x116 & ~n_984;
assign n_2446 = x117 & ~n_984;
assign n_2447 = x118 & ~n_984;
assign n_2448 = x119 & ~n_984;
assign n_2449 = x120 & ~n_984;
assign n_2450 = x121 & ~n_984;
assign n_2451 = x122 & ~n_984;
assign n_2452 = x123 & ~n_984;
assign n_2453 = x124 & ~n_984;
assign n_2454 = x125 & ~n_984;
assign n_2455 = x126 & ~n_984;
assign n_2456 = x127 & ~n_984;
assign n_2457 = n_23 & ~n_985;
assign n_2458 = x127 & ~n_985;
assign n_2459 = ~n_502 & n_986;
assign n_2460 = ~x64 & ~n_1048;
assign n_2461 = x65 & ~n_1050;
assign n_2462 = x66 & ~n_1050;
assign n_2463 = x67 & ~n_1050;
assign n_2464 = x68 & ~n_1050;
assign n_2465 = x69 & ~n_1050;
assign n_2466 = x70 & ~n_1050;
assign n_2467 = x71 & ~n_1050;
assign n_2468 = x72 & ~n_1050;
assign n_2469 = x73 & ~n_1050;
assign n_2470 = x74 & ~n_1050;
assign n_2471 = x75 & ~n_1050;
assign n_2472 = x76 & ~n_1050;
assign n_2473 = x77 & ~n_1050;
assign n_2474 = x78 & ~n_1050;
assign n_2475 = x79 & ~n_1050;
assign n_2476 = x80 & ~n_1050;
assign n_2477 = x81 & ~n_1050;
assign n_2478 = x82 & ~n_1050;
assign n_2479 = x83 & ~n_1050;
assign n_2480 = x84 & ~n_1050;
assign n_2481 = x85 & ~n_1050;
assign n_2482 = x86 & ~n_1050;
assign n_2483 = x87 & ~n_1050;
assign n_2484 = x88 & ~n_1050;
assign n_2485 = x89 & ~n_1050;
assign n_2486 = x90 & ~n_1050;
assign n_2487 = x91 & ~n_1050;
assign n_2488 = x92 & ~n_1050;
assign n_2489 = x93 & ~n_1050;
assign n_2490 = x94 & ~n_1050;
assign n_2491 = x95 & ~n_1050;
assign n_2492 = x96 & ~n_1050;
assign n_2493 = x97 & ~n_1050;
assign n_2494 = x98 & ~n_1050;
assign n_2495 = x99 & ~n_1050;
assign n_2496 = x100 & ~n_1050;
assign n_2497 = x101 & ~n_1050;
assign n_2498 = x102 & ~n_1050;
assign n_2499 = x103 & ~n_1050;
assign n_2500 = x104 & ~n_1050;
assign n_2501 = x105 & ~n_1050;
assign n_2502 = x106 & ~n_1050;
assign n_2503 = x107 & ~n_1050;
assign n_2504 = x108 & ~n_1050;
assign n_2505 = x109 & ~n_1050;
assign n_2506 = x110 & ~n_1050;
assign n_2507 = x111 & ~n_1050;
assign n_2508 = x112 & ~n_1050;
assign n_2509 = x113 & ~n_1050;
assign n_2510 = x114 & ~n_1050;
assign n_2511 = x115 & ~n_1050;
assign n_2512 = x116 & ~n_1050;
assign n_2513 = x117 & ~n_1050;
assign n_2514 = x118 & ~n_1050;
assign n_2515 = x119 & ~n_1050;
assign n_2516 = x120 & ~n_1050;
assign n_2517 = x121 & ~n_1050;
assign n_2518 = x122 & ~n_1050;
assign n_2519 = x123 & ~n_1050;
assign n_2520 = x124 & ~n_1050;
assign n_2521 = x125 & ~n_1050;
assign n_2522 = x126 & ~n_1050;
assign n_2523 = x127 & ~n_1050;
assign n_2524 = n_26 & ~n_1051;
assign n_2525 = x127 & ~n_1051;
assign n_2526 = ~n_502 & n_1052;
assign n_2527 = x65 & n_1114;
assign n_2528 = x66 & n_1114;
assign n_2529 = x67 & n_1114;
assign n_2530 = x68 & n_1114;
assign n_2531 = x69 & n_1114;
assign n_2532 = x70 & n_1114;
assign n_2533 = x71 & n_1114;
assign n_2534 = x72 & n_1114;
assign n_2535 = x73 & n_1114;
assign n_2536 = x74 & n_1114;
assign n_2537 = x75 & n_1114;
assign n_2538 = x76 & n_1114;
assign n_2539 = x77 & n_1114;
assign n_2540 = x78 & n_1114;
assign n_2541 = x79 & n_1114;
assign n_2542 = x80 & n_1114;
assign n_2543 = x81 & n_1114;
assign n_2544 = x82 & n_1114;
assign n_2545 = x83 & n_1114;
assign n_2546 = x84 & n_1114;
assign n_2547 = x85 & n_1114;
assign n_2548 = x86 & n_1114;
assign n_2549 = x87 & n_1114;
assign n_2550 = x88 & n_1114;
assign n_2551 = x89 & n_1114;
assign n_2552 = x90 & n_1114;
assign n_2553 = x91 & n_1114;
assign n_2554 = x92 & n_1114;
assign n_2555 = x93 & n_1114;
assign n_2556 = x94 & n_1114;
assign n_2557 = x95 & n_1114;
assign n_2558 = x96 & n_1114;
assign n_2559 = x97 & n_1114;
assign n_2560 = x98 & n_1114;
assign n_2561 = x99 & n_1114;
assign n_2562 = x100 & n_1114;
assign n_2563 = x101 & n_1114;
assign n_2564 = x102 & n_1114;
assign n_2565 = x103 & n_1114;
assign n_2566 = x104 & n_1114;
assign n_2567 = x105 & n_1114;
assign n_2568 = x106 & n_1114;
assign n_2569 = x107 & n_1114;
assign n_2570 = x108 & n_1114;
assign n_2571 = x109 & n_1114;
assign n_2572 = x110 & n_1114;
assign n_2573 = x111 & n_1114;
assign n_2574 = x112 & n_1114;
assign n_2575 = x113 & n_1114;
assign n_2576 = x114 & n_1114;
assign n_2577 = x115 & n_1114;
assign n_2578 = x116 & n_1114;
assign n_2579 = x117 & n_1114;
assign n_2580 = x118 & n_1114;
assign n_2581 = x119 & n_1114;
assign n_2582 = x120 & n_1114;
assign n_2583 = x121 & n_1114;
assign n_2584 = x122 & n_1114;
assign n_2585 = x123 & n_1114;
assign n_2586 = x124 & n_1114;
assign n_2587 = x125 & n_1114;
assign n_2588 = x126 & n_1114;
assign n_2589 = x127 & n_1114;
assign n_2590 = n_29 & n_1115;
assign n_2591 = ~n_502 & n_1117;
assign n_2592 = x65 & n_1178;
assign n_2593 = x66 & n_1178;
assign n_2594 = x67 & n_1178;
assign n_2595 = x68 & n_1178;
assign n_2596 = x69 & n_1178;
assign n_2597 = x70 & n_1178;
assign n_2598 = x71 & n_1178;
assign n_2599 = x72 & n_1178;
assign n_2600 = x73 & n_1178;
assign n_2601 = x74 & n_1178;
assign n_2602 = x75 & n_1178;
assign n_2603 = x76 & n_1178;
assign n_2604 = x77 & n_1178;
assign n_2605 = x78 & n_1178;
assign n_2606 = x79 & n_1178;
assign n_2607 = x80 & n_1178;
assign n_2608 = x81 & n_1178;
assign n_2609 = x82 & n_1178;
assign n_2610 = x83 & n_1178;
assign n_2611 = x84 & n_1178;
assign n_2612 = x85 & n_1178;
assign n_2613 = x86 & n_1178;
assign n_2614 = x87 & n_1178;
assign n_2615 = x88 & n_1178;
assign n_2616 = x89 & n_1178;
assign n_2617 = x90 & n_1178;
assign n_2618 = x91 & n_1178;
assign n_2619 = x92 & n_1178;
assign n_2620 = x93 & n_1178;
assign n_2621 = x94 & n_1178;
assign n_2622 = x95 & n_1178;
assign n_2623 = x96 & n_1178;
assign n_2624 = x97 & n_1178;
assign n_2625 = x98 & n_1178;
assign n_2626 = x99 & n_1178;
assign n_2627 = x100 & n_1178;
assign n_2628 = x101 & n_1178;
assign n_2629 = x102 & n_1178;
assign n_2630 = x103 & n_1178;
assign n_2631 = x104 & n_1178;
assign n_2632 = x105 & n_1178;
assign n_2633 = x106 & n_1178;
assign n_2634 = x107 & n_1178;
assign n_2635 = x108 & n_1178;
assign n_2636 = x109 & n_1178;
assign n_2637 = x110 & n_1178;
assign n_2638 = x111 & n_1178;
assign n_2639 = x112 & n_1178;
assign n_2640 = x113 & n_1178;
assign n_2641 = x114 & n_1178;
assign n_2642 = x115 & n_1178;
assign n_2643 = x116 & n_1178;
assign n_2644 = x117 & n_1178;
assign n_2645 = x118 & n_1178;
assign n_2646 = x119 & n_1178;
assign n_2647 = x120 & n_1178;
assign n_2648 = x121 & n_1178;
assign n_2649 = x122 & n_1178;
assign n_2650 = x123 & n_1178;
assign n_2651 = x124 & n_1178;
assign n_2652 = x125 & n_1178;
assign n_2653 = x126 & n_1178;
assign n_2654 = x127 & n_1178;
assign n_2655 = n_32 & n_1179;
assign n_2656 = x127 & n_1179;
assign n_2657 = ~n_502 & n_1181;
assign n_2658 = ~x64 & ~n_1243;
assign n_2659 = x65 & ~n_1245;
assign n_2660 = x66 & ~n_1245;
assign n_2661 = x67 & ~n_1245;
assign n_2662 = x68 & ~n_1245;
assign n_2663 = x69 & ~n_1245;
assign n_2664 = x70 & ~n_1245;
assign n_2665 = x71 & ~n_1245;
assign n_2666 = x72 & ~n_1245;
assign n_2667 = x73 & ~n_1245;
assign n_2668 = x74 & ~n_1245;
assign n_2669 = x75 & ~n_1245;
assign n_2670 = x76 & ~n_1245;
assign n_2671 = x77 & ~n_1245;
assign n_2672 = x78 & ~n_1245;
assign n_2673 = x79 & ~n_1245;
assign n_2674 = x80 & ~n_1245;
assign n_2675 = x81 & ~n_1245;
assign n_2676 = x82 & ~n_1245;
assign n_2677 = x83 & ~n_1245;
assign n_2678 = x84 & ~n_1245;
assign n_2679 = x85 & ~n_1245;
assign n_2680 = x86 & ~n_1245;
assign n_2681 = x87 & ~n_1245;
assign n_2682 = x88 & ~n_1245;
assign n_2683 = x89 & ~n_1245;
assign n_2684 = x90 & ~n_1245;
assign n_2685 = x91 & ~n_1245;
assign n_2686 = x92 & ~n_1245;
assign n_2687 = x93 & ~n_1245;
assign n_2688 = x94 & ~n_1245;
assign n_2689 = x95 & ~n_1245;
assign n_2690 = x96 & ~n_1245;
assign n_2691 = x97 & ~n_1245;
assign n_2692 = x98 & ~n_1245;
assign n_2693 = x99 & ~n_1245;
assign n_2694 = x100 & ~n_1245;
assign n_2695 = x101 & ~n_1245;
assign n_2696 = x102 & ~n_1245;
assign n_2697 = x103 & ~n_1245;
assign n_2698 = x104 & ~n_1245;
assign n_2699 = x105 & ~n_1245;
assign n_2700 = x106 & ~n_1245;
assign n_2701 = x107 & ~n_1245;
assign n_2702 = x108 & ~n_1245;
assign n_2703 = x109 & ~n_1245;
assign n_2704 = x110 & ~n_1245;
assign n_2705 = x111 & ~n_1245;
assign n_2706 = x112 & ~n_1245;
assign n_2707 = x113 & ~n_1245;
assign n_2708 = x114 & ~n_1245;
assign n_2709 = x115 & ~n_1245;
assign n_2710 = x116 & ~n_1245;
assign n_2711 = x117 & ~n_1245;
assign n_2712 = x118 & ~n_1245;
assign n_2713 = x119 & ~n_1245;
assign n_2714 = x120 & ~n_1245;
assign n_2715 = x121 & ~n_1245;
assign n_2716 = x122 & ~n_1245;
assign n_2717 = x123 & ~n_1245;
assign n_2718 = x124 & ~n_1245;
assign n_2719 = x125 & ~n_1245;
assign n_2720 = x126 & ~n_1245;
assign n_2721 = x127 & ~n_1245;
assign n_2722 = n_35 & ~n_1246;
assign n_2723 = x32 & n_1247;
assign n_2724 = x127 & n_1247;
assign n_2725 = ~n_502 & n_1248;
assign n_2726 = ~x64 & ~n_1310;
assign n_2727 = x65 & ~n_1312;
assign n_2728 = x66 & ~n_1312;
assign n_2729 = x67 & ~n_1312;
assign n_2730 = x68 & ~n_1312;
assign n_2731 = x69 & ~n_1312;
assign n_2732 = x70 & ~n_1312;
assign n_2733 = x71 & ~n_1312;
assign n_2734 = x72 & ~n_1312;
assign n_2735 = x73 & ~n_1312;
assign n_2736 = x74 & ~n_1312;
assign n_2737 = x75 & ~n_1312;
assign n_2738 = x76 & ~n_1312;
assign n_2739 = x77 & ~n_1312;
assign n_2740 = x78 & ~n_1312;
assign n_2741 = x79 & ~n_1312;
assign n_2742 = x80 & ~n_1312;
assign n_2743 = x81 & ~n_1312;
assign n_2744 = x82 & ~n_1312;
assign n_2745 = x83 & ~n_1312;
assign n_2746 = x84 & ~n_1312;
assign n_2747 = x85 & ~n_1312;
assign n_2748 = x86 & ~n_1312;
assign n_2749 = x87 & ~n_1312;
assign n_2750 = x88 & ~n_1312;
assign n_2751 = x89 & ~n_1312;
assign n_2752 = x90 & ~n_1312;
assign n_2753 = x91 & ~n_1312;
assign n_2754 = x92 & ~n_1312;
assign n_2755 = x93 & ~n_1312;
assign n_2756 = x94 & ~n_1312;
assign n_2757 = x95 & ~n_1312;
assign n_2758 = x96 & ~n_1312;
assign n_2759 = x97 & ~n_1312;
assign n_2760 = x98 & ~n_1312;
assign n_2761 = x99 & ~n_1312;
assign n_2762 = x100 & ~n_1312;
assign n_2763 = x101 & ~n_1312;
assign n_2764 = x102 & ~n_1312;
assign n_2765 = x103 & ~n_1312;
assign n_2766 = x104 & ~n_1312;
assign n_2767 = x105 & ~n_1312;
assign n_2768 = x106 & ~n_1312;
assign n_2769 = x107 & ~n_1312;
assign n_2770 = x108 & ~n_1312;
assign n_2771 = x109 & ~n_1312;
assign n_2772 = x110 & ~n_1312;
assign n_2773 = x111 & ~n_1312;
assign n_2774 = x112 & ~n_1312;
assign n_2775 = x113 & ~n_1312;
assign n_2776 = x114 & ~n_1312;
assign n_2777 = x115 & ~n_1312;
assign n_2778 = x116 & ~n_1312;
assign n_2779 = x117 & ~n_1312;
assign n_2780 = x118 & ~n_1312;
assign n_2781 = x119 & ~n_1312;
assign n_2782 = x120 & ~n_1312;
assign n_2783 = x121 & ~n_1312;
assign n_2784 = x122 & ~n_1312;
assign n_2785 = x123 & ~n_1312;
assign n_2786 = x124 & ~n_1312;
assign n_2787 = x125 & ~n_1312;
assign n_2788 = x126 & ~n_1312;
assign n_2789 = x127 & ~n_1312;
assign n_2790 = n_38 & ~n_1313;
assign n_2791 = x127 & ~n_1313;
assign n_2792 = ~n_502 & n_1314;
assign n_2793 = ~x64 & ~n_1376;
assign n_2794 = x65 & ~n_1378;
assign n_2795 = x66 & ~n_1378;
assign n_2796 = x67 & ~n_1378;
assign n_2797 = x68 & ~n_1378;
assign n_2798 = x69 & ~n_1378;
assign n_2799 = x70 & ~n_1378;
assign n_2800 = x71 & ~n_1378;
assign n_2801 = x72 & ~n_1378;
assign n_2802 = x73 & ~n_1378;
assign n_2803 = x74 & ~n_1378;
assign n_2804 = x75 & ~n_1378;
assign n_2805 = x76 & ~n_1378;
assign n_2806 = x77 & ~n_1378;
assign n_2807 = x78 & ~n_1378;
assign n_2808 = x79 & ~n_1378;
assign n_2809 = x80 & ~n_1378;
assign n_2810 = x81 & ~n_1378;
assign n_2811 = x82 & ~n_1378;
assign n_2812 = x83 & ~n_1378;
assign n_2813 = x84 & ~n_1378;
assign n_2814 = x85 & ~n_1378;
assign n_2815 = x86 & ~n_1378;
assign n_2816 = x87 & ~n_1378;
assign n_2817 = x88 & ~n_1378;
assign n_2818 = x89 & ~n_1378;
assign n_2819 = x90 & ~n_1378;
assign n_2820 = x91 & ~n_1378;
assign n_2821 = x92 & ~n_1378;
assign n_2822 = x93 & ~n_1378;
assign n_2823 = x94 & ~n_1378;
assign n_2824 = x95 & ~n_1378;
assign n_2825 = x96 & ~n_1378;
assign n_2826 = x97 & ~n_1378;
assign n_2827 = x98 & ~n_1378;
assign n_2828 = x99 & ~n_1378;
assign n_2829 = x100 & ~n_1378;
assign n_2830 = x101 & ~n_1378;
assign n_2831 = x102 & ~n_1378;
assign n_2832 = x103 & ~n_1378;
assign n_2833 = x104 & ~n_1378;
assign n_2834 = x105 & ~n_1378;
assign n_2835 = x106 & ~n_1378;
assign n_2836 = x107 & ~n_1378;
assign n_2837 = x108 & ~n_1378;
assign n_2838 = x109 & ~n_1378;
assign n_2839 = x110 & ~n_1378;
assign n_2840 = x111 & ~n_1378;
assign n_2841 = x112 & ~n_1378;
assign n_2842 = x113 & ~n_1378;
assign n_2843 = x114 & ~n_1378;
assign n_2844 = x115 & ~n_1378;
assign n_2845 = x116 & ~n_1378;
assign n_2846 = x117 & ~n_1378;
assign n_2847 = x118 & ~n_1378;
assign n_2848 = x119 & ~n_1378;
assign n_2849 = x120 & ~n_1378;
assign n_2850 = x121 & ~n_1378;
assign n_2851 = x122 & ~n_1378;
assign n_2852 = x123 & ~n_1378;
assign n_2853 = x124 & ~n_1378;
assign n_2854 = x125 & ~n_1378;
assign n_2855 = x126 & ~n_1378;
assign n_2856 = x127 & ~n_1378;
assign n_2857 = n_41 & ~n_1379;
assign n_2858 = x127 & ~n_1379;
assign n_2859 = ~n_502 & n_1380;
assign n_2860 = n_1442 ^ n_42;
assign n_2861 = n_1442 ^ x40;
assign n_2862 = x65 & ~n_1443;
assign n_2863 = x66 & ~n_1443;
assign n_2864 = x67 & ~n_1443;
assign n_2865 = x68 & ~n_1443;
assign n_2866 = x69 & ~n_1443;
assign n_2867 = x70 & ~n_1443;
assign n_2868 = x71 & ~n_1443;
assign n_2869 = x72 & ~n_1443;
assign n_2870 = x73 & ~n_1443;
assign n_2871 = x74 & ~n_1443;
assign n_2872 = x75 & ~n_1443;
assign n_2873 = x76 & ~n_1443;
assign n_2874 = x77 & ~n_1443;
assign n_2875 = x78 & ~n_1443;
assign n_2876 = x79 & ~n_1443;
assign n_2877 = x80 & ~n_1443;
assign n_2878 = x81 & ~n_1443;
assign n_2879 = x82 & ~n_1443;
assign n_2880 = x83 & ~n_1443;
assign n_2881 = x84 & ~n_1443;
assign n_2882 = x85 & ~n_1443;
assign n_2883 = x86 & ~n_1443;
assign n_2884 = x87 & ~n_1443;
assign n_2885 = x88 & ~n_1443;
assign n_2886 = x89 & ~n_1443;
assign n_2887 = x90 & ~n_1443;
assign n_2888 = x91 & ~n_1443;
assign n_2889 = x92 & ~n_1443;
assign n_2890 = x93 & ~n_1443;
assign n_2891 = x94 & ~n_1443;
assign n_2892 = x95 & ~n_1443;
assign n_2893 = x96 & ~n_1443;
assign n_2894 = x97 & ~n_1443;
assign n_2895 = x98 & ~n_1443;
assign n_2896 = x99 & ~n_1443;
assign n_2897 = x100 & ~n_1443;
assign n_2898 = x101 & ~n_1443;
assign n_2899 = x102 & ~n_1443;
assign n_2900 = x103 & ~n_1443;
assign n_2901 = x104 & ~n_1443;
assign n_2902 = x105 & ~n_1443;
assign n_2903 = x106 & ~n_1443;
assign n_2904 = x107 & ~n_1443;
assign n_2905 = x108 & ~n_1443;
assign n_2906 = x109 & ~n_1443;
assign n_2907 = x110 & ~n_1443;
assign n_2908 = x111 & ~n_1443;
assign n_2909 = x112 & ~n_1443;
assign n_2910 = x113 & ~n_1443;
assign n_2911 = x114 & ~n_1443;
assign n_2912 = x115 & ~n_1443;
assign n_2913 = x116 & ~n_1443;
assign n_2914 = x117 & ~n_1443;
assign n_2915 = x118 & ~n_1443;
assign n_2916 = x119 & ~n_1443;
assign n_2917 = x120 & ~n_1443;
assign n_2918 = x121 & ~n_1443;
assign n_2919 = x122 & ~n_1443;
assign n_2920 = x123 & ~n_1443;
assign n_2921 = x124 & ~n_1443;
assign n_2922 = x125 & ~n_1443;
assign n_2923 = x126 & ~n_1443;
assign n_2924 = x127 & ~n_1443;
assign n_2925 = n_44 & ~n_1444;
assign n_2926 = ~n_502 & n_1445;
assign n_2927 = ~x64 & ~n_1506;
assign n_2928 = x65 & ~n_1508;
assign n_2929 = x66 & ~n_1508;
assign n_2930 = x67 & ~n_1508;
assign n_2931 = x68 & ~n_1508;
assign n_2932 = x69 & ~n_1508;
assign n_2933 = x70 & ~n_1508;
assign n_2934 = x71 & ~n_1508;
assign n_2935 = x72 & ~n_1508;
assign n_2936 = x73 & ~n_1508;
assign n_2937 = x74 & ~n_1508;
assign n_2938 = x75 & ~n_1508;
assign n_2939 = x76 & ~n_1508;
assign n_2940 = x77 & ~n_1508;
assign n_2941 = x78 & ~n_1508;
assign n_2942 = x79 & ~n_1508;
assign n_2943 = x80 & ~n_1508;
assign n_2944 = x81 & ~n_1508;
assign n_2945 = x82 & ~n_1508;
assign n_2946 = x83 & ~n_1508;
assign n_2947 = x84 & ~n_1508;
assign n_2948 = x85 & ~n_1508;
assign n_2949 = x86 & ~n_1508;
assign n_2950 = x87 & ~n_1508;
assign n_2951 = x88 & ~n_1508;
assign n_2952 = x89 & ~n_1508;
assign n_2953 = x90 & ~n_1508;
assign n_2954 = x91 & ~n_1508;
assign n_2955 = x92 & ~n_1508;
assign n_2956 = x93 & ~n_1508;
assign n_2957 = x94 & ~n_1508;
assign n_2958 = x95 & ~n_1508;
assign n_2959 = x96 & ~n_1508;
assign n_2960 = x97 & ~n_1508;
assign n_2961 = x98 & ~n_1508;
assign n_2962 = x99 & ~n_1508;
assign n_2963 = x100 & ~n_1508;
assign n_2964 = x101 & ~n_1508;
assign n_2965 = x102 & ~n_1508;
assign n_2966 = x103 & ~n_1508;
assign n_2967 = x104 & ~n_1508;
assign n_2968 = x105 & ~n_1508;
assign n_2969 = x106 & ~n_1508;
assign n_2970 = x107 & ~n_1508;
assign n_2971 = x108 & ~n_1508;
assign n_2972 = x109 & ~n_1508;
assign n_2973 = x110 & ~n_1508;
assign n_2974 = x111 & ~n_1508;
assign n_2975 = x112 & ~n_1508;
assign n_2976 = x113 & ~n_1508;
assign n_2977 = x114 & ~n_1508;
assign n_2978 = x115 & ~n_1508;
assign n_2979 = x116 & ~n_1508;
assign n_2980 = x117 & ~n_1508;
assign n_2981 = x118 & ~n_1508;
assign n_2982 = x119 & ~n_1508;
assign n_2983 = x120 & ~n_1508;
assign n_2984 = x121 & ~n_1508;
assign n_2985 = x122 & ~n_1508;
assign n_2986 = x123 & ~n_1508;
assign n_2987 = x124 & ~n_1508;
assign n_2988 = x125 & ~n_1508;
assign n_2989 = x126 & ~n_1508;
assign n_2990 = x127 & ~n_1508;
assign n_2991 = n_47 & ~n_1509;
assign n_2992 = x127 & ~n_1509;
assign n_2993 = ~n_502 & n_1510;
assign n_2994 = ~x64 & ~n_1572;
assign n_2995 = n_50 & ~n_1573;
assign n_2996 = x127 & ~n_1573;
assign n_2997 = x65 & ~n_1574;
assign n_2998 = x66 & ~n_1574;
assign n_2999 = x67 & ~n_1574;
assign n_3000 = x68 & ~n_1574;
assign n_3001 = x69 & ~n_1574;
assign n_3002 = x70 & ~n_1574;
assign n_3003 = x71 & ~n_1574;
assign n_3004 = x72 & ~n_1574;
assign n_3005 = x73 & ~n_1574;
assign n_3006 = x74 & ~n_1574;
assign n_3007 = x75 & ~n_1574;
assign n_3008 = x76 & ~n_1574;
assign n_3009 = x77 & ~n_1574;
assign n_3010 = x78 & ~n_1574;
assign n_3011 = x79 & ~n_1574;
assign n_3012 = x80 & ~n_1574;
assign n_3013 = x81 & ~n_1574;
assign n_3014 = x82 & ~n_1574;
assign n_3015 = x83 & ~n_1574;
assign n_3016 = x84 & ~n_1574;
assign n_3017 = x85 & ~n_1574;
assign n_3018 = x86 & ~n_1574;
assign n_3019 = x87 & ~n_1574;
assign n_3020 = x88 & ~n_1574;
assign n_3021 = x89 & ~n_1574;
assign n_3022 = x90 & ~n_1574;
assign n_3023 = x91 & ~n_1574;
assign n_3024 = x92 & ~n_1574;
assign n_3025 = x93 & ~n_1574;
assign n_3026 = x94 & ~n_1574;
assign n_3027 = x95 & ~n_1574;
assign n_3028 = x96 & ~n_1574;
assign n_3029 = x97 & ~n_1574;
assign n_3030 = x98 & ~n_1574;
assign n_3031 = x99 & ~n_1574;
assign n_3032 = x100 & ~n_1574;
assign n_3033 = x101 & ~n_1574;
assign n_3034 = x102 & ~n_1574;
assign n_3035 = x103 & ~n_1574;
assign n_3036 = x104 & ~n_1574;
assign n_3037 = x105 & ~n_1574;
assign n_3038 = x106 & ~n_1574;
assign n_3039 = x107 & ~n_1574;
assign n_3040 = x108 & ~n_1574;
assign n_3041 = x109 & ~n_1574;
assign n_3042 = x110 & ~n_1574;
assign n_3043 = x111 & ~n_1574;
assign n_3044 = x112 & ~n_1574;
assign n_3045 = x113 & ~n_1574;
assign n_3046 = x114 & ~n_1574;
assign n_3047 = x115 & ~n_1574;
assign n_3048 = x116 & ~n_1574;
assign n_3049 = x117 & ~n_1574;
assign n_3050 = x118 & ~n_1574;
assign n_3051 = x119 & ~n_1574;
assign n_3052 = x120 & ~n_1574;
assign n_3053 = x121 & ~n_1574;
assign n_3054 = x122 & ~n_1574;
assign n_3055 = x123 & ~n_1574;
assign n_3056 = x124 & ~n_1574;
assign n_3057 = x125 & ~n_1574;
assign n_3058 = x126 & ~n_1574;
assign n_3059 = x127 & ~n_1574;
assign n_3060 = x64 & n_1575;
assign n_3061 = ~n_502 & n_1576;
assign n_3062 = ~x64 & ~n_1637;
assign n_3063 = x65 & ~n_1639;
assign n_3064 = x66 & ~n_1639;
assign n_3065 = x67 & ~n_1639;
assign n_3066 = x68 & ~n_1639;
assign n_3067 = x69 & ~n_1639;
assign n_3068 = x70 & ~n_1639;
assign n_3069 = x71 & ~n_1639;
assign n_3070 = x72 & ~n_1639;
assign n_3071 = x73 & ~n_1639;
assign n_3072 = x74 & ~n_1639;
assign n_3073 = x75 & ~n_1639;
assign n_3074 = x76 & ~n_1639;
assign n_3075 = x77 & ~n_1639;
assign n_3076 = x78 & ~n_1639;
assign n_3077 = x79 & ~n_1639;
assign n_3078 = x80 & ~n_1639;
assign n_3079 = x81 & ~n_1639;
assign n_3080 = x82 & ~n_1639;
assign n_3081 = x83 & ~n_1639;
assign n_3082 = x84 & ~n_1639;
assign n_3083 = x85 & ~n_1639;
assign n_3084 = x86 & ~n_1639;
assign n_3085 = x87 & ~n_1639;
assign n_3086 = x88 & ~n_1639;
assign n_3087 = x89 & ~n_1639;
assign n_3088 = x90 & ~n_1639;
assign n_3089 = x91 & ~n_1639;
assign n_3090 = x92 & ~n_1639;
assign n_3091 = x93 & ~n_1639;
assign n_3092 = x94 & ~n_1639;
assign n_3093 = x95 & ~n_1639;
assign n_3094 = x96 & ~n_1639;
assign n_3095 = x97 & ~n_1639;
assign n_3096 = x98 & ~n_1639;
assign n_3097 = x99 & ~n_1639;
assign n_3098 = x100 & ~n_1639;
assign n_3099 = x101 & ~n_1639;
assign n_3100 = x102 & ~n_1639;
assign n_3101 = x103 & ~n_1639;
assign n_3102 = x104 & ~n_1639;
assign n_3103 = x105 & ~n_1639;
assign n_3104 = x106 & ~n_1639;
assign n_3105 = x107 & ~n_1639;
assign n_3106 = x108 & ~n_1639;
assign n_3107 = x109 & ~n_1639;
assign n_3108 = x110 & ~n_1639;
assign n_3109 = x111 & ~n_1639;
assign n_3110 = x112 & ~n_1639;
assign n_3111 = x113 & ~n_1639;
assign n_3112 = x114 & ~n_1639;
assign n_3113 = x115 & ~n_1639;
assign n_3114 = x116 & ~n_1639;
assign n_3115 = x117 & ~n_1639;
assign n_3116 = x118 & ~n_1639;
assign n_3117 = x119 & ~n_1639;
assign n_3118 = x120 & ~n_1639;
assign n_3119 = x121 & ~n_1639;
assign n_3120 = x122 & ~n_1639;
assign n_3121 = x123 & ~n_1639;
assign n_3122 = x124 & ~n_1639;
assign n_3123 = x125 & ~n_1639;
assign n_3124 = x126 & ~n_1639;
assign n_3125 = x127 & ~n_1639;
assign n_3126 = n_53 & ~n_1640;
assign n_3127 = x127 & ~n_1640;
assign n_3128 = ~n_502 & n_1641;
assign n_3129 = ~x64 & ~n_1703;
assign n_3130 = n_56 & ~n_1704;
assign n_3131 = x127 & ~n_1704;
assign n_3132 = x65 & ~n_1705;
assign n_3133 = x66 & ~n_1705;
assign n_3134 = x67 & ~n_1705;
assign n_3135 = x68 & ~n_1705;
assign n_3136 = x69 & ~n_1705;
assign n_3137 = x70 & ~n_1705;
assign n_3138 = x71 & ~n_1705;
assign n_3139 = x72 & ~n_1705;
assign n_3140 = x73 & ~n_1705;
assign n_3141 = x74 & ~n_1705;
assign n_3142 = x75 & ~n_1705;
assign n_3143 = x76 & ~n_1705;
assign n_3144 = x77 & ~n_1705;
assign n_3145 = x78 & ~n_1705;
assign n_3146 = x79 & ~n_1705;
assign n_3147 = x80 & ~n_1705;
assign n_3148 = x81 & ~n_1705;
assign n_3149 = x82 & ~n_1705;
assign n_3150 = x83 & ~n_1705;
assign n_3151 = x84 & ~n_1705;
assign n_3152 = x85 & ~n_1705;
assign n_3153 = x86 & ~n_1705;
assign n_3154 = x87 & ~n_1705;
assign n_3155 = x88 & ~n_1705;
assign n_3156 = x89 & ~n_1705;
assign n_3157 = x90 & ~n_1705;
assign n_3158 = x91 & ~n_1705;
assign n_3159 = x92 & ~n_1705;
assign n_3160 = x93 & ~n_1705;
assign n_3161 = x94 & ~n_1705;
assign n_3162 = x95 & ~n_1705;
assign n_3163 = x96 & ~n_1705;
assign n_3164 = x97 & ~n_1705;
assign n_3165 = x98 & ~n_1705;
assign n_3166 = x99 & ~n_1705;
assign n_3167 = x100 & ~n_1705;
assign n_3168 = x101 & ~n_1705;
assign n_3169 = x102 & ~n_1705;
assign n_3170 = x103 & ~n_1705;
assign n_3171 = x104 & ~n_1705;
assign n_3172 = x105 & ~n_1705;
assign n_3173 = x106 & ~n_1705;
assign n_3174 = x107 & ~n_1705;
assign n_3175 = x108 & ~n_1705;
assign n_3176 = x109 & ~n_1705;
assign n_3177 = x110 & ~n_1705;
assign n_3178 = x111 & ~n_1705;
assign n_3179 = x112 & ~n_1705;
assign n_3180 = x113 & ~n_1705;
assign n_3181 = x114 & ~n_1705;
assign n_3182 = x115 & ~n_1705;
assign n_3183 = x116 & ~n_1705;
assign n_3184 = x117 & ~n_1705;
assign n_3185 = x118 & ~n_1705;
assign n_3186 = x119 & ~n_1705;
assign n_3187 = x120 & ~n_1705;
assign n_3188 = x121 & ~n_1705;
assign n_3189 = x122 & ~n_1705;
assign n_3190 = x123 & ~n_1705;
assign n_3191 = x124 & ~n_1705;
assign n_3192 = x125 & ~n_1705;
assign n_3193 = x126 & ~n_1705;
assign n_3194 = x127 & ~n_1705;
assign n_3195 = ~n_502 & n_1706;
assign n_3196 = x65 & n_1768;
assign n_3197 = x66 & n_1768;
assign n_3198 = x67 & n_1768;
assign n_3199 = x68 & n_1768;
assign n_3200 = x69 & n_1768;
assign n_3201 = x70 & n_1768;
assign n_3202 = x71 & n_1768;
assign n_3203 = x72 & n_1768;
assign n_3204 = x73 & n_1768;
assign n_3205 = x74 & n_1768;
assign n_3206 = x75 & n_1768;
assign n_3207 = x76 & n_1768;
assign n_3208 = x77 & n_1768;
assign n_3209 = x78 & n_1768;
assign n_3210 = x79 & n_1768;
assign n_3211 = x80 & n_1768;
assign n_3212 = x81 & n_1768;
assign n_3213 = x82 & n_1768;
assign n_3214 = x83 & n_1768;
assign n_3215 = x84 & n_1768;
assign n_3216 = x85 & n_1768;
assign n_3217 = x86 & n_1768;
assign n_3218 = x87 & n_1768;
assign n_3219 = x88 & n_1768;
assign n_3220 = x89 & n_1768;
assign n_3221 = x90 & n_1768;
assign n_3222 = x91 & n_1768;
assign n_3223 = x92 & n_1768;
assign n_3224 = x93 & n_1768;
assign n_3225 = x94 & n_1768;
assign n_3226 = x95 & n_1768;
assign n_3227 = x96 & n_1768;
assign n_3228 = x97 & n_1768;
assign n_3229 = x98 & n_1768;
assign n_3230 = x99 & n_1768;
assign n_3231 = x100 & n_1768;
assign n_3232 = x101 & n_1768;
assign n_3233 = x102 & n_1768;
assign n_3234 = x103 & n_1768;
assign n_3235 = x104 & n_1768;
assign n_3236 = x105 & n_1768;
assign n_3237 = x106 & n_1768;
assign n_3238 = x107 & n_1768;
assign n_3239 = x108 & n_1768;
assign n_3240 = x109 & n_1768;
assign n_3241 = x110 & n_1768;
assign n_3242 = x111 & n_1768;
assign n_3243 = x112 & n_1768;
assign n_3244 = x113 & n_1768;
assign n_3245 = x114 & n_1768;
assign n_3246 = x115 & n_1768;
assign n_3247 = x116 & n_1768;
assign n_3248 = x117 & n_1768;
assign n_3249 = x118 & n_1768;
assign n_3250 = x119 & n_1768;
assign n_3251 = x120 & n_1768;
assign n_3252 = x121 & n_1768;
assign n_3253 = x122 & n_1768;
assign n_3254 = x123 & n_1768;
assign n_3255 = x124 & n_1768;
assign n_3256 = x125 & n_1768;
assign n_3257 = x126 & n_1768;
assign n_3258 = x127 & n_1768;
assign n_3259 = n_59 & n_1769;
assign n_3260 = ~n_502 & n_1771;
assign n_3261 = x65 & n_1832;
assign n_3262 = x66 & n_1832;
assign n_3263 = x67 & n_1832;
assign n_3264 = x68 & n_1832;
assign n_3265 = x69 & n_1832;
assign n_3266 = x70 & n_1832;
assign n_3267 = x71 & n_1832;
assign n_3268 = x72 & n_1832;
assign n_3269 = x73 & n_1832;
assign n_3270 = x74 & n_1832;
assign n_3271 = x75 & n_1832;
assign n_3272 = x76 & n_1832;
assign n_3273 = x77 & n_1832;
assign n_3274 = x78 & n_1832;
assign n_3275 = x79 & n_1832;
assign n_3276 = x80 & n_1832;
assign n_3277 = x81 & n_1832;
assign n_3278 = x82 & n_1832;
assign n_3279 = x83 & n_1832;
assign n_3280 = x84 & n_1832;
assign n_3281 = x85 & n_1832;
assign n_3282 = x86 & n_1832;
assign n_3283 = x87 & n_1832;
assign n_3284 = x88 & n_1832;
assign n_3285 = x89 & n_1832;
assign n_3286 = x90 & n_1832;
assign n_3287 = x91 & n_1832;
assign n_3288 = x92 & n_1832;
assign n_3289 = x93 & n_1832;
assign n_3290 = x94 & n_1832;
assign n_3291 = x95 & n_1832;
assign n_3292 = x96 & n_1832;
assign n_3293 = x97 & n_1832;
assign n_3294 = x98 & n_1832;
assign n_3295 = x99 & n_1832;
assign n_3296 = x100 & n_1832;
assign n_3297 = x101 & n_1832;
assign n_3298 = x102 & n_1832;
assign n_3299 = x103 & n_1832;
assign n_3300 = x104 & n_1832;
assign n_3301 = x105 & n_1832;
assign n_3302 = x106 & n_1832;
assign n_3303 = x107 & n_1832;
assign n_3304 = x108 & n_1832;
assign n_3305 = x109 & n_1832;
assign n_3306 = x110 & n_1832;
assign n_3307 = x111 & n_1832;
assign n_3308 = x112 & n_1832;
assign n_3309 = x113 & n_1832;
assign n_3310 = x114 & n_1832;
assign n_3311 = x115 & n_1832;
assign n_3312 = x116 & n_1832;
assign n_3313 = x117 & n_1832;
assign n_3314 = x118 & n_1832;
assign n_3315 = x119 & n_1832;
assign n_3316 = x120 & n_1832;
assign n_3317 = x121 & n_1832;
assign n_3318 = x122 & n_1832;
assign n_3319 = x123 & n_1832;
assign n_3320 = x124 & n_1832;
assign n_3321 = x125 & n_1832;
assign n_3322 = x126 & n_1832;
assign n_3323 = x127 & n_1832;
assign n_3324 = n_62 & n_1833;
assign n_3325 = ~n_502 & n_1835;
assign n_3326 = x65 & n_1896;
assign n_3327 = x66 & n_1896;
assign n_3328 = x67 & n_1896;
assign n_3329 = x68 & n_1896;
assign n_3330 = x69 & n_1896;
assign n_3331 = x70 & n_1896;
assign n_3332 = x71 & n_1896;
assign n_3333 = x72 & n_1896;
assign n_3334 = x73 & n_1896;
assign n_3335 = x74 & n_1896;
assign n_3336 = x75 & n_1896;
assign n_3337 = x76 & n_1896;
assign n_3338 = x77 & n_1896;
assign n_3339 = x78 & n_1896;
assign n_3340 = x79 & n_1896;
assign n_3341 = x80 & n_1896;
assign n_3342 = x81 & n_1896;
assign n_3343 = x82 & n_1896;
assign n_3344 = x83 & n_1896;
assign n_3345 = x84 & n_1896;
assign n_3346 = x85 & n_1896;
assign n_3347 = x86 & n_1896;
assign n_3348 = x87 & n_1896;
assign n_3349 = x88 & n_1896;
assign n_3350 = x89 & n_1896;
assign n_3351 = x90 & n_1896;
assign n_3352 = x91 & n_1896;
assign n_3353 = x92 & n_1896;
assign n_3354 = x93 & n_1896;
assign n_3355 = x94 & n_1896;
assign n_3356 = x95 & n_1896;
assign n_3357 = x96 & n_1896;
assign n_3358 = x97 & n_1896;
assign n_3359 = x98 & n_1896;
assign n_3360 = x99 & n_1896;
assign n_3361 = x100 & n_1896;
assign n_3362 = x101 & n_1896;
assign n_3363 = x102 & n_1896;
assign n_3364 = x103 & n_1896;
assign n_3365 = x104 & n_1896;
assign n_3366 = x105 & n_1896;
assign n_3367 = x106 & n_1896;
assign n_3368 = x107 & n_1896;
assign n_3369 = x108 & n_1896;
assign n_3370 = x109 & n_1896;
assign n_3371 = x110 & n_1896;
assign n_3372 = x111 & n_1896;
assign n_3373 = x112 & n_1896;
assign n_3374 = x113 & n_1896;
assign n_3375 = x114 & n_1896;
assign n_3376 = x115 & n_1896;
assign n_3377 = x116 & n_1896;
assign n_3378 = x117 & n_1896;
assign n_3379 = x118 & n_1896;
assign n_3380 = x119 & n_1896;
assign n_3381 = x120 & n_1896;
assign n_3382 = x121 & n_1896;
assign n_3383 = x122 & n_1896;
assign n_3384 = x123 & n_1896;
assign n_3385 = x124 & n_1896;
assign n_3386 = x125 & n_1896;
assign n_3387 = x126 & n_1896;
assign n_3388 = x127 & n_1896;
assign n_3389 = n_65 & n_1897;
assign n_3390 = ~n_502 & n_1899;
assign n_3391 = n_1961 ^ n_457;
assign n_3392 = n_459 ^ n_1961;
assign n_3393 = n_1962 ^ x71;
assign n_3394 = n_1963 ^ n_460;
assign n_3395 = ~x74 & n_1963;
assign n_3396 = n_1964 ^ x82;
assign n_3397 = n_1965 ^ n_461;
assign n_3398 = n_462 ^ n_1965;
assign n_3399 = n_1966 ^ x85;
assign n_3400 = n_1967 ^ n_464;
assign n_3401 = n_1968 ^ x88;
assign n_3402 = n_1969 ^ n_465;
assign n_3403 = n_466 ^ n_1969;
assign n_3404 = n_1970 ^ x89;
assign n_3405 = n_1971 ^ x94;
assign n_3406 = n_1972 ^ n_468;
assign n_3407 = n_470 ^ n_1972;
assign n_3408 = n_1973 ^ x95;
assign n_3409 = n_1974 ^ n_471;
assign n_3410 = n_473 ^ n_1974;
assign n_3411 = n_1975 ^ x98;
assign n_3412 = n_1976 ^ n_474;
assign n_3413 = n_475 ^ n_1976;
assign n_3414 = n_1977 ^ n_476;
assign n_3415 = n_478 ^ n_1977;
assign n_3416 = n_1978 ^ x110;
assign n_3417 = n_1979 ^ n_479;
assign n_3418 = n_480 ^ n_1979;
assign n_3419 = n_1980 ^ x116;
assign n_3420 = n_1981 ^ n_483;
assign n_3421 = n_484 ^ n_1981;
assign n_3422 = n_1982 ^ x122;
assign n_3423 = n_1983 ^ n_486;
assign n_3424 = n_622 & n_1983;
assign n_3425 = n_342 & n_1993;
assign n_3426 = n_1995 ^ x65;
assign n_3427 = ~x66 & n_1996;
assign n_3428 = n_1997 ^ x64;
assign n_3429 = n_1998 ^ x4;
assign n_3430 = n_1999 ^ x10;
assign n_3431 = n_2000 ^ x13;
assign n_3432 = n_2001 ^ x16;
assign n_3433 = n_2002 ^ x19;
assign n_3434 = n_2003 ^ x22;
assign n_3435 = n_2004 ^ x25;
assign n_3436 = n_2005 ^ x28;
assign n_3437 = n_2006 ^ x31;
assign n_3438 = n_2007 ^ x34;
assign n_3439 = n_2008 ^ x37;
assign n_3440 = n_2009 ^ x40;
assign n_3441 = n_2010 ^ x43;
assign n_3442 = n_2011 ^ x46;
assign n_3443 = n_2012 ^ x49;
assign n_3444 = n_2013 ^ x52;
assign n_3445 = n_2014 ^ x55;
assign n_3446 = n_2015 ^ x58;
assign n_3447 = n_2016 ^ x61;
assign n_3448 = n_2017 ^ x66;
assign n_3449 = n_2018 ^ n_103;
assign n_3450 = ~n_2019 & ~n_80;
assign n_3451 = ~x69 & ~n_2020;
assign n_3452 = n_2021 ^ x67;
assign n_3453 = n_2022 ^ n_110;
assign n_3454 = n_2022 ^ x2;
assign n_3455 = n_2023 ^ n_112;
assign n_3456 = n_2023 ^ x2;
assign n_3457 = n_2024 ^ x68;
assign n_3458 = n_2025 ^ x70;
assign n_3459 = n_2026 ^ n_114;
assign n_3460 = n_2027 ^ n_122;
assign n_3461 = n_2028 ^ n_126;
assign n_3462 = n_2029 ^ n_131;
assign n_3463 = x63 & n_2030;
assign n_3464 = n_2031 ^ x76;
assign n_3465 = n_2032 ^ x77;
assign n_3466 = ~n_66 & n_2033;
assign n_3467 = ~x62 & ~n_2034;
assign n_3468 = n_2035 ^ n_140;
assign n_3469 = n_2036 ^ x79;
assign n_3470 = n_2037 ^ x79;
assign n_3471 = n_2038 ^ n_148;
assign n_3472 = n_2038 ^ x80;
assign n_3473 = n_2039 ^ n_150;
assign n_3474 = ~x62 & ~n_2040;
assign n_3475 = n_2041 ^ x82;
assign n_3476 = n_2042 ^ n_159;
assign n_3477 = n_2043 ^ n_165;
assign n_3478 = ~n_66 & n_2044;
assign n_3479 = n_2045 ^ n_169;
assign n_3480 = n_2046 ^ n_172;
assign n_3481 = n_2047 ^ n_176;
assign n_3482 = n_2048 ^ n_177;
assign n_3483 = n_2049 ^ n_181;
assign n_3484 = n_2050 ^ x90;
assign n_3485 = n_2051 ^ x91;
assign n_3486 = n_2052 ^ x92;
assign n_3487 = ~n_66 & n_2053;
assign n_3488 = n_2054 ^ n_195;
assign n_3489 = n_2055 ^ x93;
assign n_3490 = n_2056 ^ n_572;
assign n_3491 = n_2057 ^ n_203;
assign n_3492 = n_2058 ^ n_207;
assign n_3493 = n_2059 ^ n_210;
assign n_3494 = n_2060 ^ n_212;
assign n_3495 = n_2061 ^ x99;
assign n_3496 = n_2062 ^ x101;
assign n_3497 = n_2063 ^ n_225;
assign n_3498 = n_2064 ^ n_228;
assign n_3499 = x63 & n_2065;
assign n_3500 = n_2066 ^ x103;
assign n_3501 = n_2067 ^ n_232;
assign n_3502 = n_2068 ^ x104;
assign n_3503 = n_2069 ^ x105;
assign n_3504 = n_2070 ^ n_237;
assign n_3505 = n_2071 ^ x106;
assign n_3506 = n_2072 ^ x107;
assign n_3507 = ~n_66 & n_2073;
assign n_3508 = n_2074 ^ n_243;
assign n_3509 = n_2075 ^ x107;
assign n_3510 = n_2076 ^ x108;
assign n_3511 = n_2077 ^ n_596;
assign n_3512 = n_2077 ^ n_594;
assign n_3513 = n_2078 ^ x109;
assign n_3514 = n_2079 ^ n_251;
assign n_3515 = n_2080 ^ n_254;
assign n_3516 = n_2081 ^ x113;
assign n_3517 = n_2082 ^ n_261;
assign n_3518 = ~n_66 & n_2083;
assign n_3519 = n_2084 ^ n_264;
assign n_3520 = n_2085 ^ x114;
assign n_3521 = ~x62 & ~n_2086;
assign n_3522 = n_2087 ^ x115;
assign n_3523 = n_2088 ^ x115;
assign n_3524 = n_2089 ^ x119;
assign n_3525 = n_2090 ^ x118;
assign n_3526 = ~n_610 & n_2091;
assign n_3527 = x63 & n_2092;
assign n_3528 = n_2093 ^ x121;
assign n_3529 = n_2094 ^ x124;
assign n_3530 = n_2095 ^ n_1984;
assign n_3531 = n_2096 ^ n_298;
assign n_3532 = n_2097 ^ x125;
assign n_3533 = n_1 & ~n_2098;
assign n_3534 = x63 & n_2099;
assign n_3535 = x64 & n_2184;
assign n_3536 = x65 & n_2184;
assign n_3537 = x66 & n_2184;
assign n_3538 = x67 & n_2184;
assign n_3539 = x68 & n_2184;
assign n_3540 = x69 & n_2184;
assign n_3541 = x70 & n_2184;
assign n_3542 = x71 & n_2184;
assign n_3543 = x72 & n_2184;
assign n_3544 = x73 & n_2184;
assign n_3545 = x74 & n_2184;
assign n_3546 = x75 & n_2184;
assign n_3547 = x76 & n_2184;
assign n_3548 = x77 & n_2184;
assign n_3549 = x78 & n_2184;
assign n_3550 = x79 & n_2184;
assign n_3551 = x80 & n_2184;
assign n_3552 = x81 & n_2184;
assign n_3553 = x82 & n_2184;
assign n_3554 = x83 & n_2184;
assign n_3555 = x84 & n_2184;
assign n_3556 = x85 & n_2184;
assign n_3557 = x86 & n_2184;
assign n_3558 = x87 & n_2184;
assign n_3559 = x88 & n_2184;
assign n_3560 = x89 & n_2184;
assign n_3561 = x90 & n_2184;
assign n_3562 = x91 & n_2184;
assign n_3563 = x92 & n_2184;
assign n_3564 = x93 & n_2184;
assign n_3565 = x94 & n_2184;
assign n_3566 = x95 & n_2184;
assign n_3567 = x96 & n_2184;
assign n_3568 = x97 & n_2184;
assign n_3569 = x98 & n_2184;
assign n_3570 = x99 & n_2184;
assign n_3571 = x100 & n_2184;
assign n_3572 = x101 & n_2184;
assign n_3573 = x102 & n_2184;
assign n_3574 = x103 & n_2184;
assign n_3575 = x104 & n_2184;
assign n_3576 = x105 & n_2184;
assign n_3577 = x106 & n_2184;
assign n_3578 = x107 & n_2184;
assign n_3579 = x108 & n_2184;
assign n_3580 = x109 & n_2184;
assign n_3581 = x110 & n_2184;
assign n_3582 = x111 & n_2184;
assign n_3583 = x112 & n_2184;
assign n_3584 = x113 & n_2184;
assign n_3585 = x114 & n_2184;
assign n_3586 = x115 & n_2184;
assign n_3587 = x116 & n_2184;
assign n_3588 = x117 & n_2184;
assign n_3589 = x118 & n_2184;
assign n_3590 = x119 & n_2184;
assign n_3591 = x120 & n_2184;
assign n_3592 = x121 & n_2184;
assign n_3593 = x122 & n_2184;
assign n_3594 = x123 & n_2184;
assign n_3595 = x124 & n_2184;
assign n_3596 = x125 & n_2184;
assign n_3597 = x126 & n_2184;
assign n_3598 = ~x5 ^ ~n_2185;
assign n_3599 = n_2186 ^ n_82;
assign n_3600 = x65 & n_2188;
assign n_3601 = x66 & n_2188;
assign n_3602 = x67 & n_2188;
assign n_3603 = x68 & n_2188;
assign n_3604 = x69 & n_2188;
assign n_3605 = x70 & n_2188;
assign n_3606 = x71 & n_2188;
assign n_3607 = x72 & n_2188;
assign n_3608 = x73 & n_2188;
assign n_3609 = x74 & n_2188;
assign n_3610 = x75 & n_2188;
assign n_3611 = x76 & n_2188;
assign n_3612 = x77 & n_2188;
assign n_3613 = x78 & n_2188;
assign n_3614 = x79 & n_2188;
assign n_3615 = x80 & n_2188;
assign n_3616 = x81 & n_2188;
assign n_3617 = x82 & n_2188;
assign n_3618 = x83 & n_2188;
assign n_3619 = x84 & n_2188;
assign n_3620 = x85 & n_2188;
assign n_3621 = x86 & n_2188;
assign n_3622 = x87 & n_2188;
assign n_3623 = x88 & n_2188;
assign n_3624 = x89 & n_2188;
assign n_3625 = x90 & n_2188;
assign n_3626 = x91 & n_2188;
assign n_3627 = x92 & n_2188;
assign n_3628 = x93 & n_2188;
assign n_3629 = x94 & n_2188;
assign n_3630 = x95 & n_2188;
assign n_3631 = x96 & n_2188;
assign n_3632 = x97 & n_2188;
assign n_3633 = x98 & n_2188;
assign n_3634 = x99 & n_2188;
assign n_3635 = x100 & n_2188;
assign n_3636 = x101 & n_2188;
assign n_3637 = x102 & n_2188;
assign n_3638 = x103 & n_2188;
assign n_3639 = x104 & n_2188;
assign n_3640 = x105 & n_2188;
assign n_3641 = x106 & n_2188;
assign n_3642 = x107 & n_2188;
assign n_3643 = x108 & n_2188;
assign n_3644 = x109 & n_2188;
assign n_3645 = x110 & n_2188;
assign n_3646 = x111 & n_2188;
assign n_3647 = x112 & n_2188;
assign n_3648 = x113 & n_2188;
assign n_3649 = x114 & n_2188;
assign n_3650 = x115 & n_2188;
assign n_3651 = x116 & n_2188;
assign n_3652 = x117 & n_2188;
assign n_3653 = x118 & n_2188;
assign n_3654 = x119 & n_2188;
assign n_3655 = x120 & n_2188;
assign n_3656 = x121 & n_2188;
assign n_3657 = x122 & n_2188;
assign n_3658 = x123 & n_2188;
assign n_3659 = x124 & n_2188;
assign n_3660 = x125 & n_2188;
assign n_3661 = x126 & n_2188;
assign n_3662 = n_2189 ^ n_719;
assign n_3663 = n_2190 ^ x8;
assign n_3664 = n_340 ^ n_2191;
assign n_3665 = n_2255 ^ n_12;
assign n_3666 = x67 & ~n_2255;
assign n_3667 = x68 & ~n_2255;
assign n_3668 = x69 & ~n_2255;
assign n_3669 = x70 & ~n_2255;
assign n_3670 = x71 & ~n_2255;
assign n_3671 = x72 & ~n_2255;
assign n_3672 = x73 & ~n_2255;
assign n_3673 = x74 & ~n_2255;
assign n_3674 = x75 & ~n_2255;
assign n_3675 = x76 & ~n_2255;
assign n_3676 = x77 & ~n_2255;
assign n_3677 = x78 & ~n_2255;
assign n_3678 = x79 & ~n_2255;
assign n_3679 = x80 & ~n_2255;
assign n_3680 = x81 & ~n_2255;
assign n_3681 = x82 & ~n_2255;
assign n_3682 = x83 & ~n_2255;
assign n_3683 = x84 & ~n_2255;
assign n_3684 = x85 & ~n_2255;
assign n_3685 = x86 & ~n_2255;
assign n_3686 = x87 & ~n_2255;
assign n_3687 = x88 & ~n_2255;
assign n_3688 = x89 & ~n_2255;
assign n_3689 = x90 & ~n_2255;
assign n_3690 = x91 & ~n_2255;
assign n_3691 = x92 & ~n_2255;
assign n_3692 = x93 & ~n_2255;
assign n_3693 = x94 & ~n_2255;
assign n_3694 = x95 & ~n_2255;
assign n_3695 = x96 & ~n_2255;
assign n_3696 = x97 & ~n_2255;
assign n_3697 = x98 & ~n_2255;
assign n_3698 = x99 & ~n_2255;
assign n_3699 = x100 & ~n_2255;
assign n_3700 = x101 & ~n_2255;
assign n_3701 = x102 & ~n_2255;
assign n_3702 = x103 & ~n_2255;
assign n_3703 = x104 & ~n_2255;
assign n_3704 = x105 & ~n_2255;
assign n_3705 = x106 & ~n_2255;
assign n_3706 = x107 & ~n_2255;
assign n_3707 = x108 & ~n_2255;
assign n_3708 = x109 & ~n_2255;
assign n_3709 = x110 & ~n_2255;
assign n_3710 = x111 & ~n_2255;
assign n_3711 = x112 & ~n_2255;
assign n_3712 = x113 & ~n_2255;
assign n_3713 = x114 & ~n_2255;
assign n_3714 = x115 & ~n_2255;
assign n_3715 = x116 & ~n_2255;
assign n_3716 = x117 & ~n_2255;
assign n_3717 = x118 & ~n_2255;
assign n_3718 = x119 & ~n_2255;
assign n_3719 = x120 & ~n_2255;
assign n_3720 = x121 & ~n_2255;
assign n_3721 = x122 & ~n_2255;
assign n_3722 = x123 & ~n_2255;
assign n_3723 = x124 & ~n_2255;
assign n_3724 = x125 & ~n_2255;
assign n_3725 = x126 & ~n_2255;
assign n_3726 = x127 & ~n_2255;
assign n_3727 = x65 & n_2258;
assign n_3728 = x66 & n_2258;
assign n_3729 = x67 & n_2258;
assign n_3730 = x68 & n_2258;
assign n_3731 = x69 & n_2258;
assign n_3732 = x70 & n_2258;
assign n_3733 = x71 & n_2258;
assign n_3734 = x72 & n_2258;
assign n_3735 = x73 & n_2258;
assign n_3736 = x74 & n_2258;
assign n_3737 = x75 & n_2258;
assign n_3738 = x76 & n_2258;
assign n_3739 = x77 & n_2258;
assign n_3740 = x78 & n_2258;
assign n_3741 = x79 & n_2258;
assign n_3742 = x80 & n_2258;
assign n_3743 = x81 & n_2258;
assign n_3744 = x82 & n_2258;
assign n_3745 = x83 & n_2258;
assign n_3746 = x84 & n_2258;
assign n_3747 = x85 & n_2258;
assign n_3748 = x86 & n_2258;
assign n_3749 = x87 & n_2258;
assign n_3750 = x88 & n_2258;
assign n_3751 = x89 & n_2258;
assign n_3752 = x90 & n_2258;
assign n_3753 = x91 & n_2258;
assign n_3754 = x92 & n_2258;
assign n_3755 = x93 & n_2258;
assign n_3756 = x94 & n_2258;
assign n_3757 = x95 & n_2258;
assign n_3758 = x96 & n_2258;
assign n_3759 = x97 & n_2258;
assign n_3760 = x98 & n_2258;
assign n_3761 = x99 & n_2258;
assign n_3762 = x100 & n_2258;
assign n_3763 = x101 & n_2258;
assign n_3764 = x102 & n_2258;
assign n_3765 = x103 & n_2258;
assign n_3766 = x104 & n_2258;
assign n_3767 = x105 & n_2258;
assign n_3768 = x106 & n_2258;
assign n_3769 = x107 & n_2258;
assign n_3770 = x108 & n_2258;
assign n_3771 = x109 & n_2258;
assign n_3772 = x110 & n_2258;
assign n_3773 = x111 & n_2258;
assign n_3774 = x112 & n_2258;
assign n_3775 = x113 & n_2258;
assign n_3776 = x114 & n_2258;
assign n_3777 = x115 & n_2258;
assign n_3778 = x116 & n_2258;
assign n_3779 = x117 & n_2258;
assign n_3780 = x118 & n_2258;
assign n_3781 = x119 & n_2258;
assign n_3782 = x120 & n_2258;
assign n_3783 = x121 & n_2258;
assign n_3784 = x122 & n_2258;
assign n_3785 = x123 & n_2258;
assign n_3786 = x124 & n_2258;
assign n_3787 = x125 & n_2258;
assign n_3788 = x126 & n_2258;
assign n_3789 = n_2259 ^ x11;
assign n_3790 = x65 & n_2323;
assign n_3791 = x66 & n_2323;
assign n_3792 = x67 & n_2323;
assign n_3793 = x68 & n_2323;
assign n_3794 = x69 & n_2323;
assign n_3795 = x70 & n_2323;
assign n_3796 = x71 & n_2323;
assign n_3797 = x72 & n_2323;
assign n_3798 = x73 & n_2323;
assign n_3799 = x74 & n_2323;
assign n_3800 = x75 & n_2323;
assign n_3801 = x76 & n_2323;
assign n_3802 = x77 & n_2323;
assign n_3803 = x78 & n_2323;
assign n_3804 = x79 & n_2323;
assign n_3805 = x80 & n_2323;
assign n_3806 = x81 & n_2323;
assign n_3807 = x82 & n_2323;
assign n_3808 = x83 & n_2323;
assign n_3809 = x84 & n_2323;
assign n_3810 = x85 & n_2323;
assign n_3811 = x86 & n_2323;
assign n_3812 = x87 & n_2323;
assign n_3813 = x88 & n_2323;
assign n_3814 = x89 & n_2323;
assign n_3815 = x90 & n_2323;
assign n_3816 = x91 & n_2323;
assign n_3817 = x92 & n_2323;
assign n_3818 = x93 & n_2323;
assign n_3819 = x94 & n_2323;
assign n_3820 = x95 & n_2323;
assign n_3821 = x96 & n_2323;
assign n_3822 = x97 & n_2323;
assign n_3823 = x98 & n_2323;
assign n_3824 = x99 & n_2323;
assign n_3825 = x100 & n_2323;
assign n_3826 = x101 & n_2323;
assign n_3827 = x102 & n_2323;
assign n_3828 = x103 & n_2323;
assign n_3829 = x104 & n_2323;
assign n_3830 = x105 & n_2323;
assign n_3831 = x106 & n_2323;
assign n_3832 = x107 & n_2323;
assign n_3833 = x108 & n_2323;
assign n_3834 = x109 & n_2323;
assign n_3835 = x110 & n_2323;
assign n_3836 = x111 & n_2323;
assign n_3837 = x112 & n_2323;
assign n_3838 = x113 & n_2323;
assign n_3839 = x114 & n_2323;
assign n_3840 = x115 & n_2323;
assign n_3841 = x116 & n_2323;
assign n_3842 = x117 & n_2323;
assign n_3843 = x118 & n_2323;
assign n_3844 = x119 & n_2323;
assign n_3845 = x120 & n_2323;
assign n_3846 = x121 & n_2323;
assign n_3847 = x122 & n_2323;
assign n_3848 = x123 & n_2323;
assign n_3849 = x124 & n_2323;
assign n_3850 = x125 & n_2323;
assign n_3851 = x126 & n_2323;
assign n_3852 = ~x14 ^ ~n_2324;
assign n_3853 = n_355 ^ n_2325;
assign n_3854 = x17 & n_2390;
assign n_3855 = x65 & n_2390;
assign n_3856 = x66 & n_2390;
assign n_3857 = x67 & n_2390;
assign n_3858 = x68 & n_2390;
assign n_3859 = x69 & n_2390;
assign n_3860 = x70 & n_2390;
assign n_3861 = x71 & n_2390;
assign n_3862 = x72 & n_2390;
assign n_3863 = x73 & n_2390;
assign n_3864 = x74 & n_2390;
assign n_3865 = x75 & n_2390;
assign n_3866 = x76 & n_2390;
assign n_3867 = x77 & n_2390;
assign n_3868 = x78 & n_2390;
assign n_3869 = x79 & n_2390;
assign n_3870 = x80 & n_2390;
assign n_3871 = x81 & n_2390;
assign n_3872 = x82 & n_2390;
assign n_3873 = x83 & n_2390;
assign n_3874 = x84 & n_2390;
assign n_3875 = x85 & n_2390;
assign n_3876 = x86 & n_2390;
assign n_3877 = x87 & n_2390;
assign n_3878 = x88 & n_2390;
assign n_3879 = x89 & n_2390;
assign n_3880 = x90 & n_2390;
assign n_3881 = x91 & n_2390;
assign n_3882 = x92 & n_2390;
assign n_3883 = x93 & n_2390;
assign n_3884 = x94 & n_2390;
assign n_3885 = x95 & n_2390;
assign n_3886 = x96 & n_2390;
assign n_3887 = x97 & n_2390;
assign n_3888 = x98 & n_2390;
assign n_3889 = x99 & n_2390;
assign n_3890 = x100 & n_2390;
assign n_3891 = x101 & n_2390;
assign n_3892 = x102 & n_2390;
assign n_3893 = x103 & n_2390;
assign n_3894 = x104 & n_2390;
assign n_3895 = x105 & n_2390;
assign n_3896 = x106 & n_2390;
assign n_3897 = x107 & n_2390;
assign n_3898 = x108 & n_2390;
assign n_3899 = x109 & n_2390;
assign n_3900 = x110 & n_2390;
assign n_3901 = x111 & n_2390;
assign n_3902 = x112 & n_2390;
assign n_3903 = x113 & n_2390;
assign n_3904 = x114 & n_2390;
assign n_3905 = x115 & n_2390;
assign n_3906 = x116 & n_2390;
assign n_3907 = x117 & n_2390;
assign n_3908 = x118 & n_2390;
assign n_3909 = x119 & n_2390;
assign n_3910 = x120 & n_2390;
assign n_3911 = x121 & n_2390;
assign n_3912 = x122 & n_2390;
assign n_3913 = x123 & n_2390;
assign n_3914 = x124 & n_2390;
assign n_3915 = x125 & n_2390;
assign n_3916 = x126 & n_2390;
assign n_3917 = ~x17 ^ ~n_2391;
assign n_3918 = n_360 ^ n_2392;
assign n_3919 = x20 & n_2457;
assign n_3920 = x65 & n_2457;
assign n_3921 = x66 & n_2457;
assign n_3922 = x67 & n_2457;
assign n_3923 = x68 & n_2457;
assign n_3924 = x69 & n_2457;
assign n_3925 = x70 & n_2457;
assign n_3926 = x71 & n_2457;
assign n_3927 = x72 & n_2457;
assign n_3928 = x73 & n_2457;
assign n_3929 = x74 & n_2457;
assign n_3930 = x75 & n_2457;
assign n_3931 = x76 & n_2457;
assign n_3932 = x77 & n_2457;
assign n_3933 = x78 & n_2457;
assign n_3934 = x79 & n_2457;
assign n_3935 = x80 & n_2457;
assign n_3936 = x81 & n_2457;
assign n_3937 = x82 & n_2457;
assign n_3938 = x83 & n_2457;
assign n_3939 = x84 & n_2457;
assign n_3940 = x85 & n_2457;
assign n_3941 = x86 & n_2457;
assign n_3942 = x87 & n_2457;
assign n_3943 = x88 & n_2457;
assign n_3944 = x89 & n_2457;
assign n_3945 = x90 & n_2457;
assign n_3946 = x91 & n_2457;
assign n_3947 = x92 & n_2457;
assign n_3948 = x93 & n_2457;
assign n_3949 = x94 & n_2457;
assign n_3950 = x95 & n_2457;
assign n_3951 = x96 & n_2457;
assign n_3952 = x97 & n_2457;
assign n_3953 = x98 & n_2457;
assign n_3954 = x99 & n_2457;
assign n_3955 = x100 & n_2457;
assign n_3956 = x101 & n_2457;
assign n_3957 = x102 & n_2457;
assign n_3958 = x103 & n_2457;
assign n_3959 = x104 & n_2457;
assign n_3960 = x105 & n_2457;
assign n_3961 = x106 & n_2457;
assign n_3962 = x107 & n_2457;
assign n_3963 = x108 & n_2457;
assign n_3964 = x109 & n_2457;
assign n_3965 = x110 & n_2457;
assign n_3966 = x111 & n_2457;
assign n_3967 = x112 & n_2457;
assign n_3968 = x113 & n_2457;
assign n_3969 = x114 & n_2457;
assign n_3970 = x115 & n_2457;
assign n_3971 = x116 & n_2457;
assign n_3972 = x117 & n_2457;
assign n_3973 = x118 & n_2457;
assign n_3974 = x119 & n_2457;
assign n_3975 = x120 & n_2457;
assign n_3976 = x121 & n_2457;
assign n_3977 = x122 & n_2457;
assign n_3978 = x123 & n_2457;
assign n_3979 = x124 & n_2457;
assign n_3980 = x125 & n_2457;
assign n_3981 = x126 & n_2457;
assign n_3982 = ~x20 ^ ~n_2458;
assign n_3983 = n_366 ^ n_2459;
assign n_3984 = x23 & n_2524;
assign n_3985 = x65 & n_2524;
assign n_3986 = x66 & n_2524;
assign n_3987 = x67 & n_2524;
assign n_3988 = x68 & n_2524;
assign n_3989 = x69 & n_2524;
assign n_3990 = x70 & n_2524;
assign n_3991 = x71 & n_2524;
assign n_3992 = x72 & n_2524;
assign n_3993 = x73 & n_2524;
assign n_3994 = x74 & n_2524;
assign n_3995 = x75 & n_2524;
assign n_3996 = x76 & n_2524;
assign n_3997 = x77 & n_2524;
assign n_3998 = x78 & n_2524;
assign n_3999 = x79 & n_2524;
assign n_4000 = x80 & n_2524;
assign n_4001 = x81 & n_2524;
assign n_4002 = x82 & n_2524;
assign n_4003 = x83 & n_2524;
assign n_4004 = x84 & n_2524;
assign n_4005 = x85 & n_2524;
assign n_4006 = x86 & n_2524;
assign n_4007 = x87 & n_2524;
assign n_4008 = x88 & n_2524;
assign n_4009 = x89 & n_2524;
assign n_4010 = x90 & n_2524;
assign n_4011 = x91 & n_2524;
assign n_4012 = x92 & n_2524;
assign n_4013 = x93 & n_2524;
assign n_4014 = x94 & n_2524;
assign n_4015 = x95 & n_2524;
assign n_4016 = x96 & n_2524;
assign n_4017 = x97 & n_2524;
assign n_4018 = x98 & n_2524;
assign n_4019 = x99 & n_2524;
assign n_4020 = x100 & n_2524;
assign n_4021 = x101 & n_2524;
assign n_4022 = x102 & n_2524;
assign n_4023 = x103 & n_2524;
assign n_4024 = x104 & n_2524;
assign n_4025 = x105 & n_2524;
assign n_4026 = x106 & n_2524;
assign n_4027 = x107 & n_2524;
assign n_4028 = x108 & n_2524;
assign n_4029 = x109 & n_2524;
assign n_4030 = x110 & n_2524;
assign n_4031 = x111 & n_2524;
assign n_4032 = x112 & n_2524;
assign n_4033 = x113 & n_2524;
assign n_4034 = x114 & n_2524;
assign n_4035 = x115 & n_2524;
assign n_4036 = x116 & n_2524;
assign n_4037 = x117 & n_2524;
assign n_4038 = x118 & n_2524;
assign n_4039 = x119 & n_2524;
assign n_4040 = x120 & n_2524;
assign n_4041 = x121 & n_2524;
assign n_4042 = x122 & n_2524;
assign n_4043 = x123 & n_2524;
assign n_4044 = x124 & n_2524;
assign n_4045 = x125 & n_2524;
assign n_4046 = x126 & n_2524;
assign n_4047 = ~x23 ^ ~n_2525;
assign n_4048 = n_372 ^ n_2526;
assign n_4049 = x64 & n_2590;
assign n_4050 = x65 & n_2590;
assign n_4051 = x66 & n_2590;
assign n_4052 = x67 & n_2590;
assign n_4053 = x68 & n_2590;
assign n_4054 = x69 & n_2590;
assign n_4055 = x70 & n_2590;
assign n_4056 = x71 & n_2590;
assign n_4057 = x72 & n_2590;
assign n_4058 = x73 & n_2590;
assign n_4059 = x74 & n_2590;
assign n_4060 = x75 & n_2590;
assign n_4061 = x76 & n_2590;
assign n_4062 = x77 & n_2590;
assign n_4063 = x78 & n_2590;
assign n_4064 = x79 & n_2590;
assign n_4065 = x80 & n_2590;
assign n_4066 = x81 & n_2590;
assign n_4067 = x82 & n_2590;
assign n_4068 = x83 & n_2590;
assign n_4069 = x84 & n_2590;
assign n_4070 = x85 & n_2590;
assign n_4071 = x86 & n_2590;
assign n_4072 = x87 & n_2590;
assign n_4073 = x88 & n_2590;
assign n_4074 = x89 & n_2590;
assign n_4075 = x90 & n_2590;
assign n_4076 = x91 & n_2590;
assign n_4077 = x92 & n_2590;
assign n_4078 = x93 & n_2590;
assign n_4079 = x94 & n_2590;
assign n_4080 = x95 & n_2590;
assign n_4081 = x96 & n_2590;
assign n_4082 = x97 & n_2590;
assign n_4083 = x98 & n_2590;
assign n_4084 = x99 & n_2590;
assign n_4085 = x100 & n_2590;
assign n_4086 = x101 & n_2590;
assign n_4087 = x102 & n_2590;
assign n_4088 = x103 & n_2590;
assign n_4089 = x104 & n_2590;
assign n_4090 = x105 & n_2590;
assign n_4091 = x106 & n_2590;
assign n_4092 = x107 & n_2590;
assign n_4093 = x108 & n_2590;
assign n_4094 = x109 & n_2590;
assign n_4095 = x110 & n_2590;
assign n_4096 = x111 & n_2590;
assign n_4097 = x112 & n_2590;
assign n_4098 = x113 & n_2590;
assign n_4099 = x114 & n_2590;
assign n_4100 = x115 & n_2590;
assign n_4101 = x116 & n_2590;
assign n_4102 = x117 & n_2590;
assign n_4103 = x118 & n_2590;
assign n_4104 = x119 & n_2590;
assign n_4105 = x120 & n_2590;
assign n_4106 = x121 & n_2590;
assign n_4107 = x122 & n_2590;
assign n_4108 = x123 & n_2590;
assign n_4109 = x124 & n_2590;
assign n_4110 = x125 & n_2590;
assign n_4111 = x126 & n_2590;
assign n_4112 = x127 & n_2590;
assign n_4113 = x65 & n_2655;
assign n_4114 = x66 & n_2655;
assign n_4115 = x67 & n_2655;
assign n_4116 = x68 & n_2655;
assign n_4117 = x69 & n_2655;
assign n_4118 = x70 & n_2655;
assign n_4119 = x71 & n_2655;
assign n_4120 = x72 & n_2655;
assign n_4121 = x73 & n_2655;
assign n_4122 = x74 & n_2655;
assign n_4123 = x75 & n_2655;
assign n_4124 = x76 & n_2655;
assign n_4125 = x77 & n_2655;
assign n_4126 = x78 & n_2655;
assign n_4127 = x79 & n_2655;
assign n_4128 = x80 & n_2655;
assign n_4129 = x81 & n_2655;
assign n_4130 = x82 & n_2655;
assign n_4131 = x83 & n_2655;
assign n_4132 = x84 & n_2655;
assign n_4133 = x85 & n_2655;
assign n_4134 = x86 & n_2655;
assign n_4135 = x87 & n_2655;
assign n_4136 = x88 & n_2655;
assign n_4137 = x89 & n_2655;
assign n_4138 = x90 & n_2655;
assign n_4139 = x91 & n_2655;
assign n_4140 = x92 & n_2655;
assign n_4141 = x93 & n_2655;
assign n_4142 = x94 & n_2655;
assign n_4143 = x95 & n_2655;
assign n_4144 = x96 & n_2655;
assign n_4145 = x97 & n_2655;
assign n_4146 = x98 & n_2655;
assign n_4147 = x99 & n_2655;
assign n_4148 = x100 & n_2655;
assign n_4149 = x101 & n_2655;
assign n_4150 = x102 & n_2655;
assign n_4151 = x103 & n_2655;
assign n_4152 = x104 & n_2655;
assign n_4153 = x105 & n_2655;
assign n_4154 = x106 & n_2655;
assign n_4155 = x107 & n_2655;
assign n_4156 = x108 & n_2655;
assign n_4157 = x109 & n_2655;
assign n_4158 = x110 & n_2655;
assign n_4159 = x111 & n_2655;
assign n_4160 = x112 & n_2655;
assign n_4161 = x113 & n_2655;
assign n_4162 = x114 & n_2655;
assign n_4163 = x115 & n_2655;
assign n_4164 = x116 & n_2655;
assign n_4165 = x117 & n_2655;
assign n_4166 = x118 & n_2655;
assign n_4167 = x119 & n_2655;
assign n_4168 = x120 & n_2655;
assign n_4169 = x121 & n_2655;
assign n_4170 = x122 & n_2655;
assign n_4171 = x123 & n_2655;
assign n_4172 = x124 & n_2655;
assign n_4173 = x125 & n_2655;
assign n_4174 = x126 & n_2655;
assign n_4175 = ~x29 ^ ~n_2656;
assign n_4176 = n_384 ^ n_2657;
assign n_4177 = x65 & n_2722;
assign n_4178 = x66 & n_2722;
assign n_4179 = x67 & n_2722;
assign n_4180 = x68 & n_2722;
assign n_4181 = x69 & n_2722;
assign n_4182 = x70 & n_2722;
assign n_4183 = x71 & n_2722;
assign n_4184 = x72 & n_2722;
assign n_4185 = x73 & n_2722;
assign n_4186 = x74 & n_2722;
assign n_4187 = x75 & n_2722;
assign n_4188 = x76 & n_2722;
assign n_4189 = x77 & n_2722;
assign n_4190 = x78 & n_2722;
assign n_4191 = x79 & n_2722;
assign n_4192 = x80 & n_2722;
assign n_4193 = x81 & n_2722;
assign n_4194 = x82 & n_2722;
assign n_4195 = x83 & n_2722;
assign n_4196 = x84 & n_2722;
assign n_4197 = x85 & n_2722;
assign n_4198 = x86 & n_2722;
assign n_4199 = x87 & n_2722;
assign n_4200 = x88 & n_2722;
assign n_4201 = x89 & n_2722;
assign n_4202 = x90 & n_2722;
assign n_4203 = x91 & n_2722;
assign n_4204 = x92 & n_2722;
assign n_4205 = x93 & n_2722;
assign n_4206 = x94 & n_2722;
assign n_4207 = x95 & n_2722;
assign n_4208 = x96 & n_2722;
assign n_4209 = x97 & n_2722;
assign n_4210 = x98 & n_2722;
assign n_4211 = x99 & n_2722;
assign n_4212 = x100 & n_2722;
assign n_4213 = x101 & n_2722;
assign n_4214 = x102 & n_2722;
assign n_4215 = x103 & n_2722;
assign n_4216 = x104 & n_2722;
assign n_4217 = x105 & n_2722;
assign n_4218 = x106 & n_2722;
assign n_4219 = x107 & n_2722;
assign n_4220 = x108 & n_2722;
assign n_4221 = x109 & n_2722;
assign n_4222 = x110 & n_2722;
assign n_4223 = x111 & n_2722;
assign n_4224 = x112 & n_2722;
assign n_4225 = x113 & n_2722;
assign n_4226 = x114 & n_2722;
assign n_4227 = x115 & n_2722;
assign n_4228 = x116 & n_2722;
assign n_4229 = x117 & n_2722;
assign n_4230 = x118 & n_2722;
assign n_4231 = x119 & n_2722;
assign n_4232 = x120 & n_2722;
assign n_4233 = x121 & n_2722;
assign n_4234 = x122 & n_2722;
assign n_4235 = x123 & n_2722;
assign n_4236 = x124 & n_2722;
assign n_4237 = x125 & n_2722;
assign n_4238 = x126 & n_2722;
assign n_4239 = x64 & n_2723;
assign n_4240 = n_2724 ^ x32;
assign n_4241 = n_390 ^ n_2725;
assign n_4242 = x35 & n_2790;
assign n_4243 = x65 & n_2790;
assign n_4244 = x66 & n_2790;
assign n_4245 = x67 & n_2790;
assign n_4246 = x68 & n_2790;
assign n_4247 = x69 & n_2790;
assign n_4248 = x70 & n_2790;
assign n_4249 = x71 & n_2790;
assign n_4250 = x72 & n_2790;
assign n_4251 = x73 & n_2790;
assign n_4252 = x74 & n_2790;
assign n_4253 = x75 & n_2790;
assign n_4254 = x76 & n_2790;
assign n_4255 = x77 & n_2790;
assign n_4256 = x78 & n_2790;
assign n_4257 = x79 & n_2790;
assign n_4258 = x80 & n_2790;
assign n_4259 = x81 & n_2790;
assign n_4260 = x82 & n_2790;
assign n_4261 = x83 & n_2790;
assign n_4262 = x84 & n_2790;
assign n_4263 = x85 & n_2790;
assign n_4264 = x86 & n_2790;
assign n_4265 = x87 & n_2790;
assign n_4266 = x88 & n_2790;
assign n_4267 = x89 & n_2790;
assign n_4268 = x90 & n_2790;
assign n_4269 = x91 & n_2790;
assign n_4270 = x92 & n_2790;
assign n_4271 = x93 & n_2790;
assign n_4272 = x94 & n_2790;
assign n_4273 = x95 & n_2790;
assign n_4274 = x96 & n_2790;
assign n_4275 = x97 & n_2790;
assign n_4276 = x98 & n_2790;
assign n_4277 = x99 & n_2790;
assign n_4278 = x100 & n_2790;
assign n_4279 = x101 & n_2790;
assign n_4280 = x102 & n_2790;
assign n_4281 = x103 & n_2790;
assign n_4282 = x104 & n_2790;
assign n_4283 = x105 & n_2790;
assign n_4284 = x106 & n_2790;
assign n_4285 = x107 & n_2790;
assign n_4286 = x108 & n_2790;
assign n_4287 = x109 & n_2790;
assign n_4288 = x110 & n_2790;
assign n_4289 = x111 & n_2790;
assign n_4290 = x112 & n_2790;
assign n_4291 = x113 & n_2790;
assign n_4292 = x114 & n_2790;
assign n_4293 = x115 & n_2790;
assign n_4294 = x116 & n_2790;
assign n_4295 = x117 & n_2790;
assign n_4296 = x118 & n_2790;
assign n_4297 = x119 & n_2790;
assign n_4298 = x120 & n_2790;
assign n_4299 = x121 & n_2790;
assign n_4300 = x122 & n_2790;
assign n_4301 = x123 & n_2790;
assign n_4302 = x124 & n_2790;
assign n_4303 = x125 & n_2790;
assign n_4304 = x126 & n_2790;
assign n_4305 = ~x35 ^ ~n_2791;
assign n_4306 = n_397 ^ n_2792;
assign n_4307 = x38 & n_2857;
assign n_4308 = x65 & n_2857;
assign n_4309 = x66 & n_2857;
assign n_4310 = x67 & n_2857;
assign n_4311 = x68 & n_2857;
assign n_4312 = x69 & n_2857;
assign n_4313 = x70 & n_2857;
assign n_4314 = x71 & n_2857;
assign n_4315 = x72 & n_2857;
assign n_4316 = x73 & n_2857;
assign n_4317 = x74 & n_2857;
assign n_4318 = x75 & n_2857;
assign n_4319 = x76 & n_2857;
assign n_4320 = x77 & n_2857;
assign n_4321 = x78 & n_2857;
assign n_4322 = x79 & n_2857;
assign n_4323 = x80 & n_2857;
assign n_4324 = x81 & n_2857;
assign n_4325 = x82 & n_2857;
assign n_4326 = x83 & n_2857;
assign n_4327 = x84 & n_2857;
assign n_4328 = x85 & n_2857;
assign n_4329 = x86 & n_2857;
assign n_4330 = x87 & n_2857;
assign n_4331 = x88 & n_2857;
assign n_4332 = x89 & n_2857;
assign n_4333 = x90 & n_2857;
assign n_4334 = x91 & n_2857;
assign n_4335 = x92 & n_2857;
assign n_4336 = x93 & n_2857;
assign n_4337 = x94 & n_2857;
assign n_4338 = x95 & n_2857;
assign n_4339 = x96 & n_2857;
assign n_4340 = x97 & n_2857;
assign n_4341 = x98 & n_2857;
assign n_4342 = x99 & n_2857;
assign n_4343 = x100 & n_2857;
assign n_4344 = x101 & n_2857;
assign n_4345 = x102 & n_2857;
assign n_4346 = x103 & n_2857;
assign n_4347 = x104 & n_2857;
assign n_4348 = x105 & n_2857;
assign n_4349 = x106 & n_2857;
assign n_4350 = x107 & n_2857;
assign n_4351 = x108 & n_2857;
assign n_4352 = x109 & n_2857;
assign n_4353 = x110 & n_2857;
assign n_4354 = x111 & n_2857;
assign n_4355 = x112 & n_2857;
assign n_4356 = x113 & n_2857;
assign n_4357 = x114 & n_2857;
assign n_4358 = x115 & n_2857;
assign n_4359 = x116 & n_2857;
assign n_4360 = x117 & n_2857;
assign n_4361 = x118 & n_2857;
assign n_4362 = x119 & n_2857;
assign n_4363 = x120 & n_2857;
assign n_4364 = x121 & n_2857;
assign n_4365 = x122 & n_2857;
assign n_4366 = x123 & n_2857;
assign n_4367 = x124 & n_2857;
assign n_4368 = x125 & n_2857;
assign n_4369 = x126 & n_2857;
assign n_4370 = ~x38 ^ ~n_2858;
assign n_4371 = n_403 ^ n_2859;
assign n_4372 = n_2860 ^ n_407;
assign n_4373 = ~n_42 & ~n_2861;
assign n_4374 = x64 & n_2925;
assign n_4375 = x65 & n_2925;
assign n_4376 = x66 & n_2925;
assign n_4377 = x67 & n_2925;
assign n_4378 = x68 & n_2925;
assign n_4379 = x69 & n_2925;
assign n_4380 = x70 & n_2925;
assign n_4381 = x71 & n_2925;
assign n_4382 = x72 & n_2925;
assign n_4383 = x73 & n_2925;
assign n_4384 = x74 & n_2925;
assign n_4385 = x75 & n_2925;
assign n_4386 = x76 & n_2925;
assign n_4387 = x77 & n_2925;
assign n_4388 = x78 & n_2925;
assign n_4389 = x79 & n_2925;
assign n_4390 = x80 & n_2925;
assign n_4391 = x81 & n_2925;
assign n_4392 = x82 & n_2925;
assign n_4393 = x83 & n_2925;
assign n_4394 = x84 & n_2925;
assign n_4395 = x85 & n_2925;
assign n_4396 = x86 & n_2925;
assign n_4397 = x87 & n_2925;
assign n_4398 = x88 & n_2925;
assign n_4399 = x89 & n_2925;
assign n_4400 = x90 & n_2925;
assign n_4401 = x91 & n_2925;
assign n_4402 = x92 & n_2925;
assign n_4403 = x93 & n_2925;
assign n_4404 = x94 & n_2925;
assign n_4405 = x95 & n_2925;
assign n_4406 = x96 & n_2925;
assign n_4407 = x97 & n_2925;
assign n_4408 = x98 & n_2925;
assign n_4409 = x99 & n_2925;
assign n_4410 = x100 & n_2925;
assign n_4411 = x101 & n_2925;
assign n_4412 = x102 & n_2925;
assign n_4413 = x103 & n_2925;
assign n_4414 = x104 & n_2925;
assign n_4415 = x105 & n_2925;
assign n_4416 = x106 & n_2925;
assign n_4417 = x107 & n_2925;
assign n_4418 = x108 & n_2925;
assign n_4419 = x109 & n_2925;
assign n_4420 = x110 & n_2925;
assign n_4421 = x111 & n_2925;
assign n_4422 = x112 & n_2925;
assign n_4423 = x113 & n_2925;
assign n_4424 = x114 & n_2925;
assign n_4425 = x115 & n_2925;
assign n_4426 = x116 & n_2925;
assign n_4427 = x117 & n_2925;
assign n_4428 = x118 & n_2925;
assign n_4429 = x119 & n_2925;
assign n_4430 = x120 & n_2925;
assign n_4431 = x121 & n_2925;
assign n_4432 = x122 & n_2925;
assign n_4433 = x123 & n_2925;
assign n_4434 = x124 & n_2925;
assign n_4435 = x125 & n_2925;
assign n_4436 = x126 & n_2925;
assign n_4437 = x127 & n_2925;
assign n_4438 = x44 & n_2991;
assign n_4439 = x65 & n_2991;
assign n_4440 = x66 & n_2991;
assign n_4441 = x67 & n_2991;
assign n_4442 = x68 & n_2991;
assign n_4443 = x69 & n_2991;
assign n_4444 = x70 & n_2991;
assign n_4445 = x71 & n_2991;
assign n_4446 = x72 & n_2991;
assign n_4447 = x73 & n_2991;
assign n_4448 = x74 & n_2991;
assign n_4449 = x75 & n_2991;
assign n_4450 = x76 & n_2991;
assign n_4451 = x77 & n_2991;
assign n_4452 = x78 & n_2991;
assign n_4453 = x79 & n_2991;
assign n_4454 = x80 & n_2991;
assign n_4455 = x81 & n_2991;
assign n_4456 = x82 & n_2991;
assign n_4457 = x83 & n_2991;
assign n_4458 = x84 & n_2991;
assign n_4459 = x85 & n_2991;
assign n_4460 = x86 & n_2991;
assign n_4461 = x87 & n_2991;
assign n_4462 = x88 & n_2991;
assign n_4463 = x89 & n_2991;
assign n_4464 = x90 & n_2991;
assign n_4465 = x91 & n_2991;
assign n_4466 = x92 & n_2991;
assign n_4467 = x93 & n_2991;
assign n_4468 = x94 & n_2991;
assign n_4469 = x95 & n_2991;
assign n_4470 = x96 & n_2991;
assign n_4471 = x97 & n_2991;
assign n_4472 = x98 & n_2991;
assign n_4473 = x99 & n_2991;
assign n_4474 = x100 & n_2991;
assign n_4475 = x101 & n_2991;
assign n_4476 = x102 & n_2991;
assign n_4477 = x103 & n_2991;
assign n_4478 = x104 & n_2991;
assign n_4479 = x105 & n_2991;
assign n_4480 = x106 & n_2991;
assign n_4481 = x107 & n_2991;
assign n_4482 = x108 & n_2991;
assign n_4483 = x109 & n_2991;
assign n_4484 = x110 & n_2991;
assign n_4485 = x111 & n_2991;
assign n_4486 = x112 & n_2991;
assign n_4487 = x113 & n_2991;
assign n_4488 = x114 & n_2991;
assign n_4489 = x115 & n_2991;
assign n_4490 = x116 & n_2991;
assign n_4491 = x117 & n_2991;
assign n_4492 = x118 & n_2991;
assign n_4493 = x119 & n_2991;
assign n_4494 = x120 & n_2991;
assign n_4495 = x121 & n_2991;
assign n_4496 = x122 & n_2991;
assign n_4497 = x123 & n_2991;
assign n_4498 = x124 & n_2991;
assign n_4499 = x125 & n_2991;
assign n_4500 = x126 & n_2991;
assign n_4501 = ~x44 ^ ~n_2992;
assign n_4502 = n_416 ^ n_2993;
assign n_4503 = x47 & n_2995;
assign n_4504 = x65 & n_2995;
assign n_4505 = x66 & n_2995;
assign n_4506 = x67 & n_2995;
assign n_4507 = x68 & n_2995;
assign n_4508 = x69 & n_2995;
assign n_4509 = x70 & n_2995;
assign n_4510 = x71 & n_2995;
assign n_4511 = x72 & n_2995;
assign n_4512 = x73 & n_2995;
assign n_4513 = x74 & n_2995;
assign n_4514 = x75 & n_2995;
assign n_4515 = x76 & n_2995;
assign n_4516 = x77 & n_2995;
assign n_4517 = x78 & n_2995;
assign n_4518 = x79 & n_2995;
assign n_4519 = x80 & n_2995;
assign n_4520 = x81 & n_2995;
assign n_4521 = x82 & n_2995;
assign n_4522 = x83 & n_2995;
assign n_4523 = x84 & n_2995;
assign n_4524 = x85 & n_2995;
assign n_4525 = x86 & n_2995;
assign n_4526 = x87 & n_2995;
assign n_4527 = x88 & n_2995;
assign n_4528 = x89 & n_2995;
assign n_4529 = x90 & n_2995;
assign n_4530 = x91 & n_2995;
assign n_4531 = x92 & n_2995;
assign n_4532 = x93 & n_2995;
assign n_4533 = x94 & n_2995;
assign n_4534 = x95 & n_2995;
assign n_4535 = x96 & n_2995;
assign n_4536 = x97 & n_2995;
assign n_4537 = x98 & n_2995;
assign n_4538 = x99 & n_2995;
assign n_4539 = x100 & n_2995;
assign n_4540 = x101 & n_2995;
assign n_4541 = x102 & n_2995;
assign n_4542 = x103 & n_2995;
assign n_4543 = x104 & n_2995;
assign n_4544 = x105 & n_2995;
assign n_4545 = x106 & n_2995;
assign n_4546 = x107 & n_2995;
assign n_4547 = x108 & n_2995;
assign n_4548 = x109 & n_2995;
assign n_4549 = x110 & n_2995;
assign n_4550 = x111 & n_2995;
assign n_4551 = x112 & n_2995;
assign n_4552 = x113 & n_2995;
assign n_4553 = x114 & n_2995;
assign n_4554 = x115 & n_2995;
assign n_4555 = x116 & n_2995;
assign n_4556 = x117 & n_2995;
assign n_4557 = x118 & n_2995;
assign n_4558 = x119 & n_2995;
assign n_4559 = x120 & n_2995;
assign n_4560 = x121 & n_2995;
assign n_4561 = x122 & n_2995;
assign n_4562 = x123 & n_2995;
assign n_4563 = x124 & n_2995;
assign n_4564 = x125 & n_2995;
assign n_4565 = x126 & n_2995;
assign n_4566 = ~x47 ^ ~n_2996;
assign n_4567 = n_423 ^ n_3061;
assign n_4568 = x65 & n_3126;
assign n_4569 = x66 & n_3126;
assign n_4570 = x67 & n_3126;
assign n_4571 = x68 & n_3126;
assign n_4572 = x69 & n_3126;
assign n_4573 = x70 & n_3126;
assign n_4574 = x71 & n_3126;
assign n_4575 = x72 & n_3126;
assign n_4576 = x73 & n_3126;
assign n_4577 = x74 & n_3126;
assign n_4578 = x75 & n_3126;
assign n_4579 = x76 & n_3126;
assign n_4580 = x77 & n_3126;
assign n_4581 = x78 & n_3126;
assign n_4582 = x79 & n_3126;
assign n_4583 = x80 & n_3126;
assign n_4584 = x81 & n_3126;
assign n_4585 = x82 & n_3126;
assign n_4586 = x83 & n_3126;
assign n_4587 = x84 & n_3126;
assign n_4588 = x85 & n_3126;
assign n_4589 = x86 & n_3126;
assign n_4590 = x87 & n_3126;
assign n_4591 = x88 & n_3126;
assign n_4592 = x89 & n_3126;
assign n_4593 = x90 & n_3126;
assign n_4594 = x91 & n_3126;
assign n_4595 = x92 & n_3126;
assign n_4596 = x93 & n_3126;
assign n_4597 = x94 & n_3126;
assign n_4598 = x95 & n_3126;
assign n_4599 = x96 & n_3126;
assign n_4600 = x97 & n_3126;
assign n_4601 = x98 & n_3126;
assign n_4602 = x99 & n_3126;
assign n_4603 = x100 & n_3126;
assign n_4604 = x101 & n_3126;
assign n_4605 = x102 & n_3126;
assign n_4606 = x103 & n_3126;
assign n_4607 = x104 & n_3126;
assign n_4608 = x105 & n_3126;
assign n_4609 = x106 & n_3126;
assign n_4610 = x107 & n_3126;
assign n_4611 = x108 & n_3126;
assign n_4612 = x109 & n_3126;
assign n_4613 = x110 & n_3126;
assign n_4614 = x111 & n_3126;
assign n_4615 = x112 & n_3126;
assign n_4616 = x113 & n_3126;
assign n_4617 = x114 & n_3126;
assign n_4618 = x115 & n_3126;
assign n_4619 = x116 & n_3126;
assign n_4620 = x117 & n_3126;
assign n_4621 = x118 & n_3126;
assign n_4622 = x119 & n_3126;
assign n_4623 = x120 & n_3126;
assign n_4624 = x121 & n_3126;
assign n_4625 = x122 & n_3126;
assign n_4626 = x123 & n_3126;
assign n_4627 = x124 & n_3126;
assign n_4628 = x125 & n_3126;
assign n_4629 = x126 & n_3126;
assign n_4630 = ~x50 ^ ~n_3127;
assign n_4631 = n_428 ^ n_3128;
assign n_4632 = x52 & n_3130;
assign n_4633 = x65 & n_3130;
assign n_4634 = x66 & n_3130;
assign n_4635 = x67 & n_3130;
assign n_4636 = x68 & n_3130;
assign n_4637 = x69 & n_3130;
assign n_4638 = x70 & n_3130;
assign n_4639 = x71 & n_3130;
assign n_4640 = x72 & n_3130;
assign n_4641 = x73 & n_3130;
assign n_4642 = x74 & n_3130;
assign n_4643 = x75 & n_3130;
assign n_4644 = x76 & n_3130;
assign n_4645 = x77 & n_3130;
assign n_4646 = x78 & n_3130;
assign n_4647 = x79 & n_3130;
assign n_4648 = x80 & n_3130;
assign n_4649 = x81 & n_3130;
assign n_4650 = x82 & n_3130;
assign n_4651 = x83 & n_3130;
assign n_4652 = x84 & n_3130;
assign n_4653 = x85 & n_3130;
assign n_4654 = x86 & n_3130;
assign n_4655 = x87 & n_3130;
assign n_4656 = x88 & n_3130;
assign n_4657 = x89 & n_3130;
assign n_4658 = x90 & n_3130;
assign n_4659 = x91 & n_3130;
assign n_4660 = x92 & n_3130;
assign n_4661 = x93 & n_3130;
assign n_4662 = x94 & n_3130;
assign n_4663 = x95 & n_3130;
assign n_4664 = x96 & n_3130;
assign n_4665 = x97 & n_3130;
assign n_4666 = x98 & n_3130;
assign n_4667 = x99 & n_3130;
assign n_4668 = x100 & n_3130;
assign n_4669 = x101 & n_3130;
assign n_4670 = x102 & n_3130;
assign n_4671 = x103 & n_3130;
assign n_4672 = x104 & n_3130;
assign n_4673 = x105 & n_3130;
assign n_4674 = x106 & n_3130;
assign n_4675 = x107 & n_3130;
assign n_4676 = x108 & n_3130;
assign n_4677 = x109 & n_3130;
assign n_4678 = x110 & n_3130;
assign n_4679 = x111 & n_3130;
assign n_4680 = x112 & n_3130;
assign n_4681 = x113 & n_3130;
assign n_4682 = x114 & n_3130;
assign n_4683 = x115 & n_3130;
assign n_4684 = x116 & n_3130;
assign n_4685 = x117 & n_3130;
assign n_4686 = x118 & n_3130;
assign n_4687 = x119 & n_3130;
assign n_4688 = x120 & n_3130;
assign n_4689 = x121 & n_3130;
assign n_4690 = x122 & n_3130;
assign n_4691 = x123 & n_3130;
assign n_4692 = x124 & n_3130;
assign n_4693 = x125 & n_3130;
assign n_4694 = x126 & n_3130;
assign n_4695 = ~x53 ^ ~n_3131;
assign n_4696 = n_435 ^ n_3195;
assign n_4697 = x64 & n_3259;
assign n_4698 = x65 & n_3259;
assign n_4699 = x66 & n_3259;
assign n_4700 = x67 & n_3259;
assign n_4701 = x68 & n_3259;
assign n_4702 = x69 & n_3259;
assign n_4703 = x70 & n_3259;
assign n_4704 = x71 & n_3259;
assign n_4705 = x72 & n_3259;
assign n_4706 = x73 & n_3259;
assign n_4707 = x74 & n_3259;
assign n_4708 = x75 & n_3259;
assign n_4709 = x76 & n_3259;
assign n_4710 = x77 & n_3259;
assign n_4711 = x78 & n_3259;
assign n_4712 = x79 & n_3259;
assign n_4713 = x80 & n_3259;
assign n_4714 = x81 & n_3259;
assign n_4715 = x82 & n_3259;
assign n_4716 = x83 & n_3259;
assign n_4717 = x84 & n_3259;
assign n_4718 = x85 & n_3259;
assign n_4719 = x86 & n_3259;
assign n_4720 = x87 & n_3259;
assign n_4721 = x88 & n_3259;
assign n_4722 = x89 & n_3259;
assign n_4723 = x90 & n_3259;
assign n_4724 = x91 & n_3259;
assign n_4725 = x92 & n_3259;
assign n_4726 = x93 & n_3259;
assign n_4727 = x94 & n_3259;
assign n_4728 = x95 & n_3259;
assign n_4729 = x96 & n_3259;
assign n_4730 = x97 & n_3259;
assign n_4731 = x98 & n_3259;
assign n_4732 = x99 & n_3259;
assign n_4733 = x100 & n_3259;
assign n_4734 = x101 & n_3259;
assign n_4735 = x102 & n_3259;
assign n_4736 = x103 & n_3259;
assign n_4737 = x104 & n_3259;
assign n_4738 = x105 & n_3259;
assign n_4739 = x106 & n_3259;
assign n_4740 = x107 & n_3259;
assign n_4741 = x108 & n_3259;
assign n_4742 = x109 & n_3259;
assign n_4743 = x110 & n_3259;
assign n_4744 = x111 & n_3259;
assign n_4745 = x112 & n_3259;
assign n_4746 = x113 & n_3259;
assign n_4747 = x114 & n_3259;
assign n_4748 = x115 & n_3259;
assign n_4749 = x116 & n_3259;
assign n_4750 = x117 & n_3259;
assign n_4751 = x118 & n_3259;
assign n_4752 = x119 & n_3259;
assign n_4753 = x120 & n_3259;
assign n_4754 = x121 & n_3259;
assign n_4755 = x122 & n_3259;
assign n_4756 = x123 & n_3259;
assign n_4757 = x124 & n_3259;
assign n_4758 = x125 & n_3259;
assign n_4759 = x126 & n_3259;
assign n_4760 = x127 & n_3259;
assign n_4761 = x64 & n_3324;
assign n_4762 = x65 & n_3324;
assign n_4763 = x66 & n_3324;
assign n_4764 = x67 & n_3324;
assign n_4765 = x68 & n_3324;
assign n_4766 = x69 & n_3324;
assign n_4767 = x70 & n_3324;
assign n_4768 = x71 & n_3324;
assign n_4769 = x72 & n_3324;
assign n_4770 = x73 & n_3324;
assign n_4771 = x74 & n_3324;
assign n_4772 = x75 & n_3324;
assign n_4773 = x76 & n_3324;
assign n_4774 = x77 & n_3324;
assign n_4775 = x78 & n_3324;
assign n_4776 = x79 & n_3324;
assign n_4777 = x80 & n_3324;
assign n_4778 = x81 & n_3324;
assign n_4779 = x82 & n_3324;
assign n_4780 = x83 & n_3324;
assign n_4781 = x84 & n_3324;
assign n_4782 = x85 & n_3324;
assign n_4783 = x86 & n_3324;
assign n_4784 = x87 & n_3324;
assign n_4785 = x88 & n_3324;
assign n_4786 = x89 & n_3324;
assign n_4787 = x90 & n_3324;
assign n_4788 = x91 & n_3324;
assign n_4789 = x92 & n_3324;
assign n_4790 = x93 & n_3324;
assign n_4791 = x94 & n_3324;
assign n_4792 = x95 & n_3324;
assign n_4793 = x96 & n_3324;
assign n_4794 = x97 & n_3324;
assign n_4795 = x98 & n_3324;
assign n_4796 = x99 & n_3324;
assign n_4797 = x100 & n_3324;
assign n_4798 = x101 & n_3324;
assign n_4799 = x102 & n_3324;
assign n_4800 = x103 & n_3324;
assign n_4801 = x104 & n_3324;
assign n_4802 = x105 & n_3324;
assign n_4803 = x106 & n_3324;
assign n_4804 = x107 & n_3324;
assign n_4805 = x108 & n_3324;
assign n_4806 = x109 & n_3324;
assign n_4807 = x110 & n_3324;
assign n_4808 = x111 & n_3324;
assign n_4809 = x112 & n_3324;
assign n_4810 = x113 & n_3324;
assign n_4811 = x114 & n_3324;
assign n_4812 = x115 & n_3324;
assign n_4813 = x116 & n_3324;
assign n_4814 = x117 & n_3324;
assign n_4815 = x118 & n_3324;
assign n_4816 = x119 & n_3324;
assign n_4817 = x120 & n_3324;
assign n_4818 = x121 & n_3324;
assign n_4819 = x122 & n_3324;
assign n_4820 = x123 & n_3324;
assign n_4821 = x124 & n_3324;
assign n_4822 = x125 & n_3324;
assign n_4823 = x126 & n_3324;
assign n_4824 = x127 & n_3324;
assign n_4825 = x64 & n_3389;
assign n_4826 = x65 & n_3389;
assign n_4827 = x66 & n_3389;
assign n_4828 = x67 & n_3389;
assign n_4829 = x68 & n_3389;
assign n_4830 = x69 & n_3389;
assign n_4831 = x70 & n_3389;
assign n_4832 = x71 & n_3389;
assign n_4833 = x72 & n_3389;
assign n_4834 = x73 & n_3389;
assign n_4835 = x74 & n_3389;
assign n_4836 = x75 & n_3389;
assign n_4837 = x76 & n_3389;
assign n_4838 = x77 & n_3389;
assign n_4839 = x78 & n_3389;
assign n_4840 = x79 & n_3389;
assign n_4841 = x80 & n_3389;
assign n_4842 = x81 & n_3389;
assign n_4843 = x82 & n_3389;
assign n_4844 = x83 & n_3389;
assign n_4845 = x84 & n_3389;
assign n_4846 = x85 & n_3389;
assign n_4847 = x86 & n_3389;
assign n_4848 = x87 & n_3389;
assign n_4849 = x88 & n_3389;
assign n_4850 = x89 & n_3389;
assign n_4851 = x90 & n_3389;
assign n_4852 = x91 & n_3389;
assign n_4853 = x92 & n_3389;
assign n_4854 = x93 & n_3389;
assign n_4855 = x94 & n_3389;
assign n_4856 = x95 & n_3389;
assign n_4857 = x96 & n_3389;
assign n_4858 = x97 & n_3389;
assign n_4859 = x98 & n_3389;
assign n_4860 = x99 & n_3389;
assign n_4861 = x100 & n_3389;
assign n_4862 = x101 & n_3389;
assign n_4863 = x102 & n_3389;
assign n_4864 = x103 & n_3389;
assign n_4865 = x104 & n_3389;
assign n_4866 = x105 & n_3389;
assign n_4867 = x106 & n_3389;
assign n_4868 = x107 & n_3389;
assign n_4869 = x108 & n_3389;
assign n_4870 = x109 & n_3389;
assign n_4871 = x110 & n_3389;
assign n_4872 = x111 & n_3389;
assign n_4873 = x112 & n_3389;
assign n_4874 = x113 & n_3389;
assign n_4875 = x114 & n_3389;
assign n_4876 = x115 & n_3389;
assign n_4877 = x116 & n_3389;
assign n_4878 = x117 & n_3389;
assign n_4879 = x118 & n_3389;
assign n_4880 = x119 & n_3389;
assign n_4881 = x120 & n_3389;
assign n_4882 = x121 & n_3389;
assign n_4883 = x122 & n_3389;
assign n_4884 = x123 & n_3389;
assign n_4885 = x124 & n_3389;
assign n_4886 = x125 & n_3389;
assign n_4887 = x126 & n_3389;
assign n_4888 = x127 & n_3389;
assign n_4889 = n_1985 ^ n_3392;
assign n_4890 = x71 & n_3392;
assign n_4891 = n_3393 ^ x72;
assign n_4892 = n_3394 ^ x11;
assign n_4893 = n_3395 ^ n_1960;
assign n_4894 = n_3396 ^ x81;
assign n_4895 = x83 & n_3398;
assign n_4896 = n_1986 ^ n_3398;
assign n_4897 = n_3399 ^ x84;
assign n_4898 = n_3401 ^ x87;
assign n_4899 = x89 & n_3403;
assign n_4900 = n_1987 ^ n_3403;
assign n_4901 = n_3404 ^ x90;
assign n_4902 = n_3405 ^ x93;
assign n_4903 = n_1988 ^ n_3407;
assign n_4904 = x95 & n_3407;
assign n_4905 = n_3408 ^ x96;
assign n_4906 = n_1989 ^ n_3410;
assign n_4907 = x98 & n_3410;
assign n_4908 = n_3411 ^ x99;
assign n_4909 = n_3412 ^ x38;
assign n_4910 = x101 & n_3413;
assign n_4911 = n_1990 ^ n_3415;
assign n_4912 = x110 & n_3415;
assign n_4913 = n_3416 ^ x111;
assign n_4914 = x116 & n_3418;
assign n_4915 = n_1991 ^ n_3418;
assign n_4916 = n_3419 ^ x117;
assign n_4917 = x122 & n_3421;
assign n_4918 = n_1992 ^ n_3421;
assign n_4919 = n_3422 ^ x123;
assign n_4920 = n_3424 ^ n_629;
assign n_4921 = n_719 ^ n_3425;
assign n_4922 = n_3427 ^ n_105;
assign n_4923 = x67 & ~n_3427;
assign n_4924 = x14 & n_3428;
assign n_4925 = n_3428 ^ n_494;
assign n_4926 = n_3429 ^ n_653;
assign n_4927 = n_3430 ^ n_2256;
assign n_4928 = x64 & n_3431;
assign n_4929 = n_3432 ^ n_2326;
assign n_4930 = n_3433 ^ n_2393;
assign n_4931 = n_3434 ^ n_2460;
assign n_4932 = n_3435 ^ n_1116;
assign n_4933 = n_3436 ^ n_1180;
assign n_4934 = n_3437 ^ n_2658;
assign n_4935 = n_3438 ^ n_2726;
assign n_4936 = n_3439 ^ n_2793;
assign n_4937 = n_3441 ^ n_2927;
assign n_4938 = n_3442 ^ n_2994;
assign n_4939 = n_3443 ^ n_3062;
assign n_4940 = n_3444 ^ n_3129;
assign n_4941 = n_3445 ^ n_1770;
assign n_4942 = n_3446 ^ n_1834;
assign n_4943 = n_3447 ^ n_1898;
assign n_4944 = n_3450 ^ n_527;
assign n_4945 = x70 & ~n_3451;
assign n_4946 = n_0 & ~n_3452;
assign n_4947 = ~x62 & ~n_3453;
assign n_4948 = ~x62 & ~n_3455;
assign n_4949 = n_3457 ^ n_115;
assign n_4950 = n_3457 ^ x2;
assign n_4951 = n_3458 ^ n_7;
assign n_4952 = n_3458 ^ x5;
assign n_4953 = n_3463 ^ n_132;
assign n_4954 = n_3464 ^ n_3394;
assign n_4955 = n_3465 ^ x14;
assign n_4956 = n_3466 ^ n_547;
assign n_4957 = n_3469 ^ x14;
assign n_4958 = n_3469 ^ n_3465;
assign n_4959 = n_0 & ~n_3470;
assign n_4960 = ~x62 & ~n_3471;
assign n_4961 = n_3472 ^ n_149;
assign n_4962 = n_0 & ~n_3475;
assign n_4963 = n_3478 ^ n_171;
assign n_4964 = n_0 & ~n_3484;
assign n_4965 = n_0 & ~n_3485;
assign n_4966 = n_3487 ^ n_196;
assign n_4967 = n_0 & ~n_3489;
assign n_4968 = x63 & n_3490;
assign n_4969 = n_0 & ~n_3495;
assign n_4970 = n_3496 ^ x2;
assign n_4971 = n_3499 ^ ~n_230;
assign n_4972 = n_3500 ^ n_3412;
assign n_4973 = n_3502 ^ x41;
assign n_4974 = n_3503 ^ n_3502;
assign n_4975 = n_3505 ^ n_3502;
assign n_4976 = n_3506 ^ x44;
assign n_4977 = n_3507 ^ n_592;
assign n_4978 = n_0 & ~n_3509;
assign n_4979 = n_0 & ~n_3510;
assign n_4980 = n_3513 ^ n_3506;
assign n_4981 = n_3516 ^ x50;
assign n_4982 = n_3518 ^ n_605;
assign n_4983 = n_0 & ~n_3520;
assign n_4984 = n_3522 ^ x50;
assign n_4985 = n_3522 ^ n_3516;
assign n_4986 = n_0 & ~n_3523;
assign n_4987 = ~n_66 & n_3524;
assign n_4988 = n_66 & ~n_3525;
assign n_4989 = n_3527 ^ n_281;
assign n_4990 = n_3528 ^ x56;
assign n_4991 = n_0 & ~n_3529;
assign n_4992 = ~n_309 & ~n_3532;
assign n_4993 = n_3534 ^ n_308;
assign n_4994 = n_3535 ^ n_2187;
assign n_4995 = n_656 ^ n_3536;
assign n_4996 = n_3537 ^ n_657;
assign n_4997 = n_3538 ^ n_658;
assign n_4998 = n_659 ^ n_3539;
assign n_4999 = n_3540 ^ n_660;
assign n_5000 = n_3541 ^ n_661;
assign n_5001 = n_3542 ^ n_662;
assign n_5002 = n_663 ^ n_3543;
assign n_5003 = n_3544 ^ n_664;
assign n_5004 = n_3545 ^ n_665;
assign n_5005 = n_3546 ^ n_666;
assign n_5006 = n_3547 ^ n_667;
assign n_5007 = n_3548 ^ n_668;
assign n_5008 = n_669 ^ n_3549;
assign n_5009 = n_3550 ^ n_670;
assign n_5010 = n_3551 ^ n_671;
assign n_5011 = n_3552 ^ n_672;
assign n_5012 = n_3553 ^ n_673;
assign n_5013 = n_3554 ^ n_674;
assign n_5014 = n_3555 ^ n_675;
assign n_5015 = n_3556 ^ n_676;
assign n_5016 = n_3557 ^ n_677;
assign n_5017 = n_3558 ^ n_678;
assign n_5018 = n_3559 ^ n_679;
assign n_5019 = n_3560 ^ n_680;
assign n_5020 = n_3561 ^ n_681;
assign n_5021 = n_3562 ^ n_682;
assign n_5022 = n_3563 ^ n_683;
assign n_5023 = n_3564 ^ n_684;
assign n_5024 = n_3565 ^ n_685;
assign n_5025 = n_3566 ^ n_686;
assign n_5026 = n_3567 ^ n_687;
assign n_5027 = n_3568 ^ n_688;
assign n_5028 = n_3569 ^ n_689;
assign n_5029 = n_3570 ^ n_690;
assign n_5030 = n_3571 ^ n_691;
assign n_5031 = n_3572 ^ n_692;
assign n_5032 = n_3573 ^ n_693;
assign n_5033 = n_3574 ^ n_694;
assign n_5034 = n_3575 ^ n_695;
assign n_5035 = n_3576 ^ n_696;
assign n_5036 = n_3577 ^ n_697;
assign n_5037 = n_3578 ^ n_698;
assign n_5038 = n_3579 ^ n_699;
assign n_5039 = n_3580 ^ n_700;
assign n_5040 = n_3581 ^ n_701;
assign n_5041 = n_3582 ^ n_702;
assign n_5042 = n_3583 ^ n_703;
assign n_5043 = n_3584 ^ n_704;
assign n_5044 = n_3585 ^ n_705;
assign n_5045 = n_3586 ^ n_706;
assign n_5046 = n_3587 ^ n_707;
assign n_5047 = n_3588 ^ n_708;
assign n_5048 = n_3589 ^ n_709;
assign n_5049 = n_3590 ^ n_710;
assign n_5050 = n_3591 ^ n_711;
assign n_5051 = n_3592 ^ n_712;
assign n_5052 = n_3593 ^ n_713;
assign n_5053 = n_3594 ^ n_714;
assign n_5054 = n_3595 ^ n_715;
assign n_5055 = n_3596 ^ n_716;
assign n_5056 = ~n_3598 ^ x4;
assign n_5057 = x5 & n_3599;
assign n_5058 = n_785 ^ n_3600;
assign n_5059 = n_3601 ^ n_786;
assign n_5060 = n_3602 ^ n_787;
assign n_5061 = n_3603 ^ n_788;
assign n_5062 = n_3604 ^ n_789;
assign n_5063 = n_3605 ^ n_790;
assign n_5064 = n_3606 ^ n_791;
assign n_5065 = n_3607 ^ n_792;
assign n_5066 = n_3608 ^ n_793;
assign n_5067 = n_3609 ^ n_794;
assign n_5068 = n_3610 ^ n_795;
assign n_5069 = n_3611 ^ n_796;
assign n_5070 = n_3612 ^ n_797;
assign n_5071 = n_3613 ^ n_798;
assign n_5072 = n_3614 ^ n_799;
assign n_5073 = n_3615 ^ n_800;
assign n_5074 = n_3616 ^ n_801;
assign n_5075 = n_3617 ^ n_802;
assign n_5076 = n_3618 ^ n_803;
assign n_5077 = n_3619 ^ n_804;
assign n_5078 = n_3620 ^ n_805;
assign n_5079 = n_3621 ^ n_806;
assign n_5080 = n_3622 ^ n_807;
assign n_5081 = n_3623 ^ n_808;
assign n_5082 = n_3624 ^ n_809;
assign n_5083 = n_3625 ^ n_810;
assign n_5084 = n_3626 ^ n_811;
assign n_5085 = n_3627 ^ n_812;
assign n_5086 = n_3628 ^ n_813;
assign n_5087 = n_3629 ^ n_814;
assign n_5088 = n_3630 ^ n_815;
assign n_5089 = n_3631 ^ n_816;
assign n_5090 = n_3632 ^ n_817;
assign n_5091 = n_3633 ^ n_818;
assign n_5092 = n_3634 ^ n_819;
assign n_5093 = n_3635 ^ n_820;
assign n_5094 = n_3636 ^ n_821;
assign n_5095 = n_3637 ^ n_822;
assign n_5096 = n_3638 ^ n_823;
assign n_5097 = n_3639 ^ n_824;
assign n_5098 = n_3640 ^ n_825;
assign n_5099 = n_3641 ^ n_826;
assign n_5100 = n_3642 ^ n_827;
assign n_5101 = n_3643 ^ n_828;
assign n_5102 = n_3644 ^ n_829;
assign n_5103 = n_3645 ^ n_830;
assign n_5104 = n_3646 ^ n_831;
assign n_5105 = n_3647 ^ n_832;
assign n_5106 = n_3648 ^ n_833;
assign n_5107 = n_3649 ^ n_834;
assign n_5108 = n_3650 ^ n_835;
assign n_5109 = n_3651 ^ n_836;
assign n_5110 = n_3652 ^ n_837;
assign n_5111 = n_3653 ^ n_838;
assign n_5112 = n_3654 ^ n_839;
assign n_5113 = n_3655 ^ n_840;
assign n_5114 = n_3656 ^ n_841;
assign n_5115 = n_3657 ^ n_842;
assign n_5116 = n_3658 ^ n_843;
assign n_5117 = n_3659 ^ n_844;
assign n_5118 = n_3660 ^ n_845;
assign n_5119 = n_721 ^ n_3664;
assign n_5120 = ~n_502 & ~n_3665;
assign n_5121 = n_3666 ^ n_3727;
assign n_5122 = n_3667 ^ n_3728;
assign n_5123 = n_3668 ^ n_3729;
assign n_5124 = n_3669 ^ n_3730;
assign n_5125 = n_3670 ^ n_3731;
assign n_5126 = n_3671 ^ n_3732;
assign n_5127 = n_3733 ^ n_3672;
assign n_5128 = n_3673 ^ n_3734;
assign n_5129 = n_3735 ^ n_3674;
assign n_5130 = n_3675 ^ n_3736;
assign n_5131 = n_3676 ^ n_3737;
assign n_5132 = n_3677 ^ n_3738;
assign n_5133 = n_3739 ^ n_3678;
assign n_5134 = n_3679 ^ n_3740;
assign n_5135 = n_3741 ^ n_3680;
assign n_5136 = n_3681 ^ n_3742;
assign n_5137 = n_3682 ^ n_3743;
assign n_5138 = n_3683 ^ n_3744;
assign n_5139 = n_3745 ^ n_3684;
assign n_5140 = n_3685 ^ n_3746;
assign n_5141 = n_3747 ^ n_3686;
assign n_5142 = n_3687 ^ n_3748;
assign n_5143 = n_3749 ^ n_3688;
assign n_5144 = n_3750 ^ n_3689;
assign n_5145 = n_3690 ^ n_3751;
assign n_5146 = n_3752 ^ n_3691;
assign n_5147 = n_3692 ^ n_3753;
assign n_5148 = n_3754 ^ n_3693;
assign n_5149 = n_3755 ^ n_3694;
assign n_5150 = n_3695 ^ n_3756;
assign n_5151 = n_3696 ^ n_3757;
assign n_5152 = n_3697 ^ n_3758;
assign n_5153 = n_3759 ^ n_3698;
assign n_5154 = n_3760 ^ n_3699;
assign n_5155 = n_3761 ^ n_3700;
assign n_5156 = n_3701 ^ n_3762;
assign n_5157 = n_3763 ^ n_3702;
assign n_5158 = n_3703 ^ n_3764;
assign n_5159 = n_3704 ^ n_3765;
assign n_5160 = n_3705 ^ n_3766;
assign n_5161 = n_3706 ^ n_3767;
assign n_5162 = n_3707 ^ n_3768;
assign n_5163 = n_3708 ^ n_3769;
assign n_5164 = n_3709 ^ n_3770;
assign n_5165 = n_3771 ^ n_3710;
assign n_5166 = n_3772 ^ n_3711;
assign n_5167 = n_3712 ^ n_3773;
assign n_5168 = n_3774 ^ n_3713;
assign n_5169 = n_3714 ^ n_3775;
assign n_5170 = n_3776 ^ n_3715;
assign n_5171 = n_3777 ^ n_3716;
assign n_5172 = n_3778 ^ n_3717;
assign n_5173 = n_3718 ^ n_3779;
assign n_5174 = n_3719 ^ n_3780;
assign n_5175 = n_3781 ^ n_3720;
assign n_5176 = n_3721 ^ n_3782;
assign n_5177 = n_3722 ^ n_3783;
assign n_5178 = n_3723 ^ n_3784;
assign n_5179 = n_3724 ^ n_3785;
assign n_5180 = n_3786 ^ n_3725;
assign n_5181 = n_3726 ^ n_3787;
assign n_5182 = n_3790 ^ n_855;
assign n_5183 = n_3791 ^ n_856;
assign n_5184 = n_3792 ^ n_857;
assign n_5185 = n_3793 ^ n_858;
assign n_5186 = n_3794 ^ n_859;
assign n_5187 = n_3795 ^ n_860;
assign n_5188 = n_3796 ^ n_861;
assign n_5189 = n_3797 ^ n_862;
assign n_5190 = n_3798 ^ n_863;
assign n_5191 = n_3799 ^ n_864;
assign n_5192 = n_3800 ^ n_865;
assign n_5193 = n_3801 ^ n_866;
assign n_5194 = n_3802 ^ n_867;
assign n_5195 = n_3803 ^ n_868;
assign n_5196 = n_3804 ^ n_869;
assign n_5197 = n_3805 ^ n_870;
assign n_5198 = n_3806 ^ n_871;
assign n_5199 = n_3807 ^ n_872;
assign n_5200 = n_3808 ^ n_873;
assign n_5201 = n_3809 ^ n_874;
assign n_5202 = n_3810 ^ n_875;
assign n_5203 = n_3811 ^ n_876;
assign n_5204 = n_3812 ^ n_877;
assign n_5205 = n_3813 ^ n_878;
assign n_5206 = n_3814 ^ n_879;
assign n_5207 = n_3815 ^ n_880;
assign n_5208 = n_3816 ^ n_881;
assign n_5209 = n_3817 ^ n_882;
assign n_5210 = n_3818 ^ n_883;
assign n_5211 = n_3819 ^ n_884;
assign n_5212 = n_3820 ^ n_885;
assign n_5213 = n_3821 ^ n_886;
assign n_5214 = n_3822 ^ n_887;
assign n_5215 = n_3823 ^ n_888;
assign n_5216 = n_3824 ^ n_889;
assign n_5217 = n_3825 ^ n_890;
assign n_5218 = n_3826 ^ n_891;
assign n_5219 = n_3827 ^ n_892;
assign n_5220 = n_3828 ^ n_893;
assign n_5221 = n_3829 ^ n_894;
assign n_5222 = n_3830 ^ n_895;
assign n_5223 = n_3831 ^ n_896;
assign n_5224 = n_3832 ^ n_897;
assign n_5225 = n_3833 ^ n_898;
assign n_5226 = n_3834 ^ n_899;
assign n_5227 = n_3835 ^ n_900;
assign n_5228 = n_3836 ^ n_901;
assign n_5229 = n_3837 ^ n_902;
assign n_5230 = n_3838 ^ n_903;
assign n_5231 = n_3839 ^ n_904;
assign n_5232 = n_3840 ^ n_905;
assign n_5233 = n_3841 ^ n_906;
assign n_5234 = n_3842 ^ n_907;
assign n_5235 = n_3843 ^ n_908;
assign n_5236 = n_3844 ^ n_909;
assign n_5237 = n_3845 ^ n_910;
assign n_5238 = n_3846 ^ n_911;
assign n_5239 = n_3847 ^ n_912;
assign n_5240 = n_3848 ^ n_913;
assign n_5241 = n_3849 ^ n_914;
assign n_5242 = n_3850 ^ n_915;
assign n_5243 = ~n_3852 ^ x13;
assign n_5244 = n_2260 ^ n_3853;
assign n_5245 = x64 & n_3854;
assign n_5246 = n_921 ^ n_3855;
assign n_5247 = n_922 ^ n_3856;
assign n_5248 = n_3857 ^ n_923;
assign n_5249 = n_3858 ^ n_924;
assign n_5250 = n_3859 ^ n_925;
assign n_5251 = n_3860 ^ n_926;
assign n_5252 = n_3861 ^ n_927;
assign n_5253 = n_928 ^ n_3862;
assign n_5254 = n_929 ^ n_3863;
assign n_5255 = n_3864 ^ n_930;
assign n_5256 = n_931 ^ n_3865;
assign n_5257 = n_932 ^ n_3866;
assign n_5258 = n_933 ^ n_3867;
assign n_5259 = n_934 ^ n_3868;
assign n_5260 = n_935 ^ n_3869;
assign n_5261 = n_936 ^ n_3870;
assign n_5262 = n_937 ^ n_3871;
assign n_5263 = n_938 ^ n_3872;
assign n_5264 = n_939 ^ n_3873;
assign n_5265 = n_940 ^ n_3874;
assign n_5266 = n_941 ^ n_3875;
assign n_5267 = n_942 ^ n_3876;
assign n_5268 = n_943 ^ n_3877;
assign n_5269 = n_944 ^ n_3878;
assign n_5270 = n_945 ^ n_3879;
assign n_5271 = n_946 ^ n_3880;
assign n_5272 = n_947 ^ n_3881;
assign n_5273 = n_948 ^ n_3882;
assign n_5274 = n_949 ^ n_3883;
assign n_5275 = n_950 ^ n_3884;
assign n_5276 = n_951 ^ n_3885;
assign n_5277 = n_952 ^ n_3886;
assign n_5278 = n_953 ^ n_3887;
assign n_5279 = n_954 ^ n_3888;
assign n_5280 = n_955 ^ n_3889;
assign n_5281 = n_956 ^ n_3890;
assign n_5282 = n_957 ^ n_3891;
assign n_5283 = n_958 ^ n_3892;
assign n_5284 = n_959 ^ n_3893;
assign n_5285 = n_960 ^ n_3894;
assign n_5286 = n_961 ^ n_3895;
assign n_5287 = n_962 ^ n_3896;
assign n_5288 = n_963 ^ n_3897;
assign n_5289 = n_964 ^ n_3898;
assign n_5290 = n_965 ^ n_3899;
assign n_5291 = n_966 ^ n_3900;
assign n_5292 = n_967 ^ n_3901;
assign n_5293 = n_968 ^ n_3902;
assign n_5294 = n_969 ^ n_3903;
assign n_5295 = n_970 ^ n_3904;
assign n_5296 = n_971 ^ n_3905;
assign n_5297 = n_972 ^ n_3906;
assign n_5298 = n_973 ^ n_3907;
assign n_5299 = n_974 ^ n_3908;
assign n_5300 = n_975 ^ n_3909;
assign n_5301 = n_976 ^ n_3910;
assign n_5302 = n_977 ^ n_3911;
assign n_5303 = n_978 ^ n_3912;
assign n_5304 = n_979 ^ n_3913;
assign n_5305 = n_980 ^ n_3914;
assign n_5306 = n_981 ^ n_3915;
assign n_5307 = ~n_3917 ^ x16;
assign n_5308 = n_2327 ^ n_3918;
assign n_5309 = x64 & n_3919;
assign n_5310 = n_987 ^ n_3920;
assign n_5311 = n_3921 ^ n_988;
assign n_5312 = n_3922 ^ n_989;
assign n_5313 = n_990 ^ n_3923;
assign n_5314 = n_991 ^ n_3924;
assign n_5315 = n_3925 ^ n_992;
assign n_5316 = n_3926 ^ n_993;
assign n_5317 = n_994 ^ n_3927;
assign n_5318 = n_995 ^ n_3928;
assign n_5319 = n_996 ^ n_3929;
assign n_5320 = n_997 ^ n_3930;
assign n_5321 = n_998 ^ n_3931;
assign n_5322 = n_999 ^ n_3932;
assign n_5323 = n_1000 ^ n_3933;
assign n_5324 = n_3934 ^ n_1001;
assign n_5325 = n_1002 ^ n_3935;
assign n_5326 = n_1003 ^ n_3936;
assign n_5327 = n_1004 ^ n_3937;
assign n_5328 = n_1005 ^ n_3938;
assign n_5329 = n_3939 ^ n_1006;
assign n_5330 = n_1007 ^ n_3940;
assign n_5331 = n_1008 ^ n_3941;
assign n_5332 = n_1009 ^ n_3942;
assign n_5333 = n_1010 ^ n_3943;
assign n_5334 = n_3944 ^ n_1011;
assign n_5335 = n_1012 ^ n_3945;
assign n_5336 = n_1013 ^ n_3946;
assign n_5337 = n_1014 ^ n_3947;
assign n_5338 = n_1015 ^ n_3948;
assign n_5339 = n_1016 ^ n_3949;
assign n_5340 = n_1017 ^ n_3950;
assign n_5341 = n_3951 ^ n_1018;
assign n_5342 = n_1019 ^ n_3952;
assign n_5343 = n_1020 ^ n_3953;
assign n_5344 = n_1021 ^ n_3954;
assign n_5345 = n_1022 ^ n_3955;
assign n_5346 = n_3956 ^ n_1023;
assign n_5347 = n_1024 ^ n_3957;
assign n_5348 = n_1025 ^ n_3958;
assign n_5349 = n_1026 ^ n_3959;
assign n_5350 = n_1027 ^ n_3960;
assign n_5351 = n_1028 ^ n_3961;
assign n_5352 = n_1029 ^ n_3962;
assign n_5353 = n_1030 ^ n_3963;
assign n_5354 = n_1031 ^ n_3964;
assign n_5355 = n_1032 ^ n_3965;
assign n_5356 = n_1033 ^ n_3966;
assign n_5357 = n_1034 ^ n_3967;
assign n_5358 = n_1035 ^ n_3968;
assign n_5359 = n_1036 ^ n_3969;
assign n_5360 = n_1037 ^ n_3970;
assign n_5361 = n_1038 ^ n_3971;
assign n_5362 = n_1039 ^ n_3972;
assign n_5363 = n_1040 ^ n_3973;
assign n_5364 = n_3974 ^ n_1041;
assign n_5365 = n_1042 ^ n_3975;
assign n_5366 = n_3976 ^ n_1043;
assign n_5367 = n_1044 ^ n_3977;
assign n_5368 = n_1045 ^ n_3978;
assign n_5369 = n_1046 ^ n_3979;
assign n_5370 = n_1047 ^ n_3980;
assign n_5371 = ~n_3982 ^ x19;
assign n_5372 = n_2394 ^ n_3983;
assign n_5373 = x64 & n_3984;
assign n_5374 = n_3985 ^ n_1053;
assign n_5375 = n_3986 ^ n_1054;
assign n_5376 = n_3987 ^ n_1055;
assign n_5377 = n_3988 ^ n_1056;
assign n_5378 = n_1057 ^ n_3989;
assign n_5379 = n_3990 ^ n_1058;
assign n_5380 = n_3991 ^ n_1059;
assign n_5381 = n_1060 ^ n_3992;
assign n_5382 = n_1061 ^ n_3993;
assign n_5383 = n_3994 ^ n_1062;
assign n_5384 = n_1063 ^ n_3995;
assign n_5385 = n_3996 ^ n_1064;
assign n_5386 = n_1065 ^ n_3997;
assign n_5387 = n_1066 ^ n_3998;
assign n_5388 = n_1067 ^ n_3999;
assign n_5389 = n_1068 ^ n_4000;
assign n_5390 = n_1069 ^ n_4001;
assign n_5391 = n_1070 ^ n_4002;
assign n_5392 = n_1071 ^ n_4003;
assign n_5393 = n_1072 ^ n_4004;
assign n_5394 = n_1073 ^ n_4005;
assign n_5395 = n_1074 ^ n_4006;
assign n_5396 = n_1075 ^ n_4007;
assign n_5397 = n_1076 ^ n_4008;
assign n_5398 = n_1077 ^ n_4009;
assign n_5399 = n_1078 ^ n_4010;
assign n_5400 = n_1079 ^ n_4011;
assign n_5401 = n_1080 ^ n_4012;
assign n_5402 = n_1081 ^ n_4013;
assign n_5403 = n_1082 ^ n_4014;
assign n_5404 = n_1083 ^ n_4015;
assign n_5405 = n_1084 ^ n_4016;
assign n_5406 = n_1085 ^ n_4017;
assign n_5407 = n_1086 ^ n_4018;
assign n_5408 = n_1087 ^ n_4019;
assign n_5409 = n_1088 ^ n_4020;
assign n_5410 = n_1089 ^ n_4021;
assign n_5411 = n_1090 ^ n_4022;
assign n_5412 = n_1091 ^ n_4023;
assign n_5413 = n_1092 ^ n_4024;
assign n_5414 = n_1093 ^ n_4025;
assign n_5415 = n_4026 ^ n_1094;
assign n_5416 = n_1095 ^ n_4027;
assign n_5417 = n_1096 ^ n_4028;
assign n_5418 = n_1097 ^ n_4029;
assign n_5419 = n_1098 ^ n_4030;
assign n_5420 = n_1099 ^ n_4031;
assign n_5421 = n_1100 ^ n_4032;
assign n_5422 = n_1101 ^ n_4033;
assign n_5423 = n_1102 ^ n_4034;
assign n_5424 = n_1103 ^ n_4035;
assign n_5425 = n_1104 ^ n_4036;
assign n_5426 = n_4037 ^ n_1105;
assign n_5427 = n_1106 ^ n_4038;
assign n_5428 = n_1107 ^ n_4039;
assign n_5429 = n_1108 ^ n_4040;
assign n_5430 = n_1109 ^ n_4041;
assign n_5431 = n_1110 ^ n_4042;
assign n_5432 = n_1111 ^ n_4043;
assign n_5433 = n_1112 ^ n_4044;
assign n_5434 = n_1113 ^ n_4045;
assign n_5435 = ~n_4047 ^ x22;
assign n_5436 = n_2461 ^ n_4048;
assign n_5437 = n_4049 ^ n_2591;
assign n_5438 = n_2528 ^ n_4050;
assign n_5439 = n_4051 ^ n_1118;
assign n_5440 = n_4052 ^ n_1119;
assign n_5441 = n_4053 ^ n_1120;
assign n_5442 = n_4054 ^ n_1121;
assign n_5443 = n_4055 ^ n_1122;
assign n_5444 = n_4056 ^ n_1123;
assign n_5445 = n_4057 ^ n_1124;
assign n_5446 = n_4058 ^ n_1125;
assign n_5447 = n_4059 ^ n_1126;
assign n_5448 = n_4060 ^ n_1127;
assign n_5449 = n_4061 ^ n_1128;
assign n_5450 = n_4062 ^ n_1129;
assign n_5451 = n_1130 ^ n_4063;
assign n_5452 = n_4064 ^ n_1131;
assign n_5453 = n_4065 ^ n_1132;
assign n_5454 = n_4066 ^ n_1133;
assign n_5455 = n_4067 ^ n_1134;
assign n_5456 = n_4068 ^ n_1135;
assign n_5457 = n_4069 ^ n_1136;
assign n_5458 = n_4070 ^ n_1137;
assign n_5459 = n_4071 ^ n_1138;
assign n_5460 = n_4072 ^ n_1139;
assign n_5461 = n_4073 ^ n_1140;
assign n_5462 = n_4074 ^ n_1141;
assign n_5463 = n_4075 ^ n_1142;
assign n_5464 = n_4076 ^ n_1143;
assign n_5465 = n_4077 ^ n_1144;
assign n_5466 = n_4078 ^ n_1145;
assign n_5467 = n_4079 ^ n_1146;
assign n_5468 = n_4080 ^ n_1147;
assign n_5469 = n_4081 ^ n_1148;
assign n_5470 = n_4082 ^ n_1149;
assign n_5471 = n_4083 ^ n_1150;
assign n_5472 = n_4084 ^ n_1151;
assign n_5473 = n_4085 ^ n_1152;
assign n_5474 = n_4086 ^ n_1153;
assign n_5475 = n_4087 ^ n_1154;
assign n_5476 = n_4088 ^ n_1155;
assign n_5477 = n_4089 ^ n_1156;
assign n_5478 = n_4090 ^ n_1157;
assign n_5479 = n_4091 ^ n_1158;
assign n_5480 = n_4092 ^ n_1159;
assign n_5481 = n_4093 ^ n_1160;
assign n_5482 = n_4094 ^ n_1161;
assign n_5483 = n_4095 ^ n_1162;
assign n_5484 = n_4096 ^ n_1163;
assign n_5485 = n_4097 ^ n_1164;
assign n_5486 = n_4098 ^ n_1165;
assign n_5487 = n_4099 ^ n_1166;
assign n_5488 = n_4100 ^ n_1167;
assign n_5489 = n_4101 ^ n_1168;
assign n_5490 = n_4102 ^ n_1169;
assign n_5491 = n_4103 ^ n_1170;
assign n_5492 = n_4104 ^ n_1171;
assign n_5493 = n_4105 ^ n_1172;
assign n_5494 = n_4106 ^ n_1173;
assign n_5495 = n_4107 ^ n_1174;
assign n_5496 = n_4108 ^ n_1175;
assign n_5497 = n_4109 ^ n_1176;
assign n_5498 = n_4110 ^ n_1177;
assign n_5499 = n_4113 ^ n_1182;
assign n_5500 = n_4114 ^ n_1183;
assign n_5501 = n_4115 ^ n_1184;
assign n_5502 = n_4116 ^ n_1185;
assign n_5503 = n_4117 ^ n_1186;
assign n_5504 = n_4118 ^ n_1187;
assign n_5505 = n_4119 ^ n_1188;
assign n_5506 = n_4120 ^ n_1189;
assign n_5507 = n_4121 ^ n_1190;
assign n_5508 = n_4122 ^ n_1191;
assign n_5509 = n_4123 ^ n_1192;
assign n_5510 = n_4124 ^ n_1193;
assign n_5511 = n_4125 ^ n_1194;
assign n_5512 = n_4126 ^ n_1195;
assign n_5513 = n_4127 ^ n_1196;
assign n_5514 = n_4128 ^ n_1197;
assign n_5515 = n_4129 ^ n_1198;
assign n_5516 = n_4130 ^ n_1199;
assign n_5517 = n_4131 ^ n_1200;
assign n_5518 = n_4132 ^ n_1201;
assign n_5519 = n_4133 ^ n_1202;
assign n_5520 = n_4134 ^ n_1203;
assign n_5521 = n_4135 ^ n_1204;
assign n_5522 = n_4136 ^ n_1205;
assign n_5523 = n_4137 ^ n_1206;
assign n_5524 = n_4138 ^ n_1207;
assign n_5525 = n_4139 ^ n_1208;
assign n_5526 = n_4140 ^ n_1209;
assign n_5527 = n_4141 ^ n_1210;
assign n_5528 = n_4142 ^ n_1211;
assign n_5529 = n_4143 ^ n_1212;
assign n_5530 = n_4144 ^ n_1213;
assign n_5531 = n_4145 ^ n_1214;
assign n_5532 = n_4146 ^ n_1215;
assign n_5533 = n_4147 ^ n_1216;
assign n_5534 = n_4148 ^ n_1217;
assign n_5535 = n_4149 ^ n_1218;
assign n_5536 = n_4150 ^ n_1219;
assign n_5537 = n_4151 ^ n_1220;
assign n_5538 = n_4152 ^ n_1221;
assign n_5539 = n_4153 ^ n_1222;
assign n_5540 = n_4154 ^ n_1223;
assign n_5541 = n_4155 ^ n_1224;
assign n_5542 = n_4156 ^ n_1225;
assign n_5543 = n_4157 ^ n_1226;
assign n_5544 = n_4158 ^ n_1227;
assign n_5545 = n_4159 ^ n_1228;
assign n_5546 = n_4160 ^ n_1229;
assign n_5547 = n_4161 ^ n_1230;
assign n_5548 = n_4162 ^ n_1231;
assign n_5549 = n_4163 ^ n_1232;
assign n_5550 = n_4164 ^ n_1233;
assign n_5551 = n_4165 ^ n_1234;
assign n_5552 = n_4166 ^ n_1235;
assign n_5553 = n_4167 ^ n_1236;
assign n_5554 = n_4168 ^ n_1237;
assign n_5555 = n_4169 ^ n_1238;
assign n_5556 = n_4170 ^ n_1239;
assign n_5557 = n_4171 ^ n_1240;
assign n_5558 = n_4172 ^ n_1241;
assign n_5559 = n_4173 ^ n_1242;
assign n_5560 = ~n_4175 ^ x28;
assign n_5561 = n_2592 ^ n_4176;
assign n_5562 = n_4177 ^ n_1249;
assign n_5563 = n_1250 ^ n_4178;
assign n_5564 = n_1251 ^ n_4179;
assign n_5565 = n_4180 ^ n_1252;
assign n_5566 = n_1253 ^ n_4181;
assign n_5567 = n_4182 ^ n_1254;
assign n_5568 = n_1255 ^ n_4183;
assign n_5569 = n_4184 ^ n_1256;
assign n_5570 = n_1257 ^ n_4185;
assign n_5571 = n_1258 ^ n_4186;
assign n_5572 = n_1259 ^ n_4187;
assign n_5573 = n_1260 ^ n_4188;
assign n_5574 = n_1261 ^ n_4189;
assign n_5575 = n_1262 ^ n_4190;
assign n_5576 = n_1263 ^ n_4191;
assign n_5577 = n_1264 ^ n_4192;
assign n_5578 = n_1265 ^ n_4193;
assign n_5579 = n_1266 ^ n_4194;
assign n_5580 = n_1267 ^ n_4195;
assign n_5581 = n_1268 ^ n_4196;
assign n_5582 = n_1269 ^ n_4197;
assign n_5583 = n_1270 ^ n_4198;
assign n_5584 = n_1271 ^ n_4199;
assign n_5585 = n_1272 ^ n_4200;
assign n_5586 = n_1273 ^ n_4201;
assign n_5587 = n_1274 ^ n_4202;
assign n_5588 = n_1275 ^ n_4203;
assign n_5589 = n_1276 ^ n_4204;
assign n_5590 = n_1277 ^ n_4205;
assign n_5591 = n_1278 ^ n_4206;
assign n_5592 = n_1279 ^ n_4207;
assign n_5593 = n_1280 ^ n_4208;
assign n_5594 = n_1281 ^ n_4209;
assign n_5595 = n_1282 ^ n_4210;
assign n_5596 = n_1283 ^ n_4211;
assign n_5597 = n_4212 ^ n_1284;
assign n_5598 = n_1285 ^ n_4213;
assign n_5599 = n_1286 ^ n_4214;
assign n_5600 = n_1287 ^ n_4215;
assign n_5601 = n_1288 ^ n_4216;
assign n_5602 = n_1289 ^ n_4217;
assign n_5603 = n_1290 ^ n_4218;
assign n_5604 = n_1291 ^ n_4219;
assign n_5605 = n_1292 ^ n_4220;
assign n_5606 = n_1293 ^ n_4221;
assign n_5607 = n_1294 ^ n_4222;
assign n_5608 = n_1295 ^ n_4223;
assign n_5609 = n_1296 ^ n_4224;
assign n_5610 = n_1297 ^ n_4225;
assign n_5611 = n_1298 ^ n_4226;
assign n_5612 = n_1299 ^ n_4227;
assign n_5613 = n_1300 ^ n_4228;
assign n_5614 = n_1301 ^ n_4229;
assign n_5615 = n_1302 ^ n_4230;
assign n_5616 = n_1303 ^ n_4231;
assign n_5617 = n_1304 ^ n_4232;
assign n_5618 = n_1305 ^ n_4233;
assign n_5619 = n_1306 ^ n_4234;
assign n_5620 = n_1307 ^ n_4235;
assign n_5621 = n_1308 ^ n_4236;
assign n_5622 = n_1309 ^ n_4237;
assign n_5623 = n_2659 ^ n_4241;
assign n_5624 = x64 & n_4242;
assign n_5625 = n_4243 ^ n_1315;
assign n_5626 = n_4244 ^ n_1316;
assign n_5627 = n_1317 ^ n_4245;
assign n_5628 = n_1318 ^ n_4246;
assign n_5629 = n_1319 ^ n_4247;
assign n_5630 = n_1320 ^ n_4248;
assign n_5631 = n_1321 ^ n_4249;
assign n_5632 = n_1322 ^ n_4250;
assign n_5633 = n_4251 ^ n_1323;
assign n_5634 = n_4252 ^ n_1324;
assign n_5635 = n_1325 ^ n_4253;
assign n_5636 = n_4254 ^ n_1326;
assign n_5637 = n_1327 ^ n_4255;
assign n_5638 = n_1328 ^ n_4256;
assign n_5639 = n_4257 ^ n_1329;
assign n_5640 = n_4258 ^ n_1330;
assign n_5641 = n_1331 ^ n_4259;
assign n_5642 = n_1332 ^ n_4260;
assign n_5643 = n_4261 ^ n_1333;
assign n_5644 = n_4262 ^ n_1334;
assign n_5645 = n_1335 ^ n_4263;
assign n_5646 = n_1336 ^ n_4264;
assign n_5647 = n_4265 ^ n_1337;
assign n_5648 = n_4266 ^ n_1338;
assign n_5649 = n_1339 ^ n_4267;
assign n_5650 = n_1340 ^ n_4268;
assign n_5651 = n_4269 ^ n_1341;
assign n_5652 = n_4270 ^ n_1342;
assign n_5653 = n_1343 ^ n_4271;
assign n_5654 = n_4272 ^ n_1344;
assign n_5655 = n_1345 ^ n_4273;
assign n_5656 = n_1346 ^ n_4274;
assign n_5657 = n_1347 ^ n_4275;
assign n_5658 = n_1348 ^ n_4276;
assign n_5659 = n_1349 ^ n_4277;
assign n_5660 = n_4278 ^ n_1350;
assign n_5661 = n_4279 ^ n_1351;
assign n_5662 = n_1352 ^ n_4280;
assign n_5663 = n_1353 ^ n_4281;
assign n_5664 = n_4282 ^ n_1354;
assign n_5665 = n_1355 ^ n_4283;
assign n_5666 = n_1356 ^ n_4284;
assign n_5667 = n_4285 ^ n_1357;
assign n_5668 = n_4286 ^ n_1358;
assign n_5669 = n_4287 ^ n_1359;
assign n_5670 = n_4288 ^ n_1360;
assign n_5671 = n_4289 ^ n_1361;
assign n_5672 = n_4290 ^ n_1362;
assign n_5673 = n_1363 ^ n_4291;
assign n_5674 = n_4292 ^ n_1364;
assign n_5675 = n_1365 ^ n_4293;
assign n_5676 = n_4294 ^ n_1366;
assign n_5677 = n_1367 ^ n_4295;
assign n_5678 = n_1368 ^ n_4296;
assign n_5679 = n_1369 ^ n_4297;
assign n_5680 = n_1370 ^ n_4298;
assign n_5681 = n_4299 ^ n_1371;
assign n_5682 = n_4300 ^ n_1372;
assign n_5683 = n_4301 ^ n_1373;
assign n_5684 = n_4302 ^ n_1374;
assign n_5685 = n_1375 ^ n_4303;
assign n_5686 = ~n_4305 ^ x34;
assign n_5687 = n_2727 ^ n_4306;
assign n_5688 = x64 & n_4307;
assign n_5689 = n_1381 ^ n_4308;
assign n_5690 = n_1382 ^ n_4309;
assign n_5691 = n_1383 ^ n_4310;
assign n_5692 = n_1384 ^ n_4311;
assign n_5693 = n_1385 ^ n_4312;
assign n_5694 = n_1386 ^ n_4313;
assign n_5695 = n_4314 ^ n_1387;
assign n_5696 = n_1388 ^ n_4315;
assign n_5697 = n_1389 ^ n_4316;
assign n_5698 = n_4317 ^ n_1390;
assign n_5699 = n_1391 ^ n_4318;
assign n_5700 = n_4319 ^ n_1392;
assign n_5701 = n_1393 ^ n_4320;
assign n_5702 = n_4321 ^ n_1394;
assign n_5703 = n_1395 ^ n_4322;
assign n_5704 = n_4323 ^ n_1396;
assign n_5705 = n_1397 ^ n_4324;
assign n_5706 = n_1398 ^ n_4325;
assign n_5707 = n_4326 ^ n_1399;
assign n_5708 = n_4327 ^ n_1400;
assign n_5709 = n_1401 ^ n_4328;
assign n_5710 = n_4329 ^ n_1402;
assign n_5711 = n_4330 ^ n_1403;
assign n_5712 = n_4331 ^ n_1404;
assign n_5713 = n_4332 ^ n_1405;
assign n_5714 = n_1406 ^ n_4333;
assign n_5715 = n_4334 ^ n_1407;
assign n_5716 = n_1408 ^ n_4335;
assign n_5717 = n_4336 ^ n_1409;
assign n_5718 = n_1410 ^ n_4337;
assign n_5719 = n_4338 ^ n_1411;
assign n_5720 = n_4339 ^ n_1412;
assign n_5721 = n_4340 ^ n_1413;
assign n_5722 = n_1414 ^ n_4341;
assign n_5723 = n_1415 ^ n_4342;
assign n_5724 = n_1416 ^ n_4343;
assign n_5725 = n_4344 ^ n_1417;
assign n_5726 = n_4345 ^ n_1418;
assign n_5727 = n_4346 ^ n_1419;
assign n_5728 = n_4347 ^ n_1420;
assign n_5729 = n_1421 ^ n_4348;
assign n_5730 = n_4349 ^ n_1422;
assign n_5731 = n_1423 ^ n_4350;
assign n_5732 = n_1424 ^ n_4351;
assign n_5733 = n_4352 ^ n_1425;
assign n_5734 = n_4353 ^ n_1426;
assign n_5735 = n_4354 ^ n_1427;
assign n_5736 = n_1428 ^ n_4355;
assign n_5737 = n_4356 ^ n_1429;
assign n_5738 = n_4357 ^ n_1430;
assign n_5739 = n_4358 ^ n_1431;
assign n_5740 = n_4359 ^ n_1432;
assign n_5741 = n_4360 ^ n_1433;
assign n_5742 = n_4361 ^ n_1434;
assign n_5743 = n_4362 ^ n_1435;
assign n_5744 = n_4363 ^ n_1436;
assign n_5745 = n_1437 ^ n_4364;
assign n_5746 = n_1438 ^ n_4365;
assign n_5747 = n_4366 ^ n_1439;
assign n_5748 = n_4367 ^ n_1440;
assign n_5749 = n_4368 ^ n_1441;
assign n_5750 = ~n_4370 ^ x37;
assign n_5751 = n_2794 ^ n_4371;
assign n_5752 = n_4372 ^ n_3440;
assign n_5753 = n_4373 ^ n_412;
assign n_5754 = n_4374 ^ n_2926;
assign n_5755 = n_2863 ^ n_4375;
assign n_5756 = n_1446 ^ n_4376;
assign n_5757 = n_1447 ^ n_4377;
assign n_5758 = n_1448 ^ n_4378;
assign n_5759 = n_1449 ^ n_4379;
assign n_5760 = n_1450 ^ n_4380;
assign n_5761 = n_1451 ^ n_4381;
assign n_5762 = n_1452 ^ n_4382;
assign n_5763 = n_4383 ^ n_1453;
assign n_5764 = n_1454 ^ n_4384;
assign n_5765 = n_1455 ^ n_4385;
assign n_5766 = n_4386 ^ n_1456;
assign n_5767 = n_4387 ^ n_1457;
assign n_5768 = n_1458 ^ n_4388;
assign n_5769 = n_1459 ^ n_4389;
assign n_5770 = n_1460 ^ n_4390;
assign n_5771 = n_1461 ^ n_4391;
assign n_5772 = n_1462 ^ n_4392;
assign n_5773 = n_4393 ^ n_1463;
assign n_5774 = n_4394 ^ n_1464;
assign n_5775 = n_1465 ^ n_4395;
assign n_5776 = n_4396 ^ n_1466;
assign n_5777 = n_1467 ^ n_4397;
assign n_5778 = n_4398 ^ n_1468;
assign n_5779 = n_1469 ^ n_4399;
assign n_5780 = n_1470 ^ n_4400;
assign n_5781 = n_4401 ^ n_1471;
assign n_5782 = n_1472 ^ n_4402;
assign n_5783 = n_4403 ^ n_1473;
assign n_5784 = n_1474 ^ n_4404;
assign n_5785 = n_1475 ^ n_4405;
assign n_5786 = n_1476 ^ n_4406;
assign n_5787 = n_1477 ^ n_4407;
assign n_5788 = n_4408 ^ n_1478;
assign n_5789 = n_1479 ^ n_4409;
assign n_5790 = n_4410 ^ n_1480;
assign n_5791 = n_1481 ^ n_4411;
assign n_5792 = n_1482 ^ n_4412;
assign n_5793 = n_1483 ^ n_4413;
assign n_5794 = n_1484 ^ n_4414;
assign n_5795 = n_4415 ^ n_1485;
assign n_5796 = n_4416 ^ n_1486;
assign n_5797 = n_1487 ^ n_4417;
assign n_5798 = n_4418 ^ n_1488;
assign n_5799 = n_4419 ^ n_1489;
assign n_5800 = n_4420 ^ n_1490;
assign n_5801 = n_4421 ^ n_1491;
assign n_5802 = n_1492 ^ n_4422;
assign n_5803 = n_4423 ^ n_1493;
assign n_5804 = n_1494 ^ n_4424;
assign n_5805 = n_4425 ^ n_1495;
assign n_5806 = n_4426 ^ n_1496;
assign n_5807 = n_1497 ^ n_4427;
assign n_5808 = n_4428 ^ n_1498;
assign n_5809 = n_4429 ^ n_1499;
assign n_5810 = n_1500 ^ n_4430;
assign n_5811 = n_4431 ^ n_1501;
assign n_5812 = n_1502 ^ n_4432;
assign n_5813 = n_1503 ^ n_4433;
assign n_5814 = n_1504 ^ n_4434;
assign n_5815 = n_4435 ^ n_1505;
assign n_5816 = x64 & n_4438;
assign n_5817 = n_1511 ^ n_4439;
assign n_5818 = n_1512 ^ n_4440;
assign n_5819 = n_1513 ^ n_4441;
assign n_5820 = n_1514 ^ n_4442;
assign n_5821 = n_1515 ^ n_4443;
assign n_5822 = n_1516 ^ n_4444;
assign n_5823 = n_1517 ^ n_4445;
assign n_5824 = n_1518 ^ n_4446;
assign n_5825 = n_1519 ^ n_4447;
assign n_5826 = n_1520 ^ n_4448;
assign n_5827 = n_4449 ^ n_1521;
assign n_5828 = n_1522 ^ n_4450;
assign n_5829 = n_4451 ^ n_1523;
assign n_5830 = n_1524 ^ n_4452;
assign n_5831 = n_1525 ^ n_4453;
assign n_5832 = n_1526 ^ n_4454;
assign n_5833 = n_1527 ^ n_4455;
assign n_5834 = n_4456 ^ n_1528;
assign n_5835 = n_1529 ^ n_4457;
assign n_5836 = n_1530 ^ n_4458;
assign n_5837 = n_1531 ^ n_4459;
assign n_5838 = n_4460 ^ n_1532;
assign n_5839 = n_1533 ^ n_4461;
assign n_5840 = n_1534 ^ n_4462;
assign n_5841 = n_4463 ^ n_1535;
assign n_5842 = n_4464 ^ n_1536;
assign n_5843 = n_1537 ^ n_4465;
assign n_5844 = n_4466 ^ n_1538;
assign n_5845 = n_1539 ^ n_4467;
assign n_5846 = n_4468 ^ n_1540;
assign n_5847 = n_1541 ^ n_4469;
assign n_5848 = n_4470 ^ n_1542;
assign n_5849 = n_1543 ^ n_4471;
assign n_5850 = n_4472 ^ n_1544;
assign n_5851 = n_4473 ^ n_1545;
assign n_5852 = n_1546 ^ n_4474;
assign n_5853 = n_4475 ^ n_1547;
assign n_5854 = n_1548 ^ n_4476;
assign n_5855 = n_1549 ^ n_4477;
assign n_5856 = n_1550 ^ n_4478;
assign n_5857 = n_1551 ^ n_4479;
assign n_5858 = n_1552 ^ n_4480;
assign n_5859 = n_4481 ^ n_1553;
assign n_5860 = n_4482 ^ n_1554;
assign n_5861 = n_4483 ^ n_1555;
assign n_5862 = n_4484 ^ n_1556;
assign n_5863 = n_4485 ^ n_1557;
assign n_5864 = n_4486 ^ n_1558;
assign n_5865 = n_4487 ^ n_1559;
assign n_5866 = n_4488 ^ n_1560;
assign n_5867 = n_4489 ^ n_1561;
assign n_5868 = n_1562 ^ n_4490;
assign n_5869 = n_1563 ^ n_4491;
assign n_5870 = n_4492 ^ n_1564;
assign n_5871 = n_4493 ^ n_1565;
assign n_5872 = n_1566 ^ n_4494;
assign n_5873 = n_1567 ^ n_4495;
assign n_5874 = n_1568 ^ n_4496;
assign n_5875 = n_1569 ^ n_4497;
assign n_5876 = n_1570 ^ n_4498;
assign n_5877 = n_4499 ^ n_1571;
assign n_5878 = ~n_4501 ^ x43;
assign n_5879 = n_2928 ^ n_4502;
assign n_5880 = x64 & n_4503;
assign n_5881 = n_2998 ^ n_4504;
assign n_5882 = n_1577 ^ n_4505;
assign n_5883 = n_1578 ^ n_4506;
assign n_5884 = n_1579 ^ n_4507;
assign n_5885 = n_1580 ^ n_4508;
assign n_5886 = n_1581 ^ n_4509;
assign n_5887 = n_1582 ^ n_4510;
assign n_5888 = n_1583 ^ n_4511;
assign n_5889 = n_1584 ^ n_4512;
assign n_5890 = n_4513 ^ n_1585;
assign n_5891 = n_1586 ^ n_4514;
assign n_5892 = n_1587 ^ n_4515;
assign n_5893 = n_1588 ^ n_4516;
assign n_5894 = n_1589 ^ n_4517;
assign n_5895 = n_4518 ^ n_1590;
assign n_5896 = n_4519 ^ n_1591;
assign n_5897 = n_1592 ^ n_4520;
assign n_5898 = n_4521 ^ n_1593;
assign n_5899 = n_4522 ^ n_1594;
assign n_5900 = n_4523 ^ n_1595;
assign n_5901 = n_4524 ^ n_1596;
assign n_5902 = n_4525 ^ n_1597;
assign n_5903 = n_1598 ^ n_4526;
assign n_5904 = n_4527 ^ n_1599;
assign n_5905 = n_1600 ^ n_4528;
assign n_5906 = n_1601 ^ n_4529;
assign n_5907 = n_4530 ^ n_1602;
assign n_5908 = n_1603 ^ n_4531;
assign n_5909 = n_4532 ^ n_1604;
assign n_5910 = n_4533 ^ n_1605;
assign n_5911 = n_4534 ^ n_1606;
assign n_5912 = n_4535 ^ n_1607;
assign n_5913 = n_1608 ^ n_4536;
assign n_5914 = n_1609 ^ n_4537;
assign n_5915 = n_4538 ^ n_1610;
assign n_5916 = n_1611 ^ n_4539;
assign n_5917 = n_4540 ^ n_1612;
assign n_5918 = n_1613 ^ n_4541;
assign n_5919 = n_4542 ^ n_1614;
assign n_5920 = n_4543 ^ n_1615;
assign n_5921 = n_4544 ^ n_1616;
assign n_5922 = n_1617 ^ n_4545;
assign n_5923 = n_1618 ^ n_4546;
assign n_5924 = n_1619 ^ n_4547;
assign n_5925 = n_1620 ^ n_4548;
assign n_5926 = n_1621 ^ n_4549;
assign n_5927 = n_4550 ^ n_1622;
assign n_5928 = n_4551 ^ n_1623;
assign n_5929 = n_1624 ^ n_4552;
assign n_5930 = n_4553 ^ n_1625;
assign n_5931 = n_4554 ^ n_1626;
assign n_5932 = n_1627 ^ n_4555;
assign n_5933 = n_1628 ^ n_4556;
assign n_5934 = n_1629 ^ n_4557;
assign n_5935 = n_1630 ^ n_4558;
assign n_5936 = n_4559 ^ n_1631;
assign n_5937 = n_4560 ^ n_1632;
assign n_5938 = n_4561 ^ n_1633;
assign n_5939 = n_1634 ^ n_4562;
assign n_5940 = n_4563 ^ n_1635;
assign n_5941 = n_1636 ^ n_4564;
assign n_5942 = ~n_4566 ^ x46;
assign n_5943 = n_2997 ^ n_4567;
assign n_5944 = n_1642 ^ n_4568;
assign n_5945 = n_1643 ^ n_4569;
assign n_5946 = n_1644 ^ n_4570;
assign n_5947 = n_1645 ^ n_4571;
assign n_5948 = n_1646 ^ n_4572;
assign n_5949 = n_1647 ^ n_4573;
assign n_5950 = n_1648 ^ n_4574;
assign n_5951 = n_1649 ^ n_4575;
assign n_5952 = n_4576 ^ n_1650;
assign n_5953 = n_4577 ^ n_1651;
assign n_5954 = n_1652 ^ n_4578;
assign n_5955 = n_1653 ^ n_4579;
assign n_5956 = n_4580 ^ n_1654;
assign n_5957 = n_1655 ^ n_4581;
assign n_5958 = n_1656 ^ n_4582;
assign n_5959 = n_1657 ^ n_4583;
assign n_5960 = n_4584 ^ n_1658;
assign n_5961 = n_1659 ^ n_4585;
assign n_5962 = n_4586 ^ n_1660;
assign n_5963 = n_4587 ^ n_1661;
assign n_5964 = n_4588 ^ n_1662;
assign n_5965 = n_4589 ^ n_1663;
assign n_5966 = n_1664 ^ n_4590;
assign n_5967 = n_1665 ^ n_4591;
assign n_5968 = n_1666 ^ n_4592;
assign n_5969 = n_4593 ^ n_1667;
assign n_5970 = n_4594 ^ n_1668;
assign n_5971 = n_4595 ^ n_1669;
assign n_5972 = n_1670 ^ n_4596;
assign n_5973 = n_1671 ^ n_4597;
assign n_5974 = n_1672 ^ n_4598;
assign n_5975 = n_4599 ^ n_1673;
assign n_5976 = n_4600 ^ n_1674;
assign n_5977 = n_4601 ^ n_1675;
assign n_5978 = n_1676 ^ n_4602;
assign n_5979 = n_4603 ^ n_1677;
assign n_5980 = n_4604 ^ n_1678;
assign n_5981 = n_1679 ^ n_4605;
assign n_5982 = n_1680 ^ n_4606;
assign n_5983 = n_4607 ^ n_1681;
assign n_5984 = n_1682 ^ n_4608;
assign n_5985 = n_1683 ^ n_4609;
assign n_5986 = n_1684 ^ n_4610;
assign n_5987 = n_1685 ^ n_4611;
assign n_5988 = n_1686 ^ n_4612;
assign n_5989 = n_1687 ^ n_4613;
assign n_5990 = n_1688 ^ n_4614;
assign n_5991 = n_1689 ^ n_4615;
assign n_5992 = n_4616 ^ n_1690;
assign n_5993 = n_4617 ^ n_1691;
assign n_5994 = n_4618 ^ n_1692;
assign n_5995 = n_4619 ^ n_1693;
assign n_5996 = n_1694 ^ n_4620;
assign n_5997 = n_1695 ^ n_4621;
assign n_5998 = n_1696 ^ n_4622;
assign n_5999 = n_1697 ^ n_4623;
assign n_6000 = n_1698 ^ n_4624;
assign n_6001 = n_1699 ^ n_4625;
assign n_6002 = n_1700 ^ n_4626;
assign n_6003 = n_4627 ^ n_1701;
assign n_6004 = n_1702 ^ n_4628;
assign n_6005 = ~n_4630 ^ x49;
assign n_6006 = n_3063 ^ n_4631;
assign n_6007 = x64 & n_4632;
assign n_6008 = n_4633 ^ n_1707;
assign n_6009 = n_1708 ^ n_4634;
assign n_6010 = n_4635 ^ n_1709;
assign n_6011 = n_1710 ^ n_4636;
assign n_6012 = n_1711 ^ n_4637;
assign n_6013 = n_4638 ^ n_1712;
assign n_6014 = n_1713 ^ n_4639;
assign n_6015 = n_1714 ^ n_4640;
assign n_6016 = n_1715 ^ n_4641;
assign n_6017 = n_1716 ^ n_4642;
assign n_6018 = n_1717 ^ n_4643;
assign n_6019 = n_1718 ^ n_4644;
assign n_6020 = n_1719 ^ n_4645;
assign n_6021 = n_1720 ^ n_4646;
assign n_6022 = n_1721 ^ n_4647;
assign n_6023 = n_1722 ^ n_4648;
assign n_6024 = n_1723 ^ n_4649;
assign n_6025 = n_1724 ^ n_4650;
assign n_6026 = n_1725 ^ n_4651;
assign n_6027 = n_1726 ^ n_4652;
assign n_6028 = n_4653 ^ n_1727;
assign n_6029 = n_1728 ^ n_4654;
assign n_6030 = n_1729 ^ n_4655;
assign n_6031 = n_1730 ^ n_4656;
assign n_6032 = n_1731 ^ n_4657;
assign n_6033 = n_1732 ^ n_4658;
assign n_6034 = n_1733 ^ n_4659;
assign n_6035 = n_1734 ^ n_4660;
assign n_6036 = n_1735 ^ n_4661;
assign n_6037 = n_4662 ^ n_1736;
assign n_6038 = n_1737 ^ n_4663;
assign n_6039 = n_1738 ^ n_4664;
assign n_6040 = n_1739 ^ n_4665;
assign n_6041 = n_1740 ^ n_4666;
assign n_6042 = n_1741 ^ n_4667;
assign n_6043 = n_1742 ^ n_4668;
assign n_6044 = n_4669 ^ n_1743;
assign n_6045 = n_1744 ^ n_4670;
assign n_6046 = n_4671 ^ n_1745;
assign n_6047 = n_1746 ^ n_4672;
assign n_6048 = n_1747 ^ n_4673;
assign n_6049 = n_1748 ^ n_4674;
assign n_6050 = n_4675 ^ n_1749;
assign n_6051 = n_4676 ^ n_1750;
assign n_6052 = n_1751 ^ n_4677;
assign n_6053 = n_1752 ^ n_4678;
assign n_6054 = n_1753 ^ n_4679;
assign n_6055 = n_1754 ^ n_4680;
assign n_6056 = n_1755 ^ n_4681;
assign n_6057 = n_1756 ^ n_4682;
assign n_6058 = n_1757 ^ n_4683;
assign n_6059 = n_4684 ^ n_1758;
assign n_6060 = n_1759 ^ n_4685;
assign n_6061 = n_1760 ^ n_4686;
assign n_6062 = n_1761 ^ n_4687;
assign n_6063 = n_1762 ^ n_4688;
assign n_6064 = n_1763 ^ n_4689;
assign n_6065 = n_4690 ^ n_1764;
assign n_6066 = n_4691 ^ n_1765;
assign n_6067 = n_1766 ^ n_4692;
assign n_6068 = n_1767 ^ n_4693;
assign n_6069 = ~n_4695 ^ x52;
assign n_6070 = n_3132 ^ n_4696;
assign n_6071 = n_4697 ^ n_3260;
assign n_6072 = n_3197 ^ n_4698;
assign n_6073 = n_4699 ^ n_1772;
assign n_6074 = n_4700 ^ n_1773;
assign n_6075 = n_4701 ^ n_1774;
assign n_6076 = n_4702 ^ n_1775;
assign n_6077 = n_4703 ^ n_1776;
assign n_6078 = n_4704 ^ n_1777;
assign n_6079 = n_4705 ^ n_1778;
assign n_6080 = n_4706 ^ n_1779;
assign n_6081 = n_4707 ^ n_1780;
assign n_6082 = n_4708 ^ n_1781;
assign n_6083 = n_4709 ^ n_1782;
assign n_6084 = n_4710 ^ n_1783;
assign n_6085 = n_4711 ^ n_1784;
assign n_6086 = n_4712 ^ n_1785;
assign n_6087 = n_4713 ^ n_1786;
assign n_6088 = n_4714 ^ n_1787;
assign n_6089 = n_4715 ^ n_1788;
assign n_6090 = n_4716 ^ n_1789;
assign n_6091 = n_4717 ^ n_1790;
assign n_6092 = n_4718 ^ n_1791;
assign n_6093 = n_4719 ^ n_1792;
assign n_6094 = n_4720 ^ n_1793;
assign n_6095 = n_4721 ^ n_1794;
assign n_6096 = n_4722 ^ n_1795;
assign n_6097 = n_4723 ^ n_1796;
assign n_6098 = n_4724 ^ n_1797;
assign n_6099 = n_4725 ^ n_1798;
assign n_6100 = n_4726 ^ n_1799;
assign n_6101 = n_4727 ^ n_1800;
assign n_6102 = n_4728 ^ n_1801;
assign n_6103 = n_4729 ^ n_1802;
assign n_6104 = n_4730 ^ n_1803;
assign n_6105 = n_4731 ^ n_1804;
assign n_6106 = n_4732 ^ n_1805;
assign n_6107 = n_4733 ^ n_1806;
assign n_6108 = n_4734 ^ n_1807;
assign n_6109 = n_4735 ^ n_1808;
assign n_6110 = n_4736 ^ n_1809;
assign n_6111 = n_4737 ^ n_1810;
assign n_6112 = n_4738 ^ n_1811;
assign n_6113 = n_4739 ^ n_1812;
assign n_6114 = n_4740 ^ n_1813;
assign n_6115 = n_4741 ^ n_1814;
assign n_6116 = n_4742 ^ n_1815;
assign n_6117 = n_4743 ^ n_1816;
assign n_6118 = n_4744 ^ n_1817;
assign n_6119 = n_4745 ^ n_1818;
assign n_6120 = n_4746 ^ n_1819;
assign n_6121 = n_4747 ^ n_1820;
assign n_6122 = n_4748 ^ n_1821;
assign n_6123 = n_4749 ^ n_1822;
assign n_6124 = n_4750 ^ n_1823;
assign n_6125 = n_4751 ^ n_1824;
assign n_6126 = n_4752 ^ n_1825;
assign n_6127 = n_4753 ^ n_1826;
assign n_6128 = n_4754 ^ n_1827;
assign n_6129 = n_4755 ^ n_1828;
assign n_6130 = n_4756 ^ n_1829;
assign n_6131 = n_4757 ^ n_1830;
assign n_6132 = n_4758 ^ n_1831;
assign n_6133 = n_4761 ^ n_3325;
assign n_6134 = n_3262 ^ n_4762;
assign n_6135 = n_4763 ^ n_1836;
assign n_6136 = n_4764 ^ n_1837;
assign n_6137 = n_4765 ^ n_1838;
assign n_6138 = n_4766 ^ n_1839;
assign n_6139 = n_4767 ^ n_1840;
assign n_6140 = n_4768 ^ n_1841;
assign n_6141 = n_4769 ^ n_1842;
assign n_6142 = n_4770 ^ n_1843;
assign n_6143 = n_4771 ^ n_1844;
assign n_6144 = n_4772 ^ n_1845;
assign n_6145 = n_4773 ^ n_1846;
assign n_6146 = n_4774 ^ n_1847;
assign n_6147 = n_4775 ^ n_1848;
assign n_6148 = n_4776 ^ n_1849;
assign n_6149 = n_4777 ^ n_1850;
assign n_6150 = n_4778 ^ n_1851;
assign n_6151 = n_4779 ^ n_1852;
assign n_6152 = n_4780 ^ n_1853;
assign n_6153 = n_4781 ^ n_1854;
assign n_6154 = n_4782 ^ n_1855;
assign n_6155 = n_4783 ^ n_1856;
assign n_6156 = n_1857 ^ n_4784;
assign n_6157 = n_4785 ^ n_1858;
assign n_6158 = n_4786 ^ n_1859;
assign n_6159 = n_4787 ^ n_1860;
assign n_6160 = n_4788 ^ n_1861;
assign n_6161 = n_4789 ^ n_1862;
assign n_6162 = n_4790 ^ n_1863;
assign n_6163 = n_4791 ^ n_1864;
assign n_6164 = n_4792 ^ n_1865;
assign n_6165 = n_4793 ^ n_1866;
assign n_6166 = n_4794 ^ n_1867;
assign n_6167 = n_4795 ^ n_1868;
assign n_6168 = n_4796 ^ n_1869;
assign n_6169 = n_4797 ^ n_1870;
assign n_6170 = n_4798 ^ n_1871;
assign n_6171 = n_4799 ^ n_1872;
assign n_6172 = n_4800 ^ n_1873;
assign n_6173 = n_4801 ^ n_1874;
assign n_6174 = n_4802 ^ n_1875;
assign n_6175 = n_4803 ^ n_1876;
assign n_6176 = n_4804 ^ n_1877;
assign n_6177 = n_4805 ^ n_1878;
assign n_6178 = n_4806 ^ n_1879;
assign n_6179 = n_4807 ^ n_1880;
assign n_6180 = n_4808 ^ n_1881;
assign n_6181 = n_4809 ^ n_1882;
assign n_6182 = n_4810 ^ n_1883;
assign n_6183 = n_4811 ^ n_1884;
assign n_6184 = n_4812 ^ n_1885;
assign n_6185 = n_4813 ^ n_1886;
assign n_6186 = n_4814 ^ n_1887;
assign n_6187 = n_4815 ^ n_1888;
assign n_6188 = n_4816 ^ n_1889;
assign n_6189 = n_4817 ^ n_1890;
assign n_6190 = n_4818 ^ n_1891;
assign n_6191 = n_4819 ^ n_1892;
assign n_6192 = n_4820 ^ n_1893;
assign n_6193 = n_4821 ^ n_1894;
assign n_6194 = n_4822 ^ n_1895;
assign n_6195 = n_4825 ^ n_3390;
assign n_6196 = n_3327 ^ n_4826;
assign n_6197 = n_4827 ^ n_1900;
assign n_6198 = n_4828 ^ n_1901;
assign n_6199 = n_4829 ^ n_1902;
assign n_6200 = n_4830 ^ n_1903;
assign n_6201 = n_4831 ^ n_1904;
assign n_6202 = n_4832 ^ n_1905;
assign n_6203 = n_4833 ^ n_1906;
assign n_6204 = n_4834 ^ n_1907;
assign n_6205 = n_4835 ^ n_1908;
assign n_6206 = n_4836 ^ n_1909;
assign n_6207 = n_4837 ^ n_1910;
assign n_6208 = n_4838 ^ n_1911;
assign n_6209 = n_4839 ^ n_1912;
assign n_6210 = n_4840 ^ n_1913;
assign n_6211 = n_4841 ^ n_1914;
assign n_6212 = n_4842 ^ n_1915;
assign n_6213 = n_4843 ^ n_1916;
assign n_6214 = n_4844 ^ n_1917;
assign n_6215 = n_4845 ^ n_1918;
assign n_6216 = n_4846 ^ n_1919;
assign n_6217 = n_4847 ^ n_1920;
assign n_6218 = n_4848 ^ n_1921;
assign n_6219 = n_4849 ^ n_1922;
assign n_6220 = n_4850 ^ n_1923;
assign n_6221 = n_4851 ^ n_1924;
assign n_6222 = n_4852 ^ n_1925;
assign n_6223 = n_4853 ^ n_1926;
assign n_6224 = n_4854 ^ n_1927;
assign n_6225 = n_4855 ^ n_1928;
assign n_6226 = n_4856 ^ n_1929;
assign n_6227 = n_4857 ^ n_1930;
assign n_6228 = n_4858 ^ n_1931;
assign n_6229 = n_4859 ^ n_1932;
assign n_6230 = n_4860 ^ n_1933;
assign n_6231 = n_4861 ^ n_1934;
assign n_6232 = n_4862 ^ n_1935;
assign n_6233 = n_4863 ^ n_1936;
assign n_6234 = n_4864 ^ n_1937;
assign n_6235 = n_4865 ^ n_1938;
assign n_6236 = n_4866 ^ n_1939;
assign n_6237 = n_4867 ^ n_1940;
assign n_6238 = n_4868 ^ n_1941;
assign n_6239 = n_4869 ^ n_1942;
assign n_6240 = n_4870 ^ n_1943;
assign n_6241 = n_4871 ^ n_1944;
assign n_6242 = n_4872 ^ n_1945;
assign n_6243 = n_4873 ^ n_1946;
assign n_6244 = n_4874 ^ n_1947;
assign n_6245 = n_4875 ^ n_1948;
assign n_6246 = n_4876 ^ n_1949;
assign n_6247 = n_4877 ^ n_1950;
assign n_6248 = n_4878 ^ n_1951;
assign n_6249 = n_4879 ^ n_1952;
assign n_6250 = n_4880 ^ n_1953;
assign n_6251 = n_4881 ^ n_1954;
assign n_6252 = n_4882 ^ n_1955;
assign n_6253 = n_4883 ^ n_1956;
assign n_6254 = n_4884 ^ n_1957;
assign n_6255 = n_4885 ^ n_1958;
assign n_6256 = n_4886 ^ n_1959;
assign n_6257 = n_4889 ^ x70;
assign n_6258 = n_4890 ^ n_1961;
assign n_6259 = n_488 & n_4891;
assign n_6260 = n_4891 & ~n_124;
assign n_6261 = n_488 & n_4894;
assign n_6262 = n_4894 & ~n_152;
assign n_6263 = n_4895 ^ n_1965;
assign n_6264 = n_4896 ^ x82;
assign n_6265 = n_488 & n_4897;
assign n_6266 = n_4897 & ~n_163;
assign n_6267 = n_488 & n_4898;
assign n_6268 = n_4898 & ~n_174;
assign n_6269 = n_4899 ^ n_1969;
assign n_6270 = n_4900 ^ x88;
assign n_6271 = n_488 & n_4901;
assign n_6272 = n_4901 & ~n_184;
assign n_6273 = n_488 & n_4902;
assign n_6274 = n_4902 & ~n_197;
assign n_6275 = n_4903 ^ x94;
assign n_6276 = n_4904 ^ n_1972;
assign n_6277 = n_488 & n_4905;
assign n_6278 = n_4905 & ~n_208;
assign n_6279 = n_4906 ^ x97;
assign n_6280 = n_4907 ^ n_1974;
assign n_6281 = n_488 & n_4908;
assign n_6282 = n_4908 & ~n_219;
assign n_6283 = n_4910 ^ n_1976;
assign n_6284 = n_4911 ^ x109;
assign n_6285 = n_4912 ^ n_1977;
assign n_6286 = n_488 & n_4913;
assign n_6287 = n_4913 & ~n_256;
assign n_6288 = n_4914 ^ n_1979;
assign n_6289 = n_4915 ^ x115;
assign n_6290 = n_488 & n_4916;
assign n_6291 = n_4916 & ~n_271;
assign n_6292 = n_4917 ^ n_1981;
assign n_6293 = n_4918 ^ x121;
assign n_6294 = n_488 & n_4919;
assign n_6295 = n_4919 & ~n_288;
assign n_6296 = n_3662 ^ n_4921;
assign n_6297 = n_4922 & n_1;
assign n_6298 = n_4922 ^ n_529;
assign n_6299 = n_4922 ^ x67;
assign n_6300 = ~n_4922 & ~n_29;
assign n_6301 = ~n_4922 & ~n_44;
assign n_6302 = ~n_4922 & n_50;
assign n_6303 = ~n_4922 & n_59;
assign n_6304 = ~n_4922 & n_62;
assign n_6305 = ~n_4922 & n_65;
assign n_6306 = n_4923 ^ n_528;
assign n_6307 = ~x68 & ~n_4923;
assign n_6308 = n_4924 ^ n_494;
assign n_6309 = x14 & ~n_4925;
assign n_6310 = ~n_347 & ~n_4927;
assign n_6311 = n_4928 ^ n_1997;
assign n_6312 = ~n_358 & ~n_4929;
assign n_6313 = ~n_364 & ~n_4930;
assign n_6314 = ~n_370 & ~n_4931;
assign n_6315 = ~n_376 & ~n_4932;
assign n_6316 = ~n_382 & ~n_4933;
assign n_6317 = ~n_388 & ~n_4934;
assign n_6318 = ~n_395 & ~n_4935;
assign n_6319 = ~n_401 & ~n_4936;
assign n_6320 = ~n_414 & ~n_4937;
assign n_6321 = ~n_420 & ~n_4938;
assign n_6322 = ~n_426 & ~n_4939;
assign n_6323 = ~n_432 & ~n_4940;
assign n_6324 = ~n_438 & ~n_4941;
assign n_6325 = ~n_444 & ~n_4942;
assign n_6326 = n_4943 ^ x59;
assign n_6327 = ~n_450 & ~n_4943;
assign n_6328 = ~n_489 & ~n_4944;
assign n_6329 = ~n_4945 & n_539;
assign n_6330 = n_4946 ^ n_530;
assign n_6331 = n_4947 ^ n_2022;
assign n_6332 = n_4948 ^ n_2023;
assign n_6333 = ~x62 & ~n_4949;
assign n_6334 = n_7 & n_4952;
assign n_6335 = ~n_66 & n_4953;
assign n_6336 = n_4954 ^ x11;
assign n_6337 = ~n_4954 & ~n_4892;
assign n_6338 = n_4957 ^ n_3465;
assign n_6339 = ~n_4955 & ~n_4958;
assign n_6340 = n_4959 ^ n_551;
assign n_6341 = n_4960 ^ n_2038;
assign n_6342 = ~n_66 & n_4961;
assign n_6343 = n_4962 ^ n_556;
assign n_6344 = ~x86 & n_4963;
assign n_6345 = n_66 & n_4963;
assign n_6346 = n_4964 ^ n_565;
assign n_6347 = n_4965 ^ n_566;
assign n_6348 = n_4967 ^ n_571;
assign n_6349 = n_4968 ^ n_572;
assign n_6350 = n_4969 ^ n_577;
assign n_6351 = ~n_66 & n_4971;
assign n_6352 = n_4972 ^ x38;
assign n_6353 = ~n_4972 & ~n_4909;
assign n_6354 = n_4975 ^ x41;
assign n_6355 = ~n_4975 & ~n_4973;
assign n_6356 = n_4978 ^ n_591;
assign n_6357 = n_4979 ^ n_593;
assign n_6358 = n_4980 ^ x44;
assign n_6359 = ~n_4980 & ~n_4976;
assign n_6360 = n_4983 ^ n_604;
assign n_6361 = n_4984 ^ n_3516;
assign n_6362 = ~n_4981 & ~n_4985;
assign n_6363 = n_4986 ^ n_608;
assign n_6364 = n_4987 ^ x119;
assign n_6365 = n_4988 ^ n_609;
assign n_6366 = ~n_66 & n_4989;
assign n_6367 = n_4991 ^ n_615;
assign n_6368 = n_4992 ^ x62;
assign n_6369 = ~n_66 & n_4993;
assign n_6370 = n_334 ^ n_4994;
assign n_6371 = n_5057 ^ x5;
assign n_6372 = n_492 ^ n_5119;
assign n_6373 = n_5119 ^ n_3662;
assign n_6374 = n_349 ^ n_5120;
assign n_6375 = n_5308 ^ x17;
assign n_6376 = n_5372 ^ x20;
assign n_6377 = n_5436 ^ x23;
assign n_6378 = n_378 ^ n_5437;
assign n_6379 = n_5561 ^ x29;
assign n_6380 = n_5623 ^ x32;
assign n_6381 = n_5687 ^ x35;
assign n_6382 = n_5751 ^ x38;
assign n_6383 = n_503 & n_5753;
assign n_6384 = n_409 ^ n_5754;
assign n_6385 = n_5879 ^ x44;
assign n_6386 = n_5880 ^ n_5943;
assign n_6387 = n_5943 ^ n_3060;
assign n_6388 = n_6006 ^ x50;
assign n_6389 = n_6007 ^ n_498;
assign n_6390 = n_6070 ^ x53;
assign n_6391 = n_440 ^ n_6071;
assign n_6392 = n_446 ^ n_6133;
assign n_6393 = n_452 ^ n_6195;
assign n_6394 = n_458 & n_6257;
assign n_6395 = n_6259 ^ x8;
assign n_6396 = n_6260 ^ x72;
assign n_6397 = n_6261 ^ x17;
assign n_6398 = n_6262 ^ x81;
assign n_6399 = n_463 & n_6264;
assign n_6400 = n_6265 ^ x20;
assign n_6401 = n_6266 ^ x84;
assign n_6402 = n_6267 ^ x23;
assign n_6403 = n_6268 ^ x87;
assign n_6404 = n_467 & n_6270;
assign n_6405 = n_6271 ^ x26;
assign n_6406 = n_6272 ^ x90;
assign n_6407 = n_6273 ^ x29;
assign n_6408 = n_6274 ^ x93;
assign n_6409 = n_469 & n_6275;
assign n_6410 = n_6277 ^ x32;
assign n_6411 = n_6278 ^ x96;
assign n_6412 = n_472 & n_6279;
assign n_6413 = n_6281 ^ x35;
assign n_6414 = n_6282 ^ x99;
assign n_6415 = n_477 & n_6284;
assign n_6416 = n_6286 ^ x47;
assign n_6417 = n_6287 ^ x111;
assign n_6418 = n_481 & n_6289;
assign n_6419 = n_6290 ^ x53;
assign n_6420 = n_6291 ^ x117;
assign n_6421 = n_485 & n_6293;
assign n_6422 = n_6294 ^ x59;
assign n_6423 = n_6295 ^ x123;
assign n_6424 = ~n_339 & n_6296;
assign n_6425 = n_6297 ^ x1;
assign n_6426 = ~n_501 & ~n_6298;
assign n_6427 = n_655 & ~n_6299;
assign n_6428 = ~n_6299 & n_784;
assign n_6429 = ~n_6299 & ~n_3665;
assign n_6430 = ~n_6299 & n_854;
assign n_6431 = ~n_6299 & n_920;
assign n_6432 = ~n_6299 & n_986;
assign n_6433 = ~n_6299 & n_1052;
assign n_6434 = ~n_6299 & n_1181;
assign n_6435 = ~n_6299 & n_1248;
assign n_6436 = ~n_6299 & n_1314;
assign n_6437 = ~n_6299 & n_1380;
assign n_6438 = ~n_6299 & n_1510;
assign n_6439 = ~n_6299 & n_1641;
assign n_6440 = ~n_6299 & n_1706;
assign n_6441 = n_6300 ^ n_6299;
assign n_6442 = n_6301 ^ n_6299;
assign n_6443 = n_6302 ^ x67;
assign n_6444 = n_6303 ^ x67;
assign n_6445 = n_6304 ^ x67;
assign n_6446 = n_6305 ^ x67;
assign n_6447 = n_1 & n_6306;
assign n_6448 = n_6306 ^ x68;
assign n_6449 = n_6307 ^ n_2020;
assign n_6450 = x69 & ~n_6307;
assign n_6451 = n_6308 ^ n_5244;
assign n_6452 = ~n_5244 & n_6309;
assign n_6453 = x11 & n_6310;
assign n_6454 = x17 & n_6312;
assign n_6455 = x20 & n_6313;
assign n_6456 = x23 & n_6314;
assign n_6457 = x26 & n_6315;
assign n_6458 = n_495 ^ n_6316;
assign n_6459 = n_6316 & n_1994;
assign n_6460 = x32 & n_6317;
assign n_6461 = x35 & n_6318;
assign n_6462 = x38 & n_6319;
assign n_6463 = x44 & n_6320;
assign n_6464 = x50 & n_6322;
assign n_6465 = x53 & n_6323;
assign n_6466 = x56 & n_6324;
assign n_6467 = x59 & n_6325;
assign n_6468 = x62 & n_6327;
assign n_6469 = n_6328 ^ n_80;
assign n_6470 = ~n_6329 & n_125;
assign n_6471 = n_6330 ^ x67;
assign n_6472 = n_6331 ^ x2;
assign n_6473 = n_6332 ^ x2;
assign n_6474 = n_6333 ^ n_3457;
assign n_6475 = n_6334 ^ x2;
assign n_6476 = n_6335 ^ n_132;
assign n_6477 = n_6337 ^ x11;
assign n_6478 = n_6339 ^ x14;
assign n_6479 = n_6340 ^ x79;
assign n_6480 = n_6342 ^ n_553;
assign n_6481 = n_6343 ^ x82;
assign n_6482 = n_6346 ^ x90;
assign n_6483 = n_6347 ^ x91;
assign n_6484 = n_6348 ^ x93;
assign n_6485 = ~n_66 & n_6349;
assign n_6486 = n_6350 ^ x99;
assign n_6487 = n_6351 ^ ~n_230;
assign n_6488 = n_6353 ^ x38;
assign n_6489 = n_6355 ^ x41;
assign n_6490 = n_6356 ^ x107;
assign n_6491 = n_6357 ^ x108;
assign n_6492 = n_6359 ^ x44;
assign n_6493 = n_6360 ^ x114;
assign n_6494 = n_6362 ^ x50;
assign n_6495 = n_6363 ^ x115;
assign n_6496 = n_4990 ^ n_6364;
assign n_6497 = n_6364 ^ x56;
assign n_6498 = n_3528 ^ n_6364;
assign n_6499 = n_6365 ^ x118;
assign n_6500 = n_6366 ^ n_281;
assign n_6501 = n_6367 ^ x124;
assign n_6502 = x63 & ~n_6368;
assign n_6503 = n_6369 ^ n_628;
assign n_6504 = n_2121 ^ n_6370;
assign n_6505 = n_2192 ^ n_6374;
assign n_6506 = x64 & ~n_6375;
assign n_6507 = x64 & ~n_6376;
assign n_6508 = x64 & ~n_6377;
assign n_6509 = n_2527 ^ n_6378;
assign n_6510 = x64 & ~n_6380;
assign n_6511 = x64 & ~n_6381;
assign n_6512 = x64 & ~n_6382;
assign n_6513 = n_2862 ^ n_6384;
assign n_6514 = x64 & ~n_6385;
assign n_6515 = n_6321 ^ n_6386;
assign n_6516 = ~n_6386 & n_6321;
assign n_6517 = x64 & ~n_6388;
assign n_6518 = ~n_6389 & n_6390;
assign n_6519 = n_3196 ^ n_6391;
assign n_6520 = n_3261 ^ n_6392;
assign n_6521 = n_3326 ^ n_6393;
assign n_6522 = n_6394 ^ n_121;
assign n_6523 = n_488 & n_6396;
assign n_6524 = n_488 & n_6398;
assign n_6525 = ~n_6263 ^ ~n_6399;
assign n_6526 = n_488 & n_6401;
assign n_6527 = n_488 & n_6403;
assign n_6528 = ~n_6269 ^ ~n_6404;
assign n_6529 = n_488 & n_6406;
assign n_6530 = n_488 & n_6408;
assign n_6531 = n_6409 ^ n_205;
assign n_6532 = n_488 & n_6411;
assign n_6533 = n_6412 ^ n_216;
assign n_6534 = n_488 & n_6414;
assign n_6535 = n_6415 ^ n_255;
assign n_6536 = n_488 & n_6417;
assign n_6537 = ~n_6288 ^ ~n_6418;
assign n_6538 = n_488 & n_6420;
assign n_6539 = ~n_6292 ^ ~n_6421;
assign n_6540 = n_488 & n_6423;
assign n_6541 = n_6424 ^ n_6372;
assign n_6542 = n_6425 ^ x67;
assign n_6543 = n_490 & n_6426;
assign n_6544 = n_6427 ^ n_2122;
assign n_6545 = n_6428 ^ n_722;
assign n_6546 = n_6429 ^ n_2193;
assign n_6547 = n_6430 ^ n_2261;
assign n_6548 = n_6431 ^ n_2328;
assign n_6549 = n_6432 ^ n_2395;
assign n_6550 = n_6433 ^ n_2462;
assign n_6551 = n_6434 ^ n_2593;
assign n_6552 = n_6435 ^ n_2660;
assign n_6553 = n_6436 ^ n_2728;
assign n_6554 = n_6437 ^ n_2795;
assign n_6555 = n_6438 ^ n_2929;
assign n_6556 = n_6439 ^ n_3064;
assign n_6557 = n_6440 ^ n_3133;
assign n_6558 = n_27 & ~n_6441;
assign n_6559 = n_42 & ~n_6442;
assign n_6560 = n_48 & n_6443;
assign n_6561 = n_57 & n_6444;
assign n_6562 = n_60 & n_6445;
assign n_6563 = n_63 & n_6446;
assign n_6564 = n_6447 ^ x1;
assign n_6565 = n_655 & ~n_6448;
assign n_6566 = ~n_6448 & n_784;
assign n_6567 = ~n_6448 & ~n_3665;
assign n_6568 = ~n_6448 & n_854;
assign n_6569 = ~n_6448 & n_920;
assign n_6570 = ~n_6448 & n_986;
assign n_6571 = ~n_6448 & n_1052;
assign n_6572 = ~n_6448 & n_1117;
assign n_6573 = ~n_6448 & n_1181;
assign n_6574 = ~n_6448 & n_1248;
assign n_6575 = ~n_6448 & n_1314;
assign n_6576 = ~n_6448 & n_1380;
assign n_6577 = ~n_6448 & n_1445;
assign n_6578 = ~n_6448 & n_1510;
assign n_6579 = ~n_6448 & n_1576;
assign n_6580 = ~n_6448 & n_1641;
assign n_6581 = ~n_6448 & n_1706;
assign n_6582 = ~n_6448 & n_1771;
assign n_6583 = ~n_6448 & n_1835;
assign n_6584 = ~n_6448 & n_1899;
assign n_6585 = n_1 & n_6449;
assign n_6586 = n_6449 ^ x69;
assign n_6587 = n_6450 ^ n_3451;
assign n_6588 = ~x70 & ~n_6450;
assign n_6589 = n_6452 ^ n_358;
assign n_6590 = ~n_358 & ~n_6452;
assign n_6591 = n_6457 ^ x26;
assign n_6592 = ~n_5561 & n_6458;
assign n_6593 = ~n_5561 & n_6459;
assign n_6594 = n_6466 ^ x56;
assign n_6595 = n_6467 ^ x59;
assign n_6596 = n_6468 ^ x62;
assign n_6597 = ~n_524 ^ n_6469;
assign n_6598 = n_6470 ^ x73;
assign n_6599 = n_6474 ^ x2;
assign n_6600 = n_6475 ^ n_3391;
assign n_6601 = n_1960 ^ n_6476;
assign n_6602 = n_6477 ^ n_3465;
assign n_6603 = n_6478 ^ n_6341;
assign n_6604 = n_6485 ^ n_572;
assign n_6605 = ~n_6487 & ~n_6283;
assign n_6606 = n_6488 ^ n_3502;
assign n_6607 = n_6489 ^ n_3506;
assign n_6608 = n_6492 ^ n_3414;
assign n_6609 = n_6494 ^ n_3417;
assign n_6610 = ~n_6497 & ~n_6498;
assign n_6611 = ~n_482 & n_6499;
assign n_6612 = n_6502 ^ n_4920;
assign n_6613 = n_6371 ^ n_6504;
assign n_6614 = ~n_6504 & n_5057;
assign n_6615 = n_493 ^ n_6505;
assign n_6616 = n_6505 ^ n_2257;
assign n_6617 = n_917 & n_6506;
assign n_6618 = n_983 & n_6507;
assign n_6619 = n_1049 & n_6508;
assign n_6620 = ~n_6509 & n_6457;
assign n_6621 = n_1244 & n_6510;
assign n_6622 = n_1311 & n_6511;
assign n_6623 = n_1377 & n_6512;
assign n_6624 = n_6383 ^ n_6513;
assign n_6625 = ~n_6513 & ~n_6383;
assign n_6626 = n_1507 & n_6514;
assign n_6627 = n_6515 ^ n_6387;
assign n_6628 = x47 & n_6516;
assign n_6629 = n_1638 & n_6517;
assign n_6630 = n_6518 ^ n_6007;
assign n_6631 = ~n_6519 & n_6466;
assign n_6632 = ~n_6520 & n_6467;
assign n_6633 = ~n_6521 & n_6468;
assign n_6634 = n_6522 ^ n_6258;
assign n_6635 = n_6523 ^ n_3394;
assign n_6636 = n_6524 ^ n_3397;
assign n_6637 = n_6526 ^ n_3400;
assign n_6638 = n_6527 ^ n_3402;
assign n_6639 = n_6529 ^ n_3486;
assign n_6640 = n_6530 ^ n_3406;
assign n_6641 = n_6531 ^ n_6276;
assign n_6642 = n_6532 ^ n_3409;
assign n_6643 = n_6533 ^ n_6280;
assign n_6644 = n_6534 ^ n_3412;
assign n_6645 = n_6535 ^ n_6285;
assign n_6646 = n_6536 ^ n_3516;
assign n_6647 = n_6538 ^ n_6364;
assign n_6648 = n_6540 ^ n_3423;
assign n_6649 = n_6541 ^ n_6373;
assign n_6650 = x8 & n_6541;
assign n_6651 = n_3449 ^ n_6542;
assign n_6652 = n_6543 ^ n_490;
assign n_6653 = n_4995 ^ n_6544;
assign n_6654 = n_5058 ^ n_6545;
assign n_6655 = n_5121 ^ n_6546;
assign n_6656 = n_5182 ^ n_6547;
assign n_6657 = n_5246 ^ n_6548;
assign n_6658 = n_5310 ^ n_6549;
assign n_6659 = n_5374 ^ n_6550;
assign n_6660 = n_5499 ^ n_6551;
assign n_6661 = n_5562 ^ n_6552;
assign n_6662 = n_5625 ^ n_6553;
assign n_6663 = n_5689 ^ n_6554;
assign n_6664 = n_5817 ^ n_6555;
assign n_6665 = n_5944 ^ n_6556;
assign n_6666 = n_6008 ^ n_6557;
assign n_6667 = ~n_6558 ^ ~n_5438;
assign n_6668 = ~n_6559 ^ ~n_5755;
assign n_6669 = ~n_6560 ^ ~n_5881;
assign n_6670 = ~n_6561 ^ ~n_6072;
assign n_6671 = ~n_6562 ^ ~n_6134;
assign n_6672 = ~n_6563 ^ ~n_6196;
assign n_6673 = n_6564 ^ x68;
assign n_6674 = n_6565 ^ n_2123;
assign n_6675 = n_6566 ^ n_723;
assign n_6676 = n_6567 ^ n_2194;
assign n_6677 = n_6568 ^ n_2262;
assign n_6678 = n_6569 ^ n_2329;
assign n_6679 = n_6570 ^ n_2396;
assign n_6680 = n_6571 ^ n_2463;
assign n_6681 = n_6572 ^ n_2529;
assign n_6682 = n_6573 ^ n_2594;
assign n_6683 = n_6574 ^ n_2661;
assign n_6684 = n_6575 ^ n_2729;
assign n_6685 = n_6576 ^ n_2796;
assign n_6686 = n_6577 ^ n_2864;
assign n_6687 = n_6578 ^ n_2930;
assign n_6688 = n_6579 ^ n_2999;
assign n_6689 = n_6580 ^ n_3065;
assign n_6690 = n_6581 ^ n_3134;
assign n_6691 = n_6582 ^ n_3198;
assign n_6692 = n_6583 ^ n_3263;
assign n_6693 = n_6584 ^ n_3328;
assign n_6694 = n_6585 ^ x1;
assign n_6695 = n_655 & ~n_6586;
assign n_6696 = ~n_6586 & n_784;
assign n_6697 = ~n_6586 & ~n_3665;
assign n_6698 = ~n_6586 & n_854;
assign n_6699 = ~n_6586 & n_920;
assign n_6700 = ~n_6586 & n_986;
assign n_6701 = ~n_6586 & n_1052;
assign n_6702 = ~n_6586 & n_1117;
assign n_6703 = ~n_6586 & n_1181;
assign n_6704 = ~n_6586 & n_1248;
assign n_6705 = ~n_6586 & n_1314;
assign n_6706 = ~n_6586 & n_1380;
assign n_6707 = ~n_6586 & n_1445;
assign n_6708 = ~n_6586 & n_1510;
assign n_6709 = ~n_6586 & n_1576;
assign n_6710 = ~n_6586 & n_1641;
assign n_6711 = ~n_6586 & n_1706;
assign n_6712 = ~n_6586 & n_1771;
assign n_6713 = ~n_6586 & n_1835;
assign n_6714 = ~n_6586 & n_1899;
assign n_6715 = n_1 & n_6587;
assign n_6716 = n_6587 ^ x70;
assign n_6717 = n_6588 ^ n_4945;
assign n_6718 = ~n_6588 & n_120;
assign n_6719 = n_6591 ^ n_6509;
assign n_6720 = n_6592 ^ n_6316;
assign n_6721 = n_388 ^ n_6593;
assign n_6722 = ~n_6593 & ~n_388;
assign n_6723 = n_6594 ^ n_6519;
assign n_6724 = n_6595 ^ n_6520;
assign n_6725 = n_6596 ^ n_6521;
assign y2 = ~n_6597;
assign n_6726 = x74 & n_6598;
assign n_6727 = ~n_6604 ^ ~n_4966;
assign n_6728 = n_6610 ^ x56;
assign n_6729 = ~n_6500 ^ ~n_6611;
assign n_6730 = ~n_6614 & ~n_339;
assign n_6731 = n_6453 & ~n_6615;
assign n_6732 = n_6615 ^ n_6616;
assign n_6733 = n_6617 ^ n_6375;
assign n_6734 = n_6618 ^ n_6376;
assign n_6735 = n_6619 ^ n_6377;
assign n_6736 = n_6620 ^ n_382;
assign n_6737 = ~n_382 & ~n_6620;
assign n_6738 = n_6621 ^ n_6380;
assign n_6739 = n_6622 ^ n_6381;
assign n_6740 = n_6623 ^ n_6382;
assign n_6741 = x41 & ~n_6625;
assign n_6742 = n_6626 ^ n_6385;
assign n_6743 = ~x47 & ~n_6627;
assign n_6744 = n_6628 ^ n_426;
assign n_6745 = ~n_426 & ~n_6628;
assign n_6746 = n_6629 ^ n_6388;
assign n_6747 = n_6630 ^ n_6465;
assign n_6748 = n_6465 & n_6630;
assign n_6749 = ~n_444 & ~n_6631;
assign n_6750 = n_450 ^ n_6632;
assign n_6751 = ~n_6632 & ~n_450;
assign n_6752 = n_6634 ^ n_121;
assign n_6753 = n_6641 ^ n_205;
assign n_6754 = n_6643 ^ n_216;
assign n_6755 = n_6645 ^ n_255;
assign n_6756 = ~x8 & n_6649;
assign n_6757 = ~n_6372 & n_6650;
assign n_6758 = ~x0 & n_6651;
assign n_6759 = n_6653 ^ x5;
assign n_6760 = n_6654 ^ x8;
assign n_6761 = n_6655 ^ x11;
assign n_6762 = n_6656 ^ x14;
assign n_6763 = n_6657 ^ x17;
assign n_6764 = n_6658 ^ x20;
assign n_6765 = n_6659 ^ x23;
assign n_6766 = n_6660 ^ x29;
assign n_6767 = n_6661 ^ x32;
assign n_6768 = n_6662 ^ x35;
assign n_6769 = n_6663 ^ x38;
assign n_6770 = n_6664 ^ x44;
assign n_6771 = n_6665 ^ x50;
assign n_6772 = n_6666 ^ x53;
assign n_6773 = ~n_6667 ^ x26;
assign n_6774 = ~n_6668 ^ x41;
assign n_6775 = ~n_6669 ^ x47;
assign n_6776 = ~n_6670 ^ x56;
assign n_6777 = ~n_6671 ^ x59;
assign n_6778 = ~n_6672 ^ x62;
assign n_6779 = ~n_6672 & n_6633;
assign n_6780 = n_6673 ^ n_2100;
assign n_6781 = n_4996 ^ n_6674;
assign n_6782 = n_5059 ^ n_6675;
assign n_6783 = n_5122 ^ n_6676;
assign n_6784 = n_5183 ^ n_6677;
assign n_6785 = n_5247 ^ n_6678;
assign n_6786 = n_5311 ^ n_6679;
assign n_6787 = n_5375 ^ n_6680;
assign n_6788 = n_5439 ^ n_6681;
assign n_6789 = n_5500 ^ n_6682;
assign n_6790 = n_5563 ^ n_6683;
assign n_6791 = n_5626 ^ n_6684;
assign n_6792 = n_5690 ^ n_6685;
assign n_6793 = n_5756 ^ n_6686;
assign n_6794 = n_5818 ^ n_6687;
assign n_6795 = n_5882 ^ n_6688;
assign n_6796 = n_5945 ^ n_6689;
assign n_6797 = n_6009 ^ n_6690;
assign n_6798 = n_6073 ^ n_6691;
assign n_6799 = n_6135 ^ n_6692;
assign n_6800 = n_6197 ^ n_6693;
assign n_6801 = n_6694 ^ x69;
assign n_6802 = n_6695 ^ n_2124;
assign n_6803 = n_6696 ^ n_724;
assign n_6804 = n_6697 ^ n_2195;
assign n_6805 = n_6698 ^ n_2263;
assign n_6806 = n_6699 ^ n_2330;
assign n_6807 = n_6700 ^ n_2397;
assign n_6808 = n_6701 ^ n_2464;
assign n_6809 = n_6702 ^ n_2530;
assign n_6810 = n_6703 ^ n_2595;
assign n_6811 = n_6704 ^ n_2662;
assign n_6812 = n_6705 ^ n_2730;
assign n_6813 = n_6706 ^ n_2797;
assign n_6814 = n_6707 ^ n_2865;
assign n_6815 = n_6708 ^ n_2931;
assign n_6816 = n_6709 ^ n_3000;
assign n_6817 = n_6710 ^ n_3066;
assign n_6818 = n_6711 ^ n_3135;
assign n_6819 = n_6712 ^ n_3199;
assign n_6820 = n_6713 ^ n_3264;
assign n_6821 = n_6714 ^ n_3329;
assign n_6822 = n_6715 ^ x1;
assign n_6823 = n_655 & ~n_6716;
assign n_6824 = n_784 & ~n_6716;
assign n_6825 = ~n_6716 & ~n_3665;
assign n_6826 = ~n_6716 & n_854;
assign n_6827 = ~n_6716 & n_920;
assign n_6828 = ~n_6716 & n_986;
assign n_6829 = ~n_6716 & n_1052;
assign n_6830 = ~n_6716 & n_1117;
assign n_6831 = ~n_6716 & n_1181;
assign n_6832 = ~n_6716 & n_1248;
assign n_6833 = ~n_6716 & n_1314;
assign n_6834 = ~n_6716 & n_1380;
assign n_6835 = ~n_6716 & n_1445;
assign n_6836 = ~n_6716 & n_1510;
assign n_6837 = ~n_6716 & n_1576;
assign n_6838 = ~n_6716 & n_1641;
assign n_6839 = ~n_6716 & n_1706;
assign n_6840 = ~n_6716 & n_1771;
assign n_6841 = ~n_6716 & n_1835;
assign n_6842 = ~n_6716 & n_1899;
assign n_6843 = n_1 & n_6717;
assign n_6844 = n_6717 & n_117;
assign n_6845 = n_6717 ^ x71;
assign n_6846 = n_6718 ^ n_6329;
assign n_6847 = n_6718 ^ x72;
assign n_6848 = ~n_6379 & ~n_6720;
assign n_6849 = ~x75 & ~n_6726;
assign n_6850 = n_6728 ^ n_3420;
assign n_6851 = ~n_6731 & ~n_353;
assign n_6852 = ~x11 & ~n_6732;
assign n_6853 = n_6733 ^ n_5245;
assign n_6854 = n_6734 ^ n_5309;
assign n_6855 = n_6735 ^ n_5373;
assign n_6856 = n_6738 ^ n_4239;
assign n_6857 = n_6739 ^ n_5624;
assign n_6858 = n_6740 ^ n_5688;
assign n_6859 = n_6741 ^ ~n_6668;
assign n_6860 = n_6742 ^ n_5816;
assign n_6861 = n_6743 ^ n_6515;
assign n_6862 = ~n_497 & n_6746;
assign n_6863 = ~n_6748 & ~n_438;
assign n_6864 = n_6750 ^ n_6751;
assign n_6865 = n_6756 ^ n_6541;
assign n_6866 = ~n_6757 & ~n_347;
assign n_6867 = n_6758 ^ n_6542;
assign n_6868 = n_6759 ^ n_339;
assign n_6869 = n_6759 & ~n_6730;
assign n_6870 = n_6760 ^ n_347;
assign n_6871 = n_6761 ^ n_353;
assign n_6872 = n_6762 ^ n_6589;
assign n_6873 = n_6762 & ~n_6590;
assign n_6874 = n_6763 ^ n_364;
assign n_6875 = n_6764 ^ n_370;
assign n_6876 = n_6765 ^ n_376;
assign n_6877 = n_6766 ^ n_6721;
assign n_6878 = n_6766 & ~n_6722;
assign n_6879 = n_6767 ^ n_395;
assign n_6880 = n_6768 ^ n_401;
assign n_6881 = n_6769 ^ n_407;
assign n_6882 = n_6770 ^ n_420;
assign n_6883 = n_6771 ^ n_432;
assign n_6884 = n_6772 ^ n_438;
assign n_6885 = n_6773 ^ n_6736;
assign n_6886 = ~n_6773 & ~n_6737;
assign n_6887 = n_6744 ^ n_6775;
assign n_6888 = ~n_6775 & ~n_6745;
assign n_6889 = n_6776 ^ n_6749;
assign n_6890 = ~n_6749 & ~n_6776;
assign n_6891 = n_6751 ^ n_6777;
assign n_6892 = ~n_6777 & ~n_6751;
assign n_6893 = n_6778 ^ n_456;
assign n_6894 = n_456 & ~n_6778;
assign n_6895 = ~x0 & n_6780;
assign n_6896 = n_6781 ^ x5;
assign n_6897 = n_6782 ^ x8;
assign n_6898 = n_6783 ^ x11;
assign n_6899 = n_6784 ^ x14;
assign n_6900 = n_6785 ^ x17;
assign n_6901 = n_6786 ^ x20;
assign n_6902 = n_6787 ^ x23;
assign n_6903 = n_6788 ^ x26;
assign n_6904 = n_6789 ^ x29;
assign n_6905 = n_6790 ^ x32;
assign n_6906 = n_6791 ^ x35;
assign n_6907 = n_6792 ^ x38;
assign n_6908 = n_6793 ^ x41;
assign n_6909 = n_6794 ^ x44;
assign n_6910 = n_6795 ^ x47;
assign n_6911 = n_6796 ^ x50;
assign n_6912 = n_6797 ^ x53;
assign n_6913 = n_6798 ^ x56;
assign n_6914 = n_6799 ^ x59;
assign n_6915 = n_6326 ^ n_6799;
assign n_6916 = n_6800 ^ x62;
assign n_6917 = n_6471 ^ n_6801;
assign n_6918 = n_4997 ^ n_6802;
assign n_6919 = n_5060 ^ n_6803;
assign n_6920 = n_5123 ^ n_6804;
assign n_6921 = n_5184 ^ n_6805;
assign n_6922 = n_5248 ^ n_6806;
assign n_6923 = n_5312 ^ n_6807;
assign n_6924 = n_5376 ^ n_6808;
assign n_6925 = n_5440 ^ n_6809;
assign n_6926 = n_5501 ^ n_6810;
assign n_6927 = n_5564 ^ n_6811;
assign n_6928 = n_5627 ^ n_6812;
assign n_6929 = n_5691 ^ n_6813;
assign n_6930 = n_5757 ^ n_6814;
assign n_6931 = n_5819 ^ n_6815;
assign n_6932 = n_5883 ^ n_6816;
assign n_6933 = n_5946 ^ n_6817;
assign n_6934 = n_6010 ^ n_6818;
assign n_6935 = n_6074 ^ n_6819;
assign n_6936 = n_6136 ^ n_6820;
assign n_6937 = n_6198 ^ n_6821;
assign n_6938 = n_6822 ^ x70;
assign n_6939 = n_2125 ^ n_6823;
assign n_6940 = n_6824 ^ n_725;
assign n_6941 = n_6825 ^ n_2196;
assign n_6942 = n_6826 ^ n_2264;
assign n_6943 = n_6827 ^ n_2331;
assign n_6944 = n_6828 ^ n_2398;
assign n_6945 = n_6829 ^ n_2465;
assign n_6946 = n_6830 ^ n_2531;
assign n_6947 = n_6831 ^ n_2596;
assign n_6948 = n_6832 ^ n_2663;
assign n_6949 = n_6833 ^ n_2731;
assign n_6950 = n_6834 ^ n_2798;
assign n_6951 = n_6835 ^ n_2866;
assign n_6952 = n_6836 ^ n_2932;
assign n_6953 = n_6837 ^ n_3001;
assign n_6954 = n_6838 ^ n_3067;
assign n_6955 = n_6839 ^ n_3136;
assign n_6956 = n_6840 ^ n_3200;
assign n_6957 = n_6841 ^ n_3265;
assign n_6958 = n_6842 ^ n_3330;
assign n_6959 = n_6843 ^ x1;
assign n_6960 = n_1 & ~n_6844;
assign n_6961 = n_6844 ^ x72;
assign n_6962 = n_655 & ~n_6845;
assign n_6963 = n_784 & ~n_6845;
assign n_6964 = ~n_6845 & ~n_3665;
assign n_6965 = ~n_6845 & n_854;
assign n_6966 = ~n_6845 & n_920;
assign n_6967 = ~n_6845 & n_986;
assign n_6968 = ~n_6845 & n_1052;
assign n_6969 = ~n_6845 & n_1117;
assign n_6970 = ~n_6845 & n_1181;
assign n_6971 = ~n_6845 & n_1248;
assign n_6972 = ~n_6845 & n_1314;
assign n_6973 = ~n_6845 & n_1380;
assign n_6974 = ~n_6845 & n_1445;
assign n_6975 = ~n_6845 & n_1510;
assign n_6976 = ~n_6845 & n_1576;
assign n_6977 = ~n_6845 & n_1641;
assign n_6978 = ~n_6845 & n_1706;
assign n_6979 = ~n_6845 & n_1771;
assign n_6980 = ~n_6845 & n_1835;
assign n_6981 = ~n_6845 & n_1899;
assign n_6982 = n_1 & ~n_6846;
assign n_6983 = n_6846 ^ x73;
assign n_6984 = x73 & n_6847;
assign n_6985 = n_6848 ^ n_6593;
assign n_6986 = x76 & ~n_6849;
assign n_6987 = n_6761 & ~n_6851;
assign n_6988 = n_6852 ^ n_6615;
assign n_6989 = n_6853 ^ n_6454;
assign n_6990 = n_6454 & n_6853;
assign n_6991 = n_6854 ^ n_6455;
assign n_6992 = n_6455 & n_6854;
assign n_6993 = n_6855 ^ n_6456;
assign n_6994 = n_6456 & n_6855;
assign n_6995 = n_6856 ^ n_6460;
assign n_6996 = n_6460 & n_6856;
assign n_6997 = n_6857 ^ n_6461;
assign n_6998 = n_6461 & n_6857;
assign n_6999 = n_6858 ^ n_6462;
assign n_7000 = n_6462 & n_6858;
assign n_7001 = n_6859 ^ n_414;
assign n_7002 = ~n_414 & ~n_6859;
assign n_7003 = n_6860 ^ n_6463;
assign n_7004 = n_6463 & n_6860;
assign n_7005 = n_6464 ^ n_6862;
assign n_7006 = n_6862 & n_6464;
assign n_7007 = n_6772 & ~n_6863;
assign n_7008 = n_6760 & ~n_6866;
assign n_7009 = n_6867 ^ n_6652;
assign n_7010 = n_6652 & n_6867;
assign n_7011 = n_6868 ^ n_6614;
assign n_7012 = n_6870 ^ n_6757;
assign n_7013 = n_6871 ^ n_6731;
assign n_7014 = n_6873 ^ n_4929;
assign n_7015 = n_6884 ^ n_6748;
assign n_7016 = n_6888 ^ n_4939;
assign n_7017 = n_6889 ^ n_444;
assign n_7018 = n_6890 ^ n_4942;
assign n_7019 = n_6864 ^ n_6891;
assign n_7020 = n_6892 ^ n_4943;
assign n_7021 = n_4943 & n_6892;
assign n_7022 = n_6633 ^ n_6893;
assign n_7023 = ~n_6779 & ~n_6894;
assign n_7024 = n_6895 ^ n_6673;
assign n_7025 = n_6896 ^ n_6296;
assign n_7026 = n_4927 ^ n_6897;
assign n_7027 = n_6311 ^ n_6898;
assign n_7028 = n_4929 ^ n_6899;
assign n_7029 = n_6900 ^ n_4930;
assign n_7030 = n_6901 ^ n_4931;
assign n_7031 = n_6902 ^ n_4932;
assign n_7032 = n_6903 ^ n_4933;
assign n_7033 = n_6886 ^ n_6903;
assign n_7034 = n_6904 ^ n_4934;
assign n_7035 = n_6904 ^ n_6878;
assign n_7036 = n_6905 ^ n_4935;
assign n_7037 = n_4936 ^ n_6906;
assign n_7038 = n_5752 ^ n_6907;
assign n_7039 = n_4937 ^ n_6908;
assign n_7040 = n_6909 ^ n_4938;
assign n_7041 = n_4939 ^ n_6910;
assign n_7042 = n_4940 ^ n_6911;
assign n_7043 = n_6912 ^ n_4941;
assign n_7044 = n_4942 ^ n_6913;
assign n_7045 = n_6916 ^ n_3426;
assign n_7046 = ~x0 & ~n_6917;
assign n_7047 = n_6918 ^ x5;
assign n_7048 = n_6919 ^ x8;
assign n_7049 = n_6920 ^ x11;
assign n_7050 = n_6921 ^ x14;
assign n_7051 = n_6922 ^ x17;
assign n_7052 = n_6923 ^ x20;
assign n_7053 = n_6924 ^ x23;
assign n_7054 = n_6925 ^ x26;
assign n_7055 = n_6926 ^ x29;
assign n_7056 = n_6927 ^ x32;
assign n_7057 = n_6928 ^ x35;
assign n_7058 = n_6929 ^ x38;
assign n_7059 = n_6930 ^ x41;
assign n_7060 = n_6931 ^ x44;
assign n_7061 = n_6932 ^ x47;
assign n_7062 = n_6933 ^ x50;
assign n_7063 = n_6934 ^ x53;
assign n_7064 = n_6935 ^ x56;
assign n_7065 = n_6725 ^ n_6936;
assign n_7066 = n_6936 ^ x59;
assign n_7067 = n_6937 ^ x62;
assign n_7068 = n_6938 ^ n_2101;
assign n_7069 = n_4998 ^ n_6939;
assign n_7070 = n_5061 ^ n_6940;
assign n_7071 = n_5124 ^ n_6941;
assign n_7072 = n_5185 ^ n_6942;
assign n_7073 = n_5249 ^ n_6943;
assign n_7074 = n_5313 ^ n_6944;
assign n_7075 = n_5377 ^ n_6945;
assign n_7076 = n_5441 ^ n_6946;
assign n_7077 = n_5502 ^ n_6947;
assign n_7078 = n_5565 ^ n_6948;
assign n_7079 = n_5628 ^ n_6949;
assign n_7080 = n_5692 ^ n_6950;
assign n_7081 = n_5758 ^ n_6951;
assign n_7082 = n_5820 ^ n_6952;
assign n_7083 = n_5884 ^ n_6953;
assign n_7084 = n_5947 ^ n_6954;
assign n_7085 = n_6011 ^ n_6955;
assign n_7086 = n_6075 ^ n_6956;
assign n_7087 = n_6137 ^ n_6957;
assign n_7088 = n_6199 ^ n_6958;
assign n_7089 = n_6959 ^ x71;
assign n_7090 = n_6960 ^ x1;
assign n_7091 = n_655 & n_6961;
assign n_7092 = n_784 & n_6961;
assign n_7093 = n_6961 & ~n_3665;
assign n_7094 = n_6961 & n_854;
assign n_7095 = n_6961 & n_920;
assign n_7096 = n_6961 & n_986;
assign n_7097 = n_6961 & n_1052;
assign n_7098 = n_6961 & n_1117;
assign n_7099 = n_6961 & n_1181;
assign n_7100 = n_6961 & n_1248;
assign n_7101 = n_6961 & n_1314;
assign n_7102 = n_6961 & n_1380;
assign n_7103 = n_6961 & n_1445;
assign n_7104 = n_6961 & n_1510;
assign n_7105 = n_6961 & n_1576;
assign n_7106 = n_6961 & n_1641;
assign n_7107 = n_6961 & n_1706;
assign n_7108 = n_6961 & n_1771;
assign n_7109 = n_6961 & n_1835;
assign n_7110 = n_6961 & n_1899;
assign n_7111 = n_2126 ^ n_6962;
assign n_7112 = n_726 ^ n_6963;
assign n_7113 = n_2197 ^ n_6964;
assign n_7114 = n_2265 ^ n_6965;
assign n_7115 = n_2332 ^ n_6966;
assign n_7116 = n_2399 ^ n_6967;
assign n_7117 = n_2466 ^ n_6968;
assign n_7118 = n_2532 ^ n_6969;
assign n_7119 = n_2597 ^ n_6970;
assign n_7120 = n_2664 ^ n_6971;
assign n_7121 = n_2732 ^ n_6972;
assign n_7122 = n_2799 ^ n_6973;
assign n_7123 = n_2867 ^ n_6974;
assign n_7124 = n_2933 ^ n_6975;
assign n_7125 = n_3002 ^ n_6976;
assign n_7126 = n_3068 ^ n_6977;
assign n_7127 = n_3137 ^ n_6978;
assign n_7128 = n_3201 ^ n_6979;
assign n_7129 = n_3266 ^ n_6980;
assign n_7130 = n_3331 ^ n_6981;
assign n_7131 = n_6982 ^ x1;
assign n_7132 = n_655 & n_6983;
assign n_7133 = n_784 & n_6983;
assign n_7134 = ~n_3665 & n_6983;
assign n_7135 = n_6983 & n_854;
assign n_7136 = n_6983 & n_920;
assign n_7137 = n_6983 & n_986;
assign n_7138 = n_6983 & n_1052;
assign n_7139 = n_6983 & n_1117;
assign n_7140 = n_6983 & n_1181;
assign n_7141 = n_6983 & n_1248;
assign n_7142 = n_6983 & n_1314;
assign n_7143 = n_6983 & n_1380;
assign n_7144 = n_6983 & n_1445;
assign n_7145 = n_6983 & n_1510;
assign n_7146 = n_6983 & n_1576;
assign n_7147 = n_6983 & n_1641;
assign n_7148 = n_6983 & n_1706;
assign n_7149 = n_6983 & n_1771;
assign n_7150 = n_6983 & n_1835;
assign n_7151 = n_6983 & n_1899;
assign n_7152 = n_6984 ^ x73;
assign n_7153 = ~x74 & ~n_6984;
assign n_7154 = ~x77 & ~n_6986;
assign n_7155 = n_6987 ^ n_6311;
assign n_7156 = n_6988 ^ n_6453;
assign n_7157 = n_6990 ^ n_6874;
assign n_7158 = ~n_364 & ~n_6990;
assign n_7159 = n_6992 ^ n_6875;
assign n_7160 = ~n_370 & ~n_6992;
assign n_7161 = n_6994 ^ n_6876;
assign n_7162 = ~n_376 & ~n_6994;
assign n_7163 = n_6996 ^ n_6879;
assign n_7164 = ~n_395 & ~n_6996;
assign n_7165 = n_6998 ^ n_6880;
assign n_7166 = ~n_401 & ~n_6998;
assign n_7167 = n_7000 ^ n_6881;
assign n_7168 = ~n_407 & ~n_7000;
assign n_7169 = ~n_6774 & ~n_7002;
assign n_7170 = n_7004 ^ n_6882;
assign n_7171 = ~n_420 & ~n_7004;
assign n_7172 = n_6883 & ~n_7006;
assign n_7173 = n_7007 ^ n_6912;
assign n_7174 = n_7008 ^ n_4927;
assign y3 = n_7009;
assign n_7175 = n_4926 ^ n_7010;
assign n_7176 = n_7014 ^ n_6899;
assign n_7177 = n_7016 ^ n_6910;
assign n_7178 = n_7017 ^ n_6631;
assign n_7179 = n_7018 ^ n_6913;
assign n_7180 = n_7020 ^ n_6914;
assign n_7181 = ~n_7020 & n_6915;
assign n_7182 = n_7021 ^ n_7020;
assign n_7183 = n_7021 ^ n_6725;
assign n_7184 = n_6916 ^ n_7023;
assign n_7185 = n_7024 ^ n_4926;
assign n_7186 = n_6869 ^ n_7025;
assign n_7187 = ~n_7025 & n_6869;
assign n_7188 = n_6896 & n_7025;
assign n_7189 = n_7014 & ~n_7028;
assign n_7190 = n_6886 ^ n_7032;
assign n_7191 = ~n_7032 & n_7033;
assign n_7192 = n_7034 ^ n_6878;
assign n_7193 = ~n_7034 & n_7035;
assign n_7194 = n_7016 & ~n_7041;
assign n_7195 = n_7007 ^ n_7043;
assign n_7196 = n_7018 & ~n_7044;
assign n_7197 = n_7045 ^ n_7023;
assign n_7198 = n_7046 ^ n_6801;
assign n_7199 = n_6865 ^ n_7047;
assign n_7200 = n_7049 ^ n_6451;
assign n_7201 = n_6989 ^ n_7050;
assign n_7202 = n_6991 ^ n_7051;
assign n_7203 = n_6993 ^ n_7052;
assign n_7204 = n_7053 ^ n_6719;
assign n_7205 = n_6985 ^ n_7054;
assign n_7206 = n_6995 ^ n_7055;
assign n_7207 = n_6997 ^ n_7056;
assign n_7208 = n_6999 ^ n_7057;
assign n_7209 = n_7058 ^ n_6624;
assign n_7210 = n_7003 ^ n_7059;
assign n_7211 = n_6861 ^ n_7060;
assign n_7212 = n_7061 ^ n_6464;
assign n_7213 = n_6747 ^ n_7062;
assign n_7214 = n_7063 ^ n_6723;
assign n_7215 = n_6724 ^ n_7064;
assign n_7216 = n_7065 ^ n_6799;
assign n_7217 = n_7066 ^ n_6725;
assign n_7218 = n_3448 ^ n_7067;
assign n_7219 = ~x0 & n_7068;
assign n_7220 = n_7069 ^ x5;
assign n_7221 = n_7070 ^ x8;
assign n_7222 = n_7071 ^ x11;
assign n_7223 = n_7072 ^ x14;
assign n_7224 = n_7073 ^ x17;
assign n_7225 = n_7074 ^ x20;
assign n_7226 = n_7075 ^ x23;
assign n_7227 = n_7076 ^ x26;
assign n_7228 = n_7077 ^ x29;
assign n_7229 = n_7078 ^ x32;
assign n_7230 = n_7079 ^ x35;
assign n_7231 = n_7080 ^ x38;
assign n_7232 = n_7081 ^ x41;
assign n_7233 = n_7082 ^ x44;
assign n_7234 = n_7083 ^ x47;
assign n_7235 = n_7084 ^ x50;
assign n_7236 = n_7085 ^ x53;
assign n_7237 = n_7086 ^ x56;
assign n_7238 = n_7087 ^ x59;
assign n_7239 = n_6472 ^ n_7088;
assign n_7240 = n_7088 ^ x2;
assign n_7241 = n_7089 ^ n_3459;
assign n_7242 = n_7090 ^ x72;
assign n_7243 = n_2127 ^ n_7091;
assign n_7244 = n_727 ^ n_7092;
assign n_7245 = n_2198 ^ n_7093;
assign n_7246 = n_2266 ^ n_7094;
assign n_7247 = n_2333 ^ n_7095;
assign n_7248 = n_2400 ^ n_7096;
assign n_7249 = n_2467 ^ n_7097;
assign n_7250 = n_2533 ^ n_7098;
assign n_7251 = n_2598 ^ n_7099;
assign n_7252 = n_2665 ^ n_7100;
assign n_7253 = n_2733 ^ n_7101;
assign n_7254 = n_2800 ^ n_7102;
assign n_7255 = n_2868 ^ n_7103;
assign n_7256 = n_2934 ^ n_7104;
assign n_7257 = n_3003 ^ n_7105;
assign n_7258 = n_3069 ^ n_7106;
assign n_7259 = n_3138 ^ n_7107;
assign n_7260 = n_3202 ^ n_7108;
assign n_7261 = n_3267 ^ n_7109;
assign n_7262 = n_3332 ^ n_7110;
assign n_7263 = n_4999 ^ n_7111;
assign n_7264 = n_5062 ^ n_7112;
assign n_7265 = n_5125 ^ n_7113;
assign n_7266 = n_5186 ^ n_7114;
assign n_7267 = n_5250 ^ n_7115;
assign n_7268 = n_5314 ^ n_7116;
assign n_7269 = n_5378 ^ n_7117;
assign n_7270 = n_5442 ^ n_7118;
assign n_7271 = n_5503 ^ n_7119;
assign n_7272 = n_5566 ^ n_7120;
assign n_7273 = n_5629 ^ n_7121;
assign n_7274 = n_5693 ^ n_7122;
assign n_7275 = n_5759 ^ n_7123;
assign n_7276 = n_5821 ^ n_7124;
assign n_7277 = n_5885 ^ n_7125;
assign n_7278 = n_5948 ^ n_7126;
assign n_7279 = n_6012 ^ n_7127;
assign n_7280 = n_6076 ^ n_7128;
assign n_7281 = n_6138 ^ n_7129;
assign n_7282 = n_6200 ^ n_7130;
assign n_7283 = n_7131 ^ x73;
assign n_7284 = n_2128 ^ n_7132;
assign n_7285 = n_728 ^ n_7133;
assign n_7286 = n_2199 ^ n_7134;
assign n_7287 = n_2267 ^ n_7135;
assign n_7288 = n_2334 ^ n_7136;
assign n_7289 = n_2401 ^ n_7137;
assign n_7290 = n_2468 ^ n_7138;
assign n_7291 = n_2534 ^ n_7139;
assign n_7292 = n_2599 ^ n_7140;
assign n_7293 = n_2666 ^ n_7141;
assign n_7294 = n_2734 ^ n_7142;
assign n_7295 = n_2801 ^ n_7143;
assign n_7296 = n_2869 ^ n_7144;
assign n_7297 = n_2935 ^ n_7145;
assign n_7298 = n_3004 ^ n_7146;
assign n_7299 = n_3070 ^ n_7147;
assign n_7300 = n_3139 ^ n_7148;
assign n_7301 = n_3203 ^ n_7149;
assign n_7302 = n_3268 ^ n_7150;
assign n_7303 = n_3333 ^ n_7151;
assign n_7304 = n_7152 ^ n_6470;
assign n_7305 = n_7153 ^ n_6726;
assign n_7306 = x75 & ~n_7153;
assign n_7307 = n_7155 ^ n_6898;
assign n_7308 = n_7155 & ~n_7027;
assign n_7309 = n_7156 ^ n_7048;
assign n_7310 = n_6763 & ~n_7158;
assign n_7311 = n_6764 & ~n_7160;
assign n_7312 = n_6765 & ~n_7162;
assign n_7313 = n_6767 & ~n_7164;
assign n_7314 = n_6768 & ~n_7166;
assign n_7315 = n_6769 & ~n_7168;
assign n_7316 = n_7169 ^ n_4937;
assign n_7317 = n_6770 & ~n_7171;
assign n_7318 = n_6771 & ~n_7172;
assign n_7319 = ~n_7043 & n_7173;
assign n_7320 = n_7174 ^ n_6897;
assign n_7321 = n_7174 & ~n_7026;
assign n_7322 = n_7178 ^ n_6749;
assign n_7323 = n_7181 ^ n_6799;
assign n_7324 = ~n_7045 & ~n_7184;
assign n_7325 = n_7185 ^ n_7010;
assign n_7326 = n_7185 & ~n_7175;
assign n_7327 = n_7187 ^ n_7188;
assign n_7328 = n_7189 ^ n_6873;
assign n_7329 = n_7191 ^ n_6886;
assign n_7330 = n_7193 ^ n_6878;
assign n_7331 = n_7194 ^ n_6888;
assign n_7332 = n_7196 ^ n_6890;
assign n_7333 = n_7198 ^ n_6613;
assign n_7334 = n_7212 ^ n_6862;
assign n_7335 = n_6914 & ~n_7216;
assign n_7336 = ~n_7217 & n_7183;
assign n_7337 = n_7219 ^ n_6938;
assign n_7338 = n_7012 ^ n_7220;
assign n_7339 = n_7013 ^ n_7221;
assign n_7340 = n_6872 ^ n_7222;
assign n_7341 = n_7157 ^ n_7223;
assign n_7342 = n_7159 ^ n_7224;
assign n_7343 = n_7161 ^ n_7225;
assign n_7344 = n_6885 ^ n_7226;
assign n_7345 = n_6877 ^ n_7227;
assign n_7346 = n_7163 ^ n_7228;
assign n_7347 = n_7165 ^ n_7229;
assign n_7348 = n_7167 ^ n_7230;
assign n_7349 = n_7001 ^ n_7231;
assign n_7350 = n_7170 ^ n_7232;
assign n_7351 = n_6887 ^ n_7233;
assign n_7352 = n_6883 ^ n_7234;
assign n_7353 = n_7015 ^ n_7235;
assign n_7354 = n_7019 ^ n_7237;
assign n_7355 = n_7022 ^ n_7238;
assign n_7356 = ~n_7240 & n_3454;
assign n_7357 = n_7240 & n_532;
assign n_7358 = ~x0 & n_7241;
assign n_7359 = n_7242 ^ n_2102;
assign n_7360 = n_5000 ^ n_7243;
assign n_7361 = n_5063 ^ n_7244;
assign n_7362 = n_5126 ^ n_7245;
assign n_7363 = n_5187 ^ n_7246;
assign n_7364 = n_5251 ^ n_7247;
assign n_7365 = n_5315 ^ n_7248;
assign n_7366 = n_5379 ^ n_7249;
assign n_7367 = n_5443 ^ n_7250;
assign n_7368 = n_5504 ^ n_7251;
assign n_7369 = n_5567 ^ n_7252;
assign n_7370 = n_5630 ^ n_7253;
assign n_7371 = n_5694 ^ n_7254;
assign n_7372 = n_5760 ^ n_7255;
assign n_7373 = n_5822 ^ n_7256;
assign n_7374 = n_5886 ^ n_7257;
assign n_7375 = n_5949 ^ n_7258;
assign n_7376 = n_6013 ^ n_7259;
assign n_7377 = n_6077 ^ n_7260;
assign n_7378 = n_6139 ^ n_7261;
assign n_7379 = n_6201 ^ n_7262;
assign n_7380 = n_7263 ^ x5;
assign n_7381 = n_7264 ^ x8;
assign n_7382 = n_7265 ^ x11;
assign n_7383 = n_7266 ^ x14;
assign n_7384 = n_7267 ^ x17;
assign n_7385 = n_7268 ^ x20;
assign n_7386 = n_7269 ^ x23;
assign n_7387 = n_7270 ^ x26;
assign n_7388 = n_7271 ^ x29;
assign n_7389 = n_7272 ^ x32;
assign n_7390 = n_7273 ^ x35;
assign n_7391 = n_7274 ^ x38;
assign n_7392 = n_7275 ^ x41;
assign n_7393 = n_7276 ^ x44;
assign n_7394 = n_7277 ^ x47;
assign n_7395 = n_7278 ^ x50;
assign n_7396 = n_7279 ^ x53;
assign n_7397 = n_7280 ^ x56;
assign n_7398 = n_7281 ^ x59;
assign n_7399 = n_6473 ^ n_7282;
assign n_7400 = n_7282 ^ x2;
assign n_7401 = n_7283 ^ n_3460;
assign n_7402 = n_5001 ^ n_7284;
assign n_7403 = n_5064 ^ n_7285;
assign n_7404 = n_5127 ^ n_7286;
assign n_7405 = n_5188 ^ n_7287;
assign n_7406 = n_5252 ^ n_7288;
assign n_7407 = n_5316 ^ n_7289;
assign n_7408 = n_5380 ^ n_7290;
assign n_7409 = n_5444 ^ n_7291;
assign n_7410 = n_5505 ^ n_7292;
assign n_7411 = n_5568 ^ n_7293;
assign n_7412 = n_5631 ^ n_7294;
assign n_7413 = n_5695 ^ n_7295;
assign n_7414 = n_5761 ^ n_7296;
assign n_7415 = n_5823 ^ n_7297;
assign n_7416 = n_5887 ^ n_7298;
assign n_7417 = n_5950 ^ n_7299;
assign n_7418 = n_6014 ^ n_7300;
assign n_7419 = n_6078 ^ n_7301;
assign n_7420 = n_6140 ^ n_7302;
assign n_7421 = n_6202 ^ n_7303;
assign n_7422 = n_1 & ~n_7304;
assign n_7423 = n_7304 ^ x74;
assign n_7424 = n_1 & n_7305;
assign n_7425 = n_7305 ^ x75;
assign n_7426 = n_7306 ^ n_6849;
assign n_7427 = ~x76 & ~n_7306;
assign n_7428 = n_7308 ^ n_6987;
assign n_7429 = n_7310 ^ n_7029;
assign n_7430 = n_7310 ^ n_6900;
assign n_7431 = n_7311 ^ n_7030;
assign n_7432 = n_7311 ^ n_6901;
assign n_7433 = n_7312 ^ n_7031;
assign n_7434 = n_7312 ^ n_6902;
assign n_7435 = n_7313 ^ n_7036;
assign n_7436 = n_7313 ^ n_6905;
assign n_7437 = n_7314 ^ n_4936;
assign n_7438 = n_7315 ^ n_5752;
assign n_7439 = n_7316 ^ n_6908;
assign n_7440 = n_7316 & ~n_7039;
assign n_7441 = n_7317 ^ n_7040;
assign n_7442 = n_7317 ^ n_6909;
assign n_7443 = n_7318 ^ n_4940;
assign n_7444 = n_7319 ^ n_7007;
assign n_7445 = n_7321 ^ n_7008;
assign n_7446 = n_7322 ^ n_7236;
assign n_7447 = n_7323 ^ n_7065;
assign n_7448 = n_7324 ^ n_7023;
assign y4 = n_7325;
assign n_7449 = n_7326 ^ n_7024;
assign n_7450 = n_7199 ^ n_7327;
assign n_7451 = n_6865 ^ n_7327;
assign n_7452 = n_7328 ^ n_7201;
assign n_7453 = n_7328 ^ n_6989;
assign n_7454 = n_7329 ^ n_7205;
assign n_7455 = n_7329 ^ n_6985;
assign n_7456 = n_7330 ^ n_7206;
assign n_7457 = n_7330 ^ n_6995;
assign n_7458 = n_7061 & n_7331;
assign n_7459 = n_7332 ^ n_6724;
assign n_7460 = n_7331 ^ n_7334;
assign n_7461 = n_7335 & n_7182;
assign n_7462 = n_7336 ^ n_7021;
assign n_7463 = n_7011 ^ n_7337;
assign n_7464 = n_7356 ^ x2;
assign n_7465 = n_7357 ^ x2;
assign n_7466 = n_7358 ^ n_7089;
assign n_7467 = ~x0 & n_7359;
assign n_7468 = n_7360 ^ x5;
assign n_7469 = n_7361 ^ x8;
assign n_7470 = n_7362 ^ x11;
assign n_7471 = n_7363 ^ x14;
assign n_7472 = n_7364 ^ x17;
assign n_7473 = n_7365 ^ x20;
assign n_7474 = n_7366 ^ x23;
assign n_7475 = n_7367 ^ x26;
assign n_7476 = n_7368 ^ x29;
assign n_7477 = n_7369 ^ x32;
assign n_7478 = n_7370 ^ x35;
assign n_7479 = n_7371 ^ x38;
assign n_7480 = n_7372 ^ x41;
assign n_7481 = n_7373 ^ x44;
assign n_7482 = n_7374 ^ x47;
assign n_7483 = n_7375 ^ x50;
assign n_7484 = n_7376 ^ x53;
assign n_7485 = n_7377 ^ x56;
assign n_7486 = n_7378 ^ x59;
assign n_7487 = n_6599 ^ n_7379;
assign n_7488 = n_7379 ^ x2;
assign n_7489 = n_7320 ^ n_7380;
assign n_7490 = n_7307 ^ n_7381;
assign n_7491 = n_7176 ^ n_7382;
assign n_7492 = n_7190 ^ n_7386;
assign n_7493 = n_7387 ^ n_7192;
assign n_7494 = n_7177 ^ n_7393;
assign n_7495 = n_7195 ^ n_7395;
assign n_7496 = n_7179 ^ n_7396;
assign n_7497 = n_7180 ^ n_7397;
assign n_7498 = n_7197 ^ n_7398;
assign n_7499 = ~n_7400 & n_3456;
assign n_7500 = n_7400 & n_534;
assign n_7501 = ~x0 & n_7401;
assign n_7502 = n_7402 ^ x5;
assign n_7503 = n_7403 ^ x8;
assign n_7504 = n_7404 ^ x11;
assign n_7505 = n_7405 ^ x14;
assign n_7506 = n_7406 ^ x17;
assign n_7507 = n_7407 ^ x20;
assign n_7508 = n_7408 ^ x23;
assign n_7509 = n_7409 ^ x26;
assign n_7510 = n_7410 ^ x29;
assign n_7511 = n_7411 ^ x32;
assign n_7512 = n_7412 ^ x35;
assign n_7513 = n_7413 ^ x38;
assign n_7514 = n_7414 ^ x41;
assign n_7515 = n_7415 ^ x44;
assign n_7516 = n_7416 ^ x47;
assign n_7517 = n_7417 ^ x50;
assign n_7518 = n_7418 ^ x53;
assign n_7519 = n_7419 ^ x56;
assign n_7520 = n_7420 ^ x59;
assign n_7521 = n_7421 ^ x62;
assign n_7522 = n_7422 ^ x1;
assign n_7523 = n_655 & n_7423;
assign n_7524 = n_784 & n_7423;
assign n_7525 = ~n_3665 & n_7423;
assign n_7526 = n_7423 & n_854;
assign n_7527 = n_7423 & n_920;
assign n_7528 = n_7423 & n_986;
assign n_7529 = n_7423 & n_1052;
assign n_7530 = n_7423 & n_1117;
assign n_7531 = n_7423 & n_1181;
assign n_7532 = n_7423 & n_1248;
assign n_7533 = n_7423 & n_1314;
assign n_7534 = n_7423 & n_1380;
assign n_7535 = n_7423 & n_1445;
assign n_7536 = n_7423 & n_1510;
assign n_7537 = n_7423 & n_1576;
assign n_7538 = n_7423 & n_1641;
assign n_7539 = n_7423 & n_1706;
assign n_7540 = n_7423 & n_1771;
assign n_7541 = n_7423 & n_1835;
assign n_7542 = n_7423 & n_1899;
assign n_7543 = n_7424 ^ x1;
assign n_7544 = n_655 & ~n_7425;
assign n_7545 = n_784 & ~n_7425;
assign n_7546 = ~n_3665 & ~n_7425;
assign n_7547 = ~n_7425 & n_854;
assign n_7548 = ~n_7425 & n_920;
assign n_7549 = ~n_7425 & n_986;
assign n_7550 = ~n_7425 & n_1052;
assign n_7551 = ~n_7425 & n_1117;
assign n_7552 = ~n_7425 & n_1181;
assign n_7553 = ~n_7425 & n_1248;
assign n_7554 = ~n_7425 & n_1314;
assign n_7555 = ~n_7425 & n_1380;
assign n_7556 = ~n_7425 & n_1445;
assign n_7557 = ~n_7425 & n_1510;
assign n_7558 = ~n_7425 & n_1576;
assign n_7559 = ~n_7425 & n_1641;
assign n_7560 = ~n_7425 & n_1706;
assign n_7561 = ~n_7425 & n_1771;
assign n_7562 = ~n_7425 & n_1835;
assign n_7563 = ~n_7425 & n_1899;
assign n_7564 = n_1 & n_7426;
assign n_7565 = n_7426 ^ x76;
assign n_7566 = n_7427 ^ n_6986;
assign n_7567 = x77 & ~n_7427;
assign n_7568 = n_7428 ^ n_7200;
assign n_7569 = n_7428 ^ n_7049;
assign n_7570 = n_7429 ^ n_7383;
assign n_7571 = ~n_7029 & n_7430;
assign n_7572 = n_7431 ^ n_7384;
assign n_7573 = ~n_7030 & n_7432;
assign n_7574 = n_7433 ^ n_7385;
assign n_7575 = ~n_7031 & n_7434;
assign n_7576 = n_7435 ^ n_7388;
assign n_7577 = ~n_7036 & n_7436;
assign n_7578 = n_7437 ^ n_6906;
assign n_7579 = n_7437 & ~n_7037;
assign n_7580 = n_7438 ^ n_6907;
assign n_7581 = n_7438 & ~n_7038;
assign n_7582 = n_7439 ^ n_7391;
assign n_7583 = n_7440 ^ n_7169;
assign n_7584 = n_7392 ^ n_7441;
assign n_7585 = ~n_7040 & n_7442;
assign n_7586 = n_7443 ^ n_6911;
assign n_7587 = n_7443 & ~n_7042;
assign n_7588 = n_7444 ^ n_7214;
assign n_7589 = n_7444 ^ n_7063;
assign n_7590 = n_7445 ^ n_7309;
assign n_7591 = n_7445 ^ n_7156;
assign n_7592 = n_7448 ^ n_3448;
assign n_7593 = n_7449 ^ n_7333;
assign n_7594 = n_7449 ^ n_7198;
assign n_7595 = n_7199 & ~n_7451;
assign n_7596 = ~n_7201 & n_7453;
assign n_7597 = n_7205 & ~n_7455;
assign n_7598 = ~n_7206 & n_7457;
assign n_7599 = n_7458 ^ n_7006;
assign n_7600 = n_7459 ^ n_7064;
assign n_7601 = n_7459 & ~n_7215;
assign n_7602 = n_7460 ^ n_6862;
assign n_7603 = ~n_7461 & ~n_7462;
assign n_7604 = n_7464 ^ n_7465;
assign n_7605 = n_7186 ^ n_7466;
assign n_7606 = n_7467 ^ n_7242;
assign n_7607 = n_7452 ^ n_7470;
assign n_7608 = n_7454 ^ n_7474;
assign n_7609 = n_7456 ^ n_7475;
assign n_7610 = n_7460 ^ n_7481;
assign n_7611 = n_7447 ^ n_7485;
assign n_7612 = ~n_7488 & n_4950;
assign n_7613 = n_7488 & n_536;
assign n_7614 = n_7499 ^ x2;
assign n_7615 = n_7500 ^ x2;
assign n_7616 = n_7501 ^ n_7283;
assign n_7617 = n_7520 ^ n_7239;
assign n_7618 = n_4951 ^ n_7521;
assign n_7619 = n_7522 ^ x74;
assign n_7620 = n_2129 ^ n_7523;
assign n_7621 = n_729 ^ n_7524;
assign n_7622 = n_2200 ^ n_7525;
assign n_7623 = n_2268 ^ n_7526;
assign n_7624 = n_2335 ^ n_7527;
assign n_7625 = n_2402 ^ n_7528;
assign n_7626 = n_2469 ^ n_7529;
assign n_7627 = n_2535 ^ n_7530;
assign n_7628 = n_2600 ^ n_7531;
assign n_7629 = n_2667 ^ n_7532;
assign n_7630 = n_2735 ^ n_7533;
assign n_7631 = n_2802 ^ n_7534;
assign n_7632 = n_2870 ^ n_7535;
assign n_7633 = n_2936 ^ n_7536;
assign n_7634 = n_3005 ^ n_7537;
assign n_7635 = n_3071 ^ n_7538;
assign n_7636 = n_3140 ^ n_7539;
assign n_7637 = n_3204 ^ n_7540;
assign n_7638 = n_3269 ^ n_7541;
assign n_7639 = n_3334 ^ n_7542;
assign n_7640 = n_7543 ^ x75;
assign n_7641 = n_2130 ^ n_7544;
assign n_7642 = n_730 ^ n_7545;
assign n_7643 = n_2201 ^ n_7546;
assign n_7644 = n_2269 ^ n_7547;
assign n_7645 = n_2336 ^ n_7548;
assign n_7646 = n_2403 ^ n_7549;
assign n_7647 = n_2470 ^ n_7550;
assign n_7648 = n_2536 ^ n_7551;
assign n_7649 = n_2601 ^ n_7552;
assign n_7650 = n_2668 ^ n_7553;
assign n_7651 = n_2736 ^ n_7554;
assign n_7652 = n_2803 ^ n_7555;
assign n_7653 = n_2871 ^ n_7556;
assign n_7654 = n_2937 ^ n_7557;
assign n_7655 = n_3006 ^ n_7558;
assign n_7656 = n_3072 ^ n_7559;
assign n_7657 = n_3141 ^ n_7560;
assign n_7658 = n_3205 ^ n_7561;
assign n_7659 = n_3270 ^ n_7562;
assign n_7660 = n_3335 ^ n_7563;
assign n_7661 = n_7564 ^ x1;
assign n_7662 = n_655 & ~n_7565;
assign n_7663 = n_784 & ~n_7565;
assign n_7664 = ~n_3665 & ~n_7565;
assign n_7665 = n_854 & ~n_7565;
assign n_7666 = ~n_7565 & n_920;
assign n_7667 = ~n_7565 & n_986;
assign n_7668 = ~n_7565 & n_1052;
assign n_7669 = ~n_7565 & n_1117;
assign n_7670 = ~n_7565 & n_1181;
assign n_7671 = ~n_7565 & n_1248;
assign n_7672 = ~n_7565 & n_1314;
assign n_7673 = ~n_7565 & n_1380;
assign n_7674 = ~n_7565 & n_1445;
assign n_7675 = ~n_7565 & n_1510;
assign n_7676 = ~n_7565 & n_1576;
assign n_7677 = ~n_7565 & n_1641;
assign n_7678 = ~n_7565 & n_1706;
assign n_7679 = ~n_7565 & n_1771;
assign n_7680 = ~n_7565 & n_1835;
assign n_7681 = ~n_7565 & n_1899;
assign n_7682 = n_1 & n_7566;
assign n_7683 = n_7566 ^ x77;
assign n_7684 = n_7567 ^ n_7154;
assign n_7685 = n_7568 ^ n_7469;
assign n_7686 = ~n_7200 & n_7569;
assign n_7687 = n_7571 ^ n_7310;
assign n_7688 = n_7573 ^ n_7311;
assign n_7689 = n_7575 ^ n_7312;
assign n_7690 = n_7577 ^ n_7313;
assign n_7691 = n_7578 ^ n_7389;
assign n_7692 = n_7579 ^ n_7314;
assign n_7693 = n_7390 ^ n_7580;
assign n_7694 = n_7581 ^ n_7315;
assign n_7695 = n_7583 ^ n_7210;
assign n_7696 = n_7583 ^ n_7003;
assign n_7697 = n_7585 ^ n_7317;
assign n_7698 = n_7394 ^ n_7586;
assign n_7699 = n_7587 ^ n_7318;
assign n_7700 = n_7588 ^ n_7483;
assign n_7701 = ~n_7214 & n_7589;
assign n_7702 = n_7590 ^ n_7468;
assign n_7703 = n_7309 & ~n_7591;
assign n_7704 = n_7592 ^ n_7067;
assign n_7705 = ~n_7592 & ~n_7218;
assign y5 = n_7593;
assign n_7706 = ~n_7333 & n_7594;
assign n_7707 = n_7595 ^ n_7327;
assign n_7708 = n_7596 ^ n_7328;
assign n_7709 = n_7597 ^ n_7329;
assign n_7710 = n_7598 ^ n_7330;
assign n_7711 = n_7600 ^ n_7484;
assign n_7712 = n_7601 ^ n_7332;
assign n_7713 = n_7005 & ~n_7602;
assign n_7714 = n_7355 ^ n_7603;
assign n_7715 = n_7022 ^ n_7603;
assign n_7716 = ~x62 & n_7604;
assign n_7717 = n_7450 ^ n_7606;
assign n_7718 = n_7612 ^ x2;
assign n_7719 = n_7613 ^ x2;
assign n_7720 = n_7614 ^ n_7615;
assign n_7721 = n_7619 ^ n_3461;
assign n_7722 = n_5002 ^ n_7620;
assign n_7723 = n_5065 ^ n_7621;
assign n_7724 = n_5128 ^ n_7622;
assign n_7725 = n_5189 ^ n_7623;
assign n_7726 = n_5253 ^ n_7624;
assign n_7727 = n_5317 ^ n_7625;
assign n_7728 = n_5381 ^ n_7626;
assign n_7729 = n_5445 ^ n_7627;
assign n_7730 = n_5506 ^ n_7628;
assign n_7731 = n_5569 ^ n_7629;
assign n_7732 = n_5632 ^ n_7630;
assign n_7733 = n_5696 ^ n_7631;
assign n_7734 = n_5762 ^ n_7632;
assign n_7735 = n_5824 ^ n_7633;
assign n_7736 = n_5888 ^ n_7634;
assign n_7737 = n_5951 ^ n_7635;
assign n_7738 = n_6015 ^ n_7636;
assign n_7739 = n_6079 ^ n_7637;
assign n_7740 = n_6141 ^ n_7638;
assign n_7741 = n_6203 ^ n_7639;
assign n_7742 = n_7640 ^ n_2103;
assign n_7743 = n_5003 ^ n_7641;
assign n_7744 = n_5066 ^ n_7642;
assign n_7745 = n_5129 ^ n_7643;
assign n_7746 = n_5190 ^ n_7644;
assign n_7747 = n_5254 ^ n_7645;
assign n_7748 = n_5318 ^ n_7646;
assign n_7749 = n_5382 ^ n_7647;
assign n_7750 = n_5446 ^ n_7648;
assign n_7751 = n_5507 ^ n_7649;
assign n_7752 = n_5570 ^ n_7650;
assign n_7753 = n_5633 ^ n_7651;
assign n_7754 = n_5697 ^ n_7652;
assign n_7755 = n_5763 ^ n_7653;
assign n_7756 = n_5825 ^ n_7654;
assign n_7757 = n_5889 ^ n_7655;
assign n_7758 = n_5952 ^ n_7656;
assign n_7759 = n_6016 ^ n_7657;
assign n_7760 = n_6080 ^ n_7658;
assign n_7761 = n_6142 ^ n_7659;
assign n_7762 = n_6204 ^ n_7660;
assign n_7763 = n_7661 ^ x76;
assign n_7764 = n_2131 ^ n_7662;
assign n_7765 = n_731 ^ n_7663;
assign n_7766 = n_2202 ^ n_7664;
assign n_7767 = n_2270 ^ n_7665;
assign n_7768 = n_2337 ^ n_7666;
assign n_7769 = n_2404 ^ n_7667;
assign n_7770 = n_2471 ^ n_7668;
assign n_7771 = n_2537 ^ n_7669;
assign n_7772 = n_2602 ^ n_7670;
assign n_7773 = n_2669 ^ n_7671;
assign n_7774 = n_2737 ^ n_7672;
assign n_7775 = n_2804 ^ n_7673;
assign n_7776 = n_2872 ^ n_7674;
assign n_7777 = n_2938 ^ n_7675;
assign n_7778 = n_3007 ^ n_7676;
assign n_7779 = n_3073 ^ n_7677;
assign n_7780 = n_3142 ^ n_7678;
assign n_7781 = n_3206 ^ n_7679;
assign n_7782 = n_3271 ^ n_7680;
assign n_7783 = n_3336 ^ n_7681;
assign n_7784 = n_7682 ^ x1;
assign n_7785 = n_655 & ~n_7683;
assign n_7786 = n_784 & ~n_7683;
assign n_7787 = ~n_3665 & ~n_7683;
assign n_7788 = n_854 & ~n_7683;
assign n_7789 = ~n_7683 & n_920;
assign n_7790 = ~n_7683 & n_986;
assign n_7791 = ~n_7683 & n_1052;
assign n_7792 = ~n_7683 & n_1117;
assign n_7793 = ~n_7683 & n_1181;
assign n_7794 = ~n_7683 & n_1248;
assign n_7795 = ~n_7683 & n_1314;
assign n_7796 = ~n_7683 & n_1380;
assign n_7797 = ~n_7683 & n_1445;
assign n_7798 = ~n_7683 & n_1510;
assign n_7799 = ~n_7683 & n_1576;
assign n_7800 = ~n_7683 & n_1641;
assign n_7801 = ~n_7683 & n_1706;
assign n_7802 = ~n_7683 & n_1771;
assign n_7803 = ~n_7683 & n_1835;
assign n_7804 = ~n_7683 & n_1899;
assign n_7805 = n_1 & n_7684;
assign n_7806 = n_7684 & n_139;
assign n_7807 = ~x79 & n_7684;
assign n_7808 = n_7684 ^ x78;
assign n_7809 = n_7686 ^ n_7428;
assign n_7810 = n_7687 ^ n_7202;
assign n_7811 = n_7687 ^ n_6991;
assign n_7812 = n_7688 ^ n_7203;
assign n_7813 = n_7688 ^ n_6993;
assign n_7814 = n_7689 ^ n_7204;
assign n_7815 = n_7689 ^ n_7053;
assign n_7816 = n_7690 ^ n_7207;
assign n_7817 = n_7690 ^ n_6997;
assign n_7818 = n_7692 ^ n_7208;
assign n_7819 = n_7692 ^ n_6999;
assign n_7820 = n_7694 ^ n_7209;
assign n_7821 = n_7694 ^ n_7058;
assign n_7822 = n_7695 ^ n_7479;
assign n_7823 = ~n_7210 & n_7696;
assign n_7824 = n_7697 ^ n_6861;
assign n_7825 = n_7699 ^ n_7213;
assign n_7826 = n_7699 ^ n_6747;
assign n_7827 = n_7701 ^ n_7444;
assign n_7828 = n_7703 ^ n_7445;
assign n_7829 = n_7704 ^ n_7486;
assign n_7830 = n_7705 ^ n_7448;
assign n_7831 = n_7706 ^ n_7449;
assign n_7832 = n_7707 ^ n_7338;
assign n_7833 = n_7707 ^ n_7012;
assign n_7834 = n_7708 ^ n_7341;
assign n_7835 = n_7708 ^ n_7157;
assign n_7836 = n_7709 ^ n_7345;
assign n_7837 = n_7709 ^ n_7227;
assign n_7838 = n_7710 ^ n_7346;
assign n_7839 = n_7710 ^ n_7163;
assign n_7840 = n_7712 ^ n_7354;
assign n_7841 = n_7712 ^ n_7019;
assign n_7842 = n_7713 ^ n_6862;
assign n_7843 = n_7519 ^ n_7714;
assign n_7844 = n_7355 & n_7715;
assign n_7845 = n_7716 ^ n_7464;
assign n_7846 = n_7718 ^ n_7719;
assign n_7847 = ~x62 & n_7720;
assign n_7848 = ~x0 & n_7721;
assign n_7849 = n_7722 ^ x5;
assign n_7850 = n_7723 ^ x8;
assign n_7851 = n_7724 ^ x11;
assign n_7852 = n_7725 ^ x14;
assign n_7853 = n_7726 ^ x17;
assign n_7854 = n_7727 ^ x20;
assign n_7855 = n_7728 ^ x23;
assign n_7856 = n_7729 ^ x26;
assign n_7857 = n_7730 ^ x29;
assign n_7858 = n_7731 ^ x32;
assign n_7859 = n_7732 ^ x35;
assign n_7860 = n_7733 ^ x38;
assign n_7861 = n_7734 ^ x41;
assign n_7862 = n_7735 ^ x44;
assign n_7863 = n_7736 ^ x47;
assign n_7864 = n_7737 ^ x50;
assign n_7865 = n_7738 ^ x53;
assign n_7866 = n_7739 ^ x56;
assign n_7867 = n_7740 ^ x59;
assign n_7868 = n_7741 ^ x62;
assign n_7869 = ~x0 & n_7742;
assign n_7870 = n_7743 ^ x5;
assign n_7871 = n_7744 ^ x8;
assign n_7872 = n_7745 ^ x11;
assign n_7873 = n_7746 ^ x14;
assign n_7874 = n_7747 ^ x17;
assign n_7875 = n_7748 ^ x20;
assign n_7876 = n_7749 ^ x23;
assign n_7877 = n_7750 ^ x26;
assign n_7878 = n_7751 ^ x29;
assign n_7879 = n_7752 ^ x32;
assign n_7880 = n_7753 ^ x35;
assign n_7881 = n_7754 ^ x38;
assign n_7882 = n_7755 ^ x41;
assign n_7883 = n_7756 ^ x44;
assign n_7884 = n_7757 ^ x47;
assign n_7885 = n_7758 ^ x50;
assign n_7886 = n_7759 ^ x53;
assign n_7887 = n_7760 ^ x56;
assign n_7888 = n_7761 ^ x59;
assign n_7889 = n_7762 ^ x62;
assign n_7890 = n_7763 ^ n_3462;
assign n_7891 = n_5004 ^ n_7764;
assign n_7892 = n_5067 ^ n_7765;
assign n_7893 = n_5130 ^ n_7766;
assign n_7894 = n_5191 ^ n_7767;
assign n_7895 = n_5255 ^ n_7768;
assign n_7896 = n_5319 ^ n_7769;
assign n_7897 = n_5383 ^ n_7770;
assign n_7898 = n_5447 ^ n_7771;
assign n_7899 = n_5508 ^ n_7772;
assign n_7900 = n_5571 ^ n_7773;
assign n_7901 = n_5634 ^ n_7774;
assign n_7902 = n_5698 ^ n_7775;
assign n_7903 = n_5764 ^ n_7776;
assign n_7904 = n_5826 ^ n_7777;
assign n_7905 = n_5890 ^ n_7778;
assign n_7906 = n_5953 ^ n_7779;
assign n_7907 = n_6017 ^ n_7780;
assign n_7908 = n_6081 ^ n_7781;
assign n_7909 = n_6143 ^ n_7782;
assign n_7910 = n_6205 ^ n_7783;
assign n_7911 = n_7784 ^ x77;
assign n_7912 = n_2132 ^ n_7785;
assign n_7913 = n_732 ^ n_7786;
assign n_7914 = n_2203 ^ n_7787;
assign n_7915 = n_2271 ^ n_7788;
assign n_7916 = n_2338 ^ n_7789;
assign n_7917 = n_2405 ^ n_7790;
assign n_7918 = n_2472 ^ n_7791;
assign n_7919 = n_2538 ^ n_7792;
assign n_7920 = n_2603 ^ n_7793;
assign n_7921 = n_2670 ^ n_7794;
assign n_7922 = n_2738 ^ n_7795;
assign n_7923 = n_2805 ^ n_7796;
assign n_7924 = n_2873 ^ n_7797;
assign n_7925 = n_2939 ^ n_7798;
assign n_7926 = n_3008 ^ n_7799;
assign n_7927 = n_3074 ^ n_7800;
assign n_7928 = n_3143 ^ n_7801;
assign n_7929 = n_3207 ^ n_7802;
assign n_7930 = n_3272 ^ n_7803;
assign n_7931 = n_3337 ^ n_7804;
assign n_7932 = n_7805 ^ x1;
assign n_7933 = n_1 & ~n_7806;
assign n_7934 = n_7806 ^ x79;
assign n_7935 = n_7807 ^ n_7567;
assign n_7936 = n_655 & ~n_7808;
assign n_7937 = n_784 & ~n_7808;
assign n_7938 = ~n_3665 & ~n_7808;
assign n_7939 = n_854 & ~n_7808;
assign n_7940 = ~n_7808 & n_920;
assign n_7941 = ~n_7808 & n_986;
assign n_7942 = ~n_7808 & n_1052;
assign n_7943 = ~n_7808 & n_1117;
assign n_7944 = ~n_7808 & n_1181;
assign n_7945 = ~n_7808 & n_1248;
assign n_7946 = ~n_7808 & n_1314;
assign n_7947 = ~n_7808 & n_1380;
assign n_7948 = ~n_7808 & n_1445;
assign n_7949 = ~n_7808 & n_1510;
assign n_7950 = ~n_7808 & n_1576;
assign n_7951 = ~n_7808 & n_1641;
assign n_7952 = ~n_7808 & n_1706;
assign n_7953 = ~n_7808 & n_1771;
assign n_7954 = ~n_7808 & n_1835;
assign n_7955 = ~n_7808 & n_1899;
assign n_7956 = n_7809 ^ n_7340;
assign n_7957 = n_7809 ^ n_7222;
assign n_7958 = n_7810 ^ n_7471;
assign n_7959 = ~n_7202 & n_7811;
assign n_7960 = n_7812 ^ n_7472;
assign n_7961 = ~n_7203 & n_7813;
assign n_7962 = n_7814 ^ n_7473;
assign n_7963 = ~n_7204 & n_7815;
assign n_7964 = n_7816 ^ n_7476;
assign n_7965 = ~n_7207 & n_7817;
assign n_7966 = n_7818 ^ n_7477;
assign n_7967 = ~n_7208 & n_7819;
assign n_7968 = n_7820 ^ n_7478;
assign n_7969 = ~n_7209 & n_7821;
assign n_7970 = n_7823 ^ n_7583;
assign n_7971 = n_7824 ^ n_7060;
assign n_7972 = ~n_7824 & n_7211;
assign n_7973 = n_7825 ^ n_7482;
assign n_7974 = ~n_7213 & n_7826;
assign n_7975 = n_7827 ^ n_7236;
assign n_7976 = n_7828 ^ n_7339;
assign n_7977 = n_7828 ^ n_7221;
assign n_7978 = n_7830 ^ n_7617;
assign n_7979 = n_7830 ^ n_7520;
assign n_7980 = n_7831 ^ n_7463;
assign n_7981 = n_7831 ^ n_7011;
assign n_7982 = n_7832 ^ n_7616;
assign n_7983 = ~n_7338 & n_7833;
assign n_7984 = n_7834 ^ n_7504;
assign n_7985 = ~n_7341 & n_7835;
assign n_7986 = n_7836 ^ n_7508;
assign n_7987 = ~n_7345 & n_7837;
assign n_7988 = n_7838 ^ n_7509;
assign n_7989 = ~n_7346 & n_7839;
assign n_7990 = n_7840 ^ n_7518;
assign n_7991 = n_7354 & ~n_7841;
assign n_7992 = n_7842 ^ n_7599;
assign n_7993 = ~n_7458 & ~n_7842;
assign n_7994 = n_7458 & n_7842;
assign n_7995 = n_7844 ^ n_7603;
assign n_7996 = n_7845 ^ n_7399;
assign n_7997 = ~x62 & n_7846;
assign n_7998 = n_7847 ^ n_7614;
assign n_7999 = n_7848 ^ n_7619;
assign n_8000 = n_7399 ^ n_7867;
assign n_8001 = n_7868 ^ n_6600;
assign n_8002 = n_7868 ^ n_6475;
assign n_8003 = n_7869 ^ n_7640;
assign n_8004 = ~x0 & n_7890;
assign n_8005 = n_7891 ^ x5;
assign n_8006 = n_7892 ^ x8;
assign n_8007 = n_7893 ^ x11;
assign n_8008 = n_7894 ^ x14;
assign n_8009 = n_7895 ^ x17;
assign n_8010 = n_7896 ^ x20;
assign n_8011 = n_7897 ^ x23;
assign n_8012 = n_7898 ^ x26;
assign n_8013 = n_7899 ^ x29;
assign n_8014 = n_7900 ^ x32;
assign n_8015 = n_7901 ^ x35;
assign n_8016 = n_7902 ^ x38;
assign n_8017 = n_7903 ^ x41;
assign n_8018 = n_7904 ^ x44;
assign n_8019 = n_7905 ^ x47;
assign n_8020 = n_7906 ^ x50;
assign n_8021 = n_7907 ^ x53;
assign n_8022 = n_7908 ^ x56;
assign n_8023 = n_7909 ^ x59;
assign n_8024 = n_7910 ^ x62;
assign n_8025 = n_7911 ^ n_2104;
assign n_8026 = n_5005 ^ n_7912;
assign n_8027 = n_5068 ^ n_7913;
assign n_8028 = n_5131 ^ n_7914;
assign n_8029 = n_5192 ^ n_7915;
assign n_8030 = n_5256 ^ n_7916;
assign n_8031 = n_5320 ^ n_7917;
assign n_8032 = n_5384 ^ n_7918;
assign n_8033 = n_5448 ^ n_7919;
assign n_8034 = n_5509 ^ n_7920;
assign n_8035 = n_5572 ^ n_7921;
assign n_8036 = n_5635 ^ n_7922;
assign n_8037 = n_5699 ^ n_7923;
assign n_8038 = n_5765 ^ n_7924;
assign n_8039 = n_5827 ^ n_7925;
assign n_8040 = n_5891 ^ n_7926;
assign n_8041 = n_5954 ^ n_7927;
assign n_8042 = n_6018 ^ n_7928;
assign n_8043 = n_6082 ^ n_7929;
assign n_8044 = n_6144 ^ n_7930;
assign n_8045 = n_6206 ^ n_7931;
assign n_8046 = n_7932 ^ x78;
assign n_8047 = n_7933 ^ x1;
assign n_8048 = n_655 & n_7934;
assign n_8049 = n_784 & n_7934;
assign n_8050 = ~n_3665 & n_7934;
assign n_8051 = n_854 & n_7934;
assign n_8052 = n_920 & n_7934;
assign n_8053 = n_7934 & n_986;
assign n_8054 = n_7934 & n_1052;
assign n_8055 = n_7934 & n_1117;
assign n_8056 = n_7934 & n_1181;
assign n_8057 = n_7934 & n_1248;
assign n_8058 = n_7934 & n_1314;
assign n_8059 = n_7934 & n_1380;
assign n_8060 = n_7934 & n_1445;
assign n_8061 = n_7934 & n_1510;
assign n_8062 = n_7934 & n_1576;
assign n_8063 = n_7934 & n_1641;
assign n_8064 = n_7934 & n_1706;
assign n_8065 = n_7934 & n_1771;
assign n_8066 = n_7934 & n_1835;
assign n_8067 = n_7934 & n_1899;
assign n_8068 = n_142 & ~n_7935;
assign n_8069 = n_2133 ^ n_7936;
assign n_8070 = n_733 ^ n_7937;
assign n_8071 = n_2204 ^ n_7938;
assign n_8072 = n_2272 ^ n_7939;
assign n_8073 = n_2339 ^ n_7940;
assign n_8074 = n_2406 ^ n_7941;
assign n_8075 = n_2473 ^ n_7942;
assign n_8076 = n_2539 ^ n_7943;
assign n_8077 = n_2604 ^ n_7944;
assign n_8078 = n_2671 ^ n_7945;
assign n_8079 = n_2739 ^ n_7946;
assign n_8080 = n_2806 ^ n_7947;
assign n_8081 = n_2874 ^ n_7948;
assign n_8082 = n_2940 ^ n_7949;
assign n_8083 = n_3009 ^ n_7950;
assign n_8084 = n_3075 ^ n_7951;
assign n_8085 = n_3144 ^ n_7952;
assign n_8086 = n_3208 ^ n_7953;
assign n_8087 = n_3273 ^ n_7954;
assign n_8088 = n_3338 ^ n_7955;
assign n_8089 = n_7956 ^ n_7503;
assign n_8090 = ~n_7340 & n_7957;
assign n_8091 = n_7959 ^ n_7687;
assign n_8092 = n_7961 ^ n_7688;
assign n_8093 = n_7963 ^ n_7689;
assign n_8094 = n_7965 ^ n_7690;
assign n_8095 = n_7967 ^ n_7692;
assign n_8096 = n_7969 ^ n_7694;
assign n_8097 = n_7970 ^ n_7350;
assign n_8098 = n_7970 ^ n_7170;
assign n_8099 = n_7971 ^ n_7480;
assign n_8100 = n_7972 ^ n_7697;
assign n_8101 = n_7974 ^ n_7699;
assign n_8102 = n_7322 ^ n_7975;
assign n_8103 = n_7975 & n_7446;
assign n_8104 = n_7976 ^ n_7502;
assign n_8105 = ~n_7339 & n_7977;
assign n_8106 = n_7617 & ~n_7979;
assign y6 = n_7980;
assign n_8107 = ~n_7463 & n_7981;
assign n_8108 = n_7983 ^ n_7707;
assign n_8109 = n_7985 ^ n_7708;
assign n_8110 = n_7987 ^ n_7709;
assign n_8111 = n_7989 ^ n_7710;
assign n_8112 = n_7991 ^ n_7712;
assign n_8113 = n_7992 ^ n_7006;
assign n_8114 = n_7993 ^ n_7234;
assign n_8115 = ~n_7352 & ~n_7994;
assign n_8116 = n_7995 ^ n_7498;
assign n_8117 = n_7995 ^ n_7197;
assign n_8118 = n_7996 ^ n_7867;
assign n_8119 = n_7997 ^ n_7718;
assign n_8120 = n_7998 ^ n_7888;
assign n_8121 = n_7998 ^ n_7487;
assign n_8122 = ~n_7996 & n_8000;
assign n_8123 = ~n_6600 & ~n_8002;
assign n_8124 = n_8004 ^ n_7763;
assign n_8125 = n_7978 ^ n_8022;
assign n_8126 = n_8024 ^ n_6395;
assign n_8127 = ~x0 & n_8025;
assign n_8128 = n_8026 ^ x5;
assign n_8129 = n_8027 ^ x8;
assign n_8130 = n_8028 ^ x11;
assign n_8131 = n_8029 ^ x14;
assign n_8132 = n_8030 ^ x17;
assign n_8133 = n_8031 ^ x20;
assign n_8134 = n_8032 ^ x23;
assign n_8135 = n_8033 ^ x26;
assign n_8136 = n_8034 ^ x29;
assign n_8137 = n_8035 ^ x32;
assign n_8138 = n_8036 ^ x35;
assign n_8139 = n_8037 ^ x38;
assign n_8140 = n_8038 ^ x41;
assign n_8141 = n_8039 ^ x44;
assign n_8142 = n_8040 ^ x47;
assign n_8143 = n_8041 ^ x50;
assign n_8144 = n_8042 ^ x53;
assign n_8145 = n_8043 ^ x56;
assign n_8146 = n_8044 ^ x59;
assign n_8147 = n_8045 ^ x62;
assign n_8148 = n_8046 ^ n_2105;
assign n_8149 = n_8047 ^ x79;
assign n_8150 = n_2134 ^ n_8048;
assign n_8151 = n_734 ^ n_8049;
assign n_8152 = n_2205 ^ n_8050;
assign n_8153 = n_2273 ^ n_8051;
assign n_8154 = n_2340 ^ n_8052;
assign n_8155 = n_2407 ^ n_8053;
assign n_8156 = n_2474 ^ n_8054;
assign n_8157 = n_2540 ^ n_8055;
assign n_8158 = n_2605 ^ n_8056;
assign n_8159 = n_2672 ^ n_8057;
assign n_8160 = n_2740 ^ n_8058;
assign n_8161 = n_2807 ^ n_8059;
assign n_8162 = n_2875 ^ n_8060;
assign n_8163 = n_2941 ^ n_8061;
assign n_8164 = n_3010 ^ n_8062;
assign n_8165 = n_3076 ^ n_8063;
assign n_8166 = n_3145 ^ n_8064;
assign n_8167 = n_3209 ^ n_8065;
assign n_8168 = n_3274 ^ n_8066;
assign n_8169 = n_3339 ^ n_8067;
assign n_8170 = n_1 & ~n_8068;
assign n_8171 = ~n_8068 & n_145;
assign n_8172 = n_8068 ^ x80;
assign n_8173 = n_5006 ^ n_8069;
assign n_8174 = n_5069 ^ n_8070;
assign n_8175 = n_5132 ^ n_8071;
assign n_8176 = n_5193 ^ n_8072;
assign n_8177 = n_5257 ^ n_8073;
assign n_8178 = n_5321 ^ n_8074;
assign n_8179 = n_5385 ^ n_8075;
assign n_8180 = n_5449 ^ n_8076;
assign n_8181 = n_5510 ^ n_8077;
assign n_8182 = n_5573 ^ n_8078;
assign n_8183 = n_5636 ^ n_8079;
assign n_8184 = n_5700 ^ n_8080;
assign n_8185 = n_5766 ^ n_8081;
assign n_8186 = n_5828 ^ n_8082;
assign n_8187 = n_5892 ^ n_8083;
assign n_8188 = n_5955 ^ n_8084;
assign n_8189 = n_6019 ^ n_8085;
assign n_8190 = n_6083 ^ n_8086;
assign n_8191 = n_6145 ^ n_8087;
assign n_8192 = n_6207 ^ n_8088;
assign n_8193 = n_8090 ^ n_7809;
assign n_8194 = n_8091 ^ n_7342;
assign n_8195 = n_8091 ^ n_7159;
assign n_8196 = n_8092 ^ n_7343;
assign n_8197 = n_8092 ^ n_7161;
assign n_8198 = n_8093 ^ n_7344;
assign n_8199 = n_8093 ^ n_7226;
assign n_8200 = n_8094 ^ n_7347;
assign n_8201 = n_8094 ^ n_7165;
assign n_8202 = n_8095 ^ n_7348;
assign n_8203 = n_8095 ^ n_7167;
assign n_8204 = n_8096 ^ n_7349;
assign n_8205 = n_8096 ^ n_7001;
assign n_8206 = n_7513 ^ n_8097;
assign n_8207 = ~n_7350 & n_8098;
assign n_8208 = n_8100 ^ n_7351;
assign n_8209 = n_8100 ^ n_6887;
assign n_8210 = n_8101 ^ n_7353;
assign n_8211 = n_8101 ^ n_7015;
assign n_8212 = n_7517 ^ n_8102;
assign n_8213 = n_8103 ^ n_7827;
assign n_8214 = n_8105 ^ n_7828;
assign n_8215 = n_8106 ^ n_7830;
assign n_8216 = n_8107 ^ n_7831;
assign n_8217 = n_8108 ^ n_7489;
assign n_8218 = n_8108 ^ n_7320;
assign n_8219 = n_8109 ^ n_7570;
assign n_8220 = n_8109 ^ n_7429;
assign n_8221 = n_8110 ^ n_7387;
assign n_8222 = n_8111 ^ n_7576;
assign n_8223 = n_8111 ^ n_7435;
assign n_8224 = n_8112 ^ n_7497;
assign n_8225 = n_8112 ^ n_7397;
assign n_8226 = n_8113 ^ n_7352;
assign n_8227 = n_8114 & ~n_8115;
assign n_8228 = n_8116 ^ n_7866;
assign n_8229 = n_7498 & n_8117;
assign n_8230 = n_8119 ^ n_4951;
assign n_8231 = n_8120 ^ n_7487;
assign n_8232 = n_8120 & n_8121;
assign n_8233 = n_8122 ^ n_7845;
assign n_8234 = n_8123 ^ n_7868;
assign n_8235 = n_8127 ^ n_7911;
assign n_8236 = n_8118 ^ n_8145;
assign n_8237 = n_8146 ^ n_8001;
assign n_8238 = n_8147 ^ n_6635;
assign n_8239 = n_8147 ^ n_6523;
assign n_8240 = ~x0 & n_8148;
assign n_8241 = n_8149 ^ n_3468;
assign n_8242 = n_5007 ^ n_8150;
assign n_8243 = n_5070 ^ n_8151;
assign n_8244 = n_5133 ^ n_8152;
assign n_8245 = n_5194 ^ n_8153;
assign n_8246 = n_5258 ^ n_8154;
assign n_8247 = n_5322 ^ n_8155;
assign n_8248 = n_5386 ^ n_8156;
assign n_8249 = n_5450 ^ n_8157;
assign n_8250 = n_5511 ^ n_8158;
assign n_8251 = n_5574 ^ n_8159;
assign n_8252 = n_5637 ^ n_8160;
assign n_8253 = n_5701 ^ n_8161;
assign n_8254 = n_5767 ^ n_8162;
assign n_8255 = n_5829 ^ n_8163;
assign n_8256 = n_5893 ^ n_8164;
assign n_8257 = n_5956 ^ n_8165;
assign n_8258 = n_6020 ^ n_8166;
assign n_8259 = n_6084 ^ n_8167;
assign n_8260 = n_6146 ^ n_8168;
assign n_8261 = n_6208 ^ n_8169;
assign n_8262 = n_8170 ^ x1;
assign n_8263 = n_1 & ~n_8171;
assign n_8264 = ~n_8171 & n_149;
assign n_8265 = n_8171 ^ x81;
assign n_8266 = n_655 & n_8172;
assign n_8267 = n_784 & n_8172;
assign n_8268 = ~n_3665 & n_8172;
assign n_8269 = n_854 & n_8172;
assign n_8270 = n_920 & n_8172;
assign n_8271 = n_8172 & n_986;
assign n_8272 = n_8172 & n_1052;
assign n_8273 = n_8172 & n_1117;
assign n_8274 = n_8172 & n_1181;
assign n_8275 = n_8172 & n_1248;
assign n_8276 = n_8172 & n_1314;
assign n_8277 = n_8172 & n_1380;
assign n_8278 = n_8172 & n_1445;
assign n_8279 = n_8172 & n_1510;
assign n_8280 = n_8172 & n_1576;
assign n_8281 = n_8172 & n_1641;
assign n_8282 = n_8172 & n_1706;
assign n_8283 = n_8172 & n_1771;
assign n_8284 = n_8172 & n_1835;
assign n_8285 = n_8172 & n_1899;
assign n_8286 = n_8173 ^ x5;
assign n_8287 = n_8174 ^ x8;
assign n_8288 = n_8175 ^ x11;
assign n_8289 = n_8176 ^ x14;
assign n_8290 = n_8177 ^ x17;
assign n_8291 = n_8178 ^ x20;
assign n_8292 = n_8179 ^ x23;
assign n_8293 = n_8180 ^ x26;
assign n_8294 = n_8181 ^ x29;
assign n_8295 = n_8182 ^ x32;
assign n_8296 = n_8183 ^ x35;
assign n_8297 = n_8184 ^ x38;
assign n_8298 = n_8185 ^ x41;
assign n_8299 = n_8186 ^ x44;
assign n_8300 = n_8187 ^ x47;
assign n_8301 = n_8188 ^ x50;
assign n_8302 = n_8189 ^ x53;
assign n_8303 = n_8190 ^ x56;
assign n_8304 = n_8191 ^ x59;
assign n_8305 = n_8192 ^ x62;
assign n_8306 = n_8193 ^ n_7491;
assign n_8307 = n_8193 ^ n_7176;
assign n_8308 = n_8194 ^ n_7505;
assign n_8309 = ~n_7342 & n_8195;
assign n_8310 = n_8196 ^ n_7506;
assign n_8311 = ~n_7343 & n_8197;
assign n_8312 = n_8198 ^ n_7507;
assign n_8313 = n_7344 & n_8199;
assign n_8314 = n_8200 ^ n_7510;
assign n_8315 = ~n_7347 & n_8201;
assign n_8316 = n_8202 ^ n_7511;
assign n_8317 = ~n_7348 & n_8203;
assign n_8318 = n_8204 ^ n_7512;
assign n_8319 = n_7349 & ~n_8205;
assign n_8320 = n_8207 ^ n_7970;
assign n_8321 = n_8208 ^ n_7514;
assign n_8322 = n_7351 & ~n_8209;
assign n_8323 = n_8210 ^ n_7516;
assign n_8324 = ~n_7353 & n_8211;
assign n_8325 = n_8213 ^ n_7496;
assign n_8326 = n_8213 ^ n_7179;
assign n_8327 = n_8214 ^ n_7490;
assign n_8328 = n_8214 ^ n_7307;
assign n_8329 = n_8215 ^ n_8118;
assign n_8330 = n_8216 ^ n_7605;
assign n_8331 = n_8216 ^ n_7186;
assign n_8332 = n_8217 ^ n_7999;
assign n_8333 = ~n_7489 & n_8218;
assign n_8334 = n_8219 ^ n_7851;
assign n_8335 = ~n_7570 & n_8220;
assign n_8336 = n_8221 ^ n_7192;
assign n_8337 = n_8221 & ~n_7493;
assign n_8338 = n_8222 ^ n_7856;
assign n_8339 = ~n_7576 & n_8223;
assign n_8340 = n_8224 ^ n_7865;
assign n_8341 = ~n_7497 & n_8225;
assign n_8342 = n_8226 ^ n_7515;
assign n_8343 = n_8227 ^ n_7172;
assign n_8344 = n_8229 ^ n_7995;
assign n_8345 = n_8230 ^ n_7521;
assign n_8346 = n_8230 & ~n_7618;
assign n_8347 = n_8232 ^ n_7888;
assign n_8348 = n_8233 ^ n_8231;
assign n_8349 = n_8234 ^ n_6752;
assign n_8350 = ~n_6258 & ~n_8234;
assign n_8351 = n_8215 ^ n_8236;
assign n_8352 = n_6635 & n_8239;
assign n_8353 = n_8240 ^ n_8046;
assign n_8354 = ~x0 & n_8241;
assign n_8355 = n_8242 ^ x5;
assign n_8356 = n_8243 ^ x8;
assign n_8357 = n_8244 ^ x11;
assign n_8358 = n_8245 ^ x14;
assign n_8359 = n_8246 ^ x17;
assign n_8360 = n_8247 ^ x20;
assign n_8361 = n_8248 ^ x23;
assign n_8362 = n_8249 ^ x26;
assign n_8363 = n_8250 ^ x29;
assign n_8364 = n_8251 ^ x32;
assign n_8365 = n_8252 ^ x35;
assign n_8366 = n_8253 ^ x38;
assign n_8367 = n_8254 ^ x41;
assign n_8368 = n_8255 ^ x44;
assign n_8369 = n_8256 ^ x47;
assign n_8370 = n_8257 ^ x50;
assign n_8371 = n_8258 ^ x53;
assign n_8372 = n_8259 ^ x56;
assign n_8373 = n_8260 ^ x59;
assign n_8374 = n_8261 ^ x62;
assign n_8375 = n_8262 ^ x80;
assign n_8376 = n_8263 ^ x1;
assign n_8377 = n_1 & ~n_8264;
assign n_8378 = ~n_8264 & n_153;
assign n_8379 = n_8264 ^ x82;
assign n_8380 = n_655 & n_8265;
assign n_8381 = n_784 & n_8265;
assign n_8382 = ~n_3665 & n_8265;
assign n_8383 = n_854 & n_8265;
assign n_8384 = n_920 & n_8265;
assign n_8385 = n_8265 & n_986;
assign n_8386 = n_8265 & n_1052;
assign n_8387 = n_8265 & n_1117;
assign n_8388 = n_8265 & n_1181;
assign n_8389 = n_8265 & n_1248;
assign n_8390 = n_8265 & n_1314;
assign n_8391 = n_8265 & n_1380;
assign n_8392 = n_8265 & n_1445;
assign n_8393 = n_8265 & n_1510;
assign n_8394 = n_8265 & n_1576;
assign n_8395 = n_8265 & n_1641;
assign n_8396 = n_8265 & n_1706;
assign n_8397 = n_8265 & n_1771;
assign n_8398 = n_8265 & n_1835;
assign n_8399 = n_8265 & n_1899;
assign n_8400 = n_2135 ^ n_8266;
assign n_8401 = n_735 ^ n_8267;
assign n_8402 = n_2206 ^ n_8268;
assign n_8403 = n_2274 ^ n_8269;
assign n_8404 = n_2341 ^ n_8270;
assign n_8405 = n_2408 ^ n_8271;
assign n_8406 = n_2475 ^ n_8272;
assign n_8407 = n_2541 ^ n_8273;
assign n_8408 = n_2606 ^ n_8274;
assign n_8409 = n_2673 ^ n_8275;
assign n_8410 = n_2741 ^ n_8276;
assign n_8411 = n_2808 ^ n_8277;
assign n_8412 = n_2876 ^ n_8278;
assign n_8413 = n_2942 ^ n_8279;
assign n_8414 = n_3011 ^ n_8280;
assign n_8415 = n_3077 ^ n_8281;
assign n_8416 = n_3146 ^ n_8282;
assign n_8417 = n_3210 ^ n_8283;
assign n_8418 = n_3275 ^ n_8284;
assign n_8419 = n_3340 ^ n_8285;
assign n_8420 = n_8233 ^ n_8303;
assign n_8421 = n_8304 ^ n_7889;
assign n_8422 = n_8306 ^ n_7850;
assign n_8423 = ~n_7491 & n_8307;
assign n_8424 = n_8309 ^ n_8091;
assign n_8425 = n_8311 ^ n_8092;
assign n_8426 = n_8313 ^ n_8093;
assign n_8427 = n_8315 ^ n_8094;
assign n_8428 = n_8317 ^ n_8095;
assign n_8429 = n_8319 ^ n_8096;
assign n_8430 = n_8320 ^ n_7392;
assign n_8431 = n_8322 ^ n_8100;
assign n_8432 = n_8324 ^ n_8101;
assign n_8433 = n_8325 ^ n_7864;
assign n_8434 = ~n_7496 & n_8326;
assign n_8435 = n_8327 ^ n_7849;
assign n_8436 = ~n_7490 & n_8328;
assign n_8437 = ~n_8236 & ~n_8329;
assign y7 = ~n_8330;
assign n_8438 = n_7605 & ~n_8331;
assign n_8439 = n_8333 ^ n_8108;
assign n_8440 = n_8335 ^ n_8109;
assign n_8441 = n_8336 ^ n_7855;
assign n_8442 = n_8337 ^ n_8110;
assign n_8443 = n_8339 ^ n_8111;
assign n_8444 = n_8341 ^ n_8112;
assign n_8445 = n_7394 ^ n_8343;
assign n_8446 = n_8344 ^ n_7829;
assign n_8447 = n_8344 ^ n_7704;
assign n_8448 = n_8345 ^ n_8023;
assign n_8449 = n_8346 ^ n_8119;
assign n_8450 = n_8345 ^ n_8347;
assign n_8451 = n_7889 ^ n_8349;
assign n_8452 = ~n_6394 & ~n_8350;
assign n_8453 = n_8352 ^ n_8147;
assign n_8454 = n_8354 ^ n_8149;
assign n_8455 = n_8374 ^ n_6336;
assign n_8456 = n_8375 ^ n_2106;
assign n_8457 = n_8376 ^ x81;
assign n_8458 = n_8377 ^ x1;
assign n_8459 = n_1 & ~n_8378;
assign n_8460 = ~n_8378 & n_157;
assign n_8461 = n_8378 ^ x83;
assign n_8462 = n_655 & n_8379;
assign n_8463 = n_784 & n_8379;
assign n_8464 = ~n_3665 & n_8379;
assign n_8465 = n_854 & n_8379;
assign n_8466 = n_920 & n_8379;
assign n_8467 = n_986 & n_8379;
assign n_8468 = n_8379 & n_1052;
assign n_8469 = n_8379 & n_1117;
assign n_8470 = n_8379 & n_1181;
assign n_8471 = n_8379 & n_1248;
assign n_8472 = n_8379 & n_1314;
assign n_8473 = n_8379 & n_1380;
assign n_8474 = n_8379 & n_1445;
assign n_8475 = n_8379 & n_1510;
assign n_8476 = n_8379 & n_1576;
assign n_8477 = n_8379 & n_1641;
assign n_8478 = n_8379 & n_1706;
assign n_8479 = n_8379 & n_1771;
assign n_8480 = n_8379 & n_1835;
assign n_8481 = n_8379 & n_1899;
assign n_8482 = n_2136 ^ n_8380;
assign n_8483 = n_736 ^ n_8381;
assign n_8484 = n_2207 ^ n_8382;
assign n_8485 = n_2275 ^ n_8383;
assign n_8486 = n_2342 ^ n_8384;
assign n_8487 = n_2409 ^ n_8385;
assign n_8488 = n_2476 ^ n_8386;
assign n_8489 = n_2542 ^ n_8387;
assign n_8490 = n_2607 ^ n_8388;
assign n_8491 = n_2674 ^ n_8389;
assign n_8492 = n_2742 ^ n_8390;
assign n_8493 = n_2809 ^ n_8391;
assign n_8494 = n_2877 ^ n_8392;
assign n_8495 = n_2943 ^ n_8393;
assign n_8496 = n_3012 ^ n_8394;
assign n_8497 = n_3078 ^ n_8395;
assign n_8498 = n_3147 ^ n_8396;
assign n_8499 = n_3211 ^ n_8397;
assign n_8500 = n_3276 ^ n_8398;
assign n_8501 = n_3341 ^ n_8399;
assign n_8502 = n_5008 ^ n_8400;
assign n_8503 = n_5071 ^ n_8401;
assign n_8504 = n_5134 ^ n_8402;
assign n_8505 = n_5195 ^ n_8403;
assign n_8506 = n_5259 ^ n_8404;
assign n_8507 = n_5323 ^ n_8405;
assign n_8508 = n_5387 ^ n_8406;
assign n_8509 = n_5451 ^ n_8407;
assign n_8510 = n_5512 ^ n_8408;
assign n_8511 = n_5575 ^ n_8409;
assign n_8512 = n_5638 ^ n_8410;
assign n_8513 = n_5702 ^ n_8411;
assign n_8514 = n_5768 ^ n_8412;
assign n_8515 = n_5830 ^ n_8413;
assign n_8516 = n_5894 ^ n_8414;
assign n_8517 = n_5957 ^ n_8415;
assign n_8518 = n_6021 ^ n_8416;
assign n_8519 = n_6085 ^ n_8417;
assign n_8520 = n_6147 ^ n_8418;
assign n_8521 = n_6209 ^ n_8419;
assign n_8522 = n_8420 ^ n_8231;
assign n_8523 = n_8420 & n_8348;
assign n_8524 = n_8421 ^ n_8349;
assign n_8525 = n_8423 ^ n_8193;
assign n_8526 = n_8424 ^ n_7572;
assign n_8527 = n_8424 ^ n_7431;
assign n_8528 = n_8425 ^ n_7574;
assign n_8529 = n_8425 ^ n_7433;
assign n_8530 = n_8426 ^ n_7492;
assign n_8531 = n_8426 ^ n_7386;
assign n_8532 = n_8427 ^ n_7691;
assign n_8533 = n_8427 ^ n_7578;
assign n_8534 = n_8428 ^ n_7390;
assign n_8535 = n_8429 ^ n_7582;
assign n_8536 = n_8429 ^ n_7439;
assign n_8537 = n_8430 ^ n_7441;
assign n_8538 = n_8430 & ~n_7584;
assign n_8539 = n_8431 ^ n_7494;
assign n_8540 = n_8431 ^ n_7177;
assign n_8541 = n_8432 ^ n_7495;
assign n_8542 = n_8432 ^ n_7195;
assign n_8543 = n_8434 ^ n_8213;
assign n_8544 = n_8436 ^ n_8214;
assign n_8545 = n_8437 ^ n_8145;
assign n_8546 = n_8438 ^ n_8216;
assign n_8547 = n_8439 ^ n_7702;
assign n_8548 = n_8439 ^ n_7590;
assign n_8549 = n_8440 ^ n_7958;
assign n_8550 = n_8440 ^ n_7810;
assign n_8551 = n_8442 ^ n_7609;
assign n_8552 = n_8442 ^ n_7456;
assign n_8553 = n_8443 ^ n_7964;
assign n_8554 = n_8443 ^ n_7816;
assign n_8555 = n_8444 ^ n_7611;
assign n_8556 = n_8444 ^ n_7447;
assign n_8557 = n_8445 ^ n_7586;
assign n_8558 = n_8445 & ~n_7698;
assign n_8559 = n_7887 ^ n_8446;
assign n_8560 = n_7829 & n_8447;
assign n_8561 = n_8448 ^ n_8347;
assign n_8562 = n_8449 ^ n_8237;
assign n_8563 = n_8449 ^ n_8146;
assign n_8564 = ~n_8448 & n_8450;
assign n_8565 = n_8421 & n_8451;
assign n_8566 = n_8452 ^ n_8126;
assign n_8567 = n_8452 ^ n_8024;
assign n_8568 = n_8453 ^ n_6601;
assign n_8569 = ~n_6476 & ~n_8453;
assign n_8570 = ~x0 & n_8456;
assign n_8571 = n_8457 ^ n_6479;
assign n_8572 = n_8458 ^ x82;
assign n_8573 = n_8459 ^ x1;
assign n_8574 = n_1 & ~n_8460;
assign n_8575 = ~n_8460 & n_160;
assign n_8576 = n_8460 ^ x84;
assign n_8577 = n_655 & n_8461;
assign n_8578 = n_784 & n_8461;
assign n_8579 = ~n_3665 & n_8461;
assign n_8580 = n_854 & n_8461;
assign n_8581 = n_920 & n_8461;
assign n_8582 = n_986 & n_8461;
assign n_8583 = n_8461 & n_1052;
assign n_8584 = n_8461 & n_1117;
assign n_8585 = n_8461 & n_1181;
assign n_8586 = n_8461 & n_1248;
assign n_8587 = n_8461 & n_1314;
assign n_8588 = n_8461 & n_1380;
assign n_8589 = n_8461 & n_1445;
assign n_8590 = n_8461 & n_1510;
assign n_8591 = n_8461 & n_1576;
assign n_8592 = n_8461 & n_1641;
assign n_8593 = n_8461 & n_1706;
assign n_8594 = n_8461 & n_1771;
assign n_8595 = n_8461 & n_1835;
assign n_8596 = n_8461 & n_1899;
assign n_8597 = n_2137 ^ n_8462;
assign n_8598 = n_737 ^ n_8463;
assign n_8599 = n_2208 ^ n_8464;
assign n_8600 = n_2276 ^ n_8465;
assign n_8601 = n_2343 ^ n_8466;
assign n_8602 = n_2410 ^ n_8467;
assign n_8603 = n_2477 ^ n_8468;
assign n_8604 = n_2543 ^ n_8469;
assign n_8605 = n_2608 ^ n_8470;
assign n_8606 = n_2675 ^ n_8471;
assign n_8607 = n_2743 ^ n_8472;
assign n_8608 = n_2810 ^ n_8473;
assign n_8609 = n_2878 ^ n_8474;
assign n_8610 = n_2944 ^ n_8475;
assign n_8611 = n_3013 ^ n_8476;
assign n_8612 = n_3079 ^ n_8477;
assign n_8613 = n_3148 ^ n_8478;
assign n_8614 = n_3212 ^ n_8479;
assign n_8615 = n_3277 ^ n_8480;
assign n_8616 = n_3342 ^ n_8481;
assign n_8617 = n_5009 ^ n_8482;
assign n_8618 = n_5072 ^ n_8483;
assign n_8619 = n_5135 ^ n_8484;
assign n_8620 = n_5196 ^ n_8485;
assign n_8621 = n_5260 ^ n_8486;
assign n_8622 = n_5324 ^ n_8487;
assign n_8623 = n_5388 ^ n_8488;
assign n_8624 = n_5452 ^ n_8489;
assign n_8625 = n_5513 ^ n_8490;
assign n_8626 = n_5576 ^ n_8491;
assign n_8627 = n_5639 ^ n_8492;
assign n_8628 = n_5703 ^ n_8493;
assign n_8629 = n_5769 ^ n_8494;
assign n_8630 = n_5831 ^ n_8495;
assign n_8631 = n_5895 ^ n_8496;
assign n_8632 = n_5958 ^ n_8497;
assign n_8633 = n_6022 ^ n_8498;
assign n_8634 = n_6086 ^ n_8499;
assign n_8635 = n_6148 ^ n_8500;
assign n_8636 = n_6210 ^ n_8501;
assign n_8637 = n_8502 ^ x5;
assign n_8638 = n_8503 ^ x8;
assign n_8639 = n_8504 ^ x11;
assign n_8640 = n_8505 ^ x14;
assign n_8641 = n_8506 ^ x17;
assign n_8642 = n_8507 ^ x20;
assign n_8643 = n_8508 ^ x23;
assign n_8644 = n_8509 ^ x26;
assign n_8645 = n_8510 ^ x29;
assign n_8646 = n_8511 ^ x32;
assign n_8647 = n_8512 ^ x35;
assign n_8648 = n_8513 ^ x38;
assign n_8649 = n_8514 ^ x41;
assign n_8650 = n_8515 ^ x44;
assign n_8651 = n_8516 ^ x47;
assign n_8652 = n_8517 ^ x50;
assign n_8653 = n_8518 ^ x53;
assign n_8654 = n_8519 ^ x56;
assign n_8655 = n_8520 ^ x59;
assign n_8656 = n_8521 ^ x62;
assign n_8657 = n_8523 ^ n_8303;
assign n_8658 = n_8525 ^ n_7607;
assign n_8659 = n_8525 ^ n_7452;
assign n_8660 = n_8526 ^ n_7852;
assign n_8661 = ~n_7572 & n_8527;
assign n_8662 = n_8528 ^ n_7853;
assign n_8663 = ~n_7574 & n_8529;
assign n_8664 = n_8530 ^ n_7854;
assign n_8665 = ~n_7492 & n_8531;
assign n_8666 = n_8532 ^ n_7857;
assign n_8667 = ~n_7691 & n_8533;
assign n_8668 = n_8534 ^ n_7580;
assign n_8669 = n_8534 & ~n_7693;
assign n_8670 = n_8535 ^ n_7859;
assign n_8671 = ~n_7582 & n_8536;
assign n_8672 = n_8537 ^ n_7860;
assign n_8673 = n_8538 ^ n_8320;
assign n_8674 = n_8539 ^ n_7861;
assign n_8675 = ~n_7494 & n_8540;
assign n_8676 = n_8541 ^ n_7863;
assign n_8677 = ~n_7495 & n_8542;
assign n_8678 = n_8543 ^ n_7711;
assign n_8679 = n_8543 ^ n_7600;
assign n_8680 = n_8544 ^ n_7685;
assign n_8681 = n_8544 ^ n_7568;
assign n_8682 = n_8522 ^ n_8545;
assign n_8683 = n_8546 ^ n_7717;
assign n_8684 = n_8546 ^ n_7450;
assign n_8685 = n_8547 ^ n_8003;
assign n_8686 = n_7702 & ~n_8548;
assign n_8687 = n_8549 ^ n_7872;
assign n_8688 = ~n_7958 & n_8550;
assign n_8689 = n_8551 ^ n_7876;
assign n_8690 = ~n_7609 & n_8552;
assign n_8691 = n_8553 ^ n_7877;
assign n_8692 = ~n_7964 & n_8554;
assign n_8693 = n_7886 ^ n_8555;
assign n_8694 = ~n_7611 & n_8556;
assign n_8695 = n_8557 ^ n_7862;
assign n_8696 = n_8558 ^ n_8343;
assign n_8697 = n_8560 ^ n_8344;
assign n_8698 = n_8372 ^ n_8561;
assign n_8699 = ~n_8237 & n_8563;
assign n_8700 = n_8564 ^ n_8347;
assign n_8701 = n_8565 ^ n_8304;
assign n_8702 = n_8373 ^ n_8566;
assign n_8703 = n_8126 & n_8567;
assign n_8704 = n_8568 ^ n_8305;
assign n_8705 = ~n_4893 & ~n_8569;
assign n_8706 = n_8570 ^ n_8375;
assign n_8707 = ~x0 & ~n_8571;
assign n_8708 = n_8572 ^ n_3473;
assign n_8709 = n_8573 ^ x83;
assign n_8710 = n_8574 ^ x1;
assign n_8711 = n_1 & ~n_8575;
assign n_8712 = ~n_8575 & n_164;
assign n_8713 = n_8575 ^ x85;
assign n_8714 = n_655 & n_8576;
assign n_8715 = n_784 & n_8576;
assign n_8716 = ~n_3665 & n_8576;
assign n_8717 = n_854 & n_8576;
assign n_8718 = n_920 & n_8576;
assign n_8719 = n_986 & n_8576;
assign n_8720 = n_8576 & n_1052;
assign n_8721 = n_8576 & n_1117;
assign n_8722 = n_8576 & n_1181;
assign n_8723 = n_8576 & n_1248;
assign n_8724 = n_8576 & n_1314;
assign n_8725 = n_8576 & n_1380;
assign n_8726 = n_8576 & n_1445;
assign n_8727 = n_8576 & n_1510;
assign n_8728 = n_8576 & n_1576;
assign n_8729 = n_8576 & n_1641;
assign n_8730 = n_8576 & n_1706;
assign n_8731 = n_8576 & n_1771;
assign n_8732 = n_8576 & n_1835;
assign n_8733 = n_8576 & n_1899;
assign n_8734 = n_2138 ^ n_8577;
assign n_8735 = n_738 ^ n_8578;
assign n_8736 = n_2209 ^ n_8579;
assign n_8737 = n_2277 ^ n_8580;
assign n_8738 = n_2344 ^ n_8581;
assign n_8739 = n_2411 ^ n_8582;
assign n_8740 = n_2478 ^ n_8583;
assign n_8741 = n_2544 ^ n_8584;
assign n_8742 = n_2609 ^ n_8585;
assign n_8743 = n_2676 ^ n_8586;
assign n_8744 = n_2744 ^ n_8587;
assign n_8745 = n_2811 ^ n_8588;
assign n_8746 = n_2879 ^ n_8589;
assign n_8747 = n_2945 ^ n_8590;
assign n_8748 = n_3014 ^ n_8591;
assign n_8749 = n_3080 ^ n_8592;
assign n_8750 = n_3149 ^ n_8593;
assign n_8751 = n_3213 ^ n_8594;
assign n_8752 = n_3278 ^ n_8595;
assign n_8753 = n_3343 ^ n_8596;
assign n_8754 = n_5010 ^ n_8597;
assign n_8755 = n_5073 ^ n_8598;
assign n_8756 = n_5136 ^ n_8599;
assign n_8757 = n_5197 ^ n_8600;
assign n_8758 = n_5261 ^ n_8601;
assign n_8759 = n_5325 ^ n_8602;
assign n_8760 = n_5389 ^ n_8603;
assign n_8761 = n_5453 ^ n_8604;
assign n_8762 = n_5514 ^ n_8605;
assign n_8763 = n_5577 ^ n_8606;
assign n_8764 = n_5640 ^ n_8607;
assign n_8765 = n_5704 ^ n_8608;
assign n_8766 = n_5770 ^ n_8609;
assign n_8767 = n_5832 ^ n_8610;
assign n_8768 = n_5896 ^ n_8611;
assign n_8769 = n_5959 ^ n_8612;
assign n_8770 = n_6023 ^ n_8613;
assign n_8771 = n_6087 ^ n_8614;
assign n_8772 = n_6149 ^ n_8615;
assign n_8773 = n_6211 ^ n_8616;
assign n_8774 = n_8617 ^ x5;
assign n_8775 = n_8618 ^ x8;
assign n_8776 = n_8619 ^ x11;
assign n_8777 = n_8620 ^ x14;
assign n_8778 = n_8621 ^ x17;
assign n_8779 = n_8622 ^ x20;
assign n_8780 = n_8623 ^ x23;
assign n_8781 = n_8624 ^ x26;
assign n_8782 = n_8625 ^ x29;
assign n_8783 = n_8626 ^ x32;
assign n_8784 = n_8627 ^ x35;
assign n_8785 = n_8628 ^ x38;
assign n_8786 = n_8629 ^ x41;
assign n_8787 = n_8630 ^ x44;
assign n_8788 = n_8631 ^ x47;
assign n_8789 = n_8632 ^ x50;
assign n_8790 = n_8633 ^ x53;
assign n_8791 = n_8634 ^ x56;
assign n_8792 = n_8635 ^ x59;
assign n_8793 = n_4956 ^ n_8636;
assign n_8794 = n_8636 ^ x77;
assign n_8795 = n_8636 & ~n_548;
assign n_8796 = n_8636 ^ x78;
assign n_8797 = n_8653 ^ n_8351;
assign n_8798 = n_8654 ^ n_8562;
assign n_8799 = n_8655 ^ n_8238;
assign n_8800 = n_8656 ^ n_6602;
assign n_8801 = n_8656 ^ n_6477;
assign n_8802 = n_8657 ^ n_8372;
assign n_8803 = n_8658 ^ n_7871;
assign n_8804 = ~n_7607 & n_8659;
assign n_8805 = n_8661 ^ n_8424;
assign n_8806 = n_8663 ^ n_8425;
assign n_8807 = n_8665 ^ n_8426;
assign n_8808 = n_8667 ^ n_8427;
assign n_8809 = n_8668 ^ n_7858;
assign n_8810 = n_8669 ^ n_8428;
assign n_8811 = n_8671 ^ n_8429;
assign n_8812 = n_8673 ^ n_7971;
assign n_8813 = n_8675 ^ n_8431;
assign n_8814 = n_8677 ^ n_8432;
assign n_8815 = n_7885 ^ n_8678;
assign n_8816 = ~n_7711 & n_8679;
assign n_8817 = n_8680 ^ n_7870;
assign n_8818 = ~n_7685 & n_8681;
assign y8 = ~n_8683;
assign n_8819 = n_7717 & ~n_8684;
assign n_8820 = n_8686 ^ n_8439;
assign n_8821 = n_8688 ^ n_8440;
assign n_8822 = n_8690 ^ n_8442;
assign n_8823 = n_8692 ^ n_8443;
assign n_8824 = n_8694 ^ n_8444;
assign n_8825 = n_8696 ^ n_7973;
assign n_8826 = n_8696 ^ n_7825;
assign n_8827 = n_8697 ^ n_8125;
assign n_8828 = n_8697 ^ n_7978;
assign n_8829 = n_8699 ^ n_8449;
assign n_8830 = n_8562 ^ n_8700;
assign n_8831 = n_8701 ^ n_8373;
assign n_8832 = n_8703 ^ n_8452;
assign n_8833 = n_8705 ^ n_8455;
assign n_8834 = n_8705 ^ n_8374;
assign n_8835 = n_8707 ^ n_8457;
assign n_8836 = ~x0 & n_8708;
assign n_8837 = n_8709 ^ n_2107;
assign n_8838 = n_8710 ^ x84;
assign n_8839 = n_8711 ^ x1;
assign n_8840 = n_1 & ~n_8712;
assign n_8841 = ~n_8712 & n_168;
assign n_8842 = n_8712 ^ x86;
assign n_8843 = n_655 & n_8713;
assign n_8844 = n_784 & n_8713;
assign n_8845 = ~n_3665 & n_8713;
assign n_8846 = n_854 & n_8713;
assign n_8847 = n_920 & n_8713;
assign n_8848 = n_986 & n_8713;
assign n_8849 = n_1052 & n_8713;
assign n_8850 = n_8713 & n_1117;
assign n_8851 = n_8713 & n_1181;
assign n_8852 = n_8713 & n_1248;
assign n_8853 = n_8713 & n_1314;
assign n_8854 = n_8713 & n_1380;
assign n_8855 = n_8713 & n_1445;
assign n_8856 = n_8713 & n_1510;
assign n_8857 = n_8713 & n_1576;
assign n_8858 = n_8713 & n_1641;
assign n_8859 = n_8713 & n_1706;
assign n_8860 = n_8713 & n_1771;
assign n_8861 = n_8713 & n_1835;
assign n_8862 = n_8713 & n_1899;
assign n_8863 = n_2139 ^ n_8714;
assign n_8864 = n_739 ^ n_8715;
assign n_8865 = n_2210 ^ n_8716;
assign n_8866 = n_2278 ^ n_8717;
assign n_8867 = n_2345 ^ n_8718;
assign n_8868 = n_2412 ^ n_8719;
assign n_8869 = n_2479 ^ n_8720;
assign n_8870 = n_2545 ^ n_8721;
assign n_8871 = n_2610 ^ n_8722;
assign n_8872 = n_2677 ^ n_8723;
assign n_8873 = n_2745 ^ n_8724;
assign n_8874 = n_2812 ^ n_8725;
assign n_8875 = n_2880 ^ n_8726;
assign n_8876 = n_2946 ^ n_8727;
assign n_8877 = n_3015 ^ n_8728;
assign n_8878 = n_3081 ^ n_8729;
assign n_8879 = n_3150 ^ n_8730;
assign n_8880 = n_3214 ^ n_8731;
assign n_8881 = n_3279 ^ n_8732;
assign n_8882 = n_3344 ^ n_8733;
assign n_8883 = n_5011 ^ n_8734;
assign n_8884 = n_5074 ^ n_8735;
assign n_8885 = n_5137 ^ n_8736;
assign n_8886 = n_5198 ^ n_8737;
assign n_8887 = n_5262 ^ n_8738;
assign n_8888 = n_5326 ^ n_8739;
assign n_8889 = n_5390 ^ n_8740;
assign n_8890 = n_5454 ^ n_8741;
assign n_8891 = n_5515 ^ n_8742;
assign n_8892 = n_5578 ^ n_8743;
assign n_8893 = n_5641 ^ n_8744;
assign n_8894 = n_5705 ^ n_8745;
assign n_8895 = n_5771 ^ n_8746;
assign n_8896 = n_5833 ^ n_8747;
assign n_8897 = n_5897 ^ n_8748;
assign n_8898 = n_5960 ^ n_8749;
assign n_8899 = n_6024 ^ n_8750;
assign n_8900 = n_6088 ^ n_8751;
assign n_8901 = n_6150 ^ n_8752;
assign n_8902 = n_6212 ^ n_8753;
assign n_8903 = n_8754 ^ x5;
assign n_8904 = n_8755 ^ x8;
assign n_8905 = n_8756 ^ x11;
assign n_8906 = n_8757 ^ x14;
assign n_8907 = n_8758 ^ x17;
assign n_8908 = n_8759 ^ x20;
assign n_8909 = n_8760 ^ x23;
assign n_8910 = n_8761 ^ x26;
assign n_8911 = n_8762 ^ x29;
assign n_8912 = n_8763 ^ x32;
assign n_8913 = n_8764 ^ x35;
assign n_8914 = n_8765 ^ x38;
assign n_8915 = n_8766 ^ x41;
assign n_8916 = n_8767 ^ x44;
assign n_8917 = n_8768 ^ x47;
assign n_8918 = n_8769 ^ x50;
assign n_8919 = n_8770 ^ x53;
assign n_8920 = n_8771 ^ x56;
assign n_8921 = n_8772 ^ x59;
assign n_8922 = n_8773 ^ x62;
assign n_8923 = n_8788 ^ n_8301;
assign n_8924 = n_8790 ^ n_8522;
assign n_8925 = n_8791 ^ n_8524;
assign n_8926 = n_8792 ^ n_8704;
assign n_8927 = n_8792 ^ n_8305;
assign n_8928 = ~n_138 & ~n_8794;
assign n_8929 = n_3467 & ~n_8795;
assign n_8930 = ~n_139 & ~n_8796;
assign n_8931 = n_8798 ^ n_8700;
assign n_8932 = ~n_6602 & ~n_8801;
assign n_8933 = n_8802 ^ n_8561;
assign n_8934 = n_8802 & ~n_8698;
assign n_8935 = n_8804 ^ n_8525;
assign n_8936 = n_8805 ^ n_7960;
assign n_8937 = n_8805 ^ n_7812;
assign n_8938 = n_8806 ^ n_7962;
assign n_8939 = n_8806 ^ n_7814;
assign n_8940 = n_8807 ^ n_7608;
assign n_8941 = n_8807 ^ n_7474;
assign n_8942 = n_8808 ^ n_7966;
assign n_8943 = n_8808 ^ n_7818;
assign n_8944 = n_8810 ^ n_7968;
assign n_8945 = n_8810 ^ n_7820;
assign n_8946 = n_8811 ^ n_7822;
assign n_8947 = n_8811 ^ n_7695;
assign n_8948 = n_8812 ^ n_7480;
assign n_8949 = ~n_8812 & n_8099;
assign n_8950 = n_8813 ^ n_7460;
assign n_8951 = n_8814 ^ n_7700;
assign n_8952 = n_8814 ^ n_7588;
assign n_8953 = n_8816 ^ n_8543;
assign n_8954 = n_8818 ^ n_8544;
assign n_8955 = n_8819 ^ n_8546;
assign n_8956 = n_8820 ^ n_8104;
assign n_8957 = n_8820 ^ n_7976;
assign n_8958 = n_8821 ^ n_8308;
assign n_8959 = n_8821 ^ n_8194;
assign n_8960 = n_8822 ^ n_7988;
assign n_8961 = n_8822 ^ n_7838;
assign n_8962 = n_8823 ^ n_8314;
assign n_8963 = n_8823 ^ n_7510;
assign n_8964 = n_8824 ^ n_7519;
assign n_8965 = n_8825 ^ n_7883;
assign n_8966 = ~n_7973 & n_8826;
assign n_8967 = n_8827 ^ n_8371;
assign n_8968 = ~n_8125 & ~n_8828;
assign n_8969 = n_8791 ^ n_8829;
assign n_8970 = ~n_8798 & n_8830;
assign n_8971 = n_8831 ^ n_8566;
assign n_8972 = n_8831 & n_8702;
assign n_8973 = n_8799 ^ n_8832;
assign n_8974 = n_8655 ^ n_8832;
assign n_8975 = n_8455 & n_8834;
assign n_8976 = n_8836 ^ n_8572;
assign n_8977 = ~x0 & n_8837;
assign n_8978 = n_8838 ^ n_6481;
assign n_8979 = n_8839 ^ x85;
assign n_8980 = n_8840 ^ x1;
assign n_8981 = n_1 & ~n_8841;
assign n_8982 = ~n_8841 & n_171;
assign n_8983 = n_8841 ^ x87;
assign n_8984 = n_655 & n_8842;
assign n_8985 = n_784 & n_8842;
assign n_8986 = ~n_3665 & n_8842;
assign n_8987 = n_854 & n_8842;
assign n_8988 = n_920 & n_8842;
assign n_8989 = n_986 & n_8842;
assign n_8990 = n_1052 & n_8842;
assign n_8991 = n_8842 & n_1117;
assign n_8992 = n_8842 & n_1181;
assign n_8993 = n_8842 & n_1248;
assign n_8994 = n_8842 & n_1314;
assign n_8995 = n_8842 & n_1380;
assign n_8996 = n_8842 & n_1445;
assign n_8997 = n_8842 & n_1510;
assign n_8998 = n_8842 & n_1576;
assign n_8999 = n_8842 & n_1641;
assign n_9000 = n_8842 & n_1706;
assign n_9001 = n_8842 & n_1771;
assign n_9002 = n_8842 & n_1835;
assign n_9003 = n_8842 & n_1899;
assign n_9004 = n_2140 ^ n_8843;
assign n_9005 = n_740 ^ n_8844;
assign n_9006 = n_2211 ^ n_8845;
assign n_9007 = n_2279 ^ n_8846;
assign n_9008 = n_2346 ^ n_8847;
assign n_9009 = n_2413 ^ n_8848;
assign n_9010 = n_2480 ^ n_8849;
assign n_9011 = n_2546 ^ n_8850;
assign n_9012 = n_2611 ^ n_8851;
assign n_9013 = n_2678 ^ n_8852;
assign n_9014 = n_2746 ^ n_8853;
assign n_9015 = n_2813 ^ n_8854;
assign n_9016 = n_2881 ^ n_8855;
assign n_9017 = n_2947 ^ n_8856;
assign n_9018 = n_3016 ^ n_8857;
assign n_9019 = n_3082 ^ n_8858;
assign n_9020 = n_3151 ^ n_8859;
assign n_9021 = n_3215 ^ n_8860;
assign n_9022 = n_3280 ^ n_8861;
assign n_9023 = n_3345 ^ n_8862;
assign n_9024 = n_5012 ^ n_8863;
assign n_9025 = n_5075 ^ n_8864;
assign n_9026 = n_5138 ^ n_8865;
assign n_9027 = n_5199 ^ n_8866;
assign n_9028 = n_5263 ^ n_8867;
assign n_9029 = n_5327 ^ n_8868;
assign n_9030 = n_5391 ^ n_8869;
assign n_9031 = n_5455 ^ n_8870;
assign n_9032 = n_5516 ^ n_8871;
assign n_9033 = n_5579 ^ n_8872;
assign n_9034 = n_5642 ^ n_8873;
assign n_9035 = n_5706 ^ n_8874;
assign n_9036 = n_5772 ^ n_8875;
assign n_9037 = n_5834 ^ n_8876;
assign n_9038 = n_5898 ^ n_8877;
assign n_9039 = n_5961 ^ n_8878;
assign n_9040 = n_6025 ^ n_8879;
assign n_9041 = n_6089 ^ n_8880;
assign n_9042 = n_6151 ^ n_8881;
assign n_9043 = n_6213 ^ n_8882;
assign n_9044 = n_8883 ^ x5;
assign n_9045 = n_8884 ^ x8;
assign n_9046 = n_8885 ^ x11;
assign n_9047 = n_8886 ^ x14;
assign n_9048 = n_8887 ^ x17;
assign n_9049 = n_8888 ^ x20;
assign n_9050 = n_8889 ^ x23;
assign n_9051 = n_8890 ^ x26;
assign n_9052 = n_8891 ^ x29;
assign n_9053 = n_8892 ^ x32;
assign n_9054 = n_8893 ^ x35;
assign n_9055 = n_8894 ^ x38;
assign n_9056 = n_8895 ^ x41;
assign n_9057 = n_8896 ^ x44;
assign n_9058 = n_8897 ^ x47;
assign n_9059 = n_8898 ^ x50;
assign n_9060 = n_8899 ^ x53;
assign n_9061 = n_8900 ^ x56;
assign n_9062 = n_8901 ^ x59;
assign n_9063 = n_6603 ^ n_8902;
assign n_9064 = n_6478 ^ n_8902;
assign n_9065 = n_148 ^ n_8902;
assign n_9066 = n_2038 ^ n_8902;
assign n_9067 = n_8921 ^ n_8833;
assign n_9068 = n_8922 ^ n_6338;
assign n_9069 = n_8924 ^ n_8545;
assign n_9070 = ~n_8924 & n_8682;
assign n_9071 = n_8925 ^ n_8829;
assign n_9072 = ~n_8704 & ~n_8927;
assign n_9073 = n_8928 ^ x77;
assign n_9074 = n_8930 ^ x78;
assign n_9075 = n_8932 ^ n_8656;
assign n_9076 = n_8919 ^ n_8933;
assign n_9077 = n_8934 ^ n_8657;
assign n_9078 = n_8935 ^ n_7984;
assign n_9079 = n_8935 ^ n_7834;
assign n_9080 = n_8936 ^ n_7873;
assign n_9081 = ~n_7960 & n_8937;
assign n_9082 = n_7874 ^ n_8938;
assign n_9083 = ~n_7962 & n_8939;
assign n_9084 = n_8940 ^ n_7875;
assign n_9085 = n_7608 & n_8941;
assign n_9086 = n_7878 ^ n_8942;
assign n_9087 = ~n_7966 & n_8943;
assign n_9088 = n_8944 ^ n_7879;
assign n_9089 = ~n_7968 & n_8945;
assign n_9090 = n_7880 ^ n_8946;
assign n_9091 = ~n_7822 & n_8947;
assign n_9092 = n_8948 ^ n_7881;
assign n_9093 = n_8949 ^ n_8673;
assign n_9094 = n_8950 ^ n_7481;
assign n_9095 = n_8950 & ~n_7610;
assign n_9096 = n_8951 ^ n_7884;
assign n_9097 = ~n_7700 & n_8952;
assign n_9098 = n_8953 ^ n_7990;
assign n_9099 = n_8953 ^ n_7840;
assign n_9100 = n_8954 ^ n_8089;
assign n_9101 = n_8954 ^ n_7956;
assign n_9102 = n_8955 ^ n_7982;
assign n_9103 = n_8955 ^ n_7832;
assign n_9104 = n_8956 ^ n_8124;
assign n_9105 = ~n_8104 & n_8957;
assign n_9106 = n_8958 ^ n_8007;
assign n_9107 = ~n_8308 & n_8959;
assign n_9108 = n_8960 ^ n_8011;
assign n_9109 = ~n_7988 & n_8961;
assign n_9110 = n_8962 ^ n_8012;
assign n_9111 = n_8314 & ~n_8963;
assign n_9112 = n_8964 ^ n_7714;
assign n_9113 = n_8964 & ~n_7843;
assign n_9114 = n_8966 ^ n_8696;
assign n_9115 = n_8968 ^ n_8697;
assign n_9116 = ~n_8925 & ~n_8969;
assign n_9117 = n_8970 ^ n_8700;
assign n_9118 = n_8920 ^ n_8971;
assign n_9119 = n_8972 ^ n_8701;
assign n_9120 = n_8799 & n_8974;
assign n_9121 = n_8975 ^ n_8705;
assign n_9122 = n_8977 ^ n_8709;
assign n_9123 = ~x0 & ~n_8978;
assign n_9124 = n_8979 ^ n_3476;
assign n_9125 = n_8980 ^ x86;
assign n_9126 = n_8981 ^ x1;
assign n_9127 = n_1 & ~n_8982;
assign n_9128 = ~n_8982 & n_175;
assign n_9129 = n_8982 ^ x88;
assign n_9130 = n_655 & n_8983;
assign n_9131 = n_784 & n_8983;
assign n_9132 = ~n_3665 & n_8983;
assign n_9133 = n_854 & n_8983;
assign n_9134 = n_920 & n_8983;
assign n_9135 = n_986 & n_8983;
assign n_9136 = n_1052 & n_8983;
assign n_9137 = n_8983 & n_1117;
assign n_9138 = n_8983 & n_1181;
assign n_9139 = n_8983 & n_1248;
assign n_9140 = n_8983 & n_1314;
assign n_9141 = n_8983 & n_1380;
assign n_9142 = n_8983 & n_1445;
assign n_9143 = n_8983 & n_1510;
assign n_9144 = n_8983 & n_1576;
assign n_9145 = n_8983 & n_1641;
assign n_9146 = n_8983 & n_1706;
assign n_9147 = n_8983 & n_1771;
assign n_9148 = n_8983 & n_1835;
assign n_9149 = n_8983 & n_1899;
assign n_9150 = n_2141 ^ n_8984;
assign n_9151 = n_741 ^ n_8985;
assign n_9152 = n_2212 ^ n_8986;
assign n_9153 = n_2280 ^ n_8987;
assign n_9154 = n_2347 ^ n_8988;
assign n_9155 = n_2414 ^ n_8989;
assign n_9156 = n_2481 ^ n_8990;
assign n_9157 = n_2547 ^ n_8991;
assign n_9158 = n_2612 ^ n_8992;
assign n_9159 = n_2679 ^ n_8993;
assign n_9160 = n_2747 ^ n_8994;
assign n_9161 = n_2814 ^ n_8995;
assign n_9162 = n_2882 ^ n_8996;
assign n_9163 = n_2948 ^ n_8997;
assign n_9164 = n_3017 ^ n_8998;
assign n_9165 = n_3083 ^ n_8999;
assign n_9166 = n_3152 ^ n_9000;
assign n_9167 = n_3216 ^ n_9001;
assign n_9168 = n_3281 ^ n_9002;
assign n_9169 = n_3346 ^ n_9003;
assign n_9170 = n_5013 ^ n_9004;
assign n_9171 = n_5076 ^ n_9005;
assign n_9172 = n_5139 ^ n_9006;
assign n_9173 = n_5200 ^ n_9007;
assign n_9174 = n_5264 ^ n_9008;
assign n_9175 = n_5328 ^ n_9009;
assign n_9176 = n_5392 ^ n_9010;
assign n_9177 = n_5456 ^ n_9011;
assign n_9178 = n_5517 ^ n_9012;
assign n_9179 = n_5580 ^ n_9013;
assign n_9180 = n_5643 ^ n_9014;
assign n_9181 = n_5707 ^ n_9015;
assign n_9182 = n_5773 ^ n_9016;
assign n_9183 = n_5835 ^ n_9017;
assign n_9184 = n_5899 ^ n_9018;
assign n_9185 = n_5962 ^ n_9019;
assign n_9186 = n_6026 ^ n_9020;
assign n_9187 = n_6090 ^ n_9021;
assign n_9188 = n_6152 ^ n_9022;
assign n_9189 = n_6214 ^ n_9023;
assign n_9190 = n_9024 ^ x5;
assign n_9191 = n_9025 ^ x8;
assign n_9192 = n_9026 ^ x11;
assign n_9193 = n_9027 ^ x14;
assign n_9194 = n_9028 ^ x17;
assign n_9195 = n_9029 ^ x20;
assign n_9196 = n_9030 ^ x23;
assign n_9197 = n_9031 ^ x26;
assign n_9198 = n_9032 ^ x29;
assign n_9199 = n_9033 ^ x32;
assign n_9200 = n_9034 ^ x35;
assign n_9201 = n_9035 ^ x38;
assign n_9202 = n_9036 ^ x41;
assign n_9203 = n_9037 ^ x44;
assign n_9204 = n_9038 ^ x47;
assign n_9205 = n_9039 ^ x50;
assign n_9206 = n_9040 ^ x53;
assign n_9207 = n_9041 ^ x56;
assign n_9208 = n_9042 ^ x59;
assign n_9209 = n_6480 ^ n_9043;
assign n_9210 = n_9043 ^ x81;
assign n_9211 = ~n_9043 & n_3474;
assign n_9212 = n_9043 ^ x80;
assign n_9213 = n_9060 ^ n_8931;
assign n_9214 = n_9061 ^ n_8973;
assign n_9215 = n_9062 ^ n_8800;
assign n_9216 = ~n_9064 & ~n_9065;
assign n_9217 = n_9064 & n_9066;
assign n_9218 = n_9070 ^ n_8790;
assign n_9219 = n_9072 ^ n_8568;
assign n_9220 = n_487 & ~n_9073;
assign n_9221 = n_67 & ~n_9074;
assign n_9222 = n_9075 ^ n_8793;
assign n_9223 = n_9060 ^ n_9077;
assign n_9224 = n_9078 ^ n_8006;
assign n_9225 = ~n_7984 & n_9079;
assign n_9226 = n_9081 ^ n_8805;
assign n_9227 = n_9083 ^ n_8806;
assign n_9228 = n_9085 ^ n_8807;
assign n_9229 = n_9087 ^ n_8808;
assign n_9230 = n_9089 ^ n_8810;
assign n_9231 = n_9091 ^ n_8811;
assign n_9232 = n_9093 ^ n_8208;
assign n_9233 = n_7882 ^ n_9094;
assign n_9234 = n_9095 ^ n_8813;
assign n_9235 = n_9097 ^ n_8814;
assign n_9236 = n_9098 ^ n_8020;
assign n_9237 = n_7990 & ~n_9099;
assign n_9238 = n_9100 ^ n_8005;
assign n_9239 = ~n_8089 & n_9101;
assign y9 = n_9102;
assign n_9240 = ~n_7982 & n_9103;
assign n_9241 = n_9105 ^ n_8820;
assign n_9242 = n_9107 ^ n_8821;
assign n_9243 = n_9109 ^ n_8822;
assign n_9244 = n_9111 ^ n_8200;
assign n_9245 = n_9112 ^ n_8021;
assign n_9246 = n_9113 ^ n_8824;
assign n_9247 = n_9114 ^ n_8323;
assign n_9248 = n_9114 ^ n_8210;
assign n_9249 = n_9115 ^ n_8797;
assign n_9250 = n_9115 ^ n_8653;
assign n_9251 = n_9116 ^ n_8524;
assign n_9252 = n_9071 ^ n_9117;
assign n_9253 = n_9061 ^ n_9119;
assign n_9254 = n_9120 ^ n_8832;
assign n_9255 = n_9062 ^ n_9121;
assign n_9256 = n_9123 ^ n_8838;
assign n_9257 = ~x0 & n_9124;
assign n_9258 = n_9125 ^ n_3477;
assign n_9259 = n_9126 ^ x87;
assign n_9260 = n_9127 ^ x1;
assign n_9261 = n_1 & ~n_9128;
assign n_9262 = ~n_9128 & n_179;
assign n_9263 = n_9128 ^ x89;
assign n_9264 = n_655 & n_9129;
assign n_9265 = n_784 & n_9129;
assign n_9266 = ~n_3665 & n_9129;
assign n_9267 = n_854 & n_9129;
assign n_9268 = n_920 & n_9129;
assign n_9269 = n_986 & n_9129;
assign n_9270 = n_1052 & n_9129;
assign n_9271 = n_1117 & n_9129;
assign n_9272 = n_9129 & n_1181;
assign n_9273 = n_9129 & n_1248;
assign n_9274 = n_9129 & n_1314;
assign n_9275 = n_9129 & n_1380;
assign n_9276 = n_9129 & n_1445;
assign n_9277 = n_9129 & n_1510;
assign n_9278 = n_9129 & n_1576;
assign n_9279 = n_9129 & n_1641;
assign n_9280 = n_9129 & n_1706;
assign n_9281 = n_9129 & n_1771;
assign n_9282 = n_9129 & n_1835;
assign n_9283 = n_9129 & n_1899;
assign n_9284 = n_2142 ^ n_9130;
assign n_9285 = n_742 ^ n_9131;
assign n_9286 = n_2213 ^ n_9132;
assign n_9287 = n_2281 ^ n_9133;
assign n_9288 = n_2348 ^ n_9134;
assign n_9289 = n_2415 ^ n_9135;
assign n_9290 = n_2482 ^ n_9136;
assign n_9291 = n_2548 ^ n_9137;
assign n_9292 = n_2613 ^ n_9138;
assign n_9293 = n_2680 ^ n_9139;
assign n_9294 = n_2748 ^ n_9140;
assign n_9295 = n_2815 ^ n_9141;
assign n_9296 = n_2883 ^ n_9142;
assign n_9297 = n_2949 ^ n_9143;
assign n_9298 = n_3018 ^ n_9144;
assign n_9299 = n_3084 ^ n_9145;
assign n_9300 = n_3153 ^ n_9146;
assign n_9301 = n_3217 ^ n_9147;
assign n_9302 = n_3282 ^ n_9148;
assign n_9303 = n_3347 ^ n_9149;
assign n_9304 = n_5014 ^ n_9150;
assign n_9305 = n_5077 ^ n_9151;
assign n_9306 = n_5140 ^ n_9152;
assign n_9307 = n_5201 ^ n_9153;
assign n_9308 = n_5265 ^ n_9154;
assign n_9309 = n_5329 ^ n_9155;
assign n_9310 = n_5393 ^ n_9156;
assign n_9311 = n_5457 ^ n_9157;
assign n_9312 = n_5518 ^ n_9158;
assign n_9313 = n_5581 ^ n_9159;
assign n_9314 = n_5644 ^ n_9160;
assign n_9315 = n_5708 ^ n_9161;
assign n_9316 = n_5774 ^ n_9162;
assign n_9317 = n_5836 ^ n_9163;
assign n_9318 = n_5900 ^ n_9164;
assign n_9319 = n_5963 ^ n_9165;
assign n_9320 = n_6027 ^ n_9166;
assign n_9321 = n_6091 ^ n_9167;
assign n_9322 = n_6153 ^ n_9168;
assign n_9323 = n_6215 ^ n_9169;
assign n_9324 = n_9170 ^ x5;
assign n_9325 = n_9171 ^ x8;
assign n_9326 = n_9172 ^ x11;
assign n_9327 = n_9173 ^ x14;
assign n_9328 = n_9174 ^ x17;
assign n_9329 = n_9175 ^ x20;
assign n_9330 = n_9176 ^ x23;
assign n_9331 = n_9177 ^ x26;
assign n_9332 = n_9178 ^ x29;
assign n_9333 = n_9179 ^ x32;
assign n_9334 = n_9180 ^ x35;
assign n_9335 = n_9181 ^ x38;
assign n_9336 = n_9182 ^ x41;
assign n_9337 = n_9183 ^ x44;
assign n_9338 = n_9184 ^ x47;
assign n_9339 = n_9185 ^ x50;
assign n_9340 = n_9186 ^ x53;
assign n_9341 = n_9187 ^ x56;
assign n_9342 = n_9188 ^ x59;
assign n_9343 = n_9189 ^ x62;
assign n_9344 = n_9205 ^ n_9069;
assign n_9345 = n_9206 ^ n_9071;
assign n_9346 = n_9207 ^ n_8926;
assign n_9347 = n_9075 ^ n_9208;
assign n_9348 = ~n_149 & n_9210;
assign n_9349 = ~n_145 & n_9212;
assign n_9350 = n_9213 ^ n_9077;
assign n_9351 = n_9214 ^ n_9119;
assign n_9352 = n_9215 ^ n_9121;
assign n_9353 = n_9216 ^ n_8902;
assign n_9354 = n_9217 ^ n_8902;
assign n_9355 = n_9218 ^ n_9076;
assign n_9356 = n_9218 ^ n_8919;
assign n_9357 = n_9219 ^ n_9067;
assign n_9358 = n_9219 ^ n_8833;
assign n_9359 = n_9220 ^ n_8929;
assign n_9360 = n_9222 ^ n_9208;
assign n_9361 = ~n_9213 & n_9223;
assign n_9362 = n_9225 ^ n_8935;
assign n_9363 = n_9226 ^ n_8310;
assign n_9364 = n_9226 ^ n_8196;
assign n_9365 = n_9227 ^ n_8312;
assign n_9366 = n_9227 ^ n_8198;
assign n_9367 = n_9228 ^ n_7986;
assign n_9368 = n_9228 ^ n_7836;
assign n_9369 = n_9229 ^ n_8316;
assign n_9370 = n_9229 ^ n_8202;
assign n_9371 = n_9230 ^ n_8318;
assign n_9372 = n_9230 ^ n_8204;
assign n_9373 = n_9231 ^ n_7513;
assign n_9374 = n_9232 ^ n_7514;
assign n_9375 = ~n_9232 & n_8321;
assign n_9376 = n_9234 ^ n_8342;
assign n_9377 = n_9234 ^ n_8226;
assign n_9378 = n_9235 ^ n_7517;
assign n_9379 = n_9237 ^ n_8953;
assign n_9380 = n_9239 ^ n_8954;
assign n_9381 = n_9240 ^ n_8955;
assign n_9382 = n_9241 ^ n_8435;
assign n_9383 = n_9241 ^ n_8327;
assign n_9384 = n_9242 ^ n_8660;
assign n_9385 = n_9242 ^ n_8526;
assign n_9386 = n_9243 ^ n_8338;
assign n_9387 = n_9243 ^ n_8222;
assign n_9388 = n_9244 ^ n_8666;
assign n_9389 = n_9244 ^ n_8532;
assign n_9390 = n_9246 ^ n_8228;
assign n_9391 = n_9246 ^ n_8116;
assign n_9392 = n_9247 ^ n_8018;
assign n_9393 = ~n_8323 & n_9248;
assign n_9394 = n_9059 ^ n_9249;
assign n_9395 = ~n_8797 & ~n_9250;
assign n_9396 = n_9251 ^ n_9118;
assign n_9397 = n_9251 ^ n_8920;
assign n_9398 = n_9214 & n_9253;
assign n_9399 = n_8926 ^ n_9254;
assign n_9400 = ~n_9215 & n_9255;
assign n_9401 = n_9257 ^ n_8979;
assign n_9402 = ~x0 & n_9258;
assign n_9403 = n_9259 ^ n_3479;
assign n_9404 = n_9260 ^ x88;
assign n_9405 = n_9261 ^ x1;
assign n_9406 = n_1 & ~n_9262;
assign n_9407 = ~n_9262 & n_182;
assign n_9408 = n_9262 ^ x90;
assign n_9409 = n_655 & n_9263;
assign n_9410 = n_784 & n_9263;
assign n_9411 = ~n_3665 & n_9263;
assign n_9412 = n_854 & n_9263;
assign n_9413 = n_920 & n_9263;
assign n_9414 = n_986 & n_9263;
assign n_9415 = n_1052 & n_9263;
assign n_9416 = n_1117 & n_9263;
assign n_9417 = n_9263 & n_1181;
assign n_9418 = n_9263 & n_1248;
assign n_9419 = n_9263 & n_1314;
assign n_9420 = n_9263 & n_1380;
assign n_9421 = n_9263 & n_1445;
assign n_9422 = n_9263 & n_1510;
assign n_9423 = n_9263 & n_1576;
assign n_9424 = n_9263 & n_1641;
assign n_9425 = n_9263 & n_1706;
assign n_9426 = n_9263 & n_1771;
assign n_9427 = n_9263 & n_1835;
assign n_9428 = n_9263 & n_1899;
assign n_9429 = n_2143 ^ n_9264;
assign n_9430 = n_743 ^ n_9265;
assign n_9431 = n_2214 ^ n_9266;
assign n_9432 = n_2282 ^ n_9267;
assign n_9433 = n_2349 ^ n_9268;
assign n_9434 = n_2416 ^ n_9269;
assign n_9435 = n_2483 ^ n_9270;
assign n_9436 = n_2549 ^ n_9271;
assign n_9437 = n_2614 ^ n_9272;
assign n_9438 = n_2681 ^ n_9273;
assign n_9439 = n_2749 ^ n_9274;
assign n_9440 = n_2816 ^ n_9275;
assign n_9441 = n_2884 ^ n_9276;
assign n_9442 = n_2950 ^ n_9277;
assign n_9443 = n_3019 ^ n_9278;
assign n_9444 = n_3085 ^ n_9279;
assign n_9445 = n_3154 ^ n_9280;
assign n_9446 = n_3218 ^ n_9281;
assign n_9447 = n_3283 ^ n_9282;
assign n_9448 = n_3348 ^ n_9283;
assign n_9449 = n_5015 ^ n_9284;
assign n_9450 = n_5078 ^ n_9285;
assign n_9451 = n_5141 ^ n_9286;
assign n_9452 = n_5202 ^ n_9287;
assign n_9453 = n_5266 ^ n_9288;
assign n_9454 = n_5330 ^ n_9289;
assign n_9455 = n_5394 ^ n_9290;
assign n_9456 = n_5458 ^ n_9291;
assign n_9457 = n_5519 ^ n_9292;
assign n_9458 = n_5582 ^ n_9293;
assign n_9459 = n_5645 ^ n_9294;
assign n_9460 = n_5709 ^ n_9295;
assign n_9461 = n_5775 ^ n_9296;
assign n_9462 = n_5837 ^ n_9297;
assign n_9463 = n_5901 ^ n_9298;
assign n_9464 = n_5964 ^ n_9299;
assign n_9465 = n_6028 ^ n_9300;
assign n_9466 = n_6092 ^ n_9301;
assign n_9467 = n_6154 ^ n_9302;
assign n_9468 = n_6216 ^ n_9303;
assign n_9469 = n_9304 ^ x5;
assign n_9470 = n_9305 ^ x8;
assign n_9471 = n_9306 ^ x11;
assign n_9472 = n_9307 ^ x14;
assign n_9473 = n_9308 ^ x17;
assign n_9474 = n_9309 ^ x20;
assign n_9475 = n_9310 ^ x23;
assign n_9476 = n_9311 ^ x26;
assign n_9477 = n_9312 ^ x29;
assign n_9478 = n_9313 ^ x32;
assign n_9479 = n_9314 ^ x35;
assign n_9480 = n_9315 ^ x38;
assign n_9481 = n_9316 ^ x41;
assign n_9482 = n_9317 ^ x44;
assign n_9483 = n_9318 ^ x47;
assign n_9484 = n_9319 ^ x50;
assign n_9485 = n_9320 ^ x53;
assign n_9486 = n_9321 ^ x56;
assign n_9487 = n_9322 ^ x59;
assign n_9488 = n_9323 ^ x62;
assign n_9489 = n_9343 ^ n_6397;
assign n_9490 = n_9345 ^ n_9117;
assign n_9491 = ~n_9345 & n_9252;
assign n_9492 = n_9346 ^ n_9254;
assign n_9493 = n_9222 & n_9347;
assign n_9494 = n_9348 ^ x81;
assign n_9495 = n_9349 ^ x80;
assign n_9496 = n_9353 ^ n_9354;
assign n_9497 = n_9355 ^ n_9339;
assign n_9498 = n_9076 & ~n_9356;
assign n_9499 = n_9357 ^ n_9341;
assign n_9500 = n_9067 & n_9358;
assign n_9501 = n_9359 ^ n_9221;
assign n_9502 = n_9361 ^ n_9077;
assign n_9503 = n_9362 ^ n_8334;
assign n_9504 = n_9362 ^ n_8219;
assign n_9505 = n_9363 ^ n_8008;
assign n_9506 = ~n_8310 & n_9364;
assign n_9507 = n_9365 ^ n_8009;
assign n_9508 = n_8312 & ~n_9366;
assign n_9509 = n_9367 ^ n_8010;
assign n_9510 = ~n_7986 & n_9368;
assign n_9511 = n_9369 ^ n_8013;
assign n_9512 = ~n_8316 & n_9370;
assign n_9513 = n_9371 ^ n_8014;
assign n_9514 = n_8318 & ~n_9372;
assign n_9515 = n_9373 ^ n_8097;
assign n_9516 = n_9373 & ~n_8206;
assign n_9517 = n_9374 ^ n_8016;
assign n_9518 = n_9375 ^ n_9093;
assign n_9519 = n_9376 ^ n_8017;
assign n_9520 = ~n_8342 & n_9377;
assign n_9521 = n_9378 ^ n_8102;
assign n_9522 = n_9378 & n_8212;
assign n_9523 = n_9379 ^ n_8340;
assign n_9524 = n_9379 ^ n_8224;
assign n_9525 = n_9380 ^ n_8422;
assign n_9526 = n_9380 ^ n_8306;
assign n_9527 = n_9381 ^ n_8332;
assign n_9528 = n_9381 ^ n_8217;
assign n_9529 = n_9382 ^ n_8235;
assign n_9530 = ~n_8435 & n_9383;
assign n_9531 = n_9384 ^ n_8130;
assign n_9532 = ~n_8660 & n_9385;
assign n_9533 = n_9386 ^ n_8134;
assign n_9534 = ~n_8338 & n_9387;
assign n_9535 = n_9388 ^ n_8135;
assign n_9536 = ~n_8666 & n_9389;
assign n_9537 = n_8144 ^ n_9390;
assign n_9538 = ~n_8228 & n_9391;
assign n_9539 = n_9393 ^ n_9114;
assign n_9540 = n_9395 ^ n_9115;
assign n_9541 = n_9396 ^ n_9340;
assign n_9542 = ~n_9118 & n_9397;
assign n_9543 = n_9398 ^ n_9119;
assign n_9544 = ~n_9346 & n_9399;
assign n_9545 = n_9400 ^ n_9121;
assign n_9546 = n_9402 ^ n_9125;
assign n_9547 = ~x0 & n_9403;
assign n_9548 = n_9404 ^ n_3480;
assign n_9549 = n_9405 ^ x89;
assign n_9550 = n_9406 ^ x1;
assign n_9551 = n_1 & ~n_9407;
assign n_9552 = ~n_9407 & n_185;
assign n_9553 = n_9407 ^ x91;
assign n_9554 = n_655 & n_9408;
assign n_9555 = n_784 & n_9408;
assign n_9556 = ~n_3665 & n_9408;
assign n_9557 = n_854 & n_9408;
assign n_9558 = n_920 & n_9408;
assign n_9559 = n_986 & n_9408;
assign n_9560 = n_1052 & n_9408;
assign n_9561 = n_1117 & n_9408;
assign n_9562 = n_9408 & n_1181;
assign n_9563 = n_9408 & n_1248;
assign n_9564 = n_9408 & n_1314;
assign n_9565 = n_9408 & n_1380;
assign n_9566 = n_9408 & n_1445;
assign n_9567 = n_9408 & n_1510;
assign n_9568 = n_9408 & n_1576;
assign n_9569 = n_9408 & n_1641;
assign n_9570 = n_9408 & n_1706;
assign n_9571 = n_9408 & n_1771;
assign n_9572 = n_9408 & n_1835;
assign n_9573 = n_9408 & n_1899;
assign n_9574 = n_2144 ^ n_9409;
assign n_9575 = n_744 ^ n_9410;
assign n_9576 = n_2215 ^ n_9411;
assign n_9577 = n_2283 ^ n_9412;
assign n_9578 = n_2350 ^ n_9413;
assign n_9579 = n_2417 ^ n_9414;
assign n_9580 = n_2484 ^ n_9415;
assign n_9581 = n_2550 ^ n_9416;
assign n_9582 = n_2615 ^ n_9417;
assign n_9583 = n_2682 ^ n_9418;
assign n_9584 = n_2750 ^ n_9419;
assign n_9585 = n_2817 ^ n_9420;
assign n_9586 = n_2885 ^ n_9421;
assign n_9587 = n_2951 ^ n_9422;
assign n_9588 = n_3020 ^ n_9423;
assign n_9589 = n_3086 ^ n_9424;
assign n_9590 = n_3155 ^ n_9425;
assign n_9591 = n_3219 ^ n_9426;
assign n_9592 = n_3284 ^ n_9427;
assign n_9593 = n_3349 ^ n_9428;
assign n_9594 = n_5016 ^ n_9429;
assign n_9595 = n_5079 ^ n_9430;
assign n_9596 = n_5142 ^ n_9431;
assign n_9597 = n_5203 ^ n_9432;
assign n_9598 = n_5267 ^ n_9433;
assign n_9599 = n_5331 ^ n_9434;
assign n_9600 = n_5395 ^ n_9435;
assign n_9601 = n_5459 ^ n_9436;
assign n_9602 = n_5520 ^ n_9437;
assign n_9603 = n_5583 ^ n_9438;
assign n_9604 = n_5646 ^ n_9439;
assign n_9605 = n_5710 ^ n_9440;
assign n_9606 = n_5776 ^ n_9441;
assign n_9607 = n_5838 ^ n_9442;
assign n_9608 = n_5902 ^ n_9443;
assign n_9609 = n_5965 ^ n_9444;
assign n_9610 = n_6029 ^ n_9445;
assign n_9611 = n_6093 ^ n_9446;
assign n_9612 = n_6155 ^ n_9447;
assign n_9613 = n_6217 ^ n_9448;
assign n_9614 = n_9449 ^ x5;
assign n_9615 = n_9450 ^ x8;
assign n_9616 = n_9451 ^ x11;
assign n_9617 = n_9452 ^ x14;
assign n_9618 = n_9453 ^ x17;
assign n_9619 = n_9454 ^ x20;
assign n_9620 = n_9455 ^ x23;
assign n_9621 = n_9456 ^ x26;
assign n_9622 = n_9457 ^ x29;
assign n_9623 = n_9458 ^ x32;
assign n_9624 = n_9459 ^ x35;
assign n_9625 = n_9460 ^ x38;
assign n_9626 = n_9461 ^ x41;
assign n_9627 = n_9462 ^ x44;
assign n_9628 = n_9463 ^ x47;
assign n_9629 = n_9464 ^ x50;
assign n_9630 = n_9465 ^ x53;
assign n_9631 = n_9466 ^ x56;
assign n_9632 = n_9467 ^ x59;
assign n_9633 = n_9468 ^ x62;
assign n_9634 = n_9484 ^ n_9350;
assign n_9635 = n_9485 ^ n_9351;
assign n_9636 = n_9486 ^ n_9352;
assign n_9637 = n_9487 ^ n_9063;
assign n_9638 = n_9488 ^ n_6636;
assign n_9639 = n_9488 ^ n_6524;
assign n_9640 = n_9491 ^ n_9206;
assign n_9641 = n_9493 ^ n_9208;
assign n_9642 = n_67 & n_9494;
assign n_9643 = n_9495 ^ n_151;
assign n_9644 = x62 & ~n_9496;
assign n_9645 = n_9498 ^ n_8933;
assign n_9646 = n_9500 ^ n_9219;
assign n_9647 = n_9501 ^ n_9068;
assign n_9648 = n_9501 ^ n_8922;
assign n_9649 = n_9490 ^ n_9502;
assign n_9650 = n_9503 ^ n_8129;
assign n_9651 = ~n_8334 & n_9504;
assign n_9652 = n_9506 ^ n_9226;
assign n_9653 = n_9508 ^ n_9227;
assign n_9654 = n_9510 ^ n_9228;
assign n_9655 = n_9512 ^ n_9229;
assign n_9656 = n_9514 ^ n_9230;
assign n_9657 = n_9515 ^ n_8015;
assign n_9658 = n_9516 ^ n_9231;
assign n_9659 = n_9518 ^ n_8674;
assign n_9660 = n_9518 ^ n_8539;
assign n_9661 = n_9520 ^ n_9234;
assign n_9662 = n_9521 ^ n_8019;
assign n_9663 = n_9522 ^ n_9235;
assign n_9664 = n_8143 ^ n_9523;
assign n_9665 = ~n_8340 & n_9524;
assign n_9666 = n_9525 ^ n_8128;
assign n_9667 = ~n_8422 & n_9526;
assign y10 = n_9527;
assign n_9668 = ~n_8332 & n_9528;
assign n_9669 = n_9530 ^ n_9241;
assign n_9670 = n_9532 ^ n_9242;
assign n_9671 = n_9534 ^ n_9243;
assign n_9672 = n_9536 ^ n_9244;
assign n_9673 = n_9538 ^ n_9246;
assign n_9674 = n_9539 ^ n_8676;
assign n_9675 = n_9539 ^ n_8541;
assign n_9676 = n_9540 ^ n_9344;
assign n_9677 = n_9540 ^ n_9205;
assign n_9678 = n_9542 ^ n_8971;
assign n_9679 = n_9492 ^ n_9543;
assign n_9680 = n_9544 ^ n_9207;
assign n_9681 = n_9360 ^ n_9545;
assign n_9682 = n_9547 ^ n_9259;
assign n_9683 = ~x0 & n_9548;
assign n_9684 = n_9549 ^ n_3481;
assign n_9685 = n_9550 ^ x90;
assign n_9686 = n_9551 ^ x1;
assign n_9687 = n_1 & ~n_9552;
assign n_9688 = ~n_9552 & n_189;
assign n_9689 = ~n_9552 & ~n_194;
assign n_9690 = n_9552 ^ x92;
assign n_9691 = n_655 & n_9553;
assign n_9692 = n_784 & n_9553;
assign n_9693 = ~n_3665 & n_9553;
assign n_9694 = n_854 & n_9553;
assign n_9695 = n_920 & n_9553;
assign n_9696 = n_986 & n_9553;
assign n_9697 = n_1052 & n_9553;
assign n_9698 = n_1117 & n_9553;
assign n_9699 = n_1181 & n_9553;
assign n_9700 = n_9553 & n_1248;
assign n_9701 = n_9553 & n_1314;
assign n_9702 = n_9553 & n_1380;
assign n_9703 = n_9553 & n_1445;
assign n_9704 = n_9553 & n_1510;
assign n_9705 = n_9553 & n_1576;
assign n_9706 = n_9553 & n_1641;
assign n_9707 = n_9553 & n_1706;
assign n_9708 = n_9553 & n_1771;
assign n_9709 = n_9553 & n_1835;
assign n_9710 = n_9553 & n_1899;
assign n_9711 = n_2145 ^ n_9554;
assign n_9712 = n_745 ^ n_9555;
assign n_9713 = n_2216 ^ n_9556;
assign n_9714 = n_2284 ^ n_9557;
assign n_9715 = n_2351 ^ n_9558;
assign n_9716 = n_2418 ^ n_9559;
assign n_9717 = n_2485 ^ n_9560;
assign n_9718 = n_2551 ^ n_9561;
assign n_9719 = n_2616 ^ n_9562;
assign n_9720 = n_2683 ^ n_9563;
assign n_9721 = n_2751 ^ n_9564;
assign n_9722 = n_2818 ^ n_9565;
assign n_9723 = n_2886 ^ n_9566;
assign n_9724 = n_2952 ^ n_9567;
assign n_9725 = n_3021 ^ n_9568;
assign n_9726 = n_3087 ^ n_9569;
assign n_9727 = n_3156 ^ n_9570;
assign n_9728 = n_3220 ^ n_9571;
assign n_9729 = n_3285 ^ n_9572;
assign n_9730 = n_3350 ^ n_9573;
assign n_9731 = n_5017 ^ n_9574;
assign n_9732 = n_5080 ^ n_9575;
assign n_9733 = n_5143 ^ n_9576;
assign n_9734 = n_5204 ^ n_9577;
assign n_9735 = n_5268 ^ n_9578;
assign n_9736 = n_5332 ^ n_9579;
assign n_9737 = n_5396 ^ n_9580;
assign n_9738 = n_5460 ^ n_9581;
assign n_9739 = n_5521 ^ n_9582;
assign n_9740 = n_5584 ^ n_9583;
assign n_9741 = n_5647 ^ n_9584;
assign n_9742 = n_5711 ^ n_9585;
assign n_9743 = n_5777 ^ n_9586;
assign n_9744 = n_5839 ^ n_9587;
assign n_9745 = n_5903 ^ n_9588;
assign n_9746 = n_5966 ^ n_9589;
assign n_9747 = n_6030 ^ n_9590;
assign n_9748 = n_6094 ^ n_9591;
assign n_9749 = n_6156 ^ n_9592;
assign n_9750 = n_6218 ^ n_9593;
assign n_9751 = n_9594 ^ x5;
assign n_9752 = n_9595 ^ x8;
assign n_9753 = n_9596 ^ x11;
assign n_9754 = n_9597 ^ x14;
assign n_9755 = n_9598 ^ x17;
assign n_9756 = n_9599 ^ x20;
assign n_9757 = n_9600 ^ x23;
assign n_9758 = n_9601 ^ x26;
assign n_9759 = n_9602 ^ x29;
assign n_9760 = n_9603 ^ x32;
assign n_9761 = n_9604 ^ x35;
assign n_9762 = n_9605 ^ x38;
assign n_9763 = n_9606 ^ x41;
assign n_9764 = n_9607 ^ x44;
assign n_9765 = n_9608 ^ x47;
assign n_9766 = n_9609 ^ x50;
assign n_9767 = n_9610 ^ x53;
assign n_9768 = n_9611 ^ x56;
assign n_9769 = n_9612 ^ x59;
assign n_9770 = n_9613 ^ x62;
assign n_9771 = n_9629 ^ n_9490;
assign n_9772 = n_9630 ^ n_9492;
assign n_9773 = n_9631 ^ n_9360;
assign n_9774 = n_9633 ^ ~n_6525;
assign n_9775 = ~n_6525 & n_9633;
assign n_9776 = n_6636 & n_9639;
assign n_9777 = n_9640 ^ n_9541;
assign n_9778 = n_9640 ^ n_9396;
assign n_9779 = n_9342 ^ n_9641;
assign n_9780 = n_9642 ^ n_9211;
assign n_9781 = x62 & n_9643;
assign n_9782 = n_9644 ^ n_9353;
assign n_9783 = n_9645 ^ n_9634;
assign n_9784 = n_9645 ^ n_9484;
assign n_9785 = n_9646 ^ n_9486;
assign n_9786 = n_9647 ^ n_9342;
assign n_9787 = n_9068 & ~n_9648;
assign n_9788 = n_9651 ^ n_9362;
assign n_9789 = n_9652 ^ n_8662;
assign n_9790 = n_9652 ^ n_8528;
assign n_9791 = n_9653 ^ n_8664;
assign n_9792 = n_9653 ^ n_8530;
assign n_9793 = n_9654 ^ n_8441;
assign n_9794 = n_9654 ^ n_8336;
assign n_9795 = n_9655 ^ n_8809;
assign n_9796 = n_9655 ^ n_8668;
assign n_9797 = n_9656 ^ n_8670;
assign n_9798 = n_9656 ^ n_8535;
assign n_9799 = n_9658 ^ n_8672;
assign n_9800 = n_9658 ^ n_8537;
assign n_9801 = n_9659 ^ n_8139;
assign n_9802 = ~n_8674 & n_9660;
assign n_9803 = n_9661 ^ n_8695;
assign n_9804 = n_9661 ^ n_8557;
assign n_9805 = n_9663 ^ n_8433;
assign n_9806 = n_9663 ^ n_8325;
assign n_9807 = n_9665 ^ n_9379;
assign n_9808 = n_9667 ^ n_9380;
assign n_9809 = n_9668 ^ n_9381;
assign n_9810 = n_9669 ^ n_8817;
assign n_9811 = n_9669 ^ n_8680;
assign n_9812 = n_9670 ^ n_9080;
assign n_9813 = n_9670 ^ n_8936;
assign n_9814 = n_9671 ^ n_8691;
assign n_9815 = n_9671 ^ n_8553;
assign n_9816 = n_9672 ^ n_7878;
assign n_9817 = n_9673 ^ n_7887;
assign n_9818 = n_8141 ^ n_9674;
assign n_9819 = ~n_8676 & n_9675;
assign n_9820 = n_9676 ^ n_9628;
assign n_9821 = n_9344 & ~n_9677;
assign n_9822 = n_9678 ^ n_9485;
assign n_9823 = n_9680 ^ n_9499;
assign n_9824 = n_9680 ^ n_9357;
assign n_9825 = n_9683 ^ n_9404;
assign n_9826 = ~x0 & n_9684;
assign n_9827 = n_9685 ^ n_3482;
assign n_9828 = n_9686 ^ x91;
assign n_9829 = n_9687 ^ x1;
assign n_9830 = n_1 & ~n_9688;
assign n_9831 = n_9688 ^ x93;
assign n_9832 = n_193 & n_9689;
assign n_9833 = n_655 & n_9690;
assign n_9834 = n_784 & n_9690;
assign n_9835 = ~n_3665 & n_9690;
assign n_9836 = n_854 & n_9690;
assign n_9837 = n_920 & n_9690;
assign n_9838 = n_986 & n_9690;
assign n_9839 = n_1052 & n_9690;
assign n_9840 = n_1117 & n_9690;
assign n_9841 = n_1181 & n_9690;
assign n_9842 = n_9690 & n_1248;
assign n_9843 = n_9690 & n_1314;
assign n_9844 = n_9690 & n_1380;
assign n_9845 = n_9690 & n_1445;
assign n_9846 = n_9690 & n_1510;
assign n_9847 = n_9690 & n_1576;
assign n_9848 = n_9690 & n_1641;
assign n_9849 = n_9690 & n_1706;
assign n_9850 = n_9690 & n_1771;
assign n_9851 = n_9690 & n_1835;
assign n_9852 = n_9690 & n_1899;
assign n_9853 = n_2146 ^ n_9691;
assign n_9854 = n_746 ^ n_9692;
assign n_9855 = n_2217 ^ n_9693;
assign n_9856 = n_2285 ^ n_9694;
assign n_9857 = n_2352 ^ n_9695;
assign n_9858 = n_2419 ^ n_9696;
assign n_9859 = n_2486 ^ n_9697;
assign n_9860 = n_2552 ^ n_9698;
assign n_9861 = n_2617 ^ n_9699;
assign n_9862 = n_2684 ^ n_9700;
assign n_9863 = n_2752 ^ n_9701;
assign n_9864 = n_2819 ^ n_9702;
assign n_9865 = n_2887 ^ n_9703;
assign n_9866 = n_2953 ^ n_9704;
assign n_9867 = n_3022 ^ n_9705;
assign n_9868 = n_3088 ^ n_9706;
assign n_9869 = n_3157 ^ n_9707;
assign n_9870 = n_3221 ^ n_9708;
assign n_9871 = n_3286 ^ n_9709;
assign n_9872 = n_3351 ^ n_9710;
assign n_9873 = n_5018 ^ n_9711;
assign n_9874 = n_5081 ^ n_9712;
assign n_9875 = n_5144 ^ n_9713;
assign n_9876 = n_5205 ^ n_9714;
assign n_9877 = n_5269 ^ n_9715;
assign n_9878 = n_5333 ^ n_9716;
assign n_9879 = n_5397 ^ n_9717;
assign n_9880 = n_5461 ^ n_9718;
assign n_9881 = n_5522 ^ n_9719;
assign n_9882 = n_5585 ^ n_9720;
assign n_9883 = n_5648 ^ n_9721;
assign n_9884 = n_5712 ^ n_9722;
assign n_9885 = n_5778 ^ n_9723;
assign n_9886 = n_5840 ^ n_9724;
assign n_9887 = n_5904 ^ n_9725;
assign n_9888 = n_5967 ^ n_9726;
assign n_9889 = n_6031 ^ n_9727;
assign n_9890 = n_6095 ^ n_9728;
assign n_9891 = n_6157 ^ n_9729;
assign n_9892 = n_6219 ^ n_9730;
assign n_9893 = n_9731 ^ x5;
assign n_9894 = n_9732 ^ x8;
assign n_9895 = n_9733 ^ x11;
assign n_9896 = n_9734 ^ x14;
assign n_9897 = n_9735 ^ x17;
assign n_9898 = n_9736 ^ x20;
assign n_9899 = n_9737 ^ x23;
assign n_9900 = n_9738 ^ x26;
assign n_9901 = n_9739 ^ x29;
assign n_9902 = n_9740 ^ x32;
assign n_9903 = n_9741 ^ x35;
assign n_9904 = n_9742 ^ x38;
assign n_9905 = n_9743 ^ x41;
assign n_9906 = n_9744 ^ x44;
assign n_9907 = n_9745 ^ x47;
assign n_9908 = n_9746 ^ x50;
assign n_9909 = n_9747 ^ x53;
assign n_9910 = n_9748 ^ x56;
assign n_9911 = n_9749 ^ x59;
assign n_9912 = n_9750 ^ x62;
assign n_9913 = n_9770 ^ n_6400;
assign n_9914 = n_9771 ^ n_9502;
assign n_9915 = ~n_9771 & n_9649;
assign n_9916 = n_9772 ^ n_9543;
assign n_9917 = ~n_9772 & n_9679;
assign n_9918 = n_9773 ^ n_9545;
assign n_9919 = ~n_9773 & n_9681;
assign n_9920 = n_9775 ^ n_6263;
assign n_9921 = n_9776 ^ n_9488;
assign n_9922 = n_9777 ^ n_9766;
assign n_9923 = ~n_9541 & n_9778;
assign n_9924 = n_9781 ^ n_151;
assign n_9925 = n_9782 ^ n_9209;
assign n_9926 = n_9782 ^ n_9632;
assign n_9927 = ~n_9634 & n_9784;
assign n_9928 = n_9785 ^ n_9352;
assign n_9929 = ~n_9785 & ~n_9636;
assign n_9930 = n_9786 ^ n_9641;
assign n_9931 = ~n_9786 & n_9779;
assign n_9932 = n_9787 ^ n_9501;
assign n_9933 = n_9788 ^ n_8687;
assign n_9934 = n_9788 ^ n_8549;
assign n_9935 = n_9789 ^ n_8131;
assign n_9936 = ~n_8662 & n_9790;
assign n_9937 = n_9791 ^ n_8132;
assign n_9938 = ~n_8664 & n_9792;
assign n_9939 = n_9793 ^ n_8133;
assign n_9940 = ~n_8441 & n_9794;
assign n_9941 = n_9795 ^ n_8136;
assign n_9942 = ~n_8809 & n_9796;
assign n_9943 = n_9797 ^ n_8137;
assign n_9944 = ~n_8670 & n_9798;
assign n_9945 = n_8138 ^ n_9799;
assign n_9946 = ~n_8672 & n_9800;
assign n_9947 = n_9802 ^ n_9518;
assign n_9948 = n_8140 ^ n_9803;
assign n_9949 = ~n_8695 & n_9804;
assign n_9950 = n_9805 ^ n_8142;
assign n_9951 = ~n_8433 & n_9806;
assign n_9952 = n_9807 ^ n_7886;
assign n_9953 = n_9808 ^ n_8803;
assign n_9954 = n_9808 ^ n_8658;
assign n_9955 = n_9809 ^ n_8685;
assign n_9956 = n_9809 ^ n_8547;
assign n_9957 = n_9810 ^ n_8353;
assign n_9958 = ~n_8817 & n_9811;
assign n_9959 = n_9812 ^ n_8288;
assign n_9960 = ~n_9080 & n_9813;
assign n_9961 = n_9814 ^ n_8292;
assign n_9962 = ~n_8691 & n_9815;
assign n_9963 = n_9816 ^ n_8942;
assign n_9964 = n_9816 & ~n_9086;
assign n_9965 = n_9817 ^ n_8446;
assign n_9966 = n_9817 & ~n_8559;
assign n_9967 = n_9819 ^ n_9539;
assign n_9968 = n_9821 ^ n_9540;
assign n_9969 = n_9822 ^ n_9351;
assign n_9970 = ~n_9822 & n_9635;
assign n_9971 = n_9823 ^ n_9767;
assign n_9972 = ~n_9499 & n_9824;
assign n_9973 = n_9826 ^ n_9549;
assign n_9974 = ~x0 & n_9827;
assign n_9975 = n_9828 ^ n_3483;
assign n_9976 = n_9829 ^ x92;
assign n_9977 = n_9830 ^ x1;
assign n_9978 = n_655 & n_9831;
assign n_9979 = n_784 & n_9831;
assign n_9980 = ~n_3665 & n_9831;
assign n_9981 = n_854 & n_9831;
assign n_9982 = n_920 & n_9831;
assign n_9983 = n_986 & n_9831;
assign n_9984 = n_1052 & n_9831;
assign n_9985 = n_1117 & n_9831;
assign n_9986 = n_1181 & n_9831;
assign n_9987 = n_9831 & n_1248;
assign n_9988 = n_9831 & n_1314;
assign n_9989 = n_9831 & n_1380;
assign n_9990 = n_9831 & n_1445;
assign n_9991 = n_9831 & n_1510;
assign n_9992 = n_9831 & n_1576;
assign n_9993 = n_9831 & n_1641;
assign n_9994 = n_9831 & n_1706;
assign n_9995 = n_9831 & n_1771;
assign n_9996 = n_9831 & n_1835;
assign n_9997 = n_9831 & n_1899;
assign n_9998 = n_9832 ^ n_193;
assign n_9999 = n_2147 ^ n_9833;
assign n_10000 = n_747 ^ n_9834;
assign n_10001 = n_2218 ^ n_9835;
assign n_10002 = n_2286 ^ n_9836;
assign n_10003 = n_2353 ^ n_9837;
assign n_10004 = n_2420 ^ n_9838;
assign n_10005 = n_2487 ^ n_9839;
assign n_10006 = n_2553 ^ n_9840;
assign n_10007 = n_2618 ^ n_9841;
assign n_10008 = n_2685 ^ n_9842;
assign n_10009 = n_2753 ^ n_9843;
assign n_10010 = n_2820 ^ n_9844;
assign n_10011 = n_2888 ^ n_9845;
assign n_10012 = n_2954 ^ n_9846;
assign n_10013 = n_3023 ^ n_9847;
assign n_10014 = n_3089 ^ n_9848;
assign n_10015 = n_3158 ^ n_9849;
assign n_10016 = n_3222 ^ n_9850;
assign n_10017 = n_3287 ^ n_9851;
assign n_10018 = n_3352 ^ n_9852;
assign n_10019 = n_5019 ^ n_9853;
assign n_10020 = n_5082 ^ n_9854;
assign n_10021 = n_5145 ^ n_9855;
assign n_10022 = n_5206 ^ n_9856;
assign n_10023 = n_5270 ^ n_9857;
assign n_10024 = n_5334 ^ n_9858;
assign n_10025 = n_5398 ^ n_9859;
assign n_10026 = n_5462 ^ n_9860;
assign n_10027 = n_5523 ^ n_9861;
assign n_10028 = n_5586 ^ n_9862;
assign n_10029 = n_5649 ^ n_9863;
assign n_10030 = n_5713 ^ n_9864;
assign n_10031 = n_5779 ^ n_9865;
assign n_10032 = n_5841 ^ n_9866;
assign n_10033 = n_5905 ^ n_9867;
assign n_10034 = n_5968 ^ n_9868;
assign n_10035 = n_6032 ^ n_9869;
assign n_10036 = n_6096 ^ n_9870;
assign n_10037 = n_6158 ^ n_9871;
assign n_10038 = n_6220 ^ n_9872;
assign n_10039 = n_9873 ^ x5;
assign n_10040 = n_9874 ^ x8;
assign n_10041 = n_9875 ^ x11;
assign n_10042 = n_9876 ^ x14;
assign n_10043 = n_9877 ^ x17;
assign n_10044 = n_9878 ^ x20;
assign n_10045 = n_9879 ^ x23;
assign n_10046 = n_9880 ^ x26;
assign n_10047 = n_9881 ^ x29;
assign n_10048 = n_9882 ^ x32;
assign n_10049 = n_9883 ^ x35;
assign n_10050 = n_9884 ^ x38;
assign n_10051 = n_9885 ^ x41;
assign n_10052 = n_9886 ^ x44;
assign n_10053 = n_9887 ^ x47;
assign n_10054 = n_9888 ^ x50;
assign n_10055 = n_9889 ^ x53;
assign n_10056 = n_9890 ^ x56;
assign n_10057 = n_9891 ^ x59;
assign n_10058 = n_9892 ^ x62;
assign n_10059 = n_9907 ^ n_9783;
assign n_10060 = n_9911 ^ n_9638;
assign n_10061 = n_9912 ^ n_6526;
assign n_10062 = n_9915 ^ n_9629;
assign n_10063 = n_9917 ^ n_9630;
assign n_10064 = n_9919 ^ n_9631;
assign n_10065 = n_9920 ^ n_9913;
assign n_10066 = n_9920 ^ n_9770;
assign n_10067 = n_9921 ^ n_9774;
assign n_10068 = n_9923 ^ n_9640;
assign n_10069 = x63 & n_9924;
assign n_10070 = n_9925 ^ n_9632;
assign n_10071 = n_9925 & n_9926;
assign n_10072 = n_9927 ^ n_9645;
assign n_10073 = n_9928 ^ n_9909;
assign n_10074 = n_9929 ^ n_9646;
assign n_10075 = n_9930 ^ n_9768;
assign n_10076 = n_9931 ^ n_9641;
assign n_10077 = n_9932 ^ n_9637;
assign n_10078 = n_9932 ^ n_9063;
assign n_10079 = n_9933 ^ n_8287;
assign n_10080 = ~n_8687 & n_9934;
assign n_10081 = n_9936 ^ n_9652;
assign n_10082 = n_9938 ^ n_9653;
assign n_10083 = n_9940 ^ n_9654;
assign n_10084 = n_9942 ^ n_9655;
assign n_10085 = n_9944 ^ n_9656;
assign n_10086 = n_9946 ^ n_9658;
assign n_10087 = n_9947 ^ n_7882;
assign n_10088 = n_9949 ^ n_9661;
assign n_10089 = n_9951 ^ n_9663;
assign n_10090 = n_9952 ^ n_8555;
assign n_10091 = n_9952 & ~n_8693;
assign n_10092 = n_9953 ^ n_8286;
assign n_10093 = ~n_8803 & n_9954;
assign y11 = ~n_9955;
assign n_10094 = n_8685 & ~n_9956;
assign n_10095 = n_9958 ^ n_9669;
assign n_10096 = n_9960 ^ n_9670;
assign n_10097 = n_9962 ^ n_9671;
assign n_10098 = n_8293 ^ n_9963;
assign n_10099 = n_9964 ^ n_9672;
assign n_10100 = n_8302 ^ n_9965;
assign n_10101 = n_9966 ^ n_9673;
assign n_10102 = n_9967 ^ n_9096;
assign n_10103 = n_9967 ^ n_8951;
assign n_10104 = n_9968 ^ n_9497;
assign n_10105 = n_9968 ^ n_9355;
assign n_10106 = n_9969 ^ n_9908;
assign n_10107 = n_9970 ^ n_9678;
assign n_10108 = n_9972 ^ n_9680;
assign n_10109 = n_9974 ^ n_9685;
assign n_10110 = ~x0 & n_9975;
assign n_10111 = n_9976 ^ n_6482;
assign n_10112 = n_9977 ^ x93;
assign n_10113 = n_2148 ^ n_9978;
assign n_10114 = n_748 ^ n_9979;
assign n_10115 = n_2219 ^ n_9980;
assign n_10116 = n_2287 ^ n_9981;
assign n_10117 = n_2354 ^ n_9982;
assign n_10118 = n_2421 ^ n_9983;
assign n_10119 = n_2488 ^ n_9984;
assign n_10120 = n_2554 ^ n_9985;
assign n_10121 = n_2619 ^ n_9986;
assign n_10122 = n_2686 ^ n_9987;
assign n_10123 = n_2754 ^ n_9988;
assign n_10124 = n_2821 ^ n_9989;
assign n_10125 = n_2889 ^ n_9990;
assign n_10126 = n_2955 ^ n_9991;
assign n_10127 = n_3024 ^ n_9992;
assign n_10128 = n_3090 ^ n_9993;
assign n_10129 = n_3159 ^ n_9994;
assign n_10130 = n_3223 ^ n_9995;
assign n_10131 = n_3288 ^ n_9996;
assign n_10132 = n_3353 ^ n_9997;
assign n_10133 = n_1 & ~n_9998;
assign n_10134 = ~n_9998 & n_198;
assign n_10135 = n_9998 ^ x94;
assign n_10136 = n_5020 ^ n_9999;
assign n_10137 = n_5083 ^ n_10000;
assign n_10138 = n_5146 ^ n_10001;
assign n_10139 = n_5207 ^ n_10002;
assign n_10140 = n_5271 ^ n_10003;
assign n_10141 = n_5335 ^ n_10004;
assign n_10142 = n_5399 ^ n_10005;
assign n_10143 = n_5463 ^ n_10006;
assign n_10144 = n_5524 ^ n_10007;
assign n_10145 = n_5587 ^ n_10008;
assign n_10146 = n_5650 ^ n_10009;
assign n_10147 = n_5714 ^ n_10010;
assign n_10148 = n_5780 ^ n_10011;
assign n_10149 = n_5842 ^ n_10012;
assign n_10150 = n_5906 ^ n_10013;
assign n_10151 = n_5969 ^ n_10014;
assign n_10152 = n_6033 ^ n_10015;
assign n_10153 = n_6097 ^ n_10016;
assign n_10154 = n_6159 ^ n_10017;
assign n_10155 = n_6221 ^ n_10018;
assign n_10156 = n_10019 ^ x5;
assign n_10157 = n_10020 ^ x8;
assign n_10158 = n_10021 ^ x11;
assign n_10159 = n_10022 ^ x14;
assign n_10160 = n_10023 ^ x17;
assign n_10161 = n_10024 ^ x20;
assign n_10162 = n_10025 ^ x23;
assign n_10163 = n_10026 ^ x26;
assign n_10164 = n_10027 ^ x29;
assign n_10165 = n_10028 ^ x32;
assign n_10166 = n_10029 ^ x35;
assign n_10167 = n_10030 ^ x38;
assign n_10168 = n_10031 ^ x41;
assign n_10169 = n_10032 ^ x44;
assign n_10170 = n_10033 ^ x47;
assign n_10171 = n_10034 ^ x50;
assign n_10172 = n_10035 ^ x53;
assign n_10173 = n_10036 ^ x56;
assign n_10174 = n_10037 ^ x59;
assign n_10175 = n_10038 ^ x62;
assign n_10176 = n_9921 ^ n_10057;
assign n_10177 = n_10058 ^ n_4963;
assign n_10178 = ~n_4963 & n_10058;
assign n_10179 = n_10061 ^ n_3400;
assign n_10180 = n_10061 & n_6637;
assign n_10181 = n_10062 ^ n_9922;
assign n_10182 = n_10062 ^ n_9766;
assign n_10183 = n_10063 ^ n_9971;
assign n_10184 = n_10063 ^ n_9767;
assign n_10185 = n_9768 ^ n_10064;
assign n_10186 = n_9913 & n_10066;
assign n_10187 = n_10067 ^ n_10057;
assign n_10188 = n_9969 ^ n_10068;
assign n_10189 = ~n_9780 & ~n_10069;
assign n_10190 = n_10071 ^ n_9632;
assign n_10191 = n_10072 ^ n_10053;
assign n_10192 = n_10072 ^ n_9914;
assign n_10193 = n_10074 ^ n_10055;
assign n_10194 = n_10074 ^ n_9918;
assign n_10195 = n_10075 ^ n_10064;
assign n_10196 = n_10076 ^ n_9910;
assign n_10197 = n_10076 ^ n_10077;
assign n_10198 = ~n_9637 & ~n_10078;
assign n_10199 = n_10080 ^ n_9788;
assign n_10200 = n_10081 ^ n_7874;
assign n_10201 = n_10082 ^ n_9084;
assign n_10202 = n_10082 ^ n_8940;
assign n_10203 = n_10083 ^ n_8689;
assign n_10204 = n_10083 ^ n_8551;
assign n_10205 = n_10084 ^ n_9088;
assign n_10206 = n_10084 ^ n_8944;
assign n_10207 = n_10085 ^ n_7880;
assign n_10208 = n_10086 ^ n_8948;
assign n_10209 = n_10087 ^ n_9094;
assign n_10210 = n_10087 & ~n_9233;
assign n_10211 = n_10088 ^ n_8965;
assign n_10212 = n_10088 ^ n_8825;
assign n_10213 = n_10089 ^ n_7885;
assign n_10214 = n_10090 ^ n_8923;
assign n_10215 = n_10090 ^ n_8301;
assign n_10216 = n_10091 ^ n_9807;
assign n_10217 = n_10093 ^ n_9808;
assign n_10218 = n_10094 ^ n_9809;
assign n_10219 = n_10095 ^ n_9238;
assign n_10220 = n_10095 ^ n_9100;
assign n_10221 = n_10096 ^ n_9505;
assign n_10222 = n_10096 ^ n_9363;
assign n_10223 = n_10097 ^ n_9110;
assign n_10224 = n_10097 ^ n_8962;
assign n_10225 = n_10099 ^ n_9511;
assign n_10226 = n_10099 ^ n_9369;
assign n_10227 = n_10101 ^ n_8967;
assign n_10228 = n_10101 ^ n_8827;
assign n_10229 = n_10102 ^ n_8299;
assign n_10230 = ~n_9096 & n_10103;
assign n_10231 = n_10104 ^ n_9765;
assign n_10232 = ~n_9497 & ~n_10105;
assign n_10233 = n_10106 ^ n_10068;
assign n_10234 = n_10107 ^ n_10054;
assign n_10235 = n_10107 ^ n_9916;
assign n_10236 = n_10073 ^ n_10108;
assign n_10237 = n_9928 ^ n_10108;
assign n_10238 = n_10110 ^ n_9828;
assign n_10239 = ~x0 & ~n_10111;
assign n_10240 = n_10112 ^ n_6483;
assign n_10241 = n_5021 ^ n_10113;
assign n_10242 = n_5084 ^ n_10114;
assign n_10243 = n_5147 ^ n_10115;
assign n_10244 = n_5208 ^ n_10116;
assign n_10245 = n_5272 ^ n_10117;
assign n_10246 = n_5336 ^ n_10118;
assign n_10247 = n_5400 ^ n_10119;
assign n_10248 = n_5464 ^ n_10120;
assign n_10249 = n_5525 ^ n_10121;
assign n_10250 = n_5588 ^ n_10122;
assign n_10251 = n_5651 ^ n_10123;
assign n_10252 = n_5715 ^ n_10124;
assign n_10253 = n_5781 ^ n_10125;
assign n_10254 = n_5843 ^ n_10126;
assign n_10255 = n_5907 ^ n_10127;
assign n_10256 = n_5970 ^ n_10128;
assign n_10257 = n_6034 ^ n_10129;
assign n_10258 = n_6098 ^ n_10130;
assign n_10259 = n_6160 ^ n_10131;
assign n_10260 = n_6222 ^ n_10132;
assign n_10261 = n_10133 ^ x1;
assign n_10262 = n_1 & ~n_10134;
assign n_10263 = ~n_10134 & n_202;
assign n_10264 = n_10134 & ~n_206;
assign n_10265 = n_10134 ^ x95;
assign n_10266 = n_210 ^ n_10134;
assign n_10267 = n_655 & n_10135;
assign n_10268 = n_784 & n_10135;
assign n_10269 = ~n_3665 & n_10135;
assign n_10270 = n_854 & n_10135;
assign n_10271 = n_920 & n_10135;
assign n_10272 = n_986 & n_10135;
assign n_10273 = n_1052 & n_10135;
assign n_10274 = n_1117 & n_10135;
assign n_10275 = n_1181 & n_10135;
assign n_10276 = n_1248 & n_10135;
assign n_10277 = n_10135 & n_1314;
assign n_10278 = n_10135 & n_1380;
assign n_10279 = n_10135 & n_1445;
assign n_10280 = n_10135 & n_1510;
assign n_10281 = n_10135 & n_1576;
assign n_10282 = n_10135 & n_1641;
assign n_10283 = n_10135 & n_1706;
assign n_10284 = n_10135 & n_1771;
assign n_10285 = n_10135 & n_1835;
assign n_10286 = n_10135 & n_1899;
assign n_10287 = n_10136 ^ x5;
assign n_10288 = n_10137 ^ x8;
assign n_10289 = n_10138 ^ x11;
assign n_10290 = n_10139 ^ x14;
assign n_10291 = n_10140 ^ x17;
assign n_10292 = n_10141 ^ x20;
assign n_10293 = n_10142 ^ x23;
assign n_10294 = n_10143 ^ x26;
assign n_10295 = n_10144 ^ x29;
assign n_10296 = n_10145 ^ x32;
assign n_10297 = n_10146 ^ x35;
assign n_10298 = n_10147 ^ x38;
assign n_10299 = n_10148 ^ x41;
assign n_10300 = n_10149 ^ x44;
assign n_10301 = n_10150 ^ x47;
assign n_10302 = n_10151 ^ x50;
assign n_10303 = n_10152 ^ x53;
assign n_10304 = n_10153 ^ x56;
assign n_10305 = n_10154 ^ x59;
assign n_10306 = n_10155 ^ x62;
assign n_10307 = n_10174 ^ n_10065;
assign n_10308 = n_10175 ^ n_6402;
assign n_10309 = ~n_10067 & n_10176;
assign n_10310 = n_10178 ^ n_6344;
assign n_10311 = n_10180 ^ n_9912;
assign n_10312 = n_10181 ^ n_10170;
assign n_10313 = ~n_9922 & n_10182;
assign n_10314 = n_10183 ^ n_10171;
assign n_10315 = ~n_9971 & n_10184;
assign n_10316 = ~n_10075 & n_10185;
assign n_10317 = n_10186 ^ n_9920;
assign n_10318 = n_10106 & ~n_10188;
assign n_10319 = n_10189 ^ n_9489;
assign n_10320 = n_10189 ^ n_9343;
assign n_10321 = n_10190 ^ n_9769;
assign n_10322 = n_10191 ^ n_9914;
assign n_10323 = n_10191 & n_10192;
assign n_10324 = n_10193 ^ n_9918;
assign n_10325 = ~n_10193 & ~n_10194;
assign n_10326 = n_10195 ^ n_10172;
assign n_10327 = n_10196 ^ n_10077;
assign n_10328 = n_10196 & ~n_10197;
assign n_10329 = n_10198 ^ n_9487;
assign n_10330 = n_10199 ^ n_9106;
assign n_10331 = n_10199 ^ n_8958;
assign n_10332 = n_10200 ^ n_8938;
assign n_10333 = n_10200 & ~n_9082;
assign n_10334 = n_10201 ^ n_8290;
assign n_10335 = n_9084 & ~n_10202;
assign n_10336 = n_10203 ^ n_8291;
assign n_10337 = ~n_8689 & n_10204;
assign n_10338 = n_10205 ^ n_8294;
assign n_10339 = ~n_9088 & n_10206;
assign n_10340 = n_10207 ^ n_8946;
assign n_10341 = n_10207 & ~n_9090;
assign n_10342 = n_10208 ^ n_7881;
assign n_10343 = ~n_10208 & n_9092;
assign n_10344 = n_10209 ^ n_8297;
assign n_10345 = n_10210 ^ n_9947;
assign n_10346 = n_10211 ^ n_8298;
assign n_10347 = ~n_8965 & n_10212;
assign n_10348 = n_10213 ^ n_8678;
assign n_10349 = n_10213 & ~n_8815;
assign n_10350 = n_10216 ^ n_9245;
assign n_10351 = n_10216 ^ n_9112;
assign n_10352 = n_10217 ^ n_9224;
assign n_10353 = n_10217 ^ n_9078;
assign n_10354 = n_10218 ^ n_9104;
assign n_10355 = n_10218 ^ n_8956;
assign n_10356 = n_10219 ^ n_8454;
assign n_10357 = ~n_9238 & n_10220;
assign n_10358 = n_10221 ^ n_8357;
assign n_10359 = ~n_9505 & n_10222;
assign n_10360 = n_10223 ^ n_8361;
assign n_10361 = ~n_9110 & n_10224;
assign n_10362 = n_10225 ^ n_8362;
assign n_10363 = ~n_9511 & n_10226;
assign n_10364 = n_10227 ^ n_8918;
assign n_10365 = n_8967 & ~n_10228;
assign n_10366 = n_10229 ^ n_8786;
assign n_10367 = n_10230 ^ n_9967;
assign n_10368 = n_10232 ^ n_9968;
assign n_10369 = n_10234 ^ n_9916;
assign n_10370 = ~n_10234 & ~n_10235;
assign n_10371 = ~n_10073 & n_10237;
assign n_10372 = n_10239 ^ n_9976;
assign n_10373 = ~x0 & ~n_10240;
assign n_10374 = n_10241 ^ x5;
assign n_10375 = n_10242 ^ x8;
assign n_10376 = n_10243 ^ x11;
assign n_10377 = n_10244 ^ x14;
assign n_10378 = n_10245 ^ x17;
assign n_10379 = n_10246 ^ x20;
assign n_10380 = n_10247 ^ x23;
assign n_10381 = n_10248 ^ x26;
assign n_10382 = n_10249 ^ x29;
assign n_10383 = n_10250 ^ x32;
assign n_10384 = n_10251 ^ x35;
assign n_10385 = n_10252 ^ x38;
assign n_10386 = n_10253 ^ x41;
assign n_10387 = n_10254 ^ x44;
assign n_10388 = n_10255 ^ x47;
assign n_10389 = n_10256 ^ x50;
assign n_10390 = n_10257 ^ x53;
assign n_10391 = n_10258 ^ x56;
assign n_10392 = n_10259 ^ x59;
assign n_10393 = n_10260 ^ x62;
assign n_10394 = n_10261 ^ x94;
assign n_10395 = n_10262 ^ x1;
assign n_10396 = n_1 & ~n_10263;
assign n_10397 = n_10263 ^ x96;
assign n_10398 = n_10264 ^ x94;
assign n_10399 = n_655 & n_10265;
assign n_10400 = n_784 & n_10265;
assign n_10401 = ~n_3665 & n_10265;
assign n_10402 = n_854 & n_10265;
assign n_10403 = n_920 & n_10265;
assign n_10404 = n_986 & n_10265;
assign n_10405 = n_1052 & n_10265;
assign n_10406 = n_1117 & n_10265;
assign n_10407 = n_1181 & n_10265;
assign n_10408 = n_1248 & n_10265;
assign n_10409 = n_10265 & n_1314;
assign n_10410 = n_10265 & n_1380;
assign n_10411 = n_10265 & n_1445;
assign n_10412 = n_10265 & n_1510;
assign n_10413 = n_10265 & n_1576;
assign n_10414 = n_10265 & n_1641;
assign n_10415 = n_10265 & n_1706;
assign n_10416 = n_10265 & n_1771;
assign n_10417 = n_10265 & n_1835;
assign n_10418 = n_10265 & n_1899;
assign n_10419 = n_3493 & ~n_10266;
assign n_10420 = n_2149 ^ n_10267;
assign n_10421 = n_749 ^ n_10268;
assign n_10422 = n_2220 ^ n_10269;
assign n_10423 = n_2288 ^ n_10270;
assign n_10424 = n_2355 ^ n_10271;
assign n_10425 = n_2422 ^ n_10272;
assign n_10426 = n_2489 ^ n_10273;
assign n_10427 = n_2555 ^ n_10274;
assign n_10428 = n_2620 ^ n_10275;
assign n_10429 = n_2687 ^ n_10276;
assign n_10430 = n_2755 ^ n_10277;
assign n_10431 = n_2822 ^ n_10278;
assign n_10432 = n_2890 ^ n_10279;
assign n_10433 = n_2956 ^ n_10280;
assign n_10434 = n_3025 ^ n_10281;
assign n_10435 = n_3091 ^ n_10282;
assign n_10436 = n_3160 ^ n_10283;
assign n_10437 = n_3224 ^ n_10284;
assign n_10438 = n_3289 ^ n_10285;
assign n_10439 = n_3354 ^ n_10286;
assign n_10440 = n_10301 ^ n_10233;
assign n_10441 = n_10302 ^ n_10236;
assign n_10442 = n_10305 ^ n_10179;
assign n_10443 = n_10306 ^ n_6638;
assign n_10444 = n_10306 ^ n_6527;
assign n_10445 = n_10309 ^ n_10057;
assign n_10446 = n_10310 ^ n_6345;
assign n_10447 = n_10311 ^ n_10177;
assign n_10448 = n_10313 ^ n_10062;
assign n_10449 = n_10315 ^ n_10063;
assign n_10450 = n_10316 ^ n_10064;
assign n_10451 = n_10179 ^ n_10317;
assign n_10452 = n_10318 ^ n_9908;
assign n_10453 = n_9769 ^ n_10319;
assign n_10454 = n_9489 & n_10320;
assign n_10455 = n_10321 ^ n_10319;
assign n_10456 = n_10323 ^ n_10053;
assign n_10457 = n_10325 ^ n_10055;
assign n_10458 = n_10303 ^ n_10327;
assign n_10459 = n_10328 ^ n_9910;
assign n_10460 = n_10329 ^ n_10070;
assign n_10461 = n_10329 ^ n_10056;
assign n_10462 = n_10330 ^ n_8356;
assign n_10463 = ~n_9106 & n_10331;
assign n_10464 = n_10332 ^ n_8289;
assign n_10465 = n_10333 ^ n_10081;
assign n_10466 = n_10335 ^ n_10082;
assign n_10467 = n_10337 ^ n_10083;
assign n_10468 = n_10339 ^ n_10084;
assign n_10469 = n_10340 ^ n_8295;
assign n_10470 = n_10341 ^ n_10085;
assign n_10471 = n_10342 ^ n_8296;
assign n_10472 = n_10343 ^ n_10086;
assign n_10473 = n_10345 ^ n_9519;
assign n_10474 = n_10345 ^ n_9376;
assign n_10475 = n_10347 ^ n_10088;
assign n_10476 = n_8300 ^ n_10348;
assign n_10477 = n_10349 ^ n_10089;
assign n_10478 = n_10350 ^ n_8370;
assign n_10479 = ~n_9245 & n_10351;
assign n_10480 = n_10352 ^ n_8355;
assign n_10481 = ~n_9224 & n_10353;
assign y12 = n_10354;
assign n_10482 = ~n_9104 & n_10355;
assign n_10483 = n_10357 ^ n_10095;
assign n_10484 = n_10359 ^ n_10096;
assign n_10485 = n_10361 ^ n_10097;
assign n_10486 = n_10363 ^ n_10099;
assign n_10487 = n_10365 ^ n_10101;
assign n_10488 = n_10367 ^ n_9662;
assign n_10489 = n_10367 ^ n_9521;
assign n_10490 = n_10368 ^ n_10059;
assign n_10491 = n_10368 ^ n_9783;
assign n_10492 = n_10370 ^ n_10054;
assign n_10493 = n_10371 ^ n_9909;
assign n_10494 = n_10373 ^ n_10112;
assign n_10495 = n_10387 ^ n_10322;
assign n_10496 = n_10388 ^ n_10369;
assign n_10497 = n_10389 ^ n_10324;
assign n_10498 = n_10392 ^ n_10311;
assign n_10499 = n_10393 ^ ~n_6528;
assign n_10500 = ~n_6528 & n_10393;
assign n_10501 = n_10394 ^ n_3488;
assign n_10502 = n_10395 ^ x95;
assign n_10503 = n_10396 ^ x1;
assign n_10504 = n_655 & n_10397;
assign n_10505 = n_784 & n_10397;
assign n_10506 = ~n_3665 & n_10397;
assign n_10507 = n_854 & n_10397;
assign n_10508 = n_920 & n_10397;
assign n_10509 = n_986 & n_10397;
assign n_10510 = n_1052 & n_10397;
assign n_10511 = n_1117 & n_10397;
assign n_10512 = n_1181 & n_10397;
assign n_10513 = n_1248 & n_10397;
assign n_10514 = n_10397 & n_1314;
assign n_10515 = n_10397 & n_1380;
assign n_10516 = n_10397 & n_1445;
assign n_10517 = n_10397 & n_1510;
assign n_10518 = n_10397 & n_1576;
assign n_10519 = n_10397 & n_1641;
assign n_10520 = n_10397 & n_1706;
assign n_10521 = n_10397 & n_1771;
assign n_10522 = n_10397 & n_1835;
assign n_10523 = n_10397 & n_1899;
assign n_10524 = n_10398 ^ x96;
assign n_10525 = n_2150 ^ n_10399;
assign n_10526 = n_750 ^ n_10400;
assign n_10527 = n_2221 ^ n_10401;
assign n_10528 = n_2289 ^ n_10402;
assign n_10529 = n_2356 ^ n_10403;
assign n_10530 = n_2423 ^ n_10404;
assign n_10531 = n_2490 ^ n_10405;
assign n_10532 = n_2556 ^ n_10406;
assign n_10533 = n_2621 ^ n_10407;
assign n_10534 = n_2688 ^ n_10408;
assign n_10535 = n_2756 ^ n_10409;
assign n_10536 = n_2823 ^ n_10410;
assign n_10537 = n_2891 ^ n_10411;
assign n_10538 = n_2957 ^ n_10412;
assign n_10539 = n_3026 ^ n_10413;
assign n_10540 = n_3092 ^ n_10414;
assign n_10541 = n_3161 ^ n_10415;
assign n_10542 = n_3225 ^ n_10416;
assign n_10543 = n_3290 ^ n_10417;
assign n_10544 = n_3355 ^ n_10418;
assign n_10545 = n_10419 ^ n_2059;
assign n_10546 = n_5022 ^ n_10420;
assign n_10547 = n_5085 ^ n_10421;
assign n_10548 = n_5148 ^ n_10422;
assign n_10549 = n_5209 ^ n_10423;
assign n_10550 = n_5273 ^ n_10424;
assign n_10551 = n_5337 ^ n_10425;
assign n_10552 = n_5401 ^ n_10426;
assign n_10553 = n_5465 ^ n_10427;
assign n_10554 = n_5526 ^ n_10428;
assign n_10555 = n_5589 ^ n_10429;
assign n_10556 = n_5652 ^ n_10430;
assign n_10557 = n_5716 ^ n_10431;
assign n_10558 = n_5782 ^ n_10432;
assign n_10559 = n_5844 ^ n_10433;
assign n_10560 = n_5908 ^ n_10434;
assign n_10561 = n_5971 ^ n_10435;
assign n_10562 = n_6035 ^ n_10436;
assign n_10563 = n_6099 ^ n_10437;
assign n_10564 = n_6161 ^ n_10438;
assign n_10565 = n_6223 ^ n_10439;
assign n_10566 = n_10442 ^ n_10317;
assign n_10567 = n_6638 & n_10444;
assign n_10568 = n_10445 ^ n_10174;
assign n_10569 = n_10308 ^ n_10446;
assign n_10570 = n_10175 ^ n_10446;
assign n_10571 = n_10448 ^ n_10440;
assign n_10572 = n_10448 ^ n_10233;
assign n_10573 = n_10449 ^ n_10441;
assign n_10574 = n_10449 ^ n_10236;
assign n_10575 = n_10450 ^ n_10303;
assign n_10576 = ~n_10442 & n_10451;
assign n_10577 = n_10369 ^ n_10452;
assign n_10578 = n_10321 & n_10453;
assign n_10579 = n_10454 ^ n_10189;
assign n_10580 = n_10455 ^ n_10173;
assign n_10581 = n_10456 ^ n_10312;
assign n_10582 = n_10456 ^ n_10170;
assign n_10583 = n_10457 ^ n_10326;
assign n_10584 = n_10457 ^ n_10172;
assign n_10585 = n_10460 ^ n_10056;
assign n_10586 = n_10460 & n_10461;
assign n_10587 = n_10463 ^ n_10199;
assign n_10588 = n_10465 ^ n_9507;
assign n_10589 = n_10465 ^ n_9365;
assign n_10590 = n_10466 ^ n_9509;
assign n_10591 = n_10466 ^ n_9367;
assign n_10592 = n_10467 ^ n_9108;
assign n_10593 = n_10467 ^ n_8960;
assign n_10594 = n_10468 ^ n_9513;
assign n_10595 = n_10468 ^ n_9371;
assign n_10596 = n_10470 ^ n_9657;
assign n_10597 = n_10470 ^ n_9515;
assign n_10598 = n_10472 ^ n_9517;
assign n_10599 = n_10472 ^ n_9374;
assign n_10600 = n_8366 ^ n_10473;
assign n_10601 = ~n_9519 & n_10474;
assign n_10602 = n_10475 ^ n_9392;
assign n_10603 = n_10475 ^ n_9247;
assign n_10604 = n_10477 ^ n_9236;
assign n_10605 = n_10477 ^ n_9098;
assign n_10606 = n_10479 ^ n_10216;
assign n_10607 = n_10481 ^ n_10217;
assign n_10608 = n_10482 ^ n_10218;
assign n_10609 = n_10483 ^ n_9666;
assign n_10610 = n_10483 ^ n_9525;
assign n_10611 = n_10484 ^ n_9935;
assign n_10612 = n_10484 ^ n_9789;
assign n_10613 = n_10485 ^ n_9535;
assign n_10614 = n_10485 ^ n_9388;
assign n_10615 = n_10486 ^ n_9941;
assign n_10616 = n_10486 ^ n_9795;
assign n_10617 = n_10487 ^ n_9059;
assign n_10618 = n_8368 ^ n_10488;
assign n_10619 = n_9662 & ~n_10489;
assign n_10620 = n_10490 ^ n_10300;
assign n_10621 = n_10059 & n_10491;
assign n_10622 = n_10492 ^ n_10314;
assign n_10623 = n_10492 ^ n_10171;
assign n_10624 = n_10324 ^ n_10493;
assign n_10625 = n_10496 ^ n_10452;
assign n_10626 = n_10497 ^ n_10493;
assign n_10627 = n_10498 ^ n_10177;
assign n_10628 = n_10498 & n_10447;
assign n_10629 = n_10500 ^ n_6269;
assign n_10630 = ~x0 & n_10501;
assign n_10631 = n_10502 ^ n_6484;
assign n_10632 = n_10503 ^ x96;
assign n_10633 = n_2151 ^ n_10504;
assign n_10634 = n_751 ^ n_10505;
assign n_10635 = n_2222 ^ n_10506;
assign n_10636 = n_2290 ^ n_10507;
assign n_10637 = n_2357 ^ n_10508;
assign n_10638 = n_2424 ^ n_10509;
assign n_10639 = n_2491 ^ n_10510;
assign n_10640 = n_2557 ^ n_10511;
assign n_10641 = n_2622 ^ n_10512;
assign n_10642 = n_2689 ^ n_10513;
assign n_10643 = n_2757 ^ n_10514;
assign n_10644 = n_2824 ^ n_10515;
assign n_10645 = n_2892 ^ n_10516;
assign n_10646 = n_2958 ^ n_10517;
assign n_10647 = n_3027 ^ n_10518;
assign n_10648 = n_3093 ^ n_10519;
assign n_10649 = n_3162 ^ n_10520;
assign n_10650 = n_3226 ^ n_10521;
assign n_10651 = n_3291 ^ n_10522;
assign n_10652 = n_3356 ^ n_10523;
assign n_10653 = n_205 & n_10524;
assign n_10654 = n_5023 ^ n_10525;
assign n_10655 = n_5086 ^ n_10526;
assign n_10656 = n_5149 ^ n_10527;
assign n_10657 = n_5210 ^ n_10528;
assign n_10658 = n_5274 ^ n_10529;
assign n_10659 = n_5338 ^ n_10530;
assign n_10660 = n_5402 ^ n_10531;
assign n_10661 = n_5466 ^ n_10532;
assign n_10662 = n_5527 ^ n_10533;
assign n_10663 = n_5590 ^ n_10534;
assign n_10664 = n_5653 ^ n_10535;
assign n_10665 = n_5717 ^ n_10536;
assign n_10666 = n_5783 ^ n_10537;
assign n_10667 = n_5845 ^ n_10538;
assign n_10668 = n_5909 ^ n_10539;
assign n_10669 = n_5972 ^ n_10540;
assign n_10670 = n_6036 ^ n_10541;
assign n_10671 = n_6100 ^ n_10542;
assign n_10672 = n_6162 ^ n_10543;
assign n_10673 = n_6224 ^ n_10544;
assign n_10674 = n_10545 ^ n_210;
assign n_10675 = n_10546 ^ x5;
assign n_10676 = n_10547 ^ x8;
assign n_10677 = n_10548 ^ x11;
assign n_10678 = n_10549 ^ x14;
assign n_10679 = n_10550 ^ x17;
assign n_10680 = n_10551 ^ x20;
assign n_10681 = n_10552 ^ x23;
assign n_10682 = n_10553 ^ x26;
assign n_10683 = n_10554 ^ x29;
assign n_10684 = n_10555 ^ x32;
assign n_10685 = n_10556 ^ x35;
assign n_10686 = n_10557 ^ x38;
assign n_10687 = n_10558 ^ x41;
assign n_10688 = n_10559 ^ x44;
assign n_10689 = n_10560 ^ x47;
assign n_10690 = n_10561 ^ x50;
assign n_10691 = n_10562 ^ x53;
assign n_10692 = n_10563 ^ x56;
assign n_10693 = n_10564 ^ x59;
assign n_10694 = n_10565 ^ x62;
assign n_10695 = n_10567 ^ n_10306;
assign n_10696 = n_10568 ^ n_10065;
assign n_10697 = n_10568 & n_10307;
assign n_10698 = n_10308 & n_10570;
assign n_10699 = n_10440 & ~n_10572;
assign n_10700 = ~n_10441 & n_10574;
assign n_10701 = n_10575 ^ n_10327;
assign n_10702 = n_10575 & ~n_10458;
assign n_10703 = n_10576 ^ n_10305;
assign n_10704 = n_10496 & ~n_10577;
assign n_10705 = n_10578 ^ n_10190;
assign n_10706 = n_10579 ^ n_10060;
assign n_10707 = n_10579 ^ n_9638;
assign n_10708 = ~n_10312 & n_10582;
assign n_10709 = ~n_10326 & n_10584;
assign n_10710 = n_10585 ^ n_10390;
assign n_10711 = n_10585 ^ n_10459;
assign n_10712 = n_10586 ^ n_10056;
assign n_10713 = n_10587 ^ n_9531;
assign n_10714 = n_10587 ^ n_9384;
assign n_10715 = n_10588 ^ n_8358;
assign n_10716 = n_9507 & ~n_10589;
assign n_10717 = n_10590 ^ n_8359;
assign n_10718 = ~n_9509 & n_10591;
assign n_10719 = n_10592 ^ n_8360;
assign n_10720 = ~n_9108 & n_10593;
assign n_10721 = n_10594 ^ n_8363;
assign n_10722 = n_9513 & ~n_10595;
assign n_10723 = n_10596 ^ n_8364;
assign n_10724 = ~n_9657 & n_10597;
assign n_10725 = n_10598 ^ n_8365;
assign n_10726 = n_9517 & ~n_10599;
assign n_10727 = n_10601 ^ n_10345;
assign n_10728 = n_8367 ^ n_10602;
assign n_10729 = ~n_9392 & n_10603;
assign n_10730 = n_10604 ^ n_8369;
assign n_10731 = n_9236 & ~n_10605;
assign n_10732 = n_10606 ^ n_8144;
assign n_10733 = n_10607 ^ n_9650;
assign n_10734 = n_10607 ^ n_9503;
assign n_10735 = n_10608 ^ n_9529;
assign n_10736 = n_10608 ^ n_9382;
assign n_10737 = n_10609 ^ n_8706;
assign n_10738 = ~n_9666 & n_10610;
assign n_10739 = n_10611 ^ n_8639;
assign n_10740 = ~n_9935 & n_10612;
assign n_10741 = n_10613 ^ n_8643;
assign n_10742 = ~n_9535 & n_10614;
assign n_10743 = n_10615 ^ n_8644;
assign n_10744 = ~n_9941 & n_10616;
assign n_10745 = n_10617 ^ n_9249;
assign n_10746 = n_10617 & n_9394;
assign n_10747 = n_10619 ^ n_10367;
assign n_10748 = n_10621 ^ n_9907;
assign n_10749 = ~n_10314 & n_10623;
assign n_10750 = n_10497 & ~n_10624;
assign n_10751 = n_10628 ^ n_10392;
assign n_10752 = n_10629 ^ n_6405;
assign n_10753 = n_10630 ^ n_10394;
assign n_10754 = ~x0 & ~n_10631;
assign n_10755 = n_10632 ^ n_3491;
assign n_10756 = n_5024 ^ n_10633;
assign n_10757 = n_5087 ^ n_10634;
assign n_10758 = n_5150 ^ n_10635;
assign n_10759 = n_5211 ^ n_10636;
assign n_10760 = n_5275 ^ n_10637;
assign n_10761 = n_5339 ^ n_10638;
assign n_10762 = n_5403 ^ n_10639;
assign n_10763 = n_5467 ^ n_10640;
assign n_10764 = n_5528 ^ n_10641;
assign n_10765 = n_5591 ^ n_10642;
assign n_10766 = n_5654 ^ n_10643;
assign n_10767 = n_5718 ^ n_10644;
assign n_10768 = n_5784 ^ n_10645;
assign n_10769 = n_5846 ^ n_10646;
assign n_10770 = n_5910 ^ n_10647;
assign n_10771 = n_5973 ^ n_10648;
assign n_10772 = n_6037 ^ n_10649;
assign n_10773 = n_6101 ^ n_10650;
assign n_10774 = n_6163 ^ n_10651;
assign n_10775 = n_6225 ^ n_10652;
assign n_10776 = n_1 & ~n_10653;
assign n_10777 = n_10653 ^ x97;
assign n_10778 = n_10654 ^ x5;
assign n_10779 = n_10655 ^ x8;
assign n_10780 = n_10656 ^ x11;
assign n_10781 = n_10657 ^ x14;
assign n_10782 = n_10658 ^ x17;
assign n_10783 = n_10659 ^ x20;
assign n_10784 = n_10660 ^ x23;
assign n_10785 = n_10661 ^ x26;
assign n_10786 = n_10662 ^ x29;
assign n_10787 = n_10663 ^ x32;
assign n_10788 = n_10664 ^ x35;
assign n_10789 = n_10665 ^ x38;
assign n_10790 = n_10666 ^ x41;
assign n_10791 = n_10667 ^ x44;
assign n_10792 = n_10668 ^ x47;
assign n_10793 = n_10669 ^ x50;
assign n_10794 = n_10670 ^ x53;
assign n_10795 = n_10671 ^ x56;
assign n_10796 = n_10672 ^ x59;
assign n_10797 = n_10673 ^ x62;
assign n_10798 = n_10674 ^ n_205;
assign n_10799 = n_10581 ^ n_10688;
assign n_10800 = n_10689 ^ n_10622;
assign n_10801 = n_10690 ^ n_10583;
assign n_10802 = n_10693 ^ n_10569;
assign n_10803 = n_6405 ^ n_10694;
assign n_10804 = n_10695 ^ n_10499;
assign n_10805 = n_10696 ^ n_10692;
assign n_10806 = n_10697 ^ n_10445;
assign n_10807 = n_10698 ^ n_10446;
assign n_10808 = n_10699 ^ n_10301;
assign n_10809 = n_10700 ^ n_10302;
assign n_10810 = n_10702 ^ n_10450;
assign n_10811 = n_10703 ^ n_10627;
assign n_10812 = n_10704 ^ n_10388;
assign n_10813 = n_10705 ^ n_10304;
assign n_10814 = n_10304 ^ n_10706;
assign n_10815 = ~n_10060 & n_10707;
assign n_10816 = n_10708 ^ n_10456;
assign n_10817 = n_10709 ^ n_10457;
assign n_10818 = n_10710 ^ n_10459;
assign n_10819 = ~n_10710 & n_10711;
assign n_10820 = n_10712 ^ n_10580;
assign n_10821 = n_10712 ^ n_10173;
assign n_10822 = n_10713 ^ n_8638;
assign n_10823 = ~n_9531 & n_10714;
assign n_10824 = n_10716 ^ n_10465;
assign n_10825 = n_10718 ^ n_10466;
assign n_10826 = n_10720 ^ n_10467;
assign n_10827 = n_10722 ^ n_10468;
assign n_10828 = n_10724 ^ n_10470;
assign n_10829 = n_10726 ^ n_10472;
assign n_10830 = n_10727 ^ n_8140;
assign n_10831 = n_10729 ^ n_10475;
assign n_10832 = n_10731 ^ n_10477;
assign n_10833 = n_10732 ^ n_9390;
assign n_10834 = n_10732 & ~n_9537;
assign n_10835 = n_10733 ^ n_8637;
assign n_10836 = ~n_9650 & n_10734;
assign y13 = n_10735;
assign n_10837 = ~n_9529 & n_10736;
assign n_10838 = n_10738 ^ n_10483;
assign n_10839 = n_10740 ^ n_10484;
assign n_10840 = n_10742 ^ n_10485;
assign n_10841 = n_10744 ^ n_10486;
assign n_10842 = n_10745 ^ n_9483;
assign n_10843 = n_10746 ^ n_10487;
assign n_10844 = n_10747 ^ n_9950;
assign n_10845 = n_10747 ^ n_9805;
assign n_10846 = n_10748 ^ n_10495;
assign n_10847 = n_10748 ^ n_10322;
assign n_10848 = n_10749 ^ n_10492;
assign n_10849 = n_10750 ^ n_10389;
assign n_10850 = n_10751 ^ n_10693;
assign n_10851 = n_10752 ^ n_10694;
assign n_10852 = n_10754 ^ n_10502;
assign n_10853 = ~x0 & n_10755;
assign n_10854 = n_10756 ^ x5;
assign n_10855 = n_10757 ^ x8;
assign n_10856 = n_10758 ^ x11;
assign n_10857 = n_10759 ^ x14;
assign n_10858 = n_10760 ^ x17;
assign n_10859 = n_10761 ^ x20;
assign n_10860 = n_10762 ^ x23;
assign n_10861 = n_10763 ^ x26;
assign n_10862 = n_10764 ^ x29;
assign n_10863 = n_10765 ^ x32;
assign n_10864 = n_10766 ^ x35;
assign n_10865 = n_10767 ^ x38;
assign n_10866 = n_10768 ^ x41;
assign n_10867 = n_10769 ^ x44;
assign n_10868 = n_10770 ^ x47;
assign n_10869 = n_10771 ^ x50;
assign n_10870 = n_10772 ^ x53;
assign n_10871 = n_10773 ^ x56;
assign n_10872 = n_10774 ^ x59;
assign n_10873 = n_10775 ^ x62;
assign n_10874 = n_10776 ^ x1;
assign n_10875 = n_655 & n_10777;
assign n_10876 = n_784 & n_10777;
assign n_10877 = ~n_3665 & n_10777;
assign n_10878 = n_854 & n_10777;
assign n_10879 = n_920 & n_10777;
assign n_10880 = n_986 & n_10777;
assign n_10881 = n_1052 & n_10777;
assign n_10882 = n_1117 & n_10777;
assign n_10883 = n_1181 & n_10777;
assign n_10884 = n_1248 & n_10777;
assign n_10885 = n_1314 & n_10777;
assign n_10886 = n_10777 & n_1380;
assign n_10887 = n_10777 & n_1445;
assign n_10888 = n_10777 & n_1510;
assign n_10889 = n_10777 & n_1576;
assign n_10890 = n_10777 & n_1641;
assign n_10891 = n_10777 & n_1706;
assign n_10892 = n_10777 & n_1771;
assign n_10893 = n_10777 & n_1835;
assign n_10894 = n_10777 & n_1899;
assign n_10895 = n_10791 ^ n_10571;
assign n_10896 = n_10792 ^ n_10573;
assign n_10897 = n_10793 ^ n_10701;
assign n_10898 = n_10795 ^ n_10566;
assign n_10899 = n_10796 ^ n_10443;
assign n_10900 = n_10797 ^ n_6639;
assign n_10901 = n_10797 ^ n_6529;
assign n_10902 = n_209 & n_10798;
assign n_10903 = ~n_10752 & n_10803;
assign n_10904 = n_10566 ^ n_10806;
assign n_10905 = n_10443 ^ n_10807;
assign n_10906 = n_10625 ^ n_10808;
assign n_10907 = n_10626 ^ n_10809;
assign n_10908 = n_10812 ^ n_10689;
assign n_10909 = n_10813 ^ n_10706;
assign n_10910 = n_10813 & n_10814;
assign n_10911 = n_10815 ^ n_9911;
assign n_10912 = n_10571 ^ n_10816;
assign n_10913 = n_10701 ^ n_10817;
assign n_10914 = n_10818 ^ n_10810;
assign n_10915 = n_10819 ^ n_10390;
assign n_10916 = n_10820 ^ n_10691;
assign n_10917 = ~n_10580 & ~n_10821;
assign n_10918 = n_10823 ^ n_10587;
assign n_10919 = n_10824 ^ n_9937;
assign n_10920 = n_10824 ^ n_9791;
assign n_10921 = n_10825 ^ n_9939;
assign n_10922 = n_10825 ^ n_9793;
assign n_10923 = n_10826 ^ n_9533;
assign n_10924 = n_10826 ^ n_9386;
assign n_10925 = n_10827 ^ n_9943;
assign n_10926 = n_10827 ^ n_9797;
assign n_10927 = n_10828 ^ n_8138;
assign n_10928 = n_10829 ^ n_9801;
assign n_10929 = n_10829 ^ n_9659;
assign n_10930 = n_10830 ^ n_9803;
assign n_10931 = n_10830 & ~n_9948;
assign n_10932 = n_10831 ^ n_8141;
assign n_10933 = n_10832 ^ n_8143;
assign n_10934 = n_10833 ^ n_8652;
assign n_10935 = n_10834 ^ n_10606;
assign n_10936 = n_10836 ^ n_10607;
assign n_10937 = n_10837 ^ n_10608;
assign n_10938 = n_10838 ^ n_10092;
assign n_10939 = n_10838 ^ n_9953;
assign n_10940 = n_10839 ^ n_10464;
assign n_10941 = n_10839 ^ n_10332;
assign n_10942 = n_10840 ^ n_8293;
assign n_10943 = n_10841 ^ n_10338;
assign n_10944 = n_10841 ^ n_10205;
assign n_10945 = n_10843 ^ n_9676;
assign n_10946 = n_10844 ^ n_8650;
assign n_10947 = ~n_9950 & n_10845;
assign n_10948 = ~n_10495 & n_10847;
assign n_10949 = n_10573 ^ n_10848;
assign n_10950 = n_10849 ^ n_10801;
assign n_10951 = n_10849 ^ n_10690;
assign n_10952 = n_10850 ^ n_10569;
assign n_10953 = n_10850 & n_10802;
assign n_10954 = n_10853 ^ n_10632;
assign n_10955 = n_10846 ^ n_10866;
assign n_10956 = n_10867 ^ n_10625;
assign n_10957 = n_10868 ^ n_10626;
assign n_10958 = n_10869 ^ n_10818;
assign n_10959 = n_10871 ^ n_10703;
assign n_10960 = n_10872 ^ n_10804;
assign n_10961 = n_10872 ^ n_10695;
assign n_10962 = n_10874 ^ x97;
assign n_10963 = n_2152 ^ n_10875;
assign n_10964 = n_752 ^ n_10876;
assign n_10965 = n_2223 ^ n_10877;
assign n_10966 = n_2291 ^ n_10878;
assign n_10967 = n_2358 ^ n_10879;
assign n_10968 = n_2425 ^ n_10880;
assign n_10969 = n_2492 ^ n_10881;
assign n_10970 = n_2558 ^ n_10882;
assign n_10971 = n_2623 ^ n_10883;
assign n_10972 = n_2690 ^ n_10884;
assign n_10973 = n_2758 ^ n_10885;
assign n_10974 = n_2825 ^ n_10886;
assign n_10975 = n_2893 ^ n_10887;
assign n_10976 = n_2959 ^ n_10888;
assign n_10977 = n_3028 ^ n_10889;
assign n_10978 = n_3094 ^ n_10890;
assign n_10979 = n_3163 ^ n_10891;
assign n_10980 = n_3227 ^ n_10892;
assign n_10981 = n_3292 ^ n_10893;
assign n_10982 = n_3357 ^ n_10894;
assign n_10983 = n_10895 ^ n_10816;
assign n_10984 = n_10896 ^ n_10848;
assign n_10985 = n_10897 ^ n_10817;
assign n_10986 = n_10898 ^ n_10806;
assign n_10987 = n_10899 ^ n_10807;
assign n_10988 = n_6639 & n_10901;
assign n_10989 = n_10902 ^ x96;
assign n_10990 = n_10903 ^ n_10629;
assign n_10991 = ~n_10898 & n_10904;
assign n_10992 = ~n_10899 & n_10905;
assign n_10993 = n_10908 ^ n_10622;
assign n_10994 = n_10908 & ~n_10800;
assign n_10995 = n_10910 ^ n_10705;
assign n_10996 = n_10911 ^ n_10391;
assign n_10997 = n_10911 ^ n_10187;
assign n_10998 = n_10895 & ~n_10912;
assign n_10999 = n_10897 & ~n_10913;
assign n_11000 = n_10691 ^ n_10915;
assign n_11001 = n_10916 ^ n_10915;
assign n_11002 = n_10917 ^ n_10455;
assign n_11003 = n_10918 ^ n_9959;
assign n_11004 = n_10918 ^ n_9812;
assign n_11005 = n_10919 ^ n_8640;
assign n_11006 = ~n_9937 & n_10920;
assign n_11007 = n_10921 ^ n_8641;
assign n_11008 = ~n_9939 & n_10922;
assign n_11009 = n_10923 ^ n_8642;
assign n_11010 = ~n_9533 & n_10924;
assign n_11011 = n_10925 ^ n_8645;
assign n_11012 = ~n_9943 & n_10926;
assign n_11013 = n_10927 ^ n_9799;
assign n_11014 = n_10927 & ~n_9945;
assign n_11015 = n_10928 ^ n_8647;
assign n_11016 = ~n_9801 & n_10929;
assign n_11017 = n_10930 ^ n_8648;
assign n_11018 = n_10931 ^ n_10727;
assign n_11019 = n_10932 ^ n_9674;
assign n_11020 = n_10932 & ~n_9818;
assign n_11021 = n_10933 ^ n_9523;
assign n_11022 = n_10933 & ~n_9664;
assign n_11023 = n_10935 ^ n_8302;
assign n_11024 = n_10936 ^ n_10079;
assign n_11025 = n_10936 ^ n_9933;
assign n_11026 = n_10937 ^ n_9957;
assign n_11027 = n_10937 ^ n_9810;
assign n_11028 = n_10938 ^ n_8835;
assign n_11029 = ~n_10092 & n_10939;
assign n_11030 = n_10940 ^ n_8776;
assign n_11031 = ~n_10464 & n_10941;
assign n_11032 = n_10942 ^ n_9963;
assign n_11033 = n_10942 & ~n_10098;
assign n_11034 = n_10943 ^ n_8781;
assign n_11035 = ~n_10338 & n_10944;
assign n_11036 = n_10945 ^ n_9628;
assign n_11037 = n_10945 & ~n_9820;
assign n_11038 = n_10947 ^ n_10747;
assign n_11039 = n_10948 ^ n_10387;
assign n_11040 = ~n_10896 & n_10949;
assign n_11041 = ~n_10801 & n_10951;
assign n_11042 = n_10953 ^ n_10751;
assign n_11043 = n_10956 ^ n_10808;
assign n_11044 = n_10956 & ~n_10906;
assign n_11045 = n_10957 ^ n_10809;
assign n_11046 = n_10957 & ~n_10907;
assign n_11047 = n_10958 ^ n_10810;
assign n_11048 = ~n_10958 & n_10914;
assign n_11049 = n_10959 ^ n_10627;
assign n_11050 = n_10959 & n_10811;
assign n_11051 = ~n_10804 & n_10961;
assign n_11052 = n_10962 ^ n_3492;
assign n_11053 = n_5025 ^ n_10963;
assign n_11054 = n_5088 ^ n_10964;
assign n_11055 = n_5151 ^ n_10965;
assign n_11056 = n_5212 ^ n_10966;
assign n_11057 = n_5276 ^ n_10967;
assign n_11058 = n_5340 ^ n_10968;
assign n_11059 = n_5404 ^ n_10969;
assign n_11060 = n_5468 ^ n_10970;
assign n_11061 = n_5529 ^ n_10971;
assign n_11062 = n_5592 ^ n_10972;
assign n_11063 = n_5655 ^ n_10973;
assign n_11064 = n_5719 ^ n_10974;
assign n_11065 = n_5785 ^ n_10975;
assign n_11066 = n_5847 ^ n_10976;
assign n_11067 = n_5911 ^ n_10977;
assign n_11068 = n_5974 ^ n_10978;
assign n_11069 = n_6038 ^ n_10979;
assign n_11070 = n_6102 ^ n_10980;
assign n_11071 = n_6164 ^ n_10981;
assign n_11072 = n_6226 ^ n_10982;
assign n_11073 = n_10988 ^ n_10797;
assign n_11074 = n_10989 ^ x97;
assign n_11075 = n_214 ^ n_10989;
assign n_11076 = n_10900 ^ n_10990;
assign n_11077 = n_10991 ^ n_10795;
assign n_11078 = n_10992 ^ n_10796;
assign n_11079 = n_10994 ^ n_10812;
assign n_11080 = n_10996 ^ n_10187;
assign n_11081 = n_10996 & ~n_10997;
assign n_11082 = n_10998 ^ n_10791;
assign n_11083 = n_10999 ^ n_10793;
assign n_11084 = n_10916 & n_11000;
assign n_11085 = n_11002 ^ n_10909;
assign n_11086 = n_11002 ^ n_10794;
assign n_11087 = n_11003 ^ n_8775;
assign n_11088 = ~n_9959 & n_11004;
assign n_11089 = n_11006 ^ n_10824;
assign n_11090 = n_11008 ^ n_10825;
assign n_11091 = n_11010 ^ n_10826;
assign n_11092 = n_11012 ^ n_10827;
assign n_11093 = n_11013 ^ n_8646;
assign n_11094 = n_11014 ^ n_10828;
assign n_11095 = n_11016 ^ n_10829;
assign n_11096 = n_11018 ^ n_10346;
assign n_11097 = n_11018 ^ n_10211;
assign n_11098 = n_11019 ^ n_8649;
assign n_11099 = n_11020 ^ n_10831;
assign n_11100 = n_11021 ^ n_8651;
assign n_11101 = n_11022 ^ n_10832;
assign n_11102 = n_11023 ^ n_9965;
assign n_11103 = n_11023 & ~n_10100;
assign n_11104 = n_11024 ^ n_8774;
assign n_11105 = ~n_10079 & n_11025;
assign y14 = n_11026;
assign n_11106 = ~n_9957 & n_11027;
assign n_11107 = n_11029 ^ n_10838;
assign n_11108 = n_11031 ^ n_10839;
assign n_11109 = n_8780 ^ n_11032;
assign n_11110 = n_11033 ^ n_10840;
assign n_11111 = n_11035 ^ n_10841;
assign n_11112 = n_11036 ^ n_10052;
assign n_11113 = n_11037 ^ n_10843;
assign n_11114 = n_11038 ^ n_8300;
assign n_11115 = n_11039 ^ n_10581;
assign n_11116 = n_11040 ^ n_10792;
assign n_11117 = n_11041 ^ n_10849;
assign n_11118 = n_10987 ^ n_11042;
assign n_11119 = n_11044 ^ n_10867;
assign n_11120 = n_11046 ^ n_10868;
assign n_11121 = n_11048 ^ n_10869;
assign n_11122 = n_11050 ^ n_10871;
assign n_11123 = n_11051 ^ n_10872;
assign n_11124 = ~x0 & n_11052;
assign n_11125 = n_11053 ^ x5;
assign n_11126 = n_11054 ^ x8;
assign n_11127 = n_11055 ^ x11;
assign n_11128 = n_11056 ^ x14;
assign n_11129 = n_11057 ^ x17;
assign n_11130 = n_11058 ^ x20;
assign n_11131 = n_11059 ^ x23;
assign n_11132 = n_11060 ^ x26;
assign n_11133 = n_11061 ^ x29;
assign n_11134 = n_11062 ^ x32;
assign n_11135 = n_11063 ^ x35;
assign n_11136 = n_11064 ^ x38;
assign n_11137 = n_11065 ^ x41;
assign n_11138 = n_11066 ^ x44;
assign n_11139 = n_11067 ^ x47;
assign n_11140 = n_11068 ^ x50;
assign n_11141 = n_11069 ^ x53;
assign n_11142 = n_11070 ^ x56;
assign n_11143 = n_11071 ^ x59;
assign n_11144 = n_11072 ^ x62;
assign n_11145 = n_11073 ^ ~n_6727;
assign n_11146 = ~n_6727 & ~n_11073;
assign n_11147 = n_1 & ~n_11074;
assign n_11148 = ~n_11074 & n_214;
assign n_11149 = n_655 & n_11075;
assign n_11150 = n_784 & n_11075;
assign n_11151 = ~n_3665 & n_11075;
assign n_11152 = n_854 & n_11075;
assign n_11153 = n_920 & n_11075;
assign n_11154 = n_986 & n_11075;
assign n_11155 = n_1052 & n_11075;
assign n_11156 = n_1117 & n_11075;
assign n_11157 = n_1181 & n_11075;
assign n_11158 = n_1248 & n_11075;
assign n_11159 = n_1314 & n_11075;
assign n_11160 = n_11075 & n_1380;
assign n_11161 = n_11075 & n_1445;
assign n_11162 = n_11075 & n_1510;
assign n_11163 = n_11075 & n_1576;
assign n_11164 = n_11075 & n_1641;
assign n_11165 = n_11075 & n_1706;
assign n_11166 = n_11075 & n_1771;
assign n_11167 = n_11075 & n_1835;
assign n_11168 = n_11075 & n_1899;
assign n_11169 = n_11077 ^ n_11049;
assign n_11170 = n_10960 ^ n_11078;
assign n_11171 = n_10984 ^ n_11079;
assign n_11172 = n_11080 ^ n_10870;
assign n_11173 = n_11080 ^ n_10995;
assign n_11174 = n_11081 ^ n_10391;
assign n_11175 = n_11082 ^ n_11043;
assign n_11176 = n_11083 ^ n_11047;
assign n_11177 = n_11084 ^ n_10915;
assign n_11178 = n_11085 ^ n_10794;
assign n_11179 = ~n_11085 & ~n_11086;
assign n_11180 = n_11088 ^ n_10918;
assign n_11181 = n_11089 ^ n_10334;
assign n_11182 = n_11089 ^ n_10201;
assign n_11183 = n_11090 ^ n_10336;
assign n_11184 = n_11090 ^ n_10203;
assign n_11185 = n_11091 ^ n_9961;
assign n_11186 = n_11091 ^ n_9814;
assign n_11187 = n_11092 ^ n_10469;
assign n_11188 = n_11092 ^ n_10340;
assign n_11189 = n_11094 ^ n_10471;
assign n_11190 = n_11094 ^ n_10342;
assign n_11191 = n_11095 ^ n_10344;
assign n_11192 = n_11095 ^ n_10209;
assign n_11193 = n_11096 ^ n_8785;
assign n_11194 = ~n_10346 & n_11097;
assign n_11195 = n_11099 ^ n_10366;
assign n_11196 = n_11099 ^ n_10102;
assign n_11197 = n_11101 ^ n_10214;
assign n_11198 = n_11101 ^ n_10090;
assign n_11199 = n_11102 ^ n_8789;
assign n_11200 = n_11103 ^ n_10935;
assign n_11201 = n_11105 ^ n_10936;
assign n_11202 = n_11106 ^ n_10937;
assign n_11203 = n_11107 ^ n_10480;
assign n_11204 = n_11107 ^ n_10352;
assign n_11205 = n_11108 ^ n_10715;
assign n_11206 = n_11108 ^ n_10588;
assign n_11207 = n_11110 ^ n_10362;
assign n_11208 = n_11110 ^ n_10225;
assign n_11209 = n_11111 ^ n_10721;
assign n_11210 = n_11111 ^ n_10594;
assign n_11211 = n_11113 ^ n_10104;
assign n_11212 = n_11114 ^ n_10348;
assign n_11213 = n_11114 & ~n_10476;
assign n_11214 = n_11115 ^ n_10688;
assign n_11215 = n_11115 & ~n_10799;
assign n_11216 = n_11045 ^ n_11116;
assign n_11217 = n_10985 ^ n_11117;
assign n_11218 = n_10952 ^ n_11122;
assign n_11219 = n_10851 ^ n_11123;
assign n_11220 = n_11124 ^ n_10962;
assign n_11221 = n_11138 ^ n_10993;
assign n_11222 = n_11138 ^ n_11119;
assign n_11223 = n_11139 ^ n_10950;
assign n_11224 = n_11139 ^ n_11120;
assign n_11225 = n_11140 ^ n_11001;
assign n_11226 = n_11140 ^ n_11121;
assign n_11227 = n_11142 ^ n_10952;
assign n_11228 = n_11143 ^ n_10851;
assign n_11229 = n_11144 ^ n_6407;
assign n_11230 = n_11145 ^ n_10873;
assign n_11231 = n_11146 ^ n_4966;
assign n_11232 = n_11147 ^ x1;
assign n_11233 = n_1 & ~n_11148;
assign n_11234 = ~n_11148 & n_216;
assign n_11235 = n_11148 ^ x99;
assign n_11236 = n_225 ^ n_11148;
assign n_11237 = n_2153 ^ n_11149;
assign n_11238 = n_753 ^ n_11150;
assign n_11239 = n_2224 ^ n_11151;
assign n_11240 = n_2292 ^ n_11152;
assign n_11241 = n_2359 ^ n_11153;
assign n_11242 = n_2426 ^ n_11154;
assign n_11243 = n_2493 ^ n_11155;
assign n_11244 = n_2559 ^ n_11156;
assign n_11245 = n_2624 ^ n_11157;
assign n_11246 = n_2691 ^ n_11158;
assign n_11247 = n_2759 ^ n_11159;
assign n_11248 = n_2826 ^ n_11160;
assign n_11249 = n_2894 ^ n_11161;
assign n_11250 = n_2960 ^ n_11162;
assign n_11251 = n_3029 ^ n_11163;
assign n_11252 = n_3095 ^ n_11164;
assign n_11253 = n_3164 ^ n_11165;
assign n_11254 = n_3228 ^ n_11166;
assign n_11255 = n_3293 ^ n_11167;
assign n_11256 = n_3358 ^ n_11168;
assign n_11257 = n_11172 ^ n_10995;
assign n_11258 = n_11172 & ~n_11173;
assign n_11259 = n_11174 ^ n_10805;
assign n_11260 = n_11174 ^ n_10692;
assign n_11261 = n_11178 ^ n_11177;
assign n_11262 = n_11179 ^ n_10794;
assign n_11263 = n_11180 ^ n_10358;
assign n_11264 = n_11180 ^ n_10221;
assign n_11265 = n_11181 ^ n_8777;
assign n_11266 = n_10334 & ~n_11182;
assign n_11267 = n_11183 ^ n_8778;
assign n_11268 = ~n_10336 & n_11184;
assign n_11269 = n_11185 ^ n_8779;
assign n_11270 = ~n_9961 & n_11186;
assign n_11271 = n_11187 ^ n_8782;
assign n_11272 = ~n_10469 & n_11188;
assign n_11273 = n_11189 ^ n_8783;
assign n_11274 = n_10471 & ~n_11190;
assign n_11275 = n_11191 ^ n_8784;
assign n_11276 = ~n_10344 & n_11192;
assign n_11277 = n_11194 ^ n_11018;
assign n_11278 = ~n_10229 & n_11196;
assign n_11279 = ~n_10215 & n_11198;
assign n_11280 = n_11200 ^ n_10364;
assign n_11281 = n_11200 ^ n_10227;
assign n_11282 = n_11201 ^ n_10462;
assign n_11283 = n_11201 ^ n_10330;
assign n_11284 = n_11202 ^ n_10356;
assign n_11285 = n_11202 ^ n_10219;
assign n_11286 = n_11203 ^ n_8976;
assign n_11287 = ~n_10480 & n_11204;
assign n_11288 = n_11205 ^ n_8905;
assign n_11289 = n_10715 & ~n_11206;
assign n_11290 = n_11207 ^ n_8909;
assign n_11291 = ~n_10362 & n_11208;
assign n_11292 = n_11209 ^ n_8910;
assign n_11293 = n_10721 & ~n_11210;
assign n_11294 = n_11211 ^ n_9765;
assign n_11295 = ~n_11211 & n_10231;
assign n_11296 = n_11212 ^ n_8787;
assign n_11297 = n_11213 ^ n_11038;
assign n_11298 = n_11137 ^ n_11214;
assign n_11299 = n_11215 ^ n_11039;
assign n_11300 = n_11221 ^ n_11119;
assign n_11301 = ~n_11221 & n_11222;
assign n_11302 = n_11223 ^ n_11120;
assign n_11303 = ~n_11223 & n_11224;
assign n_11304 = n_11225 ^ n_11121;
assign n_11305 = n_11225 & n_11226;
assign n_11306 = n_11227 ^ n_11122;
assign n_11307 = n_11227 & ~n_11218;
assign n_11308 = n_11228 ^ n_11123;
assign n_11309 = ~n_11228 & n_11219;
assign n_11310 = n_11229 ^ n_11231;
assign n_11311 = n_11144 ^ n_11231;
assign n_11312 = n_11232 ^ x98;
assign n_11313 = n_11233 ^ x1;
assign n_11314 = n_1 & ~n_11234;
assign n_11315 = n_11234 & n_220;
assign n_11316 = n_11234 ^ x100;
assign n_11317 = n_655 & n_11235;
assign n_11318 = n_784 & n_11235;
assign n_11319 = ~n_3665 & n_11235;
assign n_11320 = n_854 & n_11235;
assign n_11321 = n_920 & n_11235;
assign n_11322 = n_986 & n_11235;
assign n_11323 = n_1052 & n_11235;
assign n_11324 = n_1117 & n_11235;
assign n_11325 = n_1181 & n_11235;
assign n_11326 = n_1248 & n_11235;
assign n_11327 = n_1314 & n_11235;
assign n_11328 = n_11235 & n_1380;
assign n_11329 = n_11235 & n_1445;
assign n_11330 = n_11235 & n_1510;
assign n_11331 = n_11235 & n_1576;
assign n_11332 = n_11235 & n_1641;
assign n_11333 = n_11235 & n_1706;
assign n_11334 = n_11235 & n_1771;
assign n_11335 = n_11235 & n_1835;
assign n_11336 = n_11235 & n_1899;
assign n_11337 = ~n_11236 & n_3497;
assign n_11338 = n_5026 ^ n_11237;
assign n_11339 = n_5089 ^ n_11238;
assign n_11340 = n_5152 ^ n_11239;
assign n_11341 = n_5213 ^ n_11240;
assign n_11342 = n_5277 ^ n_11241;
assign n_11343 = n_5341 ^ n_11242;
assign n_11344 = n_5405 ^ n_11243;
assign n_11345 = n_5469 ^ n_11244;
assign n_11346 = n_5530 ^ n_11245;
assign n_11347 = n_5593 ^ n_11246;
assign n_11348 = n_5656 ^ n_11247;
assign n_11349 = n_5720 ^ n_11248;
assign n_11350 = n_5786 ^ n_11249;
assign n_11351 = n_5848 ^ n_11250;
assign n_11352 = n_5912 ^ n_11251;
assign n_11353 = n_5975 ^ n_11252;
assign n_11354 = n_6039 ^ n_11253;
assign n_11355 = n_6103 ^ n_11254;
assign n_11356 = n_6165 ^ n_11255;
assign n_11357 = n_6227 ^ n_11256;
assign n_11358 = n_11258 ^ n_10870;
assign n_11359 = n_11141 ^ n_11259;
assign n_11360 = n_10805 & n_11260;
assign n_11361 = n_11262 ^ n_11257;
assign n_11362 = n_11263 ^ n_8904;
assign n_11363 = ~n_10358 & n_11264;
assign n_11364 = n_11266 ^ n_11089;
assign n_11365 = n_11268 ^ n_11090;
assign n_11366 = n_11270 ^ n_11091;
assign n_11367 = n_11272 ^ n_11092;
assign n_11368 = n_11274 ^ n_11094;
assign n_11369 = n_11276 ^ n_11095;
assign n_11370 = n_11277 ^ n_8367;
assign n_11371 = n_11278 ^ n_11099;
assign n_11372 = n_11279 ^ n_11101;
assign n_11373 = n_11280 ^ n_9338;
assign n_11374 = n_10364 & ~n_11281;
assign n_11375 = n_11282 ^ n_8903;
assign n_11376 = ~n_10462 & n_11283;
assign y15 = n_11284;
assign n_11377 = ~n_10356 & n_11285;
assign n_11378 = n_11287 ^ n_11107;
assign n_11379 = n_11289 ^ n_11108;
assign n_11380 = n_11291 ^ n_11110;
assign n_11381 = n_11293 ^ n_11111;
assign n_11382 = n_11294 ^ n_10169;
assign n_11383 = n_11295 ^ n_11113;
assign n_11384 = n_11297 ^ n_10730;
assign n_11385 = n_11297 ^ n_10604;
assign n_11386 = n_11299 ^ n_10983;
assign n_11387 = n_11301 ^ n_11119;
assign n_11388 = n_11303 ^ n_11120;
assign n_11389 = n_11305 ^ n_11121;
assign n_11390 = n_11307 ^ n_11122;
assign n_11391 = n_11309 ^ n_11143;
assign n_11392 = n_11229 & ~n_11311;
assign n_11393 = n_11312 ^ n_2108;
assign n_11394 = n_11313 ^ x99;
assign n_11395 = n_11314 ^ x1;
assign n_11396 = n_11315 ^ n_220;
assign n_11397 = n_655 & n_11316;
assign n_11398 = n_784 & n_11316;
assign n_11399 = ~n_3665 & n_11316;
assign n_11400 = n_854 & n_11316;
assign n_11401 = n_920 & n_11316;
assign n_11402 = n_986 & n_11316;
assign n_11403 = n_1052 & n_11316;
assign n_11404 = n_1117 & n_11316;
assign n_11405 = n_1181 & n_11316;
assign n_11406 = n_1248 & n_11316;
assign n_11407 = n_1314 & n_11316;
assign n_11408 = n_1380 & n_11316;
assign n_11409 = n_11316 & n_1445;
assign n_11410 = n_11316 & n_1510;
assign n_11411 = n_11316 & n_1576;
assign n_11412 = n_11316 & n_1641;
assign n_11413 = n_11316 & n_1706;
assign n_11414 = n_11316 & n_1771;
assign n_11415 = n_11316 & n_1835;
assign n_11416 = n_11316 & n_1899;
assign n_11417 = n_2154 ^ n_11317;
assign n_11418 = n_754 ^ n_11318;
assign n_11419 = n_2225 ^ n_11319;
assign n_11420 = n_2293 ^ n_11320;
assign n_11421 = n_2360 ^ n_11321;
assign n_11422 = n_2427 ^ n_11322;
assign n_11423 = n_2494 ^ n_11323;
assign n_11424 = n_2560 ^ n_11324;
assign n_11425 = n_2625 ^ n_11325;
assign n_11426 = n_2692 ^ n_11326;
assign n_11427 = n_2760 ^ n_11327;
assign n_11428 = n_2827 ^ n_11328;
assign n_11429 = n_2895 ^ n_11329;
assign n_11430 = n_2961 ^ n_11330;
assign n_11431 = n_3030 ^ n_11331;
assign n_11432 = n_3096 ^ n_11332;
assign n_11433 = n_3165 ^ n_11333;
assign n_11434 = n_3229 ^ n_11334;
assign n_11435 = n_3294 ^ n_11335;
assign n_11436 = n_3359 ^ n_11336;
assign n_11437 = n_11337 ^ n_2063;
assign n_11438 = n_11338 ^ x5;
assign n_11439 = n_11339 ^ x8;
assign n_11440 = n_11340 ^ x11;
assign n_11441 = n_11341 ^ x14;
assign n_11442 = n_11342 ^ x17;
assign n_11443 = n_11343 ^ x20;
assign n_11444 = n_11344 ^ x23;
assign n_11445 = n_11345 ^ x26;
assign n_11446 = n_11346 ^ x29;
assign n_11447 = n_11347 ^ x32;
assign n_11448 = n_11348 ^ x35;
assign n_11449 = n_11349 ^ x38;
assign n_11450 = n_11350 ^ x41;
assign n_11451 = n_11351 ^ x44;
assign n_11452 = n_11352 ^ x47;
assign n_11453 = n_11353 ^ x50;
assign n_11454 = n_11354 ^ x53;
assign n_11455 = n_11355 ^ x56;
assign n_11456 = n_11356 ^ x59;
assign n_11457 = n_11357 ^ x62;
assign n_11458 = n_11141 ^ n_11358;
assign n_11459 = n_11359 ^ n_11358;
assign n_11460 = n_11360 ^ n_11174;
assign n_11461 = n_11363 ^ n_11180;
assign n_11462 = n_11364 ^ n_10717;
assign n_11463 = n_11364 ^ n_10590;
assign n_11464 = n_11365 ^ n_10719;
assign n_11465 = n_11365 ^ n_10592;
assign n_11466 = n_11366 ^ n_10360;
assign n_11467 = n_11366 ^ n_10223;
assign n_11468 = n_11367 ^ n_10723;
assign n_11469 = n_11367 ^ n_10596;
assign n_11470 = n_11368 ^ n_10598;
assign n_11471 = n_11369 ^ n_8366;
assign n_11472 = n_11370 ^ n_10602;
assign n_11473 = n_11370 & ~n_10728;
assign n_11474 = n_11371 ^ n_8368;
assign n_11475 = n_11372 ^ n_10350;
assign n_11476 = n_11374 ^ n_11200;
assign n_11477 = n_11376 ^ n_11201;
assign n_11478 = n_11377 ^ n_11202;
assign n_11479 = n_11378 ^ n_10835;
assign n_11480 = n_11378 ^ n_10733;
assign n_11481 = n_11379 ^ n_11005;
assign n_11482 = n_11379 ^ n_10919;
assign n_11483 = n_11380 ^ n_10743;
assign n_11484 = n_11380 ^ n_10615;
assign n_11485 = n_11381 ^ n_11011;
assign n_11486 = n_11381 ^ n_10925;
assign n_11487 = n_11383 ^ n_10620;
assign n_11488 = n_11383 ^ n_10300;
assign n_11489 = n_11384 ^ n_8916;
assign n_11490 = n_10730 & ~n_11385;
assign n_11491 = n_11392 ^ n_11231;
assign n_11492 = ~x0 & n_11393;
assign n_11493 = n_11394 ^ n_3494;
assign n_11494 = n_11395 ^ x100;
assign n_11495 = n_1 & ~n_11396;
assign n_11496 = n_11396 ^ x101;
assign n_11497 = n_2155 ^ n_11397;
assign n_11498 = n_755 ^ n_11398;
assign n_11499 = n_2226 ^ n_11399;
assign n_11500 = n_2294 ^ n_11400;
assign n_11501 = n_2361 ^ n_11401;
assign n_11502 = n_2428 ^ n_11402;
assign n_11503 = n_2495 ^ n_11403;
assign n_11504 = n_2561 ^ n_11404;
assign n_11505 = n_2626 ^ n_11405;
assign n_11506 = n_2693 ^ n_11406;
assign n_11507 = n_2761 ^ n_11407;
assign n_11508 = n_2828 ^ n_11408;
assign n_11509 = n_2896 ^ n_11409;
assign n_11510 = n_2962 ^ n_11410;
assign n_11511 = n_3031 ^ n_11411;
assign n_11512 = n_3097 ^ n_11412;
assign n_11513 = n_3166 ^ n_11413;
assign n_11514 = n_3230 ^ n_11414;
assign n_11515 = n_3295 ^ n_11415;
assign n_11516 = n_3360 ^ n_11416;
assign n_11517 = n_5027 ^ n_11417;
assign n_11518 = n_5090 ^ n_11418;
assign n_11519 = n_5153 ^ n_11419;
assign n_11520 = n_5214 ^ n_11420;
assign n_11521 = n_5278 ^ n_11421;
assign n_11522 = n_5342 ^ n_11422;
assign n_11523 = n_5406 ^ n_11423;
assign n_11524 = n_5470 ^ n_11424;
assign n_11525 = n_5531 ^ n_11425;
assign n_11526 = n_5594 ^ n_11426;
assign n_11527 = n_5657 ^ n_11427;
assign n_11528 = n_5721 ^ n_11428;
assign n_11529 = n_5787 ^ n_11429;
assign n_11530 = n_5849 ^ n_11430;
assign n_11531 = n_5913 ^ n_11431;
assign n_11532 = n_5976 ^ n_11432;
assign n_11533 = n_6040 ^ n_11433;
assign n_11534 = n_6104 ^ n_11434;
assign n_11535 = n_6166 ^ n_11435;
assign n_11536 = n_6228 ^ n_11436;
assign n_11537 = n_11437 ^ n_225;
assign n_11538 = n_11450 ^ n_10983;
assign n_11539 = n_11451 ^ n_10984;
assign n_11540 = n_11452 ^ n_10985;
assign n_11541 = n_11453 ^ n_11261;
assign n_11542 = n_11453 ^ n_11177;
assign n_11543 = n_11454 ^ n_10986;
assign n_11544 = n_11455 ^ n_10987;
assign n_11545 = n_11456 ^ n_10900;
assign n_11546 = n_11457 ^ n_6530;
assign n_11547 = n_11359 & n_11458;
assign n_11548 = n_10986 ^ n_11460;
assign n_11549 = n_11461 ^ n_10739;
assign n_11550 = n_11461 ^ n_10611;
assign n_11551 = n_11462 ^ n_8906;
assign n_11552 = ~n_10717 & n_11463;
assign n_11553 = n_11464 ^ n_8907;
assign n_11554 = ~n_10719 & n_11465;
assign n_11555 = n_11466 ^ n_8908;
assign n_11556 = ~n_10360 & n_11467;
assign n_11557 = n_11468 ^ n_8911;
assign n_11558 = ~n_10723 & n_11469;
assign n_11559 = n_11470 ^ n_8365;
assign n_11560 = ~n_11470 & n_10725;
assign n_11561 = n_11471 ^ n_10473;
assign n_11562 = n_11471 & ~n_10600;
assign n_11563 = n_11472 ^ n_8914;
assign n_11564 = n_11473 ^ n_11277;
assign n_11565 = n_11474 ^ n_10488;
assign n_11566 = n_11474 & n_10618;
assign n_11567 = n_11475 ^ n_8370;
assign n_11568 = n_11475 & ~n_10478;
assign n_11569 = n_11476 ^ n_10842;
assign n_11570 = n_11476 ^ n_10745;
assign n_11571 = n_11477 ^ n_10822;
assign n_11572 = n_11477 ^ n_10713;
assign n_11573 = n_11478 ^ n_10737;
assign n_11574 = n_11478 ^ n_10609;
assign n_11575 = n_11479 ^ n_9122;
assign n_11576 = ~n_10835 & n_11480;
assign n_11577 = n_11481 ^ n_9046;
assign n_11578 = ~n_11005 & n_11482;
assign n_11579 = n_11483 ^ n_9050;
assign n_11580 = ~n_10743 & n_11484;
assign n_11581 = n_11485 ^ n_9051;
assign n_11582 = ~n_11011 & n_11486;
assign n_11583 = n_11487 ^ n_10790;
assign n_11584 = n_10620 & n_11488;
assign n_11585 = n_11490 ^ n_11297;
assign n_11586 = n_11492 ^ n_11312;
assign n_11587 = ~x0 & n_11493;
assign n_11588 = n_11494 ^ n_2109;
assign n_11589 = n_11495 ^ x1;
assign n_11590 = n_655 & n_11496;
assign n_11591 = n_784 & n_11496;
assign n_11592 = ~n_3665 & n_11496;
assign n_11593 = n_854 & n_11496;
assign n_11594 = n_920 & n_11496;
assign n_11595 = n_986 & n_11496;
assign n_11596 = n_1052 & n_11496;
assign n_11597 = n_1117 & n_11496;
assign n_11598 = n_1181 & n_11496;
assign n_11599 = n_1248 & n_11496;
assign n_11600 = n_1314 & n_11496;
assign n_11601 = n_1380 & n_11496;
assign n_11602 = n_11496 & n_1445;
assign n_11603 = n_11496 & n_1510;
assign n_11604 = n_11496 & n_1576;
assign n_11605 = n_11496 & n_1641;
assign n_11606 = n_11496 & n_1706;
assign n_11607 = n_11496 & n_1771;
assign n_11608 = n_11496 & n_1835;
assign n_11609 = n_11496 & n_1899;
assign n_11610 = n_5028 ^ n_11497;
assign n_11611 = n_5091 ^ n_11498;
assign n_11612 = n_5154 ^ n_11499;
assign n_11613 = n_5215 ^ n_11500;
assign n_11614 = n_5279 ^ n_11501;
assign n_11615 = n_5343 ^ n_11502;
assign n_11616 = n_5407 ^ n_11503;
assign n_11617 = n_5471 ^ n_11504;
assign n_11618 = n_5532 ^ n_11505;
assign n_11619 = n_5595 ^ n_11506;
assign n_11620 = n_5658 ^ n_11507;
assign n_11621 = n_5722 ^ n_11508;
assign n_11622 = n_5788 ^ n_11509;
assign n_11623 = n_5850 ^ n_11510;
assign n_11624 = n_5914 ^ n_11511;
assign n_11625 = n_5977 ^ n_11512;
assign n_11626 = n_6041 ^ n_11513;
assign n_11627 = n_6105 ^ n_11514;
assign n_11628 = n_6167 ^ n_11515;
assign n_11629 = n_6229 ^ n_11516;
assign n_11630 = n_11517 ^ x5;
assign n_11631 = n_11518 ^ x8;
assign n_11632 = n_11519 ^ x11;
assign n_11633 = n_11520 ^ x14;
assign n_11634 = n_11521 ^ x17;
assign n_11635 = n_11522 ^ x20;
assign n_11636 = n_11523 ^ x23;
assign n_11637 = n_11524 ^ x26;
assign n_11638 = n_11525 ^ x29;
assign n_11639 = n_11526 ^ x32;
assign n_11640 = n_11527 ^ x35;
assign n_11641 = n_11528 ^ x38;
assign n_11642 = n_11529 ^ x41;
assign n_11643 = n_11530 ^ x44;
assign n_11644 = n_11531 ^ x47;
assign n_11645 = n_11532 ^ x50;
assign n_11646 = n_11533 ^ x53;
assign n_11647 = n_11534 ^ x56;
assign n_11648 = n_11535 ^ x59;
assign n_11649 = n_11536 ^ x62;
assign n_11650 = n_11537 ^ n_220;
assign n_11651 = n_11299 ^ n_11538;
assign n_11652 = n_11538 & ~n_11386;
assign n_11653 = n_11539 ^ n_11079;
assign n_11654 = ~n_11539 & n_11171;
assign n_11655 = n_11540 ^ n_11117;
assign n_11656 = n_11540 & ~n_11217;
assign n_11657 = n_11389 ^ n_11541;
assign n_11658 = ~n_11261 & n_11542;
assign n_11659 = n_11543 ^ n_11460;
assign n_11660 = n_11544 ^ n_11042;
assign n_11661 = ~n_11544 & n_11118;
assign n_11662 = n_11545 ^ n_10990;
assign n_11663 = ~n_11545 & n_11076;
assign n_11664 = n_11546 ^ n_3406;
assign n_11665 = n_11546 & n_6640;
assign n_11666 = n_11547 ^ n_11358;
assign n_11667 = ~n_11543 & n_11548;
assign n_11668 = n_11549 ^ n_9045;
assign n_11669 = ~n_10739 & n_11550;
assign n_11670 = n_11552 ^ n_11364;
assign n_11671 = n_11554 ^ n_11365;
assign n_11672 = n_11556 ^ n_11366;
assign n_11673 = n_11558 ^ n_11367;
assign n_11674 = n_11559 ^ n_8912;
assign n_11675 = n_11560 ^ n_11368;
assign n_11676 = n_11561 ^ n_8913;
assign n_11677 = n_11562 ^ n_11369;
assign n_11678 = n_11564 ^ n_11098;
assign n_11679 = n_11564 ^ n_11019;
assign n_11680 = n_11565 ^ n_8915;
assign n_11681 = n_11566 ^ n_11371;
assign n_11682 = n_11567 ^ n_8917;
assign n_11683 = n_11568 ^ n_11372;
assign n_11684 = n_11569 ^ n_9906;
assign n_11685 = n_10842 & ~n_11570;
assign n_11686 = n_11571 ^ n_9044;
assign n_11687 = ~n_10822 & n_11572;
assign y16 = n_11573;
assign n_11688 = ~n_10737 & n_11574;
assign n_11689 = n_11576 ^ n_11378;
assign n_11690 = n_11578 ^ n_11379;
assign n_11691 = n_11580 ^ n_11380;
assign n_11692 = n_11582 ^ n_11381;
assign n_11693 = n_11584 ^ n_11383;
assign n_11694 = n_11585 ^ n_11100;
assign n_11695 = n_11585 ^ n_11021;
assign n_11696 = n_11587 ^ n_11394;
assign n_11697 = ~x0 & n_11588;
assign n_11698 = n_11589 ^ x101;
assign n_11699 = n_2156 ^ n_11590;
assign n_11700 = n_756 ^ n_11591;
assign n_11701 = n_2227 ^ n_11592;
assign n_11702 = n_2295 ^ n_11593;
assign n_11703 = n_2362 ^ n_11594;
assign n_11704 = n_2429 ^ n_11595;
assign n_11705 = n_2496 ^ n_11596;
assign n_11706 = n_2562 ^ n_11597;
assign n_11707 = n_2627 ^ n_11598;
assign n_11708 = n_2694 ^ n_11599;
assign n_11709 = n_2762 ^ n_11600;
assign n_11710 = n_2829 ^ n_11601;
assign n_11711 = n_2897 ^ n_11602;
assign n_11712 = n_2963 ^ n_11603;
assign n_11713 = n_3032 ^ n_11604;
assign n_11714 = n_3098 ^ n_11605;
assign n_11715 = n_3167 ^ n_11606;
assign n_11716 = n_3231 ^ n_11607;
assign n_11717 = n_3296 ^ n_11608;
assign n_11718 = n_3361 ^ n_11609;
assign n_11719 = n_11610 ^ x5;
assign n_11720 = n_11611 ^ x8;
assign n_11721 = n_11612 ^ x11;
assign n_11722 = n_11613 ^ x14;
assign n_11723 = n_11614 ^ x17;
assign n_11724 = n_11615 ^ x20;
assign n_11725 = n_11616 ^ x23;
assign n_11726 = n_11617 ^ x26;
assign n_11727 = n_11618 ^ x29;
assign n_11728 = n_11619 ^ x32;
assign n_11729 = n_11620 ^ x35;
assign n_11730 = n_11621 ^ x38;
assign n_11731 = n_11622 ^ x41;
assign n_11732 = n_11623 ^ x44;
assign n_11733 = n_11624 ^ x47;
assign n_11734 = n_11625 ^ x50;
assign n_11735 = n_11626 ^ x53;
assign n_11736 = n_11627 ^ x56;
assign n_11737 = n_11628 ^ x59;
assign n_11738 = n_11629 ^ x62;
assign n_11739 = n_11642 ^ n_11175;
assign n_11740 = n_11642 ^ n_11043;
assign n_11741 = n_11643 ^ n_11045;
assign n_11742 = n_11644 ^ n_11083;
assign n_11743 = n_11645 ^ n_11262;
assign n_11744 = n_11646 ^ n_11077;
assign n_11745 = n_11647 ^ n_10960;
assign n_11746 = n_11648 ^ n_11230;
assign n_11747 = n_11648 ^ n_11145;
assign n_11748 = n_224 & n_11650;
assign n_11749 = n_11652 ^ n_11450;
assign n_11750 = n_11387 ^ n_11653;
assign n_11751 = n_11654 ^ n_11451;
assign n_11752 = n_11388 ^ n_11655;
assign n_11753 = n_11656 ^ n_11452;
assign n_11754 = n_11658 ^ n_11453;
assign n_11755 = n_11390 ^ n_11660;
assign n_11756 = n_11661 ^ n_11455;
assign n_11757 = n_11391 ^ n_11662;
assign n_11758 = n_11663 ^ n_11456;
assign n_11759 = n_11664 ^ n_11491;
assign n_11760 = n_11665 ^ n_11457;
assign n_11761 = n_11659 ^ n_11666;
assign n_11762 = n_11667 ^ n_11454;
assign n_11763 = n_11669 ^ n_11461;
assign n_11764 = n_11670 ^ n_11007;
assign n_11765 = n_11670 ^ n_10921;
assign n_11766 = n_11671 ^ n_11009;
assign n_11767 = n_11671 ^ n_10923;
assign n_11768 = n_11672 ^ n_10741;
assign n_11769 = n_11672 ^ n_10613;
assign n_11770 = n_11673 ^ n_11093;
assign n_11771 = n_11673 ^ n_11013;
assign n_11772 = n_11675 ^ n_11015;
assign n_11773 = n_11675 ^ n_10928;
assign n_11774 = n_11677 ^ n_11017;
assign n_11775 = n_11677 ^ n_10930;
assign n_11776 = n_11678 ^ n_9055;
assign n_11777 = ~n_11098 & n_11679;
assign n_11778 = n_11681 ^ n_10946;
assign n_11779 = n_11681 ^ n_10844;
assign n_11780 = n_11683 ^ n_10934;
assign n_11781 = n_11683 ^ n_10833;
assign n_11782 = n_11685 ^ n_11476;
assign n_11783 = n_11687 ^ n_11477;
assign n_11784 = n_11688 ^ n_11478;
assign n_11785 = n_11689 ^ n_11104;
assign n_11786 = n_11689 ^ n_11024;
assign n_11787 = n_11690 ^ n_11265;
assign n_11788 = n_11690 ^ n_11181;
assign n_11789 = n_11691 ^ n_11034;
assign n_11790 = n_11691 ^ n_10943;
assign n_11791 = n_11692 ^ n_11271;
assign n_11792 = n_11692 ^ n_11187;
assign n_11793 = n_11693 ^ n_10955;
assign n_11794 = n_11693 ^ n_10866;
assign n_11795 = n_11694 ^ n_9057;
assign n_11796 = ~n_11100 & n_11695;
assign n_11797 = n_11697 ^ n_11494;
assign n_11798 = n_11698 ^ n_6486;
assign n_11799 = n_5029 ^ n_11699;
assign n_11800 = n_5092 ^ n_11700;
assign n_11801 = n_5155 ^ n_11701;
assign n_11802 = n_5216 ^ n_11702;
assign n_11803 = n_5280 ^ n_11703;
assign n_11804 = n_5344 ^ n_11704;
assign n_11805 = n_5408 ^ n_11705;
assign n_11806 = n_5472 ^ n_11706;
assign n_11807 = n_5533 ^ n_11707;
assign n_11808 = n_5596 ^ n_11708;
assign n_11809 = n_5659 ^ n_11709;
assign n_11810 = n_5723 ^ n_11710;
assign n_11811 = n_5789 ^ n_11711;
assign n_11812 = n_5851 ^ n_11712;
assign n_11813 = n_5915 ^ n_11713;
assign n_11814 = n_5978 ^ n_11714;
assign n_11815 = n_6042 ^ n_11715;
assign n_11816 = n_6106 ^ n_11716;
assign n_11817 = n_6168 ^ n_11717;
assign n_11818 = n_6230 ^ n_11718;
assign n_11819 = n_11731 ^ n_11300;
assign n_11820 = n_11732 ^ n_11302;
assign n_11821 = n_11733 ^ n_11304;
assign n_11822 = n_11734 ^ n_11459;
assign n_11823 = n_11735 ^ n_11306;
assign n_11824 = n_11736 ^ n_11308;
assign n_11825 = n_11737 ^ n_11310;
assign n_11826 = n_11738 ^ n_6410;
assign n_11827 = ~n_11175 & n_11740;
assign n_11828 = n_11741 ^ n_11116;
assign n_11829 = n_11741 & ~n_11216;
assign n_11830 = n_11742 ^ n_11047;
assign n_11831 = n_11742 & n_11176;
assign n_11832 = n_11743 ^ n_11257;
assign n_11833 = n_11743 & ~n_11361;
assign n_11834 = n_11744 ^ n_11049;
assign n_11835 = n_11744 & n_11169;
assign n_11836 = n_11745 ^ n_11078;
assign n_11837 = n_11745 & ~n_11170;
assign n_11838 = ~n_11230 & n_11747;
assign n_11839 = n_11748 ^ x100;
assign n_11840 = n_11749 ^ n_11739;
assign n_11841 = n_11758 ^ n_11746;
assign n_11842 = n_11760 ^ n_6753;
assign n_11843 = ~n_6276 & ~n_11760;
assign n_11844 = n_11763 ^ n_11030;
assign n_11845 = n_11763 ^ n_10940;
assign n_11846 = n_11764 ^ n_9047;
assign n_11847 = ~n_11007 & n_11765;
assign n_11848 = n_11766 ^ n_9048;
assign n_11849 = ~n_11009 & n_11767;
assign n_11850 = n_11768 ^ n_9049;
assign n_11851 = ~n_10741 & n_11769;
assign n_11852 = n_11770 ^ n_9052;
assign n_11853 = ~n_11093 & n_11771;
assign n_11854 = n_11772 ^ n_9053;
assign n_11855 = ~n_11015 & n_11773;
assign n_11856 = n_11774 ^ n_9054;
assign n_11857 = ~n_11017 & n_11775;
assign n_11858 = n_11777 ^ n_11564;
assign n_11859 = n_11778 ^ n_9056;
assign n_11860 = ~n_10946 & n_11779;
assign n_11861 = n_11780 ^ n_9058;
assign n_11862 = ~n_10934 & n_11781;
assign n_11863 = n_11782 ^ n_11112;
assign n_11864 = n_11782 ^ n_11036;
assign n_11865 = n_11783 ^ n_11087;
assign n_11866 = n_11783 ^ n_11003;
assign n_11867 = n_11784 ^ n_11028;
assign n_11868 = n_11784 ^ n_10938;
assign n_11869 = n_11785 ^ n_9256;
assign n_11870 = ~n_11104 & n_11786;
assign n_11871 = n_11787 ^ n_9192;
assign n_11872 = n_11265 & ~n_11788;
assign n_11873 = n_11789 ^ n_9196;
assign n_11874 = ~n_11034 & n_11790;
assign n_11875 = n_11791 ^ n_9197;
assign n_11876 = ~n_11271 & n_11792;
assign n_11877 = n_11793 ^ n_11641;
assign n_11878 = n_10955 & n_11794;
assign n_11879 = n_11796 ^ n_11585;
assign n_11880 = ~x0 & ~n_11798;
assign n_11881 = n_11799 ^ x5;
assign n_11882 = n_11800 ^ x8;
assign n_11883 = n_11801 ^ x11;
assign n_11884 = n_11802 ^ x14;
assign n_11885 = n_11803 ^ x17;
assign n_11886 = n_11804 ^ x20;
assign n_11887 = n_11805 ^ x23;
assign n_11888 = n_11806 ^ x26;
assign n_11889 = n_11807 ^ x29;
assign n_11890 = n_11808 ^ x32;
assign n_11891 = n_11809 ^ x35;
assign n_11892 = n_11810 ^ x38;
assign n_11893 = n_11811 ^ x41;
assign n_11894 = n_11812 ^ x44;
assign n_11895 = n_11813 ^ x47;
assign n_11896 = n_11814 ^ x50;
assign n_11897 = n_11815 ^ x53;
assign n_11898 = n_11816 ^ x56;
assign n_11899 = n_11817 ^ x59;
assign n_11900 = n_11818 ^ x62;
assign n_11901 = n_11827 ^ n_11642;
assign n_11902 = n_11828 ^ n_11751;
assign n_11903 = n_11829 ^ n_11643;
assign n_11904 = n_11830 ^ n_11753;
assign n_11905 = n_11831 ^ n_11644;
assign n_11906 = n_11832 ^ n_11754;
assign n_11907 = n_11833 ^ n_11645;
assign n_11908 = n_11762 ^ n_11834;
assign n_11909 = n_11835 ^ n_11646;
assign n_11910 = n_11836 ^ n_11756;
assign n_11911 = n_11837 ^ n_11647;
assign n_11912 = n_11838 ^ n_11648;
assign n_11913 = n_11839 ^ x101;
assign n_11914 = ~x101 & ~n_11839;
assign n_11915 = n_11842 ^ n_11649;
assign n_11916 = ~n_6409 & ~n_11843;
assign n_11917 = n_11844 ^ n_9191;
assign n_11918 = ~n_11030 & n_11845;
assign n_11919 = n_11847 ^ n_11670;
assign n_11920 = n_11849 ^ n_11671;
assign n_11921 = n_11851 ^ n_11672;
assign n_11922 = n_11853 ^ n_11673;
assign n_11923 = n_11855 ^ n_11675;
assign n_11924 = n_11857 ^ n_11677;
assign n_11925 = n_11858 ^ n_11195;
assign n_11926 = n_11858 ^ n_8786;
assign n_11927 = n_11860 ^ n_11681;
assign n_11928 = n_11862 ^ n_11683;
assign n_11929 = n_11863 ^ n_10386;
assign n_11930 = ~n_11112 & n_11864;
assign n_11931 = n_11865 ^ n_9190;
assign n_11932 = ~n_11087 & n_11866;
assign y17 = n_11867;
assign n_11933 = ~n_11028 & n_11868;
assign n_11934 = n_11870 ^ n_11689;
assign n_11935 = n_11872 ^ n_11690;
assign n_11936 = n_11874 ^ n_11691;
assign n_11937 = n_11876 ^ n_11692;
assign n_11938 = n_11878 ^ n_11693;
assign n_11939 = n_11879 ^ n_11197;
assign n_11940 = n_11879 ^ n_8788;
assign n_11941 = n_11880 ^ n_11698;
assign n_11942 = n_11892 ^ n_11651;
assign n_11943 = n_11893 ^ n_11750;
assign n_11944 = n_11893 ^ n_11387;
assign n_11945 = n_11894 ^ n_11388;
assign n_11946 = n_11895 ^ n_11657;
assign n_11947 = n_11895 ^ n_11389;
assign n_11948 = n_11896 ^ n_11659;
assign n_11949 = n_11897 ^ n_11390;
assign n_11950 = n_11898 ^ n_11391;
assign n_11951 = n_11899 ^ n_11664;
assign n_11952 = n_11900 ^ n_6532;
assign n_11953 = n_11901 ^ n_11819;
assign n_11954 = n_11901 ^ n_11731;
assign n_11955 = n_11903 ^ n_11820;
assign n_11956 = n_11903 ^ n_11732;
assign n_11957 = n_11905 ^ n_11821;
assign n_11958 = n_11905 ^ n_11733;
assign n_11959 = n_11907 ^ n_11734;
assign n_11960 = n_11909 ^ n_11735;
assign n_11961 = n_11911 ^ n_11824;
assign n_11962 = n_11911 ^ n_11736;
assign n_11963 = n_11912 ^ n_11737;
assign n_11964 = n_1 & ~n_11913;
assign n_11965 = n_11913 ^ x102;
assign n_11966 = x102 & ~n_11914;
assign n_11967 = n_11914 ^ n_11913;
assign n_11968 = n_11916 ^ n_11826;
assign n_11969 = n_11916 ^ n_11738;
assign n_11970 = n_11918 ^ n_11763;
assign n_11971 = n_11919 ^ n_11267;
assign n_11972 = n_11919 ^ n_11183;
assign n_11973 = n_11920 ^ n_11269;
assign n_11974 = n_11920 ^ n_11185;
assign n_11975 = n_11921 ^ n_8780;
assign n_11976 = n_11922 ^ n_11273;
assign n_11977 = n_11922 ^ n_11189;
assign n_11978 = n_11923 ^ n_11275;
assign n_11979 = n_11923 ^ n_11191;
assign n_11980 = n_11924 ^ n_11096;
assign n_11981 = n_11925 ^ n_9201;
assign n_11982 = ~n_11195 & n_11926;
assign n_11983 = n_11927 ^ n_11296;
assign n_11984 = n_11927 ^ n_11212;
assign n_11985 = n_11928 ^ n_11199;
assign n_11986 = n_11928 ^ n_11102;
assign n_11987 = n_11930 ^ n_11782;
assign n_11988 = n_11932 ^ n_11783;
assign n_11989 = n_11933 ^ n_11784;
assign n_11990 = n_11934 ^ n_11375;
assign n_11991 = n_11934 ^ n_11282;
assign n_11992 = n_11935 ^ n_11551;
assign n_11993 = n_11935 ^ n_11462;
assign n_11994 = n_11936 ^ n_11292;
assign n_11995 = n_11936 ^ n_11209;
assign n_11996 = n_11937 ^ n_11557;
assign n_11997 = n_11937 ^ n_11468;
assign n_11998 = n_11938 ^ n_11298;
assign n_11999 = n_11938 ^ n_11137;
assign n_12000 = n_11939 ^ n_9203;
assign n_12001 = ~n_11197 & n_11940;
assign n_12002 = n_11750 & n_11944;
assign n_12003 = n_11945 ^ n_11655;
assign n_12004 = n_11945 & ~n_11752;
assign n_12005 = ~n_11657 & n_11947;
assign n_12006 = n_11948 ^ n_11666;
assign n_12007 = ~n_11948 & n_11761;
assign n_12008 = n_11949 ^ n_11660;
assign n_12009 = n_11949 & n_11755;
assign n_12010 = n_11950 ^ n_11662;
assign n_12011 = n_11950 & n_11757;
assign n_12012 = n_11951 ^ n_11491;
assign n_12013 = ~n_11951 & ~n_11759;
assign n_12014 = n_11952 ^ n_3409;
assign n_12015 = n_11952 & n_6642;
assign n_12016 = ~n_11819 & n_11954;
assign n_12017 = ~n_11820 & n_11956;
assign n_12018 = n_11821 & n_11958;
assign n_12019 = n_11959 ^ n_11459;
assign n_12020 = n_11959 & n_11822;
assign n_12021 = n_11960 ^ n_11306;
assign n_12022 = n_11960 & n_11823;
assign n_12023 = n_11824 & n_11962;
assign n_12024 = n_11963 ^ n_11310;
assign n_12025 = n_11963 & ~n_11825;
assign n_12026 = n_11964 ^ x1;
assign n_12027 = n_655 & n_11965;
assign n_12028 = n_784 & n_11965;
assign n_12029 = ~n_3665 & n_11965;
assign n_12030 = n_854 & n_11965;
assign n_12031 = n_920 & n_11965;
assign n_12032 = n_986 & n_11965;
assign n_12033 = n_1052 & n_11965;
assign n_12034 = n_1117 & n_11965;
assign n_12035 = n_1181 & n_11965;
assign n_12036 = n_1248 & n_11965;
assign n_12037 = n_1314 & n_11965;
assign n_12038 = n_1380 & n_11965;
assign n_12039 = n_11965 & n_1445;
assign n_12040 = n_11965 & n_1510;
assign n_12041 = n_11965 & n_1576;
assign n_12042 = n_11965 & n_1641;
assign n_12043 = n_11965 & n_1706;
assign n_12044 = n_11965 & n_1771;
assign n_12045 = n_11965 & n_1835;
assign n_12046 = n_11965 & n_1899;
assign n_12047 = ~x103 & ~n_11966;
assign n_12048 = ~x102 & n_11967;
assign n_12049 = n_11826 & n_11969;
assign n_12050 = n_11970 ^ n_11288;
assign n_12051 = n_11970 ^ n_11205;
assign n_12052 = n_11971 ^ n_9193;
assign n_12053 = ~n_11267 & n_11972;
assign n_12054 = n_11973 ^ n_9194;
assign n_12055 = ~n_11269 & n_11974;
assign n_12056 = n_11975 ^ n_11032;
assign n_12057 = n_11975 & ~n_11109;
assign n_12058 = n_11976 ^ n_9198;
assign n_12059 = n_11273 & ~n_11977;
assign n_12060 = n_11978 ^ n_9199;
assign n_12061 = ~n_11275 & n_11979;
assign n_12062 = n_11980 ^ n_8785;
assign n_12063 = n_11980 & ~n_11193;
assign n_12064 = n_11982 ^ n_11858;
assign n_12065 = n_11983 ^ n_9202;
assign n_12066 = ~n_11296 & n_11984;
assign n_12067 = n_11985 ^ n_9204;
assign n_12068 = ~n_11199 & n_11986;
assign n_12069 = n_11987 ^ n_11382;
assign n_12070 = n_11987 ^ n_11294;
assign n_12071 = n_11988 ^ n_11362;
assign n_12072 = n_11988 ^ n_11263;
assign n_12073 = n_11989 ^ n_11286;
assign n_12074 = n_11989 ^ n_11203;
assign n_12075 = n_11990 ^ n_9401;
assign n_12076 = ~n_11375 & n_11991;
assign n_12077 = n_11992 ^ n_9326;
assign n_12078 = ~n_11551 & n_11993;
assign n_12079 = n_11994 ^ n_9330;
assign n_12080 = n_11292 & ~n_11995;
assign n_12081 = n_11996 ^ n_9331;
assign n_12082 = ~n_11557 & n_11997;
assign n_12083 = n_11998 ^ n_11730;
assign n_12084 = ~n_11298 & n_11999;
assign n_12085 = n_12001 ^ n_11879;
assign n_12086 = n_12002 ^ n_11893;
assign n_12087 = n_12004 ^ n_11894;
assign n_12088 = n_12005 ^ n_11895;
assign n_12089 = n_12007 ^ n_11896;
assign n_12090 = n_12009 ^ n_11897;
assign n_12091 = n_12011 ^ n_11898;
assign n_12092 = n_12013 ^ n_11899;
assign n_12093 = n_12015 ^ n_11900;
assign n_12094 = n_12016 ^ n_11901;
assign n_12095 = n_12017 ^ n_11903;
assign n_12096 = n_12018 ^ n_11905;
assign n_12097 = n_12020 ^ n_11907;
assign n_12098 = n_12022 ^ n_11909;
assign n_12099 = n_12023 ^ n_11911;
assign n_12100 = n_12025 ^ n_11912;
assign n_12101 = n_12026 ^ x102;
assign n_12102 = n_2157 ^ n_12027;
assign n_12103 = n_757 ^ n_12028;
assign n_12104 = n_2228 ^ n_12029;
assign n_12105 = n_2296 ^ n_12030;
assign n_12106 = n_2363 ^ n_12031;
assign n_12107 = n_2430 ^ n_12032;
assign n_12108 = n_2497 ^ n_12033;
assign n_12109 = n_2563 ^ n_12034;
assign n_12110 = n_2628 ^ n_12035;
assign n_12111 = n_2695 ^ n_12036;
assign n_12112 = n_2763 ^ n_12037;
assign n_12113 = n_2830 ^ n_12038;
assign n_12114 = n_2898 ^ n_12039;
assign n_12115 = n_2964 ^ n_12040;
assign n_12116 = n_3033 ^ n_12041;
assign n_12117 = n_3099 ^ n_12042;
assign n_12118 = n_3168 ^ n_12043;
assign n_12119 = n_3232 ^ n_12044;
assign n_12120 = n_3297 ^ n_12045;
assign n_12121 = n_3362 ^ n_12046;
assign n_12122 = x104 & ~n_12047;
assign n_12123 = n_11966 ^ n_12048;
assign n_12124 = x103 & ~n_12048;
assign n_12125 = n_12049 ^ n_11916;
assign n_12126 = n_12050 ^ n_9325;
assign n_12127 = n_11288 & ~n_12051;
assign n_12128 = n_12053 ^ n_11919;
assign n_12129 = n_12055 ^ n_11920;
assign n_12130 = n_12056 ^ n_9195;
assign n_12131 = n_12057 ^ n_11921;
assign n_12132 = n_12059 ^ n_11922;
assign n_12133 = n_12061 ^ n_11923;
assign n_12134 = n_12062 ^ n_9200;
assign n_12135 = n_12063 ^ n_11924;
assign n_12136 = n_12064 ^ n_11680;
assign n_12137 = n_12064 ^ n_11565;
assign n_12138 = n_12066 ^ n_11927;
assign n_12139 = n_12068 ^ n_11928;
assign n_12140 = n_12069 ^ n_10687;
assign n_12141 = n_11382 & ~n_12070;
assign n_12142 = n_12071 ^ n_9324;
assign n_12143 = ~n_11362 & n_12072;
assign y18 = n_12073;
assign n_12144 = ~n_11286 & n_12074;
assign n_12145 = n_12076 ^ n_11934;
assign n_12146 = n_12078 ^ n_11935;
assign n_12147 = n_12080 ^ n_11936;
assign n_12148 = n_12082 ^ n_11937;
assign n_12149 = n_12084 ^ n_11938;
assign n_12150 = n_12085 ^ n_11682;
assign n_12151 = n_12085 ^ n_11567;
assign n_12152 = n_12093 ^ n_6754;
assign n_12153 = ~n_6280 & ~n_12093;
assign n_12154 = n_12094 ^ n_11943;
assign n_12155 = n_12095 ^ n_12003;
assign n_12156 = n_12096 ^ n_11946;
assign n_12157 = n_12097 ^ n_12006;
assign n_12158 = n_12098 ^ n_12008;
assign n_12159 = n_12010 ^ n_12099;
assign n_12160 = n_12012 ^ n_12100;
assign n_12161 = n_12101 ^ n_4970;
assign n_12162 = n_5030 ^ n_12102;
assign n_12163 = n_5093 ^ n_12103;
assign n_12164 = n_5156 ^ n_12104;
assign n_12165 = n_5217 ^ n_12105;
assign n_12166 = n_5281 ^ n_12106;
assign n_12167 = n_5345 ^ n_12107;
assign n_12168 = n_5409 ^ n_12108;
assign n_12169 = n_5473 ^ n_12109;
assign n_12170 = n_5534 ^ n_12110;
assign n_12171 = n_5597 ^ n_12111;
assign n_12172 = n_5660 ^ n_12112;
assign n_12173 = n_5724 ^ n_12113;
assign n_12174 = n_5790 ^ n_12114;
assign n_12175 = n_5852 ^ n_12115;
assign n_12176 = n_5916 ^ n_12116;
assign n_12177 = n_5979 ^ n_12117;
assign n_12178 = n_6043 ^ n_12118;
assign n_12179 = n_6107 ^ n_12119;
assign n_12180 = n_6169 ^ n_12120;
assign n_12181 = n_6231 ^ n_12121;
assign n_12182 = ~x105 & ~n_12122;
assign n_12183 = n_1 & n_12123;
assign n_12184 = n_12123 ^ x103;
assign n_12185 = n_12047 ^ n_12124;
assign n_12186 = ~x104 & ~n_12124;
assign n_12187 = n_12014 ^ n_12125;
assign n_12188 = n_12127 ^ n_11970;
assign n_12189 = n_12128 ^ n_11553;
assign n_12190 = n_12128 ^ n_11464;
assign n_12191 = n_12129 ^ n_11555;
assign n_12192 = n_12129 ^ n_11466;
assign n_12193 = n_12131 ^ n_11290;
assign n_12194 = n_12131 ^ n_11207;
assign n_12195 = n_12132 ^ n_11674;
assign n_12196 = n_12132 ^ n_11559;
assign n_12197 = n_12133 ^ n_11676;
assign n_12198 = n_12133 ^ n_11561;
assign n_12199 = n_12135 ^ n_11563;
assign n_12200 = n_12135 ^ n_11472;
assign n_12201 = n_12136 ^ n_9335;
assign n_12202 = n_11680 & ~n_12137;
assign n_12203 = n_12138 ^ n_11489;
assign n_12204 = n_12138 ^ n_11384;
assign n_12205 = n_12139 ^ n_11373;
assign n_12206 = n_12139 ^ n_11280;
assign n_12207 = n_12141 ^ n_11987;
assign n_12208 = n_12143 ^ n_11988;
assign n_12209 = n_12144 ^ n_11989;
assign n_12210 = n_12145 ^ n_11686;
assign n_12211 = n_12145 ^ n_11571;
assign n_12212 = n_12146 ^ n_11846;
assign n_12213 = n_12146 ^ n_11764;
assign n_12214 = n_12147 ^ n_11581;
assign n_12215 = n_12147 ^ n_11485;
assign n_12216 = n_12148 ^ n_11852;
assign n_12217 = n_12148 ^ n_11770;
assign n_12218 = n_12149 ^ n_11942;
assign n_12219 = n_12149 ^ n_11892;
assign n_12220 = n_12150 ^ n_9337;
assign n_12221 = ~n_11682 & n_12151;
assign n_12222 = ~n_6412 & ~n_12153;
assign n_12223 = ~x0 & n_12161;
assign n_12224 = n_12162 ^ x5;
assign n_12225 = n_12163 ^ x8;
assign n_12226 = n_12164 ^ x11;
assign n_12227 = n_12165 ^ x14;
assign n_12228 = n_12166 ^ x17;
assign n_12229 = n_12167 ^ x20;
assign n_12230 = n_12168 ^ x23;
assign n_12231 = n_12169 ^ x26;
assign n_12232 = n_12170 ^ x29;
assign n_12233 = n_12171 ^ x32;
assign n_12234 = n_12172 ^ x35;
assign n_12235 = n_12173 ^ x38;
assign n_12236 = n_12174 ^ x41;
assign n_12237 = n_12175 ^ x44;
assign n_12238 = n_12176 ^ x47;
assign n_12239 = n_12177 ^ x50;
assign n_12240 = n_12178 ^ x53;
assign n_12241 = n_12179 ^ x56;
assign n_12242 = n_12180 ^ x59;
assign n_12243 = n_12181 ^ x62;
assign n_12244 = x106 & ~n_12182;
assign n_12245 = n_12183 ^ x1;
assign n_12246 = n_655 & ~n_12184;
assign n_12247 = n_784 & ~n_12184;
assign n_12248 = ~n_3665 & ~n_12184;
assign n_12249 = n_854 & ~n_12184;
assign n_12250 = n_920 & ~n_12184;
assign n_12251 = n_986 & ~n_12184;
assign n_12252 = n_1052 & ~n_12184;
assign n_12253 = n_1117 & ~n_12184;
assign n_12254 = n_1181 & ~n_12184;
assign n_12255 = n_1248 & ~n_12184;
assign n_12256 = n_1314 & ~n_12184;
assign n_12257 = n_1380 & ~n_12184;
assign n_12258 = n_1445 & ~n_12184;
assign n_12259 = ~n_12184 & n_1510;
assign n_12260 = ~n_12184 & n_1576;
assign n_12261 = ~n_12184 & n_1641;
assign n_12262 = ~n_12184 & n_1706;
assign n_12263 = ~n_12184 & n_1771;
assign n_12264 = ~n_12184 & n_1835;
assign n_12265 = ~n_12184 & n_1899;
assign n_12266 = n_1 & n_12185;
assign n_12267 = n_12185 ^ x104;
assign n_12268 = n_12122 ^ n_12186;
assign n_12269 = x105 & ~n_12186;
assign n_12270 = n_12188 ^ n_11577;
assign n_12271 = n_12188 ^ n_11481;
assign n_12272 = n_12189 ^ n_9327;
assign n_12273 = ~n_11553 & n_12190;
assign n_12274 = n_12191 ^ n_9328;
assign n_12275 = ~n_11555 & n_12192;
assign n_12276 = n_12193 ^ n_9329;
assign n_12277 = ~n_11290 & n_12194;
assign n_12278 = n_12195 ^ n_9332;
assign n_12279 = n_11674 & ~n_12196;
assign n_12280 = n_12197 ^ n_9333;
assign n_12281 = ~n_11676 & n_12198;
assign n_12282 = n_12199 ^ n_9334;
assign n_12283 = ~n_11563 & n_12200;
assign n_12284 = n_12202 ^ n_12064;
assign n_12285 = n_12203 ^ n_9336;
assign n_12286 = n_11489 & ~n_12204;
assign n_12287 = n_12205 ^ n_9764;
assign n_12288 = n_11373 & ~n_12206;
assign n_12289 = n_12207 ^ n_11583;
assign n_12290 = n_12207 ^ n_11487;
assign n_12291 = n_12208 ^ n_11668;
assign n_12292 = n_12208 ^ n_11549;
assign n_12293 = n_12209 ^ n_11575;
assign n_12294 = n_12209 ^ n_11479;
assign n_12295 = n_12210 ^ n_9546;
assign n_12296 = ~n_11686 & n_12211;
assign n_12297 = n_12212 ^ n_9471;
assign n_12298 = ~n_11846 & n_12213;
assign n_12299 = n_12214 ^ n_9475;
assign n_12300 = ~n_11581 & n_12215;
assign n_12301 = n_12216 ^ n_9476;
assign n_12302 = ~n_11852 & n_12217;
assign n_12303 = ~n_11942 & n_12219;
assign n_12304 = n_12221 ^ n_12085;
assign n_12305 = n_12223 ^ n_12101;
assign n_12306 = n_12235 ^ n_11840;
assign n_12307 = n_12235 ^ n_11749;
assign n_12308 = n_12236 ^ n_11902;
assign n_12309 = n_12236 ^ n_11828;
assign n_12310 = n_12237 ^ n_11830;
assign n_12311 = n_12238 ^ n_11906;
assign n_12312 = n_12238 ^ n_11754;
assign n_12313 = n_12239 ^ n_11762;
assign n_12314 = n_12240 ^ n_11836;
assign n_12315 = n_12241 ^ n_11758;
assign n_12316 = n_12242 ^ n_11915;
assign n_12317 = n_12242 ^ n_11649;
assign n_12318 = n_12152 ^ n_12243;
assign n_12319 = n_12245 ^ x103;
assign n_12320 = n_2158 ^ n_12246;
assign n_12321 = n_758 ^ n_12247;
assign n_12322 = n_2229 ^ n_12248;
assign n_12323 = n_2297 ^ n_12249;
assign n_12324 = n_2364 ^ n_12250;
assign n_12325 = n_2431 ^ n_12251;
assign n_12326 = n_2498 ^ n_12252;
assign n_12327 = n_2564 ^ n_12253;
assign n_12328 = n_2629 ^ n_12254;
assign n_12329 = n_2696 ^ n_12255;
assign n_12330 = n_2764 ^ n_12256;
assign n_12331 = n_2831 ^ n_12257;
assign n_12332 = n_2899 ^ n_12258;
assign n_12333 = n_2965 ^ n_12259;
assign n_12334 = n_3034 ^ n_12260;
assign n_12335 = n_3100 ^ n_12261;
assign n_12336 = n_3169 ^ n_12262;
assign n_12337 = n_3233 ^ n_12263;
assign n_12338 = n_3298 ^ n_12264;
assign n_12339 = n_3363 ^ n_12265;
assign n_12340 = n_12266 ^ x1;
assign n_12341 = n_655 & ~n_12267;
assign n_12342 = n_784 & ~n_12267;
assign n_12343 = ~n_3665 & ~n_12267;
assign n_12344 = n_854 & ~n_12267;
assign n_12345 = n_920 & ~n_12267;
assign n_12346 = n_986 & ~n_12267;
assign n_12347 = n_1052 & ~n_12267;
assign n_12348 = n_1117 & ~n_12267;
assign n_12349 = n_1181 & ~n_12267;
assign n_12350 = n_1248 & ~n_12267;
assign n_12351 = n_1314 & ~n_12267;
assign n_12352 = n_1380 & ~n_12267;
assign n_12353 = n_1445 & ~n_12267;
assign n_12354 = ~n_12267 & n_1510;
assign n_12355 = ~n_12267 & n_1576;
assign n_12356 = ~n_12267 & n_1641;
assign n_12357 = ~n_12267 & n_1706;
assign n_12358 = ~n_12267 & n_1771;
assign n_12359 = ~n_12267 & n_1835;
assign n_12360 = ~n_12267 & n_1899;
assign n_12361 = n_1 & n_12268;
assign n_12362 = n_12268 ^ x105;
assign n_12363 = n_12182 ^ n_12269;
assign n_12364 = ~x106 & ~n_12269;
assign n_12365 = n_12270 ^ n_9470;
assign n_12366 = ~n_11577 & n_12271;
assign n_12367 = n_12273 ^ n_12128;
assign n_12368 = n_12275 ^ n_12129;
assign n_12369 = n_12277 ^ n_12131;
assign n_12370 = n_12279 ^ n_12132;
assign n_12371 = n_12281 ^ n_12133;
assign n_12372 = n_12283 ^ n_12135;
assign n_12373 = n_12284 ^ n_11859;
assign n_12374 = n_12284 ^ n_11778;
assign n_12375 = n_12286 ^ n_12138;
assign n_12376 = n_12288 ^ n_12139;
assign n_12377 = n_12289 ^ n_11449;
assign n_12378 = n_11583 & ~n_12290;
assign n_12379 = n_12291 ^ n_9469;
assign n_12380 = ~n_11668 & n_12292;
assign y19 = n_12293;
assign n_12381 = ~n_11575 & n_12294;
assign n_12382 = n_12296 ^ n_12145;
assign n_12383 = n_12298 ^ n_12146;
assign n_12384 = n_12300 ^ n_12147;
assign n_12385 = n_12302 ^ n_12148;
assign n_12386 = n_12303 ^ n_12149;
assign n_12387 = n_12304 ^ n_11861;
assign n_12388 = n_12304 ^ n_11780;
assign n_12389 = ~n_11840 & n_12307;
assign n_12390 = n_12308 ^ n_12086;
assign n_12391 = ~n_11902 & n_12309;
assign n_12392 = n_12310 ^ n_11753;
assign n_12393 = ~n_12310 & n_11904;
assign n_12394 = n_12311 ^ n_12088;
assign n_12395 = n_11906 & ~n_12312;
assign n_12396 = n_12313 ^ n_11834;
assign n_12397 = n_12313 & n_11908;
assign n_12398 = n_12314 ^ n_11756;
assign n_12399 = n_12314 & ~n_11910;
assign n_12400 = n_12315 ^ n_11746;
assign n_12401 = n_12315 & ~n_11841;
assign n_12402 = n_12092 ^ n_12316;
assign n_12403 = ~n_11915 & ~n_12317;
assign n_12404 = n_12319 ^ n_3498;
assign n_12405 = n_5031 ^ n_12320;
assign n_12406 = n_5094 ^ n_12321;
assign n_12407 = n_5157 ^ n_12322;
assign n_12408 = n_5218 ^ n_12323;
assign n_12409 = n_5282 ^ n_12324;
assign n_12410 = n_5346 ^ n_12325;
assign n_12411 = n_5410 ^ n_12326;
assign n_12412 = n_5474 ^ n_12327;
assign n_12413 = n_5535 ^ n_12328;
assign n_12414 = n_5598 ^ n_12329;
assign n_12415 = n_5661 ^ n_12330;
assign n_12416 = n_5725 ^ n_12331;
assign n_12417 = n_5791 ^ n_12332;
assign n_12418 = n_5853 ^ n_12333;
assign n_12419 = n_5917 ^ n_12334;
assign n_12420 = n_5980 ^ n_12335;
assign n_12421 = n_6044 ^ n_12336;
assign n_12422 = n_6108 ^ n_12337;
assign n_12423 = n_6170 ^ n_12338;
assign n_12424 = n_6232 ^ n_12339;
assign n_12425 = n_12340 ^ x104;
assign n_12426 = n_2159 ^ n_12341;
assign n_12427 = n_759 ^ n_12342;
assign n_12428 = n_2230 ^ n_12343;
assign n_12429 = n_2298 ^ n_12344;
assign n_12430 = n_2365 ^ n_12345;
assign n_12431 = n_2432 ^ n_12346;
assign n_12432 = n_2499 ^ n_12347;
assign n_12433 = n_2565 ^ n_12348;
assign n_12434 = n_2630 ^ n_12349;
assign n_12435 = n_2697 ^ n_12350;
assign n_12436 = n_2765 ^ n_12351;
assign n_12437 = n_2832 ^ n_12352;
assign n_12438 = n_2900 ^ n_12353;
assign n_12439 = n_2966 ^ n_12354;
assign n_12440 = n_3035 ^ n_12355;
assign n_12441 = n_3101 ^ n_12356;
assign n_12442 = n_3170 ^ n_12357;
assign n_12443 = n_3234 ^ n_12358;
assign n_12444 = n_3299 ^ n_12359;
assign n_12445 = n_3364 ^ n_12360;
assign n_12446 = n_12361 ^ x1;
assign n_12447 = n_655 & ~n_12362;
assign n_12448 = n_784 & ~n_12362;
assign n_12449 = ~n_3665 & ~n_12362;
assign n_12450 = n_854 & ~n_12362;
assign n_12451 = n_920 & ~n_12362;
assign n_12452 = n_986 & ~n_12362;
assign n_12453 = n_1052 & ~n_12362;
assign n_12454 = n_1117 & ~n_12362;
assign n_12455 = n_1181 & ~n_12362;
assign n_12456 = n_1248 & ~n_12362;
assign n_12457 = n_1314 & ~n_12362;
assign n_12458 = n_1380 & ~n_12362;
assign n_12459 = n_1445 & ~n_12362;
assign n_12460 = ~n_12362 & n_1510;
assign n_12461 = ~n_12362 & n_1576;
assign n_12462 = ~n_12362 & n_1641;
assign n_12463 = ~n_12362 & n_1706;
assign n_12464 = ~n_12362 & n_1771;
assign n_12465 = ~n_12362 & n_1835;
assign n_12466 = ~n_12362 & n_1899;
assign n_12467 = n_1 & n_12363;
assign n_12468 = ~x107 & n_12363;
assign n_12469 = n_12363 ^ x106;
assign n_12470 = n_12244 ^ n_12364;
assign n_12471 = n_12366 ^ n_12188;
assign n_12472 = n_12367 ^ n_11848;
assign n_12473 = n_12367 ^ n_11766;
assign n_12474 = n_12368 ^ n_11850;
assign n_12475 = n_12368 ^ n_11768;
assign n_12476 = n_12369 ^ n_11579;
assign n_12477 = n_12369 ^ n_11483;
assign n_12478 = n_12370 ^ n_11854;
assign n_12479 = n_12370 ^ n_11772;
assign n_12480 = n_12371 ^ n_11856;
assign n_12481 = n_12371 ^ n_11774;
assign n_12482 = n_12372 ^ n_11776;
assign n_12483 = n_12372 ^ n_11678;
assign n_12484 = n_12373 ^ n_9480;
assign n_12485 = ~n_11859 & n_12374;
assign n_12486 = n_12375 ^ n_11795;
assign n_12487 = n_12375 ^ n_11694;
assign n_12488 = n_12376 ^ n_11684;
assign n_12489 = n_12376 ^ n_11569;
assign n_12490 = n_12378 ^ n_12207;
assign n_12491 = n_12380 ^ n_12208;
assign n_12492 = n_12381 ^ n_12209;
assign n_12493 = n_12382 ^ n_11931;
assign n_12494 = n_12382 ^ n_11865;
assign n_12495 = n_12383 ^ n_12052;
assign n_12496 = n_12383 ^ n_11971;
assign n_12497 = n_12384 ^ n_11875;
assign n_12498 = n_12384 ^ n_11791;
assign n_12499 = n_12385 ^ n_12058;
assign n_12500 = n_12385 ^ n_11976;
assign n_12501 = n_12387 ^ n_9482;
assign n_12502 = ~n_11861 & n_12388;
assign n_12503 = n_12389 ^ n_12235;
assign n_12504 = n_12391 ^ n_12236;
assign n_12505 = n_12392 ^ n_12087;
assign n_12506 = n_12393 ^ n_12237;
assign n_12507 = n_12395 ^ n_11832;
assign n_12508 = n_12089 ^ n_12396;
assign n_12509 = n_12397 ^ n_12239;
assign n_12510 = n_12398 ^ n_12090;
assign n_12511 = n_12399 ^ n_12240;
assign n_12512 = n_12091 ^ n_12400;
assign n_12513 = n_12401 ^ n_12241;
assign n_12514 = n_12403 ^ n_11842;
assign n_12515 = ~x0 & n_12404;
assign n_12516 = n_12405 ^ x5;
assign n_12517 = n_12406 ^ x8;
assign n_12518 = n_12407 ^ x11;
assign n_12519 = n_12408 ^ x14;
assign n_12520 = n_12409 ^ x17;
assign n_12521 = n_12410 ^ x20;
assign n_12522 = n_12411 ^ x23;
assign n_12523 = n_12412 ^ x26;
assign n_12524 = n_12413 ^ x29;
assign n_12525 = n_12414 ^ x32;
assign n_12526 = n_12415 ^ x35;
assign n_12527 = n_12416 ^ x38;
assign n_12528 = n_12417 ^ x41;
assign n_12529 = n_12418 ^ x44;
assign n_12530 = n_12419 ^ x47;
assign n_12531 = n_12420 ^ x50;
assign n_12532 = n_12421 ^ x53;
assign n_12533 = n_12422 ^ x56;
assign n_12534 = n_12423 ^ x59;
assign n_12535 = n_12424 ^ x62;
assign n_12536 = n_12425 ^ n_3501;
assign n_12537 = n_5032 ^ n_12426;
assign n_12538 = n_5095 ^ n_12427;
assign n_12539 = n_5158 ^ n_12428;
assign n_12540 = n_5219 ^ n_12429;
assign n_12541 = n_5283 ^ n_12430;
assign n_12542 = n_5347 ^ n_12431;
assign n_12543 = n_5411 ^ n_12432;
assign n_12544 = n_5475 ^ n_12433;
assign n_12545 = n_5536 ^ n_12434;
assign n_12546 = n_5599 ^ n_12435;
assign n_12547 = n_5662 ^ n_12436;
assign n_12548 = n_5726 ^ n_12437;
assign n_12549 = n_5792 ^ n_12438;
assign n_12550 = n_5854 ^ n_12439;
assign n_12551 = n_5918 ^ n_12440;
assign n_12552 = n_5981 ^ n_12441;
assign n_12553 = n_6045 ^ n_12442;
assign n_12554 = n_6109 ^ n_12443;
assign n_12555 = n_6171 ^ n_12444;
assign n_12556 = n_6233 ^ n_12445;
assign n_12557 = n_12446 ^ x105;
assign n_12558 = n_2160 ^ n_12447;
assign n_12559 = n_760 ^ n_12448;
assign n_12560 = n_2231 ^ n_12449;
assign n_12561 = n_2299 ^ n_12450;
assign n_12562 = n_2366 ^ n_12451;
assign n_12563 = n_2433 ^ n_12452;
assign n_12564 = n_2500 ^ n_12453;
assign n_12565 = n_2566 ^ n_12454;
assign n_12566 = n_2631 ^ n_12455;
assign n_12567 = n_2698 ^ n_12456;
assign n_12568 = n_2766 ^ n_12457;
assign n_12569 = n_2833 ^ n_12458;
assign n_12570 = n_2901 ^ n_12459;
assign n_12571 = n_2967 ^ n_12460;
assign n_12572 = n_3036 ^ n_12461;
assign n_12573 = n_3102 ^ n_12462;
assign n_12574 = n_3171 ^ n_12463;
assign n_12575 = n_3235 ^ n_12464;
assign n_12576 = n_3300 ^ n_12465;
assign n_12577 = n_3365 ^ n_12466;
assign n_12578 = n_12467 ^ x1;
assign n_12579 = n_12468 ^ n_12269;
assign n_12580 = n_655 & ~n_12469;
assign n_12581 = n_784 & ~n_12469;
assign n_12582 = ~n_3665 & ~n_12469;
assign n_12583 = n_854 & ~n_12469;
assign n_12584 = n_920 & ~n_12469;
assign n_12585 = n_986 & ~n_12469;
assign n_12586 = n_1052 & ~n_12469;
assign n_12587 = n_1117 & ~n_12469;
assign n_12588 = n_1181 & ~n_12469;
assign n_12589 = n_1248 & ~n_12469;
assign n_12590 = n_1314 & ~n_12469;
assign n_12591 = n_1380 & ~n_12469;
assign n_12592 = n_1445 & ~n_12469;
assign n_12593 = n_1510 & ~n_12469;
assign n_12594 = ~n_12469 & n_1576;
assign n_12595 = ~n_12469 & n_1641;
assign n_12596 = ~n_12469 & n_1706;
assign n_12597 = ~n_12469 & n_1771;
assign n_12598 = ~n_12469 & n_1835;
assign n_12599 = ~n_12469 & n_1899;
assign n_12600 = n_1 & n_12470;
assign n_12601 = x108 & n_12470;
assign n_12602 = n_12470 ^ x107;
assign n_12603 = n_12471 ^ n_11871;
assign n_12604 = n_12471 ^ n_11787;
assign n_12605 = n_12472 ^ n_9472;
assign n_12606 = ~n_11848 & n_12473;
assign n_12607 = n_12474 ^ n_9473;
assign n_12608 = ~n_11850 & n_12475;
assign n_12609 = n_12476 ^ n_9474;
assign n_12610 = ~n_11579 & n_12477;
assign n_12611 = n_12478 ^ n_9477;
assign n_12612 = ~n_11854 & n_12479;
assign n_12613 = n_12480 ^ n_9478;
assign n_12614 = ~n_11856 & n_12481;
assign n_12615 = n_12482 ^ n_9479;
assign n_12616 = ~n_11776 & n_12483;
assign n_12617 = n_12485 ^ n_12284;
assign n_12618 = n_12486 ^ n_9481;
assign n_12619 = ~n_11795 & n_12487;
assign n_12620 = n_12488 ^ n_10299;
assign n_12621 = n_11684 & ~n_12489;
assign n_12622 = n_12490 ^ n_11877;
assign n_12623 = n_12490 ^ n_11793;
assign n_12624 = n_12491 ^ n_11917;
assign n_12625 = n_12491 ^ n_11844;
assign n_12626 = n_12492 ^ n_11869;
assign n_12627 = n_12492 ^ n_11785;
assign n_12628 = n_12493 ^ n_9682;
assign n_12629 = ~n_11931 & n_12494;
assign n_12630 = n_12495 ^ n_9616;
assign n_12631 = ~n_12052 & n_12496;
assign n_12632 = n_12497 ^ n_9620;
assign n_12633 = ~n_11875 & n_12498;
assign n_12634 = n_12499 ^ n_9621;
assign n_12635 = n_12058 & ~n_12500;
assign n_12636 = n_12502 ^ n_12304;
assign n_12637 = n_12503 ^ n_11953;
assign n_12638 = n_11955 ^ n_12504;
assign n_12639 = n_12507 ^ n_12019;
assign n_12640 = n_12514 ^ n_11968;
assign n_12641 = n_12515 ^ n_12319;
assign n_12642 = n_11953 ^ n_12527;
assign n_12643 = n_12528 ^ n_11955;
assign n_12644 = n_12529 ^ n_11957;
assign n_12645 = n_12529 ^ n_12506;
assign n_12646 = n_12019 ^ n_12530;
assign n_12647 = n_12509 ^ n_12531;
assign n_12648 = n_12531 ^ n_12021;
assign n_12649 = n_12511 ^ n_12532;
assign n_12650 = n_12532 ^ n_11961;
assign n_12651 = n_12513 ^ n_12533;
assign n_12652 = n_12533 ^ n_12024;
assign n_12653 = n_12514 ^ n_12534;
assign n_12654 = n_12535 ^ n_6413;
assign n_12655 = n_12535 ^ n_12222;
assign n_12656 = ~x0 & n_12536;
assign n_12657 = n_12537 ^ x5;
assign n_12658 = n_12538 ^ x8;
assign n_12659 = n_12539 ^ x11;
assign n_12660 = n_12540 ^ x14;
assign n_12661 = n_12541 ^ x17;
assign n_12662 = n_12542 ^ x20;
assign n_12663 = n_12543 ^ x23;
assign n_12664 = n_12544 ^ x26;
assign n_12665 = n_12545 ^ x29;
assign n_12666 = n_12546 ^ x32;
assign n_12667 = n_12547 ^ x35;
assign n_12668 = n_12548 ^ x38;
assign n_12669 = n_12549 ^ x41;
assign n_12670 = n_12550 ^ x44;
assign n_12671 = n_12551 ^ x47;
assign n_12672 = n_12552 ^ x50;
assign n_12673 = n_12553 ^ x53;
assign n_12674 = n_12554 ^ x56;
assign n_12675 = n_12555 ^ x59;
assign n_12676 = n_12556 ^ x62;
assign n_12677 = n_12557 ^ n_2110;
assign n_12678 = n_5033 ^ n_12558;
assign n_12679 = n_5096 ^ n_12559;
assign n_12680 = n_5159 ^ n_12560;
assign n_12681 = n_5220 ^ n_12561;
assign n_12682 = n_5284 ^ n_12562;
assign n_12683 = n_5348 ^ n_12563;
assign n_12684 = n_5412 ^ n_12564;
assign n_12685 = n_5476 ^ n_12565;
assign n_12686 = n_5537 ^ n_12566;
assign n_12687 = n_5600 ^ n_12567;
assign n_12688 = n_5663 ^ n_12568;
assign n_12689 = n_5727 ^ n_12569;
assign n_12690 = n_5793 ^ n_12570;
assign n_12691 = n_5855 ^ n_12571;
assign n_12692 = n_5919 ^ n_12572;
assign n_12693 = n_5982 ^ n_12573;
assign n_12694 = n_6046 ^ n_12574;
assign n_12695 = n_6110 ^ n_12575;
assign n_12696 = n_6172 ^ n_12576;
assign n_12697 = n_6234 ^ n_12577;
assign n_12698 = n_12578 ^ x106;
assign n_12699 = n_242 & ~n_12579;
assign n_12700 = n_2161 ^ n_12580;
assign n_12701 = n_761 ^ n_12581;
assign n_12702 = n_2232 ^ n_12582;
assign n_12703 = n_2300 ^ n_12583;
assign n_12704 = n_2367 ^ n_12584;
assign n_12705 = n_2434 ^ n_12585;
assign n_12706 = n_2501 ^ n_12586;
assign n_12707 = n_2567 ^ n_12587;
assign n_12708 = n_2632 ^ n_12588;
assign n_12709 = n_2699 ^ n_12589;
assign n_12710 = n_2767 ^ n_12590;
assign n_12711 = n_2834 ^ n_12591;
assign n_12712 = n_2902 ^ n_12592;
assign n_12713 = n_2968 ^ n_12593;
assign n_12714 = n_3037 ^ n_12594;
assign n_12715 = n_3103 ^ n_12595;
assign n_12716 = n_3172 ^ n_12596;
assign n_12717 = n_3236 ^ n_12597;
assign n_12718 = n_3301 ^ n_12598;
assign n_12719 = n_3366 ^ n_12599;
assign n_12720 = n_12600 ^ x1;
assign n_12721 = n_12601 ^ n_12364;
assign n_12722 = n_655 & ~n_12602;
assign n_12723 = n_784 & ~n_12602;
assign n_12724 = ~n_3665 & ~n_12602;
assign n_12725 = n_854 & ~n_12602;
assign n_12726 = n_920 & ~n_12602;
assign n_12727 = n_986 & ~n_12602;
assign n_12728 = n_1052 & ~n_12602;
assign n_12729 = n_1117 & ~n_12602;
assign n_12730 = n_1181 & ~n_12602;
assign n_12731 = n_1248 & ~n_12602;
assign n_12732 = n_1314 & ~n_12602;
assign n_12733 = n_1380 & ~n_12602;
assign n_12734 = n_1445 & ~n_12602;
assign n_12735 = n_1510 & ~n_12602;
assign n_12736 = ~n_12602 & n_1576;
assign n_12737 = ~n_12602 & n_1641;
assign n_12738 = ~n_12602 & n_1706;
assign n_12739 = ~n_12602 & n_1771;
assign n_12740 = ~n_12602 & n_1835;
assign n_12741 = ~n_12602 & n_1899;
assign n_12742 = n_12603 ^ n_9615;
assign n_12743 = n_11871 & ~n_12604;
assign n_12744 = n_12606 ^ n_12367;
assign n_12745 = n_12608 ^ n_12368;
assign n_12746 = n_12610 ^ n_12369;
assign n_12747 = n_12612 ^ n_12370;
assign n_12748 = n_12614 ^ n_12371;
assign n_12749 = n_12616 ^ n_12372;
assign n_12750 = n_12617 ^ n_12065;
assign n_12751 = n_12617 ^ n_11983;
assign n_12752 = n_12619 ^ n_12375;
assign n_12753 = n_12621 ^ n_12376;
assign n_12754 = n_12622 ^ n_12234;
assign n_12755 = n_11877 & ~n_12623;
assign n_12756 = n_12624 ^ n_9614;
assign n_12757 = ~n_11917 & n_12625;
assign y20 = n_12626;
assign n_12758 = ~n_11869 & n_12627;
assign n_12759 = n_12629 ^ n_12382;
assign n_12760 = n_12631 ^ n_12383;
assign n_12761 = n_12633 ^ n_12384;
assign n_12762 = n_12635 ^ n_12385;
assign n_12763 = n_12636 ^ n_12067;
assign n_12764 = n_12636 ^ n_11985;
assign n_12765 = n_12637 ^ n_12527;
assign n_12766 = n_12639 ^ n_12530;
assign n_12767 = n_12637 & ~n_12642;
assign n_12768 = n_12643 ^ n_12504;
assign n_12769 = n_12643 & ~n_12638;
assign n_12770 = n_12644 ^ n_12506;
assign n_12771 = n_12644 & n_12645;
assign n_12772 = ~n_12639 & n_12646;
assign n_12773 = n_12647 ^ n_12021;
assign n_12774 = n_12647 & n_12648;
assign n_12775 = n_12649 ^ n_11961;
assign n_12776 = n_12649 & n_12650;
assign n_12777 = n_12651 ^ n_12024;
assign n_12778 = n_12651 & ~n_12652;
assign n_12779 = n_12653 ^ n_11968;
assign n_12780 = ~n_12653 & ~n_12640;
assign n_12781 = n_12654 ^ n_12222;
assign n_12782 = n_12654 & n_12655;
assign n_12783 = n_12656 ^ n_12425;
assign n_12784 = n_12218 ^ n_12667;
assign n_12785 = n_12668 ^ n_12154;
assign n_12786 = n_12668 ^ n_12094;
assign n_12787 = n_12669 ^ n_12155;
assign n_12788 = n_12669 ^ n_12095;
assign n_12789 = n_12670 ^ n_12156;
assign n_12790 = n_12670 ^ n_11946;
assign n_12791 = n_12671 ^ n_12097;
assign n_12792 = n_12672 ^ n_12098;
assign n_12793 = n_12673 ^ n_12010;
assign n_12794 = n_12674 ^ n_12012;
assign n_12795 = n_12675 ^ n_12014;
assign n_12796 = n_12676 ^ n_6644;
assign n_12797 = n_12676 ^ n_6534;
assign n_12798 = ~x0 & n_12677;
assign n_12799 = n_12678 ^ x5;
assign n_12800 = n_12679 ^ x8;
assign n_12801 = n_12680 ^ x11;
assign n_12802 = n_12681 ^ x14;
assign n_12803 = n_12682 ^ x17;
assign n_12804 = n_12683 ^ x20;
assign n_12805 = n_12684 ^ x23;
assign n_12806 = n_12685 ^ x26;
assign n_12807 = n_12686 ^ x29;
assign n_12808 = n_12687 ^ x32;
assign n_12809 = n_12688 ^ x35;
assign n_12810 = n_12689 ^ x38;
assign n_12811 = n_12690 ^ x41;
assign n_12812 = n_12691 ^ x44;
assign n_12813 = n_12692 ^ x47;
assign n_12814 = n_12693 ^ x50;
assign n_12815 = n_12694 ^ x53;
assign n_12816 = n_12695 ^ x56;
assign n_12817 = n_12696 ^ x59;
assign n_12818 = n_12697 ^ x62;
assign n_12819 = n_12698 ^ n_3504;
assign n_12820 = n_1 & ~n_12699;
assign n_12821 = n_12699 ^ x108;
assign n_12822 = n_5034 ^ n_12700;
assign n_12823 = n_5097 ^ n_12701;
assign n_12824 = n_5160 ^ n_12702;
assign n_12825 = n_5221 ^ n_12703;
assign n_12826 = n_5285 ^ n_12704;
assign n_12827 = n_5349 ^ n_12705;
assign n_12828 = n_5413 ^ n_12706;
assign n_12829 = n_5477 ^ n_12707;
assign n_12830 = n_5538 ^ n_12708;
assign n_12831 = n_5601 ^ n_12709;
assign n_12832 = n_5664 ^ n_12710;
assign n_12833 = n_5728 ^ n_12711;
assign n_12834 = n_5794 ^ n_12712;
assign n_12835 = n_5856 ^ n_12713;
assign n_12836 = n_5920 ^ n_12714;
assign n_12837 = n_5983 ^ n_12715;
assign n_12838 = n_6047 ^ n_12716;
assign n_12839 = n_6111 ^ n_12717;
assign n_12840 = n_6173 ^ n_12718;
assign n_12841 = n_6235 ^ n_12719;
assign n_12842 = n_12720 ^ x107;
assign n_12843 = n_244 & ~n_12721;
assign n_12844 = n_2162 ^ n_12722;
assign n_12845 = n_762 ^ n_12723;
assign n_12846 = n_2233 ^ n_12724;
assign n_12847 = n_2301 ^ n_12725;
assign n_12848 = n_2368 ^ n_12726;
assign n_12849 = n_2435 ^ n_12727;
assign n_12850 = n_2502 ^ n_12728;
assign n_12851 = n_2568 ^ n_12729;
assign n_12852 = n_2633 ^ n_12730;
assign n_12853 = n_2700 ^ n_12731;
assign n_12854 = n_2768 ^ n_12732;
assign n_12855 = n_2835 ^ n_12733;
assign n_12856 = n_2903 ^ n_12734;
assign n_12857 = n_2969 ^ n_12735;
assign n_12858 = n_3038 ^ n_12736;
assign n_12859 = n_3104 ^ n_12737;
assign n_12860 = n_3173 ^ n_12738;
assign n_12861 = n_3237 ^ n_12739;
assign n_12862 = n_3302 ^ n_12740;
assign n_12863 = n_3367 ^ n_12741;
assign n_12864 = n_12743 ^ n_12471;
assign n_12865 = n_12744 ^ n_12054;
assign n_12866 = n_12744 ^ n_11973;
assign n_12867 = n_12745 ^ n_12130;
assign n_12868 = n_12745 ^ n_12056;
assign n_12869 = n_12746 ^ n_11873;
assign n_12870 = n_12746 ^ n_11789;
assign n_12871 = n_12747 ^ n_12060;
assign n_12872 = n_12747 ^ n_9199;
assign n_12873 = n_12748 ^ n_12134;
assign n_12874 = n_12748 ^ n_12062;
assign n_12875 = n_12749 ^ n_11981;
assign n_12876 = n_12749 ^ n_11925;
assign n_12877 = n_12750 ^ n_9625;
assign n_12878 = ~n_12065 & n_12751;
assign n_12879 = n_12752 ^ n_12000;
assign n_12880 = n_12752 ^ n_11939;
assign n_12881 = n_12753 ^ n_11929;
assign n_12882 = n_12753 ^ n_11863;
assign n_12883 = n_12755 ^ n_12490;
assign n_12884 = n_12757 ^ n_12491;
assign n_12885 = n_12758 ^ n_12492;
assign n_12886 = n_12759 ^ n_12142;
assign n_12887 = n_12759 ^ n_12071;
assign n_12888 = n_12760 ^ n_12272;
assign n_12889 = n_12760 ^ n_12189;
assign n_12890 = n_12761 ^ n_12081;
assign n_12891 = n_12761 ^ n_11996;
assign n_12892 = n_12762 ^ n_12278;
assign n_12893 = n_12762 ^ n_12195;
assign n_12894 = n_12763 ^ n_9627;
assign n_12895 = ~n_12067 & n_12764;
assign n_12896 = n_12767 ^ n_12503;
assign n_12897 = n_12769 ^ n_12528;
assign n_12898 = n_12771 ^ n_12506;
assign n_12899 = n_12772 ^ n_12507;
assign n_12900 = n_12774 ^ n_12509;
assign n_12901 = n_12776 ^ n_12511;
assign n_12902 = n_12778 ^ n_12513;
assign n_12903 = n_12780 ^ n_12534;
assign n_12904 = n_12782 ^ n_12222;
assign n_12905 = n_12154 & n_12786;
assign n_12906 = ~n_12155 & n_12788;
assign n_12907 = n_12156 & ~n_12790;
assign n_12908 = n_12791 ^ n_12006;
assign n_12909 = n_12791 & n_12157;
assign n_12910 = n_12792 ^ n_12008;
assign n_12911 = n_12792 & n_12158;
assign n_12912 = n_12793 ^ n_12099;
assign n_12913 = ~n_12793 & n_12159;
assign n_12914 = n_12794 ^ n_12100;
assign n_12915 = n_12794 & ~n_12160;
assign n_12916 = n_12795 ^ n_12125;
assign n_12917 = ~n_12795 & n_12187;
assign n_12918 = n_6644 & n_12797;
assign n_12919 = n_12798 ^ n_12557;
assign n_12920 = n_12809 ^ n_12306;
assign n_12921 = n_12386 ^ n_12809;
assign n_12922 = n_12810 ^ n_12390;
assign n_12923 = n_12810 ^ n_12308;
assign n_12924 = n_12811 ^ n_12505;
assign n_12925 = n_12811 ^ n_12087;
assign n_12926 = n_12812 ^ n_12394;
assign n_12927 = n_12812 ^ n_12311;
assign n_12928 = n_12813 ^ n_12089;
assign n_12929 = n_12814 ^ n_12510;
assign n_12930 = n_12814 ^ n_12398;
assign n_12931 = n_12815 ^ n_12091;
assign n_12932 = n_12816 ^ n_12092;
assign n_12933 = n_12817 ^ n_12318;
assign n_12934 = n_12817 ^ n_12152;
assign n_12935 = ~x0 & n_12819;
assign n_12936 = n_12820 ^ x1;
assign n_12937 = n_655 & n_12821;
assign n_12938 = n_784 & n_12821;
assign n_12939 = ~n_3665 & n_12821;
assign n_12940 = n_854 & n_12821;
assign n_12941 = n_920 & n_12821;
assign n_12942 = n_986 & n_12821;
assign n_12943 = n_1052 & n_12821;
assign n_12944 = n_1117 & n_12821;
assign n_12945 = n_1181 & n_12821;
assign n_12946 = n_1248 & n_12821;
assign n_12947 = n_1314 & n_12821;
assign n_12948 = n_1380 & n_12821;
assign n_12949 = n_1445 & n_12821;
assign n_12950 = n_1510 & n_12821;
assign n_12951 = n_12821 & n_1576;
assign n_12952 = n_12821 & n_1641;
assign n_12953 = n_12821 & n_1706;
assign n_12954 = n_12821 & n_1771;
assign n_12955 = n_12821 & n_1835;
assign n_12956 = n_12821 & n_1899;
assign n_12957 = n_12822 ^ x5;
assign n_12958 = n_12823 ^ x8;
assign n_12959 = n_12824 ^ x11;
assign n_12960 = n_12825 ^ x14;
assign n_12961 = n_12826 ^ x17;
assign n_12962 = n_12827 ^ x20;
assign n_12963 = n_12828 ^ x23;
assign n_12964 = n_12829 ^ x26;
assign n_12965 = n_12830 ^ x29;
assign n_12966 = n_12831 ^ x32;
assign n_12967 = n_12832 ^ x35;
assign n_12968 = n_12833 ^ x38;
assign n_12969 = n_12834 ^ x41;
assign n_12970 = n_12835 ^ x44;
assign n_12971 = n_12836 ^ x47;
assign n_12972 = n_12837 ^ x50;
assign n_12973 = n_12838 ^ x53;
assign n_12974 = n_12839 ^ x56;
assign n_12975 = n_12840 ^ x59;
assign n_12976 = n_12841 ^ x62;
assign n_12977 = n_12842 ^ n_2111;
assign n_12978 = n_1 & ~n_12843;
assign n_12979 = n_12843 & n_248;
assign n_12980 = n_12843 ^ x109;
assign n_12981 = n_5035 ^ n_12844;
assign n_12982 = n_5098 ^ n_12845;
assign n_12983 = n_5161 ^ n_12846;
assign n_12984 = n_5222 ^ n_12847;
assign n_12985 = n_5286 ^ n_12848;
assign n_12986 = n_5350 ^ n_12849;
assign n_12987 = n_5414 ^ n_12850;
assign n_12988 = n_5478 ^ n_12851;
assign n_12989 = n_5539 ^ n_12852;
assign n_12990 = n_5602 ^ n_12853;
assign n_12991 = n_5665 ^ n_12854;
assign n_12992 = n_5729 ^ n_12855;
assign n_12993 = n_5795 ^ n_12856;
assign n_12994 = n_5857 ^ n_12857;
assign n_12995 = n_5921 ^ n_12858;
assign n_12996 = n_5984 ^ n_12859;
assign n_12997 = n_6048 ^ n_12860;
assign n_12998 = n_6112 ^ n_12861;
assign n_12999 = n_6174 ^ n_12862;
assign n_13000 = n_6236 ^ n_12863;
assign n_13001 = n_12864 ^ n_12077;
assign n_13002 = n_12864 ^ n_11992;
assign n_13003 = n_12865 ^ n_9617;
assign n_13004 = ~n_12054 & n_12866;
assign n_13005 = n_12867 ^ n_9618;
assign n_13006 = ~n_12130 & n_12868;
assign n_13007 = n_12869 ^ n_9619;
assign n_13008 = ~n_11873 & n_12870;
assign n_13009 = n_12871 ^ n_9622;
assign n_13010 = n_12060 & ~n_12872;
assign n_13011 = n_12873 ^ n_9623;
assign n_13012 = ~n_12134 & n_12874;
assign n_13013 = n_12875 ^ n_9624;
assign n_13014 = ~n_11981 & n_12876;
assign n_13015 = n_12878 ^ n_12617;
assign n_13016 = n_12879 ^ n_9626;
assign n_13017 = ~n_12000 & n_12880;
assign n_13018 = n_12881 ^ n_10865;
assign n_13019 = ~n_11929 & n_12882;
assign n_13020 = n_12883 ^ n_12083;
assign n_13021 = n_12883 ^ n_11998;
assign n_13022 = n_12884 ^ n_12126;
assign n_13023 = n_12884 ^ n_12050;
assign n_13024 = n_12885 ^ n_12075;
assign n_13025 = n_12885 ^ n_11990;
assign n_13026 = n_12886 ^ n_9825;
assign n_13027 = ~n_12142 & n_12887;
assign n_13028 = n_12888 ^ n_9753;
assign n_13029 = ~n_12272 & n_12889;
assign n_13030 = n_12890 ^ n_9757;
assign n_13031 = ~n_12081 & n_12891;
assign n_13032 = n_12892 ^ n_9758;
assign n_13033 = n_12278 & ~n_12893;
assign n_13034 = n_12895 ^ n_12636;
assign n_13035 = n_12896 ^ n_12785;
assign n_13036 = n_12897 ^ n_12787;
assign n_13037 = n_12898 ^ n_12789;
assign n_13038 = n_12905 ^ n_12668;
assign n_13039 = n_12906 ^ n_12669;
assign n_13040 = n_12907 ^ n_12096;
assign n_13041 = n_12899 ^ n_12908;
assign n_13042 = n_12909 ^ n_12671;
assign n_13043 = n_12900 ^ n_12910;
assign n_13044 = n_12911 ^ n_12672;
assign n_13045 = n_12901 ^ n_12912;
assign n_13046 = n_12913 ^ n_12673;
assign n_13047 = n_12915 ^ n_12674;
assign n_13048 = n_12903 ^ n_12916;
assign n_13049 = n_12917 ^ n_12675;
assign n_13050 = n_12918 ^ n_12676;
assign n_13051 = n_12386 ^ n_12920;
assign n_13052 = ~n_12920 & n_12921;
assign n_13053 = ~n_12390 & n_12923;
assign n_13054 = n_12505 & n_12925;
assign n_13055 = ~n_12394 & n_12927;
assign n_13056 = n_12928 ^ n_12396;
assign n_13057 = n_12928 & n_12508;
assign n_13058 = ~n_12510 & n_12930;
assign n_13059 = n_12931 ^ n_12400;
assign n_13060 = n_12931 & ~n_12512;
assign n_13061 = n_12932 ^ n_12316;
assign n_13062 = n_12932 & n_12402;
assign n_13063 = n_12318 & ~n_12934;
assign n_13064 = n_12935 ^ n_12698;
assign n_13065 = n_12936 ^ x108;
assign n_13066 = n_2163 ^ n_12937;
assign n_13067 = n_763 ^ n_12938;
assign n_13068 = n_2234 ^ n_12939;
assign n_13069 = n_2302 ^ n_12940;
assign n_13070 = n_2369 ^ n_12941;
assign n_13071 = n_2436 ^ n_12942;
assign n_13072 = n_2503 ^ n_12943;
assign n_13073 = n_2569 ^ n_12944;
assign n_13074 = n_2634 ^ n_12945;
assign n_13075 = n_2701 ^ n_12946;
assign n_13076 = n_2769 ^ n_12947;
assign n_13077 = n_2836 ^ n_12948;
assign n_13078 = n_2904 ^ n_12949;
assign n_13079 = n_2970 ^ n_12950;
assign n_13080 = n_3039 ^ n_12951;
assign n_13081 = n_3105 ^ n_12952;
assign n_13082 = n_3174 ^ n_12953;
assign n_13083 = n_3238 ^ n_12954;
assign n_13084 = n_3303 ^ n_12955;
assign n_13085 = n_3368 ^ n_12956;
assign n_13086 = n_12967 ^ n_12765;
assign n_13087 = n_12968 ^ n_12768;
assign n_13088 = n_12969 ^ n_12770;
assign n_13089 = n_12970 ^ n_12766;
assign n_13090 = n_12773 ^ n_12971;
assign n_13091 = n_12972 ^ n_12775;
assign n_13092 = n_12973 ^ n_12777;
assign n_13093 = n_12974 ^ n_12779;
assign n_13094 = n_12975 ^ n_12781;
assign n_13095 = n_12976 ^ n_6352;
assign n_13096 = ~x0 & n_12977;
assign n_13097 = n_12978 ^ x1;
assign n_13098 = n_12979 ^ x108;
assign n_13099 = n_655 & n_12980;
assign n_13100 = n_784 & n_12980;
assign n_13101 = ~n_3665 & n_12980;
assign n_13102 = n_854 & n_12980;
assign n_13103 = n_920 & n_12980;
assign n_13104 = n_986 & n_12980;
assign n_13105 = n_1052 & n_12980;
assign n_13106 = n_1117 & n_12980;
assign n_13107 = n_1181 & n_12980;
assign n_13108 = n_1248 & n_12980;
assign n_13109 = n_1314 & n_12980;
assign n_13110 = n_1380 & n_12980;
assign n_13111 = n_1445 & n_12980;
assign n_13112 = n_1510 & n_12980;
assign n_13113 = n_1576 & n_12980;
assign n_13114 = n_12980 & n_1641;
assign n_13115 = n_12980 & n_1706;
assign n_13116 = n_12980 & n_1771;
assign n_13117 = n_12980 & n_1835;
assign n_13118 = n_12980 & n_1899;
assign n_13119 = n_12981 ^ x5;
assign n_13120 = n_12982 ^ x8;
assign n_13121 = n_12983 ^ x11;
assign n_13122 = n_12984 ^ x14;
assign n_13123 = n_12985 ^ x17;
assign n_13124 = n_12986 ^ x20;
assign n_13125 = n_12987 ^ x23;
assign n_13126 = n_12988 ^ x26;
assign n_13127 = n_12989 ^ x29;
assign n_13128 = n_12990 ^ x32;
assign n_13129 = n_12991 ^ x35;
assign n_13130 = n_12992 ^ x38;
assign n_13131 = n_12993 ^ x41;
assign n_13132 = n_12994 ^ x44;
assign n_13133 = n_12995 ^ x47;
assign n_13134 = n_12996 ^ x50;
assign n_13135 = n_12997 ^ x53;
assign n_13136 = n_12998 ^ x56;
assign n_13137 = n_12999 ^ x59;
assign n_13138 = n_13000 ^ x62;
assign n_13139 = n_13001 ^ n_9752;
assign n_13140 = ~n_12077 & n_13002;
assign n_13141 = n_13004 ^ n_12744;
assign n_13142 = n_13006 ^ n_12745;
assign n_13143 = n_13008 ^ n_12746;
assign n_13144 = n_13010 ^ n_11978;
assign n_13145 = n_13012 ^ n_12748;
assign n_13146 = n_13014 ^ n_12749;
assign n_13147 = n_13015 ^ n_12285;
assign n_13148 = n_13015 ^ n_12203;
assign n_13149 = n_13017 ^ n_12752;
assign n_13150 = n_13019 ^ n_12753;
assign n_13151 = n_13020 ^ n_12526;
assign n_13152 = ~n_12083 & n_13021;
assign n_13153 = n_13022 ^ n_9751;
assign n_13154 = n_12126 & ~n_13023;
assign y21 = n_13024;
assign n_13155 = ~n_12075 & n_13025;
assign n_13156 = n_13027 ^ n_12759;
assign n_13157 = n_13029 ^ n_12760;
assign n_13158 = n_13031 ^ n_12761;
assign n_13159 = n_13033 ^ n_12762;
assign n_13160 = n_13034 ^ n_12287;
assign n_13161 = n_13034 ^ n_12205;
assign n_13162 = n_13038 ^ n_12922;
assign n_13163 = n_13039 ^ n_12924;
assign n_13164 = n_13040 ^ n_12926;
assign n_13165 = n_12929 ^ n_13044;
assign n_13166 = n_13050 ^ n_6605;
assign n_13167 = n_6605 & ~n_13050;
assign n_13168 = n_13052 ^ n_12386;
assign n_13169 = n_13053 ^ n_12810;
assign n_13170 = n_13054 ^ n_12811;
assign n_13171 = n_13055 ^ n_12812;
assign n_13172 = n_13056 ^ n_13042;
assign n_13173 = n_13057 ^ n_12813;
assign n_13174 = n_13058 ^ n_12814;
assign n_13175 = n_13046 ^ n_13059;
assign n_13176 = n_13060 ^ n_12815;
assign n_13177 = n_13062 ^ n_12816;
assign n_13178 = n_13063 ^ n_12817;
assign n_13179 = n_13065 ^ n_3508;
assign n_13180 = n_5036 ^ n_13066;
assign n_13181 = n_5099 ^ n_13067;
assign n_13182 = n_5162 ^ n_13068;
assign n_13183 = n_5223 ^ n_13069;
assign n_13184 = n_5287 ^ n_13070;
assign n_13185 = n_5351 ^ n_13071;
assign n_13186 = n_5415 ^ n_13072;
assign n_13187 = n_5479 ^ n_13073;
assign n_13188 = n_5540 ^ n_13074;
assign n_13189 = n_5603 ^ n_13075;
assign n_13190 = n_5666 ^ n_13076;
assign n_13191 = n_5730 ^ n_13077;
assign n_13192 = n_5796 ^ n_13078;
assign n_13193 = n_5858 ^ n_13079;
assign n_13194 = n_5922 ^ n_13080;
assign n_13195 = n_5985 ^ n_13081;
assign n_13196 = n_6049 ^ n_13082;
assign n_13197 = n_6113 ^ n_13083;
assign n_13198 = n_6175 ^ n_13084;
assign n_13199 = n_6237 ^ n_13085;
assign n_13200 = n_13096 ^ n_12842;
assign n_13201 = n_13097 ^ x109;
assign n_13202 = n_13098 ^ x109;
assign n_13203 = ~x109 & ~n_13098;
assign n_13204 = n_253 ^ n_13098;
assign n_13205 = n_2164 ^ n_13099;
assign n_13206 = n_764 ^ n_13100;
assign n_13207 = n_2235 ^ n_13101;
assign n_13208 = n_2303 ^ n_13102;
assign n_13209 = n_2370 ^ n_13103;
assign n_13210 = n_2437 ^ n_13104;
assign n_13211 = n_2504 ^ n_13105;
assign n_13212 = n_2570 ^ n_13106;
assign n_13213 = n_2635 ^ n_13107;
assign n_13214 = n_2702 ^ n_13108;
assign n_13215 = n_2770 ^ n_13109;
assign n_13216 = n_2837 ^ n_13110;
assign n_13217 = n_2905 ^ n_13111;
assign n_13218 = n_2971 ^ n_13112;
assign n_13219 = n_3040 ^ n_13113;
assign n_13220 = n_3106 ^ n_13114;
assign n_13221 = n_3175 ^ n_13115;
assign n_13222 = n_3239 ^ n_13116;
assign n_13223 = n_3304 ^ n_13117;
assign n_13224 = n_3369 ^ n_13118;
assign n_13225 = n_13035 ^ n_13129;
assign n_13226 = n_12896 ^ n_13129;
assign n_13227 = n_13036 ^ n_13130;
assign n_13228 = n_12897 ^ n_13130;
assign n_13229 = n_13037 ^ n_13131;
assign n_13230 = n_12789 ^ n_13131;
assign n_13231 = n_13041 ^ n_13132;
assign n_13232 = n_12908 ^ n_13132;
assign n_13233 = n_13043 ^ n_13133;
assign n_13234 = n_12910 ^ n_13133;
assign n_13235 = n_13045 ^ n_13134;
assign n_13236 = n_12912 ^ n_13134;
assign n_13237 = n_13135 ^ n_12902;
assign n_13238 = n_13135 ^ n_12914;
assign n_13239 = n_13136 ^ n_12903;
assign n_13240 = n_13137 ^ n_12904;
assign n_13241 = n_13137 ^ n_12796;
assign n_13242 = n_13138 ^ n_6606;
assign n_13243 = n_13138 ^ n_6488;
assign n_13244 = n_13140 ^ n_12864;
assign n_13245 = n_13141 ^ n_12274;
assign n_13246 = n_13141 ^ n_12191;
assign n_13247 = n_13142 ^ n_12276;
assign n_13248 = n_13142 ^ n_12193;
assign n_13249 = n_13143 ^ n_12079;
assign n_13250 = n_13143 ^ n_11994;
assign n_13251 = n_13144 ^ n_12280;
assign n_13252 = n_13144 ^ n_9333;
assign n_13253 = n_13145 ^ n_12282;
assign n_13254 = n_13145 ^ n_12199;
assign n_13255 = n_13146 ^ n_12201;
assign n_13256 = n_13146 ^ n_12136;
assign n_13257 = n_13147 ^ n_9762;
assign n_13258 = n_12285 & ~n_13148;
assign n_13259 = n_13149 ^ n_12220;
assign n_13260 = n_13149 ^ n_12150;
assign n_13261 = n_13150 ^ n_12140;
assign n_13262 = n_13150 ^ n_12069;
assign n_13263 = n_13152 ^ n_12883;
assign n_13264 = n_13154 ^ n_12884;
assign n_13265 = n_13155 ^ n_12885;
assign n_13266 = n_13156 ^ n_12379;
assign n_13267 = n_13156 ^ n_12291;
assign n_13268 = n_13157 ^ n_12605;
assign n_13269 = n_13157 ^ n_12472;
assign n_13270 = n_13158 ^ n_12301;
assign n_13271 = n_13158 ^ n_12216;
assign n_13272 = n_13159 ^ n_12611;
assign n_13273 = n_13159 ^ n_12478;
assign n_13274 = n_13160 ^ n_10168;
assign n_13275 = n_12287 & ~n_13161;
assign n_13276 = n_13166 ^ n_12818;
assign n_13277 = n_13167 ^ n_6283;
assign n_13278 = n_13168 ^ n_13086;
assign n_13279 = n_13168 ^ n_12967;
assign n_13280 = n_13169 ^ n_13087;
assign n_13281 = n_13169 ^ n_12968;
assign n_13282 = n_13170 ^ n_13088;
assign n_13283 = n_13170 ^ n_12969;
assign n_13284 = n_13171 ^ n_13089;
assign n_13285 = n_13171 ^ n_12970;
assign n_13286 = n_13173 ^ n_12773;
assign n_13287 = n_13174 ^ n_12972;
assign n_13288 = n_13176 ^ n_12973;
assign n_13289 = n_13177 ^ n_12974;
assign n_13290 = n_13178 ^ n_12975;
assign n_13291 = ~x0 & n_13179;
assign n_13292 = n_13180 ^ x5;
assign n_13293 = n_13181 ^ x8;
assign n_13294 = n_13182 ^ x11;
assign n_13295 = n_13183 ^ x14;
assign n_13296 = n_13184 ^ x17;
assign n_13297 = n_13185 ^ x20;
assign n_13298 = n_13186 ^ x23;
assign n_13299 = n_13187 ^ x26;
assign n_13300 = n_13188 ^ x29;
assign n_13301 = n_13189 ^ x32;
assign n_13302 = n_13190 ^ x35;
assign n_13303 = n_13191 ^ x38;
assign n_13304 = n_13192 ^ x41;
assign n_13305 = n_13193 ^ x44;
assign n_13306 = n_13194 ^ x47;
assign n_13307 = n_13195 ^ x50;
assign n_13308 = n_13196 ^ x53;
assign n_13309 = n_13197 ^ x56;
assign n_13310 = n_13198 ^ x59;
assign n_13311 = n_13199 ^ x62;
assign n_13312 = n_13201 ^ n_6490;
assign n_13313 = n_1 & ~n_13202;
assign n_13314 = x110 & ~n_13203;
assign n_13315 = n_13203 ^ n_13202;
assign n_13316 = n_655 & n_13204;
assign n_13317 = n_784 & n_13204;
assign n_13318 = ~n_3665 & n_13204;
assign n_13319 = n_854 & n_13204;
assign n_13320 = n_920 & n_13204;
assign n_13321 = n_986 & n_13204;
assign n_13322 = n_1052 & n_13204;
assign n_13323 = n_1117 & n_13204;
assign n_13324 = n_1181 & n_13204;
assign n_13325 = n_1248 & n_13204;
assign n_13326 = n_1314 & n_13204;
assign n_13327 = n_1380 & n_13204;
assign n_13328 = n_1445 & n_13204;
assign n_13329 = n_1510 & n_13204;
assign n_13330 = n_1576 & n_13204;
assign n_13331 = n_13204 & n_1641;
assign n_13332 = n_13204 & n_1706;
assign n_13333 = n_13204 & n_1771;
assign n_13334 = n_13204 & n_1835;
assign n_13335 = n_13204 & n_1899;
assign n_13336 = n_5037 ^ n_13205;
assign n_13337 = n_5100 ^ n_13206;
assign n_13338 = n_5163 ^ n_13207;
assign n_13339 = n_5224 ^ n_13208;
assign n_13340 = n_5288 ^ n_13209;
assign n_13341 = n_5352 ^ n_13210;
assign n_13342 = n_5416 ^ n_13211;
assign n_13343 = n_5480 ^ n_13212;
assign n_13344 = n_5541 ^ n_13213;
assign n_13345 = n_5604 ^ n_13214;
assign n_13346 = n_5667 ^ n_13215;
assign n_13347 = n_5731 ^ n_13216;
assign n_13348 = n_5797 ^ n_13217;
assign n_13349 = n_5859 ^ n_13218;
assign n_13350 = n_5923 ^ n_13219;
assign n_13351 = n_5986 ^ n_13220;
assign n_13352 = n_6050 ^ n_13221;
assign n_13353 = n_6114 ^ n_13222;
assign n_13354 = n_6176 ^ n_13223;
assign n_13355 = n_6238 ^ n_13224;
assign n_13356 = n_13035 & n_13226;
assign n_13357 = ~n_13036 & n_13228;
assign n_13358 = n_13037 & ~n_13230;
assign n_13359 = n_13041 & ~n_13232;
assign n_13360 = ~n_13043 & n_13234;
assign n_13361 = ~n_13045 & n_13236;
assign n_13362 = n_13237 ^ n_12914;
assign n_13363 = n_13237 & ~n_13238;
assign n_13364 = n_13239 ^ n_12916;
assign n_13365 = n_13239 & n_13048;
assign n_13366 = n_13240 ^ n_12796;
assign n_13367 = n_13240 & n_13241;
assign n_13368 = n_6606 & n_13243;
assign n_13369 = n_13244 ^ n_12297;
assign n_13370 = n_13244 ^ n_12212;
assign n_13371 = n_13245 ^ n_9754;
assign n_13372 = ~n_12274 & n_13246;
assign n_13373 = n_13247 ^ n_9755;
assign n_13374 = ~n_12276 & n_13248;
assign n_13375 = n_13249 ^ n_9756;
assign n_13376 = n_12079 & ~n_13250;
assign n_13377 = n_13251 ^ n_9759;
assign n_13378 = n_12280 & ~n_13252;
assign n_13379 = n_13253 ^ n_9760;
assign n_13380 = ~n_12282 & n_13254;
assign n_13381 = n_13255 ^ n_9761;
assign n_13382 = n_12201 & ~n_13256;
assign n_13383 = n_13258 ^ n_13015;
assign n_13384 = n_13259 ^ n_9763;
assign n_13385 = ~n_12220 & n_13260;
assign n_13386 = n_13261 ^ n_11136;
assign n_13387 = n_12140 & ~n_13262;
assign n_13388 = n_13263 ^ n_12784;
assign n_13389 = n_13263 ^ n_12218;
assign n_13390 = n_13264 ^ n_12365;
assign n_13391 = n_13264 ^ n_12270;
assign n_13392 = n_13265 ^ n_12295;
assign n_13393 = n_13265 ^ n_12210;
assign n_13394 = n_13266 ^ n_9973;
assign n_13395 = ~n_12379 & n_13267;
assign n_13396 = n_13268 ^ n_9895;
assign n_13397 = ~n_12605 & n_13269;
assign n_13398 = n_13270 ^ n_9899;
assign n_13399 = ~n_12301 & n_13271;
assign n_13400 = n_13272 ^ n_9900;
assign n_13401 = ~n_12611 & n_13273;
assign n_13402 = n_13275 ^ n_13034;
assign n_13403 = n_13277 ^ n_13095;
assign n_13404 = n_13277 ^ n_12976;
assign n_13405 = ~n_13086 & n_13279;
assign n_13406 = ~n_13087 & n_13281;
assign n_13407 = n_13088 & n_13283;
assign n_13408 = n_13089 & n_13285;
assign n_13409 = n_13286 ^ n_12971;
assign n_13410 = ~n_13286 & n_13090;
assign n_13411 = n_13287 ^ n_12775;
assign n_13412 = n_13287 & n_13091;
assign n_13413 = n_13288 ^ n_12777;
assign n_13414 = n_13288 & ~n_13092;
assign n_13415 = n_13289 ^ n_12779;
assign n_13416 = n_13289 & ~n_13093;
assign n_13417 = n_13290 ^ n_12781;
assign n_13418 = n_13290 & n_13094;
assign n_13419 = n_13291 ^ n_13065;
assign n_13420 = n_13301 ^ n_13051;
assign n_13421 = n_13302 ^ n_13162;
assign n_13422 = n_13302 ^ n_12922;
assign n_13423 = n_13303 ^ n_13163;
assign n_13424 = n_13303 ^ n_12924;
assign n_13425 = n_13304 ^ n_13164;
assign n_13426 = n_13304 ^ n_13040;
assign n_13427 = n_13305 ^ n_13172;
assign n_13428 = n_13305 ^ n_13056;
assign n_13429 = n_13306 ^ n_12929;
assign n_13430 = n_13307 ^ n_13046;
assign n_13431 = n_13308 ^ n_13047;
assign n_13432 = n_13308 ^ n_13061;
assign n_13433 = n_13309 ^ n_13049;
assign n_13434 = n_13309 ^ n_12933;
assign n_13435 = n_13310 ^ n_13166;
assign n_13436 = ~x0 & ~n_13312;
assign n_13437 = n_13313 ^ x1;
assign n_13438 = ~x111 & ~n_13314;
assign n_13439 = ~x110 & n_13315;
assign n_13440 = n_2165 ^ n_13316;
assign n_13441 = n_765 ^ n_13317;
assign n_13442 = n_2236 ^ n_13318;
assign n_13443 = n_2304 ^ n_13319;
assign n_13444 = n_2371 ^ n_13320;
assign n_13445 = n_2438 ^ n_13321;
assign n_13446 = n_2505 ^ n_13322;
assign n_13447 = n_2571 ^ n_13323;
assign n_13448 = n_2636 ^ n_13324;
assign n_13449 = n_2703 ^ n_13325;
assign n_13450 = n_2771 ^ n_13326;
assign n_13451 = n_2838 ^ n_13327;
assign n_13452 = n_2906 ^ n_13328;
assign n_13453 = n_2972 ^ n_13329;
assign n_13454 = n_3041 ^ n_13330;
assign n_13455 = n_3107 ^ n_13331;
assign n_13456 = n_3176 ^ n_13332;
assign n_13457 = n_3240 ^ n_13333;
assign n_13458 = n_3305 ^ n_13334;
assign n_13459 = n_3370 ^ n_13335;
assign n_13460 = n_13336 ^ x5;
assign n_13461 = n_13337 ^ x8;
assign n_13462 = n_13338 ^ x11;
assign n_13463 = n_13339 ^ x14;
assign n_13464 = n_13340 ^ x17;
assign n_13465 = n_13341 ^ x20;
assign n_13466 = n_13342 ^ x23;
assign n_13467 = n_13343 ^ x26;
assign n_13468 = n_13344 ^ x29;
assign n_13469 = n_13345 ^ x32;
assign n_13470 = n_13346 ^ x35;
assign n_13471 = n_13347 ^ x38;
assign n_13472 = n_13348 ^ x41;
assign n_13473 = n_13349 ^ x44;
assign n_13474 = n_13350 ^ x47;
assign n_13475 = n_13351 ^ x50;
assign n_13476 = n_13352 ^ x53;
assign n_13477 = n_13353 ^ x56;
assign n_13478 = n_13354 ^ x59;
assign n_13479 = n_13355 ^ x62;
assign n_13480 = n_13356 ^ n_13129;
assign n_13481 = n_13357 ^ n_13130;
assign n_13482 = n_13358 ^ n_12898;
assign n_13483 = n_13359 ^ n_13132;
assign n_13484 = n_13360 ^ n_12900;
assign n_13485 = n_13361 ^ n_12901;
assign n_13486 = n_13363 ^ n_12902;
assign n_13487 = n_13365 ^ n_13136;
assign n_13488 = n_13367 ^ n_12904;
assign n_13489 = n_13368 ^ n_3503;
assign n_13490 = n_13368 & ~n_4974;
assign n_13491 = n_13369 ^ n_9894;
assign n_13492 = ~n_12297 & n_13370;
assign n_13493 = n_13372 ^ n_13141;
assign n_13494 = n_13374 ^ n_13142;
assign n_13495 = n_13376 ^ n_13143;
assign n_13496 = n_13378 ^ n_12197;
assign n_13497 = n_13380 ^ n_13145;
assign n_13498 = n_13382 ^ n_13146;
assign n_13499 = n_13383 ^ n_12618;
assign n_13500 = n_13383 ^ n_12486;
assign n_13501 = n_13385 ^ n_13149;
assign n_13502 = n_13387 ^ n_13150;
assign n_13503 = n_13388 ^ n_13128;
assign n_13504 = ~n_12784 & n_13389;
assign n_13505 = n_13390 ^ n_9893;
assign n_13506 = ~n_12365 & n_13391;
assign y22 = n_13392;
assign n_13507 = ~n_12295 & n_13393;
assign n_13508 = n_13395 ^ n_13156;
assign n_13509 = n_13397 ^ n_13157;
assign n_13510 = n_13399 ^ n_13158;
assign n_13511 = n_13401 ^ n_13159;
assign n_13512 = n_13402 ^ n_12620;
assign n_13513 = n_13402 ^ n_12488;
assign n_13514 = n_13095 & ~n_13404;
assign n_13515 = n_13405 ^ n_13168;
assign n_13516 = n_13406 ^ n_13169;
assign n_13517 = n_13407 ^ n_13170;
assign n_13518 = n_13408 ^ n_13171;
assign n_13519 = n_13410 ^ n_13173;
assign n_13520 = n_13412 ^ n_13174;
assign n_13521 = n_13414 ^ n_13176;
assign n_13522 = n_13416 ^ n_13177;
assign n_13523 = n_13418 ^ n_13178;
assign n_13524 = ~n_13162 & n_13422;
assign n_13525 = n_13163 & ~n_13424;
assign n_13526 = ~n_13164 & n_13426;
assign n_13527 = ~n_13172 & n_13428;
assign n_13528 = n_13429 ^ n_13044;
assign n_13529 = n_13429 & ~n_13165;
assign n_13530 = n_13430 ^ n_13059;
assign n_13531 = n_13430 & ~n_13175;
assign n_13532 = n_13431 ^ n_13061;
assign n_13533 = n_13431 & n_13432;
assign n_13534 = n_13433 ^ n_12933;
assign n_13535 = n_13433 & n_13434;
assign n_13536 = n_13435 ^ n_12818;
assign n_13537 = n_13435 & ~n_13276;
assign n_13538 = n_13436 ^ n_13201;
assign n_13539 = n_13437 ^ x110;
assign n_13540 = x112 & ~n_13438;
assign n_13541 = n_13314 ^ n_13439;
assign n_13542 = x111 & ~n_13439;
assign n_13543 = n_5038 ^ n_13440;
assign n_13544 = n_5101 ^ n_13441;
assign n_13545 = n_5164 ^ n_13442;
assign n_13546 = n_5225 ^ n_13443;
assign n_13547 = n_5289 ^ n_13444;
assign n_13548 = n_5353 ^ n_13445;
assign n_13549 = n_5417 ^ n_13446;
assign n_13550 = n_5481 ^ n_13447;
assign n_13551 = n_5542 ^ n_13448;
assign n_13552 = n_5605 ^ n_13449;
assign n_13553 = n_5668 ^ n_13450;
assign n_13554 = n_5732 ^ n_13451;
assign n_13555 = n_5798 ^ n_13452;
assign n_13556 = n_5860 ^ n_13453;
assign n_13557 = n_5924 ^ n_13454;
assign n_13558 = n_5987 ^ n_13455;
assign n_13559 = n_6051 ^ n_13456;
assign n_13560 = n_6115 ^ n_13457;
assign n_13561 = n_6177 ^ n_13458;
assign n_13562 = n_6239 ^ n_13459;
assign n_13563 = n_13278 ^ n_13469;
assign n_13564 = n_13470 ^ n_13280;
assign n_13565 = n_13471 ^ n_13282;
assign n_13566 = n_13472 ^ n_13284;
assign n_13567 = n_13473 ^ n_13409;
assign n_13568 = n_13474 ^ n_13411;
assign n_13569 = n_13475 ^ n_13413;
assign n_13570 = n_13476 ^ n_13415;
assign n_13571 = n_13477 ^ n_13417;
assign n_13572 = n_13478 ^ n_13403;
assign n_13573 = n_13479 ^ n_6354;
assign n_13574 = n_13421 ^ n_13480;
assign n_13575 = n_13423 ^ n_13481;
assign n_13576 = n_13425 ^ n_13482;
assign n_13577 = n_13427 ^ n_13483;
assign n_13578 = n_13489 ^ n_13311;
assign n_13579 = n_13490 ^ n_3502;
assign n_13580 = n_13492 ^ n_13244;
assign n_13581 = n_13493 ^ n_12607;
assign n_13582 = n_13493 ^ n_12474;
assign n_13583 = n_13494 ^ n_12609;
assign n_13584 = n_13494 ^ n_12476;
assign n_13585 = n_13495 ^ n_12299;
assign n_13586 = n_13495 ^ n_12214;
assign n_13587 = n_13496 ^ n_12613;
assign n_13588 = n_13496 ^ n_9478;
assign n_13589 = n_13497 ^ n_12615;
assign n_13590 = n_13497 ^ n_12482;
assign n_13591 = n_13498 ^ n_12484;
assign n_13592 = n_13498 ^ n_12373;
assign n_13593 = n_13499 ^ n_9904;
assign n_13594 = ~n_12618 & n_13500;
assign n_13595 = n_13501 ^ n_12501;
assign n_13596 = n_13501 ^ n_12387;
assign n_13597 = n_13502 ^ n_12377;
assign n_13598 = n_13502 ^ n_12289;
assign n_13599 = n_13504 ^ n_13263;
assign n_13600 = n_13506 ^ n_13264;
assign n_13601 = n_13507 ^ n_13265;
assign n_13602 = n_13508 ^ n_12756;
assign n_13603 = n_13508 ^ n_12624;
assign n_13604 = n_13509 ^ n_13003;
assign n_13605 = n_13509 ^ n_12865;
assign n_13606 = n_13510 ^ n_12634;
assign n_13607 = n_13510 ^ n_12499;
assign n_13608 = n_13511 ^ n_13009;
assign n_13609 = n_13511 ^ n_12871;
assign n_13610 = n_13512 ^ n_10789;
assign n_13611 = n_12620 & ~n_13513;
assign n_13612 = n_13514 ^ n_13277;
assign n_13613 = n_13517 ^ n_13229;
assign n_13614 = n_13520 ^ n_13235;
assign n_13615 = n_13524 ^ n_13302;
assign n_13616 = n_13525 ^ n_13303;
assign n_13617 = n_13526 ^ n_13304;
assign n_13618 = n_13527 ^ n_13042;
assign n_13619 = n_13528 ^ n_13484;
assign n_13620 = n_13529 ^ n_13306;
assign n_13621 = n_13530 ^ n_13485;
assign n_13622 = n_13531 ^ n_13307;
assign n_13623 = n_13532 ^ n_13486;
assign n_13624 = n_13533 ^ n_13047;
assign n_13625 = n_13487 ^ n_13534;
assign n_13626 = n_13535 ^ n_13049;
assign n_13627 = n_13488 ^ n_13536;
assign n_13628 = n_13537 ^ n_13310;
assign n_13629 = n_13539 ^ n_6491;
assign n_13630 = ~x113 & ~n_13540;
assign n_13631 = n_1 & n_13541;
assign n_13632 = n_13541 ^ x111;
assign n_13633 = n_13438 ^ n_13542;
assign n_13634 = ~x112 & ~n_13542;
assign n_13635 = n_13543 ^ x5;
assign n_13636 = n_13544 ^ x8;
assign n_13637 = n_13545 ^ x11;
assign n_13638 = n_13546 ^ x14;
assign n_13639 = n_13547 ^ x17;
assign n_13640 = n_13548 ^ x20;
assign n_13641 = n_13549 ^ x23;
assign n_13642 = n_13550 ^ x26;
assign n_13643 = n_13551 ^ x29;
assign n_13644 = n_13552 ^ x32;
assign n_13645 = n_13553 ^ x35;
assign n_13646 = n_13554 ^ x38;
assign n_13647 = n_13555 ^ x41;
assign n_13648 = n_13556 ^ x44;
assign n_13649 = n_13557 ^ x47;
assign n_13650 = n_13558 ^ x50;
assign n_13651 = n_13559 ^ x53;
assign n_13652 = n_13560 ^ x56;
assign n_13653 = n_13561 ^ x59;
assign n_13654 = n_13562 ^ x62;
assign n_13655 = n_13579 ^ n_13479;
assign n_13656 = n_13580 ^ n_12630;
assign n_13657 = n_13580 ^ n_12495;
assign n_13658 = n_13581 ^ n_9896;
assign n_13659 = ~n_12607 & n_13582;
assign n_13660 = n_13583 ^ n_9897;
assign n_13661 = ~n_12609 & n_13584;
assign n_13662 = n_13585 ^ n_9898;
assign n_13663 = ~n_12299 & n_13586;
assign n_13664 = n_13587 ^ n_9901;
assign n_13665 = n_12613 & ~n_13588;
assign n_13666 = n_13589 ^ n_9902;
assign n_13667 = ~n_12615 & n_13590;
assign n_13668 = n_13591 ^ n_9903;
assign n_13669 = ~n_12484 & n_13592;
assign n_13670 = n_13594 ^ n_13383;
assign n_13671 = n_13595 ^ n_9905;
assign n_13672 = ~n_12501 & n_13596;
assign n_13673 = n_13597 ^ n_11891;
assign n_13674 = n_12377 & ~n_13598;
assign n_13675 = n_13599 ^ n_13420;
assign n_13676 = n_13599 ^ n_13051;
assign n_13677 = n_13600 ^ n_12742;
assign n_13678 = n_13600 ^ n_12603;
assign n_13679 = n_13601 ^ n_12628;
assign n_13680 = n_13601 ^ n_12493;
assign n_13681 = n_13602 ^ n_10109;
assign n_13682 = ~n_12756 & n_13603;
assign n_13683 = n_13604 ^ n_10041;
assign n_13684 = ~n_13003 & n_13605;
assign n_13685 = n_13606 ^ n_10045;
assign n_13686 = n_12634 & ~n_13607;
assign n_13687 = n_13608 ^ n_10046;
assign n_13688 = ~n_13009 & n_13609;
assign n_13689 = n_13611 ^ n_13402;
assign n_13690 = n_13615 ^ n_13564;
assign n_13691 = n_13615 ^ n_13470;
assign n_13692 = n_13616 ^ n_13565;
assign n_13693 = n_13616 ^ n_13471;
assign n_13694 = n_13617 ^ n_13566;
assign n_13695 = n_13617 ^ n_13284;
assign n_13696 = n_13618 ^ n_13567;
assign n_13697 = n_13618 ^ n_13473;
assign n_13698 = n_13620 ^ n_13568;
assign n_13699 = n_13620 ^ n_13474;
assign n_13700 = n_13622 ^ n_13475;
assign n_13701 = n_13624 ^ n_13476;
assign n_13702 = n_13626 ^ n_13477;
assign n_13703 = n_13628 ^ n_13478;
assign n_13704 = ~x0 & ~n_13629;
assign n_13705 = x114 & ~n_13630;
assign n_13706 = n_13631 ^ x1;
assign n_13707 = n_655 & ~n_13632;
assign n_13708 = n_784 & ~n_13632;
assign n_13709 = ~n_3665 & ~n_13632;
assign n_13710 = n_854 & ~n_13632;
assign n_13711 = n_920 & ~n_13632;
assign n_13712 = n_986 & ~n_13632;
assign n_13713 = n_1052 & ~n_13632;
assign n_13714 = n_1117 & ~n_13632;
assign n_13715 = n_1181 & ~n_13632;
assign n_13716 = n_1248 & ~n_13632;
assign n_13717 = n_1314 & ~n_13632;
assign n_13718 = n_1380 & ~n_13632;
assign n_13719 = n_1445 & ~n_13632;
assign n_13720 = n_1510 & ~n_13632;
assign n_13721 = n_1576 & ~n_13632;
assign n_13722 = ~n_13632 & n_1641;
assign n_13723 = ~n_13632 & n_1706;
assign n_13724 = ~n_13632 & n_1771;
assign n_13725 = ~n_13632 & n_1835;
assign n_13726 = ~n_13632 & n_1899;
assign n_13727 = n_1 & n_13633;
assign n_13728 = n_13633 ^ x112;
assign n_13729 = n_13540 ^ n_13634;
assign n_13730 = x113 & ~n_13634;
assign n_13731 = n_13644 ^ n_13225;
assign n_13732 = n_13644 ^ n_13515;
assign n_13733 = n_13645 ^ n_13516;
assign n_13734 = n_13645 ^ n_13227;
assign n_13735 = n_13646 ^ n_13613;
assign n_13736 = n_13646 ^ n_13229;
assign n_13737 = n_13647 ^ n_13231;
assign n_13738 = n_13647 ^ n_13518;
assign n_13739 = n_13648 ^ n_13233;
assign n_13740 = n_13648 ^ n_13519;
assign n_13741 = n_13649 ^ n_13614;
assign n_13742 = n_13649 ^ n_13235;
assign n_13743 = n_13650 ^ n_13521;
assign n_13744 = n_13650 ^ n_13362;
assign n_13745 = n_13651 ^ n_13522;
assign n_13746 = n_13651 ^ n_13364;
assign n_13747 = n_13652 ^ n_13523;
assign n_13748 = n_13652 ^ n_13366;
assign n_13749 = n_13653 ^ n_13242;
assign n_13750 = n_13653 ^ n_13612;
assign n_13751 = n_13654 ^ n_6607;
assign n_13752 = n_13654 ^ n_6489;
assign n_13753 = n_13655 ^ n_6354;
assign n_13754 = ~n_13655 & n_13573;
assign n_13755 = n_13656 ^ n_10040;
assign n_13756 = ~n_12630 & n_13657;
assign n_13757 = n_13659 ^ n_13493;
assign n_13758 = n_13661 ^ n_13494;
assign n_13759 = n_13663 ^ n_13495;
assign n_13760 = n_13665 ^ n_12480;
assign n_13761 = n_13667 ^ n_13497;
assign n_13762 = n_13669 ^ n_13498;
assign n_13763 = n_13670 ^ n_13016;
assign n_13764 = n_13670 ^ n_12879;
assign n_13765 = n_13672 ^ n_13501;
assign n_13766 = n_13674 ^ n_13502;
assign n_13767 = ~n_13420 & n_13676;
assign n_13768 = n_13677 ^ n_10039;
assign n_13769 = n_12742 & ~n_13678;
assign y23 = n_13679;
assign n_13770 = ~n_12628 & n_13680;
assign n_13771 = n_13682 ^ n_13508;
assign n_13772 = n_13684 ^ n_13509;
assign n_13773 = n_13686 ^ n_13510;
assign n_13774 = n_13688 ^ n_13511;
assign n_13775 = n_13689 ^ n_13018;
assign n_13776 = n_13689 ^ n_12881;
assign n_13777 = ~n_13564 & n_13691;
assign n_13778 = n_13565 & n_13693;
assign n_13779 = ~n_13566 & n_13695;
assign n_13780 = ~n_13567 & ~n_13697;
assign n_13781 = ~n_13568 & ~n_13699;
assign n_13782 = n_13700 ^ n_13413;
assign n_13783 = n_13700 & ~n_13569;
assign n_13784 = n_13701 ^ n_13415;
assign n_13785 = n_13701 & ~n_13570;
assign n_13786 = n_13702 ^ n_13417;
assign n_13787 = n_13702 & n_13571;
assign n_13788 = n_13703 ^ n_13403;
assign n_13789 = n_13703 & ~n_13572;
assign n_13790 = n_13704 ^ n_13539;
assign n_13791 = ~x115 & ~n_13705;
assign n_13792 = n_13706 ^ x111;
assign n_13793 = n_2166 ^ n_13707;
assign n_13794 = n_766 ^ n_13708;
assign n_13795 = n_2237 ^ n_13709;
assign n_13796 = n_2305 ^ n_13710;
assign n_13797 = n_2372 ^ n_13711;
assign n_13798 = n_2439 ^ n_13712;
assign n_13799 = n_2506 ^ n_13713;
assign n_13800 = n_2572 ^ n_13714;
assign n_13801 = n_2637 ^ n_13715;
assign n_13802 = n_2704 ^ n_13716;
assign n_13803 = n_2772 ^ n_13717;
assign n_13804 = n_2839 ^ n_13718;
assign n_13805 = n_2907 ^ n_13719;
assign n_13806 = n_2973 ^ n_13720;
assign n_13807 = n_3042 ^ n_13721;
assign n_13808 = n_3108 ^ n_13722;
assign n_13809 = n_3177 ^ n_13723;
assign n_13810 = n_3241 ^ n_13724;
assign n_13811 = n_3306 ^ n_13725;
assign n_13812 = n_3371 ^ n_13726;
assign n_13813 = n_13727 ^ x1;
assign n_13814 = n_655 & ~n_13728;
assign n_13815 = n_784 & ~n_13728;
assign n_13816 = ~n_3665 & ~n_13728;
assign n_13817 = n_854 & ~n_13728;
assign n_13818 = n_920 & ~n_13728;
assign n_13819 = n_986 & ~n_13728;
assign n_13820 = n_1052 & ~n_13728;
assign n_13821 = n_1117 & ~n_13728;
assign n_13822 = n_1181 & ~n_13728;
assign n_13823 = n_1248 & ~n_13728;
assign n_13824 = n_1314 & ~n_13728;
assign n_13825 = n_1380 & ~n_13728;
assign n_13826 = n_1445 & ~n_13728;
assign n_13827 = n_1510 & ~n_13728;
assign n_13828 = n_1576 & ~n_13728;
assign n_13829 = n_1641 & ~n_13728;
assign n_13830 = ~n_13728 & n_1706;
assign n_13831 = ~n_13728 & n_1771;
assign n_13832 = ~n_13728 & n_1835;
assign n_13833 = ~n_13728 & n_1899;
assign n_13834 = n_1 & n_13729;
assign n_13835 = n_13729 ^ x113;
assign n_13836 = n_13630 ^ n_13730;
assign n_13837 = ~x114 & ~n_13730;
assign n_13838 = n_13731 ^ n_13515;
assign n_13839 = n_13731 & n_13732;
assign n_13840 = n_13733 ^ n_13227;
assign n_13841 = n_13733 & ~n_13734;
assign n_13842 = n_13613 & ~n_13736;
assign n_13843 = n_13737 ^ n_13518;
assign n_13844 = n_13737 & n_13738;
assign n_13845 = n_13739 ^ n_13519;
assign n_13846 = n_13739 & n_13740;
assign n_13847 = ~n_13614 & n_13742;
assign n_13848 = n_13743 ^ n_13362;
assign n_13849 = n_13743 & ~n_13744;
assign n_13850 = n_13745 ^ n_13364;
assign n_13851 = n_13745 & n_13746;
assign n_13852 = n_13747 ^ n_13366;
assign n_13853 = n_13747 & n_13748;
assign n_13854 = n_13749 ^ n_13612;
assign n_13855 = ~n_13749 & ~n_13750;
assign n_13856 = ~n_6607 & ~n_13752;
assign n_13857 = n_13754 ^ n_13579;
assign n_13858 = n_13756 ^ n_13580;
assign n_13859 = n_13757 ^ n_13005;
assign n_13860 = n_13757 ^ n_12867;
assign n_13861 = n_13758 ^ n_13007;
assign n_13862 = n_13758 ^ n_12869;
assign n_13863 = n_13759 ^ n_12632;
assign n_13864 = n_13759 ^ n_12497;
assign n_13865 = n_13760 ^ n_13011;
assign n_13866 = n_13760 ^ n_12873;
assign n_13867 = n_13761 ^ n_13013;
assign n_13868 = n_13761 ^ n_12875;
assign n_13869 = n_13762 ^ n_12877;
assign n_13870 = n_13762 ^ n_12750;
assign n_13871 = n_13763 ^ n_10050;
assign n_13872 = ~n_13016 & n_13764;
assign n_13873 = n_13765 ^ n_12894;
assign n_13874 = n_13765 ^ n_12763;
assign n_13875 = n_13766 ^ n_12754;
assign n_13876 = n_13766 ^ n_12622;
assign n_13877 = n_13767 ^ n_13599;
assign n_13878 = n_13769 ^ n_13600;
assign n_13879 = n_13770 ^ n_13601;
assign n_13880 = n_13771 ^ n_13153;
assign n_13881 = n_13771 ^ n_13022;
assign n_13882 = n_13772 ^ n_13371;
assign n_13883 = n_13772 ^ n_13245;
assign n_13884 = n_13773 ^ n_13032;
assign n_13885 = n_13773 ^ n_12892;
assign n_13886 = n_13774 ^ n_13377;
assign n_13887 = n_13774 ^ n_13251;
assign n_13888 = n_13775 ^ n_11640;
assign n_13889 = ~n_13018 & n_13776;
assign n_13890 = n_13777 ^ n_13615;
assign n_13891 = n_13778 ^ n_13616;
assign n_13892 = n_13779 ^ n_13472;
assign n_13893 = n_13780 ^ n_13409;
assign n_13894 = n_13781 ^ n_13411;
assign n_13895 = n_13783 ^ n_13622;
assign n_13896 = n_13785 ^ n_13624;
assign n_13897 = n_13787 ^ n_13626;
assign n_13898 = n_13789 ^ n_13628;
assign n_13899 = x116 & ~n_13791;
assign n_13900 = n_13792 ^ n_3514;
assign n_13901 = n_5039 ^ n_13793;
assign n_13902 = n_5102 ^ n_13794;
assign n_13903 = n_5165 ^ n_13795;
assign n_13904 = n_5226 ^ n_13796;
assign n_13905 = n_5290 ^ n_13797;
assign n_13906 = n_5354 ^ n_13798;
assign n_13907 = n_5418 ^ n_13799;
assign n_13908 = n_5482 ^ n_13800;
assign n_13909 = n_5543 ^ n_13801;
assign n_13910 = n_5606 ^ n_13802;
assign n_13911 = n_5669 ^ n_13803;
assign n_13912 = n_5733 ^ n_13804;
assign n_13913 = n_5799 ^ n_13805;
assign n_13914 = n_5861 ^ n_13806;
assign n_13915 = n_5925 ^ n_13807;
assign n_13916 = n_5988 ^ n_13808;
assign n_13917 = n_6052 ^ n_13809;
assign n_13918 = n_6116 ^ n_13810;
assign n_13919 = n_6178 ^ n_13811;
assign n_13920 = n_6240 ^ n_13812;
assign n_13921 = n_13813 ^ x112;
assign n_13922 = n_2167 ^ n_13814;
assign n_13923 = n_767 ^ n_13815;
assign n_13924 = n_2238 ^ n_13816;
assign n_13925 = n_2306 ^ n_13817;
assign n_13926 = n_2373 ^ n_13818;
assign n_13927 = n_2440 ^ n_13819;
assign n_13928 = n_2507 ^ n_13820;
assign n_13929 = n_2573 ^ n_13821;
assign n_13930 = n_2638 ^ n_13822;
assign n_13931 = n_2705 ^ n_13823;
assign n_13932 = n_2773 ^ n_13824;
assign n_13933 = n_2840 ^ n_13825;
assign n_13934 = n_2908 ^ n_13826;
assign n_13935 = n_2974 ^ n_13827;
assign n_13936 = n_3043 ^ n_13828;
assign n_13937 = n_3109 ^ n_13829;
assign n_13938 = n_3178 ^ n_13830;
assign n_13939 = n_3242 ^ n_13831;
assign n_13940 = n_3307 ^ n_13832;
assign n_13941 = n_3372 ^ n_13833;
assign n_13942 = n_13834 ^ x1;
assign n_13943 = n_655 & ~n_13835;
assign n_13944 = n_784 & ~n_13835;
assign n_13945 = ~n_3665 & ~n_13835;
assign n_13946 = n_854 & ~n_13835;
assign n_13947 = n_920 & ~n_13835;
assign n_13948 = n_986 & ~n_13835;
assign n_13949 = n_1052 & ~n_13835;
assign n_13950 = n_1117 & ~n_13835;
assign n_13951 = n_1181 & ~n_13835;
assign n_13952 = n_1248 & ~n_13835;
assign n_13953 = n_1314 & ~n_13835;
assign n_13954 = n_1380 & ~n_13835;
assign n_13955 = n_1445 & ~n_13835;
assign n_13956 = n_1510 & ~n_13835;
assign n_13957 = n_1576 & ~n_13835;
assign n_13958 = n_1641 & ~n_13835;
assign n_13959 = ~n_13835 & n_1706;
assign n_13960 = ~n_13835 & n_1771;
assign n_13961 = ~n_13835 & n_1835;
assign n_13962 = ~n_13835 & n_1899;
assign n_13963 = n_1 & n_13836;
assign n_13964 = n_13836 ^ x114;
assign n_13965 = n_13705 ^ n_13837;
assign n_13966 = x115 & ~n_13837;
assign n_13967 = n_13839 ^ n_13515;
assign n_13968 = n_13841 ^ n_13516;
assign n_13969 = n_13842 ^ n_13517;
assign n_13970 = n_13844 ^ n_13518;
assign n_13971 = n_13846 ^ n_13519;
assign n_13972 = n_13847 ^ n_13520;
assign n_13973 = n_13849 ^ n_13521;
assign n_13974 = n_13851 ^ n_13522;
assign n_13975 = n_13853 ^ n_13523;
assign n_13976 = n_13855 ^ n_13612;
assign n_13977 = n_13856 ^ n_13654;
assign n_13978 = n_13857 ^ n_13751;
assign n_13979 = n_13858 ^ n_13028;
assign n_13980 = n_13858 ^ n_12888;
assign n_13981 = n_13859 ^ n_10042;
assign n_13982 = ~n_13005 & n_13860;
assign n_13983 = n_13861 ^ n_10043;
assign n_13984 = ~n_13007 & n_13862;
assign n_13985 = n_13863 ^ n_10044;
assign n_13986 = ~n_12632 & n_13864;
assign n_13987 = n_13865 ^ n_10047;
assign n_13988 = ~n_13011 & n_13866;
assign n_13989 = n_13867 ^ n_10048;
assign n_13990 = ~n_13013 & n_13868;
assign n_13991 = n_13869 ^ n_10049;
assign n_13992 = ~n_12877 & n_13870;
assign n_13993 = n_13872 ^ n_13670;
assign n_13994 = n_13873 ^ n_10051;
assign n_13995 = ~n_12894 & n_13874;
assign n_13996 = n_13875 ^ n_12808;
assign n_13997 = n_12754 & ~n_13876;
assign n_13998 = n_13877 ^ n_13563;
assign n_13999 = n_13877 ^ n_13278;
assign n_14000 = n_13878 ^ n_13139;
assign n_14001 = n_13878 ^ n_13001;
assign n_14002 = n_13879 ^ n_13026;
assign n_14003 = n_13879 ^ n_12886;
assign n_14004 = n_13880 ^ n_10238;
assign n_14005 = n_13153 & ~n_13881;
assign n_14006 = n_13882 ^ n_10158;
assign n_14007 = ~n_13371 & n_13883;
assign n_14008 = n_13884 ^ n_10162;
assign n_14009 = n_13032 & ~n_13885;
assign n_14010 = n_13886 ^ n_10163;
assign n_14011 = ~n_13377 & n_13887;
assign n_14012 = n_13889 ^ n_13689;
assign n_14013 = n_13840 ^ n_13890;
assign n_14014 = n_13735 ^ n_13891;
assign n_14015 = n_13843 ^ n_13892;
assign n_14016 = n_13845 ^ n_13893;
assign n_14017 = n_13741 ^ n_13894;
assign n_14018 = n_13848 ^ n_13895;
assign n_14019 = n_13896 ^ n_13850;
assign n_14020 = n_13897 ^ n_13852;
assign n_14021 = n_13898 ^ n_13854;
assign n_14022 = ~x117 & ~n_13899;
assign n_14023 = ~x0 & n_13900;
assign n_14024 = n_13901 ^ x5;
assign n_14025 = n_13902 ^ x8;
assign n_14026 = n_13903 ^ x11;
assign n_14027 = n_13904 ^ x14;
assign n_14028 = n_13905 ^ x17;
assign n_14029 = n_13906 ^ x20;
assign n_14030 = n_13907 ^ x23;
assign n_14031 = n_13908 ^ x26;
assign n_14032 = n_13909 ^ x29;
assign n_14033 = n_13910 ^ x32;
assign n_14034 = n_13911 ^ x35;
assign n_14035 = n_13912 ^ x38;
assign n_14036 = n_13913 ^ x41;
assign n_14037 = n_13914 ^ x44;
assign n_14038 = n_13915 ^ x47;
assign n_14039 = n_13916 ^ x50;
assign n_14040 = n_13917 ^ x53;
assign n_14041 = n_13918 ^ x56;
assign n_14042 = n_13919 ^ x59;
assign n_14043 = n_4977 ^ n_13920;
assign n_14044 = n_13920 ^ x107;
assign n_14045 = n_2077 ^ n_13920;
assign n_14046 = n_13921 ^ n_3515;
assign n_14047 = n_5040 ^ n_13922;
assign n_14048 = n_5103 ^ n_13923;
assign n_14049 = n_5166 ^ n_13924;
assign n_14050 = n_5227 ^ n_13925;
assign n_14051 = n_5291 ^ n_13926;
assign n_14052 = n_5355 ^ n_13927;
assign n_14053 = n_5419 ^ n_13928;
assign n_14054 = n_5483 ^ n_13929;
assign n_14055 = n_5544 ^ n_13930;
assign n_14056 = n_5607 ^ n_13931;
assign n_14057 = n_5670 ^ n_13932;
assign n_14058 = n_5734 ^ n_13933;
assign n_14059 = n_5800 ^ n_13934;
assign n_14060 = n_5862 ^ n_13935;
assign n_14061 = n_5926 ^ n_13936;
assign n_14062 = n_5989 ^ n_13937;
assign n_14063 = n_6053 ^ n_13938;
assign n_14064 = n_6117 ^ n_13939;
assign n_14065 = n_6179 ^ n_13940;
assign n_14066 = n_6241 ^ n_13941;
assign n_14067 = n_13942 ^ x113;
assign n_14068 = n_2168 ^ n_13943;
assign n_14069 = n_768 ^ n_13944;
assign n_14070 = n_2239 ^ n_13945;
assign n_14071 = n_2307 ^ n_13946;
assign n_14072 = n_2374 ^ n_13947;
assign n_14073 = n_2441 ^ n_13948;
assign n_14074 = n_2508 ^ n_13949;
assign n_14075 = n_2574 ^ n_13950;
assign n_14076 = n_2639 ^ n_13951;
assign n_14077 = n_2706 ^ n_13952;
assign n_14078 = n_2774 ^ n_13953;
assign n_14079 = n_2841 ^ n_13954;
assign n_14080 = n_2909 ^ n_13955;
assign n_14081 = n_2975 ^ n_13956;
assign n_14082 = n_3044 ^ n_13957;
assign n_14083 = n_3110 ^ n_13958;
assign n_14084 = n_3179 ^ n_13959;
assign n_14085 = n_3243 ^ n_13960;
assign n_14086 = n_3308 ^ n_13961;
assign n_14087 = n_3373 ^ n_13962;
assign n_14088 = n_13963 ^ x1;
assign n_14089 = n_655 & ~n_13964;
assign n_14090 = n_784 & ~n_13964;
assign n_14091 = ~n_3665 & ~n_13964;
assign n_14092 = n_854 & ~n_13964;
assign n_14093 = n_920 & ~n_13964;
assign n_14094 = n_986 & ~n_13964;
assign n_14095 = n_1052 & ~n_13964;
assign n_14096 = n_1117 & ~n_13964;
assign n_14097 = n_1181 & ~n_13964;
assign n_14098 = n_1248 & ~n_13964;
assign n_14099 = n_1314 & ~n_13964;
assign n_14100 = n_1380 & ~n_13964;
assign n_14101 = n_1445 & ~n_13964;
assign n_14102 = n_1510 & ~n_13964;
assign n_14103 = n_1576 & ~n_13964;
assign n_14104 = n_1641 & ~n_13964;
assign n_14105 = ~n_13964 & n_1706;
assign n_14106 = ~n_13964 & n_1771;
assign n_14107 = ~n_13964 & n_1835;
assign n_14108 = ~n_13964 & n_1899;
assign n_14109 = n_1 & n_13965;
assign n_14110 = n_13965 ^ x115;
assign n_14111 = n_13791 ^ n_13966;
assign n_14112 = ~x116 & ~n_13966;
assign n_14113 = n_13979 ^ n_10157;
assign n_14114 = ~n_13028 & n_13980;
assign n_14115 = n_13982 ^ n_13757;
assign n_14116 = n_13984 ^ n_13758;
assign n_14117 = n_13986 ^ n_13759;
assign n_14118 = n_13988 ^ n_13760;
assign n_14119 = n_13990 ^ n_13761;
assign n_14120 = n_13992 ^ n_13762;
assign n_14121 = n_13993 ^ n_13384;
assign n_14122 = n_13993 ^ n_13259;
assign n_14123 = n_13995 ^ n_13765;
assign n_14124 = n_13997 ^ n_13766;
assign n_14125 = ~n_13563 & n_13999;
assign n_14126 = n_14000 ^ n_10156;
assign n_14127 = ~n_13139 & n_14001;
assign y24 = n_14002;
assign n_14128 = ~n_13026 & n_14003;
assign n_14129 = n_14005 ^ n_13771;
assign n_14130 = n_14007 ^ n_13772;
assign n_14131 = n_14009 ^ n_13773;
assign n_14132 = n_14011 ^ n_13774;
assign n_14133 = n_14012 ^ n_13386;
assign n_14134 = n_14012 ^ n_13261;
assign n_14135 = n_14023 ^ n_13792;
assign n_14136 = n_13675 ^ n_14032;
assign n_14137 = n_14033 ^ n_13574;
assign n_14138 = n_14033 ^ n_13480;
assign n_14139 = n_14034 ^ n_13575;
assign n_14140 = n_14034 ^ n_13481;
assign n_14141 = n_14035 ^ n_13576;
assign n_14142 = n_14035 ^ n_13482;
assign n_14143 = n_14036 ^ n_13577;
assign n_14144 = n_14036 ^ n_13483;
assign n_14145 = n_14037 ^ n_13619;
assign n_14146 = n_14037 ^ n_13484;
assign n_14147 = n_14038 ^ n_13621;
assign n_14148 = n_14038 ^ n_13485;
assign n_14149 = n_14039 ^ n_13623;
assign n_14150 = n_14039 ^ n_13486;
assign n_14151 = n_14040 ^ n_13487;
assign n_14152 = n_14041 ^ n_13488;
assign n_14153 = n_14042 ^ n_13578;
assign n_14154 = n_14042 ^ n_13489;
assign n_14155 = n_13977 ^ n_14043;
assign n_14156 = ~n_242 & ~n_14044;
assign n_14157 = ~n_2077 & n_14045;
assign n_14158 = ~x0 & n_14046;
assign n_14159 = n_14047 ^ x5;
assign n_14160 = n_14048 ^ x8;
assign n_14161 = n_14049 ^ x11;
assign n_14162 = n_14050 ^ x14;
assign n_14163 = n_14051 ^ x17;
assign n_14164 = n_14052 ^ x20;
assign n_14165 = n_14053 ^ x23;
assign n_14166 = n_14054 ^ x26;
assign n_14167 = n_14055 ^ x29;
assign n_14168 = n_14056 ^ x32;
assign n_14169 = n_14057 ^ x35;
assign n_14170 = n_14058 ^ x38;
assign n_14171 = n_14059 ^ x41;
assign n_14172 = n_14060 ^ x44;
assign n_14173 = n_14061 ^ x47;
assign n_14174 = n_14062 ^ x50;
assign n_14175 = n_14063 ^ x53;
assign n_14176 = n_14064 ^ x56;
assign n_14177 = n_14065 ^ x59;
assign n_14178 = n_14066 ^ x62;
assign n_14179 = n_14067 ^ n_2112;
assign n_14180 = n_5041 ^ n_14068;
assign n_14181 = n_5104 ^ n_14069;
assign n_14182 = n_5167 ^ n_14070;
assign n_14183 = n_5228 ^ n_14071;
assign n_14184 = n_5292 ^ n_14072;
assign n_14185 = n_5356 ^ n_14073;
assign n_14186 = n_5420 ^ n_14074;
assign n_14187 = n_5484 ^ n_14075;
assign n_14188 = n_5545 ^ n_14076;
assign n_14189 = n_5608 ^ n_14077;
assign n_14190 = n_5671 ^ n_14078;
assign n_14191 = n_5735 ^ n_14079;
assign n_14192 = n_5801 ^ n_14080;
assign n_14193 = n_5863 ^ n_14081;
assign n_14194 = n_5927 ^ n_14082;
assign n_14195 = n_5990 ^ n_14083;
assign n_14196 = n_6054 ^ n_14084;
assign n_14197 = n_6118 ^ n_14085;
assign n_14198 = n_6180 ^ n_14086;
assign n_14199 = n_6242 ^ n_14087;
assign n_14200 = n_14088 ^ x114;
assign n_14201 = n_2169 ^ n_14089;
assign n_14202 = n_769 ^ n_14090;
assign n_14203 = n_2240 ^ n_14091;
assign n_14204 = n_2308 ^ n_14092;
assign n_14205 = n_2375 ^ n_14093;
assign n_14206 = n_2442 ^ n_14094;
assign n_14207 = n_2509 ^ n_14095;
assign n_14208 = n_2575 ^ n_14096;
assign n_14209 = n_2640 ^ n_14097;
assign n_14210 = n_2707 ^ n_14098;
assign n_14211 = n_2775 ^ n_14099;
assign n_14212 = n_2842 ^ n_14100;
assign n_14213 = n_2910 ^ n_14101;
assign n_14214 = n_2976 ^ n_14102;
assign n_14215 = n_3045 ^ n_14103;
assign n_14216 = n_3111 ^ n_14104;
assign n_14217 = n_3180 ^ n_14105;
assign n_14218 = n_3244 ^ n_14106;
assign n_14219 = n_3309 ^ n_14107;
assign n_14220 = n_3374 ^ n_14108;
assign n_14221 = n_14109 ^ x1;
assign n_14222 = n_655 & ~n_14110;
assign n_14223 = n_784 & ~n_14110;
assign n_14224 = ~n_3665 & ~n_14110;
assign n_14225 = n_854 & ~n_14110;
assign n_14226 = n_920 & ~n_14110;
assign n_14227 = n_986 & ~n_14110;
assign n_14228 = n_1052 & ~n_14110;
assign n_14229 = n_1117 & ~n_14110;
assign n_14230 = n_1181 & ~n_14110;
assign n_14231 = n_1248 & ~n_14110;
assign n_14232 = n_1314 & ~n_14110;
assign n_14233 = n_1380 & ~n_14110;
assign n_14234 = n_1445 & ~n_14110;
assign n_14235 = n_1510 & ~n_14110;
assign n_14236 = n_1576 & ~n_14110;
assign n_14237 = n_1641 & ~n_14110;
assign n_14238 = n_1706 & ~n_14110;
assign n_14239 = ~n_14110 & n_1771;
assign n_14240 = ~n_14110 & n_1835;
assign n_14241 = ~n_14110 & n_1899;
assign n_14242 = n_1 & n_14111;
assign n_14243 = n_14111 ^ x116;
assign n_14244 = n_13899 ^ n_14112;
assign n_14245 = x117 & ~n_14112;
assign n_14246 = n_14114 ^ n_13858;
assign n_14247 = n_14115 ^ n_13373;
assign n_14248 = n_14115 ^ n_13247;
assign n_14249 = n_14116 ^ n_13375;
assign n_14250 = n_14116 ^ n_13249;
assign n_14251 = n_14117 ^ n_13030;
assign n_14252 = n_14117 ^ n_12890;
assign n_14253 = n_14118 ^ n_13379;
assign n_14254 = n_14118 ^ n_13253;
assign n_14255 = n_14119 ^ n_13381;
assign n_14256 = n_14119 ^ n_13255;
assign n_14257 = n_14120 ^ n_13257;
assign n_14258 = n_14120 ^ n_13147;
assign n_14259 = n_14121 ^ n_10167;
assign n_14260 = ~n_13384 & n_14122;
assign n_14261 = n_14123 ^ n_13274;
assign n_14262 = n_14123 ^ n_13160;
assign n_14263 = n_14124 ^ n_13151;
assign n_14264 = n_14124 ^ n_13020;
assign n_14265 = n_14125 ^ n_13877;
assign n_14266 = n_14127 ^ n_13878;
assign n_14267 = n_14128 ^ n_13879;
assign n_14268 = n_14129 ^ n_13505;
assign n_14269 = n_14129 ^ n_13390;
assign n_14270 = n_14130 ^ n_13658;
assign n_14271 = n_14130 ^ n_13581;
assign n_14272 = n_14131 ^ n_13400;
assign n_14273 = n_14131 ^ n_13272;
assign n_14274 = n_14132 ^ n_13664;
assign n_14275 = n_14132 ^ n_13587;
assign n_14276 = n_14133 ^ n_11729;
assign n_14277 = n_13386 & ~n_14134;
assign n_14278 = n_14137 ^ n_13967;
assign n_14279 = ~n_13574 & n_14138;
assign n_14280 = n_14139 ^ n_13968;
assign n_14281 = n_13575 & n_14140;
assign n_14282 = n_14141 ^ n_13969;
assign n_14283 = ~n_13576 & n_14142;
assign n_14284 = n_14143 ^ n_13970;
assign n_14285 = n_13577 & n_14144;
assign n_14286 = n_14145 ^ n_13971;
assign n_14287 = ~n_13619 & n_14146;
assign n_14288 = n_14147 ^ n_13972;
assign n_14289 = ~n_13621 & n_14148;
assign n_14290 = n_14149 ^ n_13973;
assign n_14291 = n_13623 & n_14150;
assign n_14292 = n_14151 ^ n_13534;
assign n_14293 = n_14151 & n_13625;
assign n_14294 = n_14152 ^ n_13536;
assign n_14295 = n_14152 & ~n_13627;
assign n_14296 = n_13976 ^ n_14153;
assign n_14297 = ~n_13578 & n_14154;
assign n_14298 = n_14156 ^ x107;
assign n_14299 = n_14157 ^ n_2077;
assign n_14300 = n_14158 ^ n_13921;
assign n_14301 = n_13998 ^ n_14167;
assign n_14302 = n_14168 ^ n_13690;
assign n_14303 = n_14169 ^ n_13692;
assign n_14304 = n_14170 ^ n_13694;
assign n_14305 = n_14171 ^ n_13696;
assign n_14306 = n_14172 ^ n_13698;
assign n_14307 = n_14173 ^ n_13782;
assign n_14308 = n_14174 ^ n_13784;
assign n_14309 = n_14175 ^ n_13786;
assign n_14310 = n_14176 ^ n_13788;
assign n_14311 = n_14177 ^ n_13753;
assign n_14312 = n_14178 ^ n_6358;
assign n_14313 = ~x0 & n_14179;
assign n_14314 = n_14180 ^ x5;
assign n_14315 = n_14181 ^ x8;
assign n_14316 = n_14182 ^ x11;
assign n_14317 = n_14183 ^ x14;
assign n_14318 = n_14184 ^ x17;
assign n_14319 = n_14185 ^ x20;
assign n_14320 = n_14186 ^ x23;
assign n_14321 = n_14187 ^ x26;
assign n_14322 = n_14188 ^ x29;
assign n_14323 = n_14189 ^ x32;
assign n_14324 = n_14190 ^ x35;
assign n_14325 = n_14191 ^ x38;
assign n_14326 = n_14192 ^ x41;
assign n_14327 = n_14193 ^ x44;
assign n_14328 = n_14194 ^ x47;
assign n_14329 = n_14195 ^ x50;
assign n_14330 = n_14196 ^ x53;
assign n_14331 = n_14197 ^ x56;
assign n_14332 = n_14198 ^ x59;
assign n_14333 = n_14199 ^ x62;
assign n_14334 = n_14200 ^ n_3517;
assign n_14335 = n_5042 ^ n_14201;
assign n_14336 = n_5105 ^ n_14202;
assign n_14337 = n_5168 ^ n_14203;
assign n_14338 = n_5229 ^ n_14204;
assign n_14339 = n_5293 ^ n_14205;
assign n_14340 = n_5357 ^ n_14206;
assign n_14341 = n_5421 ^ n_14207;
assign n_14342 = n_5485 ^ n_14208;
assign n_14343 = n_5546 ^ n_14209;
assign n_14344 = n_5609 ^ n_14210;
assign n_14345 = n_5672 ^ n_14211;
assign n_14346 = n_5736 ^ n_14212;
assign n_14347 = n_5802 ^ n_14213;
assign n_14348 = n_5864 ^ n_14214;
assign n_14349 = n_5928 ^ n_14215;
assign n_14350 = n_5991 ^ n_14216;
assign n_14351 = n_6055 ^ n_14217;
assign n_14352 = n_6119 ^ n_14218;
assign n_14353 = n_6181 ^ n_14219;
assign n_14354 = n_6243 ^ n_14220;
assign n_14355 = n_14221 ^ x115;
assign n_14356 = n_2170 ^ n_14222;
assign n_14357 = n_770 ^ n_14223;
assign n_14358 = n_2241 ^ n_14224;
assign n_14359 = n_2309 ^ n_14225;
assign n_14360 = n_2376 ^ n_14226;
assign n_14361 = n_2443 ^ n_14227;
assign n_14362 = n_2510 ^ n_14228;
assign n_14363 = n_2576 ^ n_14229;
assign n_14364 = n_2641 ^ n_14230;
assign n_14365 = n_2708 ^ n_14231;
assign n_14366 = n_2776 ^ n_14232;
assign n_14367 = n_2843 ^ n_14233;
assign n_14368 = n_2911 ^ n_14234;
assign n_14369 = n_2977 ^ n_14235;
assign n_14370 = n_3046 ^ n_14236;
assign n_14371 = n_3112 ^ n_14237;
assign n_14372 = n_3181 ^ n_14238;
assign n_14373 = n_3245 ^ n_14239;
assign n_14374 = n_3310 ^ n_14240;
assign n_14375 = n_3375 ^ n_14241;
assign n_14376 = n_14242 ^ x1;
assign n_14377 = n_655 & ~n_14243;
assign n_14378 = n_784 & ~n_14243;
assign n_14379 = ~n_3665 & ~n_14243;
assign n_14380 = n_854 & ~n_14243;
assign n_14381 = n_920 & ~n_14243;
assign n_14382 = n_986 & ~n_14243;
assign n_14383 = n_1052 & ~n_14243;
assign n_14384 = n_1117 & ~n_14243;
assign n_14385 = n_1181 & ~n_14243;
assign n_14386 = n_1248 & ~n_14243;
assign n_14387 = n_1314 & ~n_14243;
assign n_14388 = n_1380 & ~n_14243;
assign n_14389 = n_1445 & ~n_14243;
assign n_14390 = n_1510 & ~n_14243;
assign n_14391 = n_1576 & ~n_14243;
assign n_14392 = n_1641 & ~n_14243;
assign n_14393 = n_1706 & ~n_14243;
assign n_14394 = ~n_14243 & n_1771;
assign n_14395 = ~n_14243 & n_1835;
assign n_14396 = ~n_14243 & n_1899;
assign n_14397 = n_1 & n_14244;
assign n_14398 = n_14244 ^ x117;
assign n_14399 = n_14022 ^ n_14245;
assign n_14400 = n_14246 ^ n_13396;
assign n_14401 = n_14246 ^ n_13268;
assign n_14402 = n_14247 ^ n_10159;
assign n_14403 = ~n_13373 & n_14248;
assign n_14404 = n_14249 ^ n_10160;
assign n_14405 = n_13375 & ~n_14250;
assign n_14406 = n_14251 ^ n_10161;
assign n_14407 = ~n_13030 & n_14252;
assign n_14408 = n_14253 ^ n_10164;
assign n_14409 = ~n_13379 & n_14254;
assign n_14410 = n_14255 ^ n_10165;
assign n_14411 = n_13381 & ~n_14256;
assign n_14412 = n_14257 ^ n_10166;
assign n_14413 = n_13257 & ~n_14258;
assign n_14414 = n_14260 ^ n_13993;
assign n_14415 = n_14261 ^ n_10686;
assign n_14416 = n_13274 & ~n_14262;
assign n_14417 = n_14263 ^ n_12966;
assign n_14418 = ~n_13151 & n_14264;
assign n_14419 = n_14265 ^ n_13838;
assign n_14420 = n_14266 ^ n_13491;
assign n_14421 = n_14266 ^ n_13369;
assign n_14422 = n_14267 ^ n_13394;
assign n_14423 = n_14267 ^ n_13266;
assign n_14424 = n_14268 ^ n_10372;
assign n_14425 = ~n_13505 & n_14269;
assign n_14426 = n_14270 ^ n_10289;
assign n_14427 = ~n_13658 & n_14271;
assign n_14428 = n_14272 ^ n_10293;
assign n_14429 = ~n_13400 & n_14273;
assign n_14430 = n_14274 ^ n_10294;
assign n_14431 = ~n_13664 & n_14275;
assign n_14432 = n_14277 ^ n_14012;
assign n_14433 = n_14279 ^ n_14033;
assign n_14434 = n_14281 ^ n_14034;
assign n_14435 = n_14283 ^ n_14035;
assign n_14436 = n_14285 ^ n_14036;
assign n_14437 = n_14287 ^ n_14037;
assign n_14438 = n_14289 ^ n_14038;
assign n_14439 = n_14291 ^ n_14039;
assign n_14440 = n_13974 ^ n_14292;
assign n_14441 = n_14293 ^ n_14040;
assign n_14442 = n_14294 ^ n_13975;
assign n_14443 = n_14295 ^ n_14041;
assign n_14444 = n_14297 ^ n_14042;
assign n_14445 = n_594 ^ n_14298;
assign n_14446 = ~n_3512 & ~n_14299;
assign n_14447 = n_14313 ^ n_14067;
assign n_14448 = n_13838 ^ n_14322;
assign n_14449 = n_14323 ^ n_14013;
assign n_14450 = n_14323 ^ n_13840;
assign n_14451 = n_14324 ^ n_14014;
assign n_14452 = n_14324 ^ n_13735;
assign n_14453 = n_14325 ^ n_14015;
assign n_14454 = n_14325 ^ n_13892;
assign n_14455 = n_14326 ^ n_14016;
assign n_14456 = n_14326 ^ n_13893;
assign n_14457 = n_14327 ^ n_14017;
assign n_14458 = n_14327 ^ n_13741;
assign n_14459 = n_14328 ^ n_14018;
assign n_14460 = n_14328 ^ n_13848;
assign n_14461 = n_14329 ^ n_13896;
assign n_14462 = n_14330 ^ n_13897;
assign n_14463 = n_14331 ^ n_13898;
assign n_14464 = n_14332 ^ n_13857;
assign n_14465 = n_14333 ^ n_6492;
assign n_14466 = ~x0 & n_14334;
assign n_14467 = n_14335 ^ x5;
assign n_14468 = n_14336 ^ x8;
assign n_14469 = n_14337 ^ x11;
assign n_14470 = n_14338 ^ x14;
assign n_14471 = n_14339 ^ x17;
assign n_14472 = n_14340 ^ x20;
assign n_14473 = n_14341 ^ x23;
assign n_14474 = n_14342 ^ x26;
assign n_14475 = n_14343 ^ x29;
assign n_14476 = n_14344 ^ x32;
assign n_14477 = n_14345 ^ x35;
assign n_14478 = n_14346 ^ x38;
assign n_14479 = n_14347 ^ x41;
assign n_14480 = n_14348 ^ x44;
assign n_14481 = n_14349 ^ x47;
assign n_14482 = n_14350 ^ x50;
assign n_14483 = n_14351 ^ x53;
assign n_14484 = n_14352 ^ x56;
assign n_14485 = n_14353 ^ x59;
assign n_14486 = n_14354 ^ x62;
assign n_14487 = n_14355 ^ n_3519;
assign n_14488 = n_5043 ^ n_14356;
assign n_14489 = n_5106 ^ n_14357;
assign n_14490 = n_5169 ^ n_14358;
assign n_14491 = n_5230 ^ n_14359;
assign n_14492 = n_5294 ^ n_14360;
assign n_14493 = n_5358 ^ n_14361;
assign n_14494 = n_5422 ^ n_14362;
assign n_14495 = n_5486 ^ n_14363;
assign n_14496 = n_5547 ^ n_14364;
assign n_14497 = n_5610 ^ n_14365;
assign n_14498 = n_5673 ^ n_14366;
assign n_14499 = n_5737 ^ n_14367;
assign n_14500 = n_5803 ^ n_14368;
assign n_14501 = n_5865 ^ n_14369;
assign n_14502 = n_5929 ^ n_14370;
assign n_14503 = n_5992 ^ n_14371;
assign n_14504 = n_6056 ^ n_14372;
assign n_14505 = n_6120 ^ n_14373;
assign n_14506 = n_6182 ^ n_14374;
assign n_14507 = n_6244 ^ n_14375;
assign n_14508 = n_14376 ^ x116;
assign n_14509 = n_2171 ^ n_14377;
assign n_14510 = n_771 ^ n_14378;
assign n_14511 = n_2242 ^ n_14379;
assign n_14512 = n_2310 ^ n_14380;
assign n_14513 = n_2377 ^ n_14381;
assign n_14514 = n_2444 ^ n_14382;
assign n_14515 = n_2511 ^ n_14383;
assign n_14516 = n_2577 ^ n_14384;
assign n_14517 = n_2642 ^ n_14385;
assign n_14518 = n_2709 ^ n_14386;
assign n_14519 = n_2777 ^ n_14387;
assign n_14520 = n_2844 ^ n_14388;
assign n_14521 = n_2912 ^ n_14389;
assign n_14522 = n_2978 ^ n_14390;
assign n_14523 = n_3047 ^ n_14391;
assign n_14524 = n_3113 ^ n_14392;
assign n_14525 = n_3182 ^ n_14393;
assign n_14526 = n_3246 ^ n_14394;
assign n_14527 = n_3311 ^ n_14395;
assign n_14528 = n_3376 ^ n_14396;
assign n_14529 = n_14397 ^ x1;
assign n_14530 = n_655 & ~n_14398;
assign n_14531 = n_784 & ~n_14398;
assign n_14532 = ~n_3665 & ~n_14398;
assign n_14533 = n_854 & ~n_14398;
assign n_14534 = n_920 & ~n_14398;
assign n_14535 = n_986 & ~n_14398;
assign n_14536 = n_1052 & ~n_14398;
assign n_14537 = n_1117 & ~n_14398;
assign n_14538 = n_1181 & ~n_14398;
assign n_14539 = n_1248 & ~n_14398;
assign n_14540 = n_1314 & ~n_14398;
assign n_14541 = n_1380 & ~n_14398;
assign n_14542 = n_1445 & ~n_14398;
assign n_14543 = n_1510 & ~n_14398;
assign n_14544 = n_1576 & ~n_14398;
assign n_14545 = n_1641 & ~n_14398;
assign n_14546 = n_1706 & ~n_14398;
assign n_14547 = ~n_14398 & n_1771;
assign n_14548 = ~n_14398 & n_1835;
assign n_14549 = ~n_14398 & n_1899;
assign n_14550 = n_1 & n_14399;
assign n_14551 = n_14399 & n_272;
assign n_14552 = ~x119 & n_14399;
assign n_14553 = n_14399 ^ x117;
assign n_14554 = n_14400 ^ n_10288;
assign n_14555 = ~n_13396 & n_14401;
assign n_14556 = n_14403 ^ n_14115;
assign n_14557 = n_14405 ^ n_14116;
assign n_14558 = n_14407 ^ n_14117;
assign n_14559 = n_14409 ^ n_14118;
assign n_14560 = n_14411 ^ n_14119;
assign n_14561 = n_14413 ^ n_14120;
assign n_14562 = n_14414 ^ n_13671;
assign n_14563 = n_14414 ^ n_13595;
assign n_14564 = n_14416 ^ n_14123;
assign n_14565 = n_14418 ^ n_14124;
assign n_14566 = n_14419 ^ n_14322;
assign n_14567 = n_14420 ^ n_10287;
assign n_14568 = ~n_13491 & n_14421;
assign y25 = n_14422;
assign n_14569 = ~n_13394 & n_14423;
assign n_14570 = n_14425 ^ n_14129;
assign n_14571 = n_14427 ^ n_14130;
assign n_14572 = n_14429 ^ n_14131;
assign n_14573 = n_14431 ^ n_14132;
assign n_14574 = n_14432 ^ n_13673;
assign n_14575 = n_14432 ^ n_13597;
assign n_14576 = n_14433 ^ n_14302;
assign n_14577 = n_14433 ^ n_14168;
assign n_14578 = n_14434 ^ n_14303;
assign n_14579 = n_14434 ^ n_13692;
assign n_14580 = n_14435 ^ n_14304;
assign n_14581 = n_14435 ^ n_13694;
assign n_14582 = n_14436 ^ n_14305;
assign n_14583 = n_14436 ^ n_13696;
assign n_14584 = n_14437 ^ n_14306;
assign n_14585 = n_14437 ^ n_13698;
assign n_14586 = n_14438 ^ n_14307;
assign n_14587 = n_14438 ^ n_14173;
assign n_14588 = n_14439 ^ n_14174;
assign n_14589 = n_14441 ^ n_14309;
assign n_14590 = n_14441 ^ n_14175;
assign n_14591 = n_14443 ^ n_14176;
assign n_14592 = n_14444 ^ n_14311;
assign n_14593 = n_14444 ^ n_14177;
assign n_14594 = x62 & ~n_14445;
assign n_14595 = n_14446 ^ n_14157;
assign n_14596 = ~n_14419 & n_14448;
assign n_14597 = ~n_14013 & n_14450;
assign n_14598 = ~n_14014 & n_14452;
assign n_14599 = n_14015 & n_14454;
assign n_14600 = ~n_14016 & ~n_14456;
assign n_14601 = n_14017 & n_14458;
assign n_14602 = ~n_14018 & n_14460;
assign n_14603 = n_14461 ^ n_13850;
assign n_14604 = n_14461 & n_14019;
assign n_14605 = n_14462 ^ n_13852;
assign n_14606 = n_14462 & n_14020;
assign n_14607 = n_14463 ^ n_13854;
assign n_14608 = n_14463 & n_14021;
assign n_14609 = n_14464 ^ n_13751;
assign n_14610 = ~n_14464 & n_13978;
assign n_14611 = n_14465 ^ n_3414;
assign n_14612 = ~n_14465 & ~n_6608;
assign n_14613 = n_14466 ^ n_14200;
assign n_14614 = n_14475 ^ n_14278;
assign n_14615 = n_14475 ^ n_14137;
assign n_14616 = n_14476 ^ n_14280;
assign n_14617 = n_14476 ^ n_14139;
assign n_14618 = n_14477 ^ n_14282;
assign n_14619 = n_14477 ^ n_14141;
assign n_14620 = n_14478 ^ n_14284;
assign n_14621 = n_14478 ^ n_13970;
assign n_14622 = n_14479 ^ n_14286;
assign n_14623 = n_14479 ^ n_14145;
assign n_14624 = n_14480 ^ n_14288;
assign n_14625 = n_14480 ^ n_14147;
assign n_14626 = n_14481 ^ n_14290;
assign n_14627 = n_14481 ^ n_13973;
assign n_14628 = n_14482 ^ n_13974;
assign n_14629 = n_14483 ^ n_14442;
assign n_14630 = n_14483 ^ n_13975;
assign n_14631 = n_14484 ^ n_13976;
assign n_14632 = n_14485 ^ n_14155;
assign n_14633 = n_14485 ^ n_13977;
assign n_14634 = ~x0 & n_14487;
assign n_14635 = n_14488 ^ x5;
assign n_14636 = n_14489 ^ x8;
assign n_14637 = n_14490 ^ x11;
assign n_14638 = n_14491 ^ x14;
assign n_14639 = n_14492 ^ x17;
assign n_14640 = n_14493 ^ x20;
assign n_14641 = n_14494 ^ x23;
assign n_14642 = n_14495 ^ x26;
assign n_14643 = n_14496 ^ x29;
assign n_14644 = n_14497 ^ x32;
assign n_14645 = n_14498 ^ x35;
assign n_14646 = n_14499 ^ x38;
assign n_14647 = n_14500 ^ x41;
assign n_14648 = n_14501 ^ x44;
assign n_14649 = n_14502 ^ x47;
assign n_14650 = n_14503 ^ x50;
assign n_14651 = n_14504 ^ x53;
assign n_14652 = n_14505 ^ x56;
assign n_14653 = n_14506 ^ x59;
assign n_14654 = n_14507 ^ x62;
assign n_14655 = n_14508 ^ n_6493;
assign n_14656 = n_5044 ^ n_14509;
assign n_14657 = n_5107 ^ n_14510;
assign n_14658 = n_5170 ^ n_14511;
assign n_14659 = n_5231 ^ n_14512;
assign n_14660 = n_5295 ^ n_14513;
assign n_14661 = n_5359 ^ n_14514;
assign n_14662 = n_5423 ^ n_14515;
assign n_14663 = n_5487 ^ n_14516;
assign n_14664 = n_5548 ^ n_14517;
assign n_14665 = n_5611 ^ n_14518;
assign n_14666 = n_5674 ^ n_14519;
assign n_14667 = n_5738 ^ n_14520;
assign n_14668 = n_5804 ^ n_14521;
assign n_14669 = n_5866 ^ n_14522;
assign n_14670 = n_5930 ^ n_14523;
assign n_14671 = n_5993 ^ n_14524;
assign n_14672 = n_6057 ^ n_14525;
assign n_14673 = n_6121 ^ n_14526;
assign n_14674 = n_6183 ^ n_14527;
assign n_14675 = n_6245 ^ n_14528;
assign n_14676 = n_14529 ^ x117;
assign n_14677 = n_2172 ^ n_14530;
assign n_14678 = n_772 ^ n_14531;
assign n_14679 = n_2243 ^ n_14532;
assign n_14680 = n_2311 ^ n_14533;
assign n_14681 = n_2378 ^ n_14534;
assign n_14682 = n_2445 ^ n_14535;
assign n_14683 = n_2512 ^ n_14536;
assign n_14684 = n_2578 ^ n_14537;
assign n_14685 = n_2643 ^ n_14538;
assign n_14686 = n_2710 ^ n_14539;
assign n_14687 = n_2778 ^ n_14540;
assign n_14688 = n_2845 ^ n_14541;
assign n_14689 = n_2913 ^ n_14542;
assign n_14690 = n_2979 ^ n_14543;
assign n_14691 = n_3048 ^ n_14544;
assign n_14692 = n_3114 ^ n_14545;
assign n_14693 = n_3183 ^ n_14546;
assign n_14694 = n_3247 ^ n_14547;
assign n_14695 = n_3312 ^ n_14548;
assign n_14696 = n_3377 ^ n_14549;
assign n_14697 = n_14550 ^ x1;
assign n_14698 = n_1 & ~n_14551;
assign n_14699 = n_14551 ^ x119;
assign n_14700 = n_14552 ^ n_14245;
assign n_14701 = n_14553 ^ n_272;
assign n_14702 = n_14553 & n_611;
assign n_14703 = n_14555 ^ n_14246;
assign n_14704 = n_14556 ^ n_13660;
assign n_14705 = n_14556 ^ n_13583;
assign n_14706 = n_14557 ^ n_13662;
assign n_14707 = n_14557 ^ n_13585;
assign n_14708 = n_14558 ^ n_13398;
assign n_14709 = n_14558 ^ n_13270;
assign n_14710 = n_14559 ^ n_13666;
assign n_14711 = n_14559 ^ n_13589;
assign n_14712 = n_14560 ^ n_13668;
assign n_14713 = n_14560 ^ n_13591;
assign n_14714 = n_14561 ^ n_13593;
assign n_14715 = n_14561 ^ n_13499;
assign n_14716 = n_14562 ^ n_10298;
assign n_14717 = ~n_13671 & n_14563;
assign n_14718 = n_14564 ^ n_13610;
assign n_14719 = n_14564 ^ n_13512;
assign n_14720 = n_14565 ^ n_13503;
assign n_14721 = n_14565 ^ n_13388;
assign n_14722 = n_14568 ^ n_14266;
assign n_14723 = n_14569 ^ n_14267;
assign n_14724 = n_14570 ^ n_13768;
assign n_14725 = n_14570 ^ n_13677;
assign n_14726 = n_14571 ^ n_13981;
assign n_14727 = n_14571 ^ n_13859;
assign n_14728 = n_14572 ^ n_13687;
assign n_14729 = n_14572 ^ n_13608;
assign n_14730 = n_14573 ^ n_13987;
assign n_14731 = n_14573 ^ n_13865;
assign n_14732 = n_14574 ^ n_12666;
assign n_14733 = n_13673 & ~n_14575;
assign n_14734 = ~n_14302 & n_14577;
assign n_14735 = ~n_14303 & n_14579;
assign n_14736 = ~n_14304 & n_14581;
assign n_14737 = ~n_14305 & n_14583;
assign n_14738 = ~n_14306 & n_14585;
assign n_14739 = ~n_14307 & n_14587;
assign n_14740 = n_14588 ^ n_13784;
assign n_14741 = n_14588 & ~n_14308;
assign n_14742 = n_14309 & n_14590;
assign n_14743 = n_14591 ^ n_13788;
assign n_14744 = n_14591 & ~n_14310;
assign n_14745 = ~n_14311 & n_14593;
assign n_14746 = n_14594 ^ n_594;
assign n_14747 = n_14595 ^ n_2077;
assign n_14748 = n_14596 ^ n_14265;
assign n_14749 = n_14597 ^ n_14323;
assign n_14750 = n_14598 ^ n_14324;
assign n_14751 = n_14599 ^ n_14325;
assign n_14752 = n_14600 ^ n_14326;
assign n_14753 = n_14601 ^ n_13894;
assign n_14754 = n_14602 ^ n_14328;
assign n_14755 = n_14604 ^ n_14329;
assign n_14756 = n_14606 ^ n_14330;
assign n_14757 = n_14608 ^ n_14331;
assign n_14758 = n_14610 ^ n_14332;
assign n_14759 = n_14612 ^ n_14333;
assign n_14760 = n_14278 & ~n_14615;
assign n_14761 = n_14280 & ~n_14617;
assign n_14762 = ~n_14282 & n_14619;
assign n_14763 = n_14284 & n_14621;
assign n_14764 = ~n_14286 & n_14623;
assign n_14765 = n_14288 & ~n_14625;
assign n_14766 = n_14290 & n_14627;
assign n_14767 = n_14628 ^ n_14292;
assign n_14768 = n_14628 & n_14440;
assign n_14769 = ~n_14442 & n_14630;
assign n_14770 = n_14631 ^ n_14153;
assign n_14771 = ~n_14631 & n_14296;
assign n_14772 = n_14155 & n_14633;
assign n_14773 = n_14634 ^ n_14355;
assign n_14774 = n_14643 ^ n_14576;
assign n_14775 = n_14644 ^ n_14578;
assign n_14776 = n_14645 ^ n_14580;
assign n_14777 = n_14646 ^ n_14582;
assign n_14778 = n_14647 ^ n_14584;
assign n_14779 = n_14648 ^ n_14586;
assign n_14780 = n_14589 ^ n_14650;
assign n_14781 = n_14652 ^ n_14592;
assign n_14782 = n_14654 ^ n_6416;
assign n_14783 = ~x0 & ~n_14655;
assign n_14784 = n_14656 ^ x5;
assign n_14785 = n_14657 ^ x8;
assign n_14786 = n_14658 ^ x11;
assign n_14787 = n_14659 ^ x14;
assign n_14788 = n_14660 ^ x17;
assign n_14789 = n_14661 ^ x20;
assign n_14790 = n_14662 ^ x23;
assign n_14791 = n_14663 ^ x26;
assign n_14792 = n_14664 ^ x29;
assign n_14793 = n_14665 ^ x32;
assign n_14794 = n_14666 ^ x35;
assign n_14795 = n_14667 ^ x38;
assign n_14796 = n_14668 ^ x41;
assign n_14797 = n_14669 ^ x44;
assign n_14798 = n_14670 ^ x47;
assign n_14799 = n_14671 ^ x50;
assign n_14800 = n_14672 ^ x53;
assign n_14801 = n_14673 ^ x56;
assign n_14802 = n_14674 ^ x59;
assign n_14803 = n_14675 ^ x62;
assign n_14804 = n_14676 ^ n_6495;
assign n_14805 = n_5045 ^ n_14677;
assign n_14806 = n_5108 ^ n_14678;
assign n_14807 = n_5171 ^ n_14679;
assign n_14808 = n_5232 ^ n_14680;
assign n_14809 = n_5296 ^ n_14681;
assign n_14810 = n_5360 ^ n_14682;
assign n_14811 = n_5424 ^ n_14683;
assign n_14812 = n_5488 ^ n_14684;
assign n_14813 = n_5549 ^ n_14685;
assign n_14814 = n_5612 ^ n_14686;
assign n_14815 = n_5675 ^ n_14687;
assign n_14816 = n_5739 ^ n_14688;
assign n_14817 = n_5805 ^ n_14689;
assign n_14818 = n_5867 ^ n_14690;
assign n_14819 = n_5931 ^ n_14691;
assign n_14820 = n_5994 ^ n_14692;
assign n_14821 = n_6058 ^ n_14693;
assign n_14822 = n_6122 ^ n_14694;
assign n_14823 = n_6184 ^ n_14695;
assign n_14824 = n_6246 ^ n_14696;
assign n_14825 = n_14697 ^ x118;
assign n_14826 = n_14698 ^ x1;
assign n_14827 = n_655 & n_14699;
assign n_14828 = n_784 & n_14699;
assign n_14829 = ~n_3665 & n_14699;
assign n_14830 = n_854 & n_14699;
assign n_14831 = n_920 & n_14699;
assign n_14832 = n_986 & n_14699;
assign n_14833 = n_1052 & n_14699;
assign n_14834 = n_1117 & n_14699;
assign n_14835 = n_1181 & n_14699;
assign n_14836 = n_1248 & n_14699;
assign n_14837 = n_1314 & n_14699;
assign n_14838 = n_1380 & n_14699;
assign n_14839 = n_1445 & n_14699;
assign n_14840 = n_1510 & n_14699;
assign n_14841 = n_1576 & n_14699;
assign n_14842 = n_1641 & n_14699;
assign n_14843 = n_1706 & n_14699;
assign n_14844 = n_1771 & n_14699;
assign n_14845 = n_14699 & n_1835;
assign n_14846 = n_14699 & n_1899;
assign n_14847 = n_276 & ~n_14700;
assign n_14848 = n_655 & ~n_14701;
assign n_14849 = n_784 & ~n_14701;
assign n_14850 = ~n_3665 & ~n_14701;
assign n_14851 = n_854 & ~n_14701;
assign n_14852 = n_920 & ~n_14701;
assign n_14853 = n_986 & ~n_14701;
assign n_14854 = n_1052 & ~n_14701;
assign n_14855 = n_1117 & ~n_14701;
assign n_14856 = n_1181 & ~n_14701;
assign n_14857 = n_1248 & ~n_14701;
assign n_14858 = n_1314 & ~n_14701;
assign n_14859 = n_1380 & ~n_14701;
assign n_14860 = n_1445 & ~n_14701;
assign n_14861 = n_1510 & ~n_14701;
assign n_14862 = n_1576 & ~n_14701;
assign n_14863 = n_1641 & ~n_14701;
assign n_14864 = n_1706 & ~n_14701;
assign n_14865 = n_1771 & ~n_14701;
assign n_14866 = ~n_14701 & n_1835;
assign n_14867 = ~n_14701 & n_1899;
assign n_14868 = n_3526 & ~n_14702;
assign n_14869 = n_14703 ^ n_13683;
assign n_14870 = n_14703 ^ n_13604;
assign n_14871 = n_14704 ^ n_10290;
assign n_14872 = ~n_13660 & n_14705;
assign n_14873 = n_14706 ^ n_10291;
assign n_14874 = ~n_13662 & n_14707;
assign n_14875 = n_14708 ^ n_10292;
assign n_14876 = ~n_13398 & n_14709;
assign n_14877 = n_14710 ^ n_10295;
assign n_14878 = ~n_13666 & n_14711;
assign n_14879 = n_14712 ^ n_10296;
assign n_14880 = ~n_13668 & n_14713;
assign n_14881 = n_14714 ^ n_10297;
assign n_14882 = ~n_13593 & n_14715;
assign n_14883 = n_14717 ^ n_14414;
assign n_14884 = n_14718 ^ n_11448;
assign n_14885 = n_13610 & ~n_14719;
assign n_14886 = n_14720 ^ n_13643;
assign n_14887 = ~n_13503 & n_14721;
assign n_14888 = n_14722 ^ n_13755;
assign n_14889 = n_14722 ^ n_13656;
assign n_14890 = n_14723 ^ n_13681;
assign n_14891 = n_14723 ^ n_13602;
assign n_14892 = n_14724 ^ n_10494;
assign n_14893 = n_13768 & ~n_14725;
assign n_14894 = n_14726 ^ n_10376;
assign n_14895 = ~n_13981 & n_14727;
assign n_14896 = n_14728 ^ n_10380;
assign n_14897 = ~n_13687 & n_14729;
assign n_14898 = n_14730 ^ n_10381;
assign n_14899 = ~n_13987 & n_14731;
assign n_14900 = n_14733 ^ n_14432;
assign n_14901 = n_14734 ^ n_14433;
assign n_14902 = n_14735 ^ n_14169;
assign n_14903 = n_14736 ^ n_14170;
assign n_14904 = n_14737 ^ n_14171;
assign n_14905 = n_14738 ^ n_14172;
assign n_14906 = n_14739 ^ n_14438;
assign n_14907 = n_14740 ^ n_14649;
assign n_14908 = n_14741 ^ n_14439;
assign n_14909 = n_14742 ^ n_14441;
assign n_14910 = n_14651 ^ n_14743;
assign n_14911 = n_14744 ^ n_14443;
assign n_14912 = n_14745 ^ n_14444;
assign n_14913 = x63 & n_14746;
assign n_14914 = n_14747 ^ n_13920;
assign n_14915 = n_14748 ^ n_14614;
assign n_14916 = n_14749 ^ n_14616;
assign n_14917 = n_14750 ^ n_14618;
assign n_14918 = n_14751 ^ n_14620;
assign n_14919 = n_14752 ^ n_14622;
assign n_14920 = n_14753 ^ n_14624;
assign n_14921 = n_14754 ^ n_14626;
assign n_14922 = n_14629 ^ n_14756;
assign n_14923 = n_14632 ^ n_14758;
assign n_14924 = n_14759 ^ n_6755;
assign n_14925 = ~n_6285 & ~n_14759;
assign n_14926 = n_14760 ^ n_13967;
assign n_14927 = n_14761 ^ n_14476;
assign n_14928 = n_14762 ^ n_14477;
assign n_14929 = n_14763 ^ n_14478;
assign n_14930 = n_14764 ^ n_14479;
assign n_14931 = n_14765 ^ n_13972;
assign n_14932 = n_14766 ^ n_14481;
assign n_14933 = n_14767 ^ n_14755;
assign n_14934 = n_14768 ^ n_14482;
assign n_14935 = n_14769 ^ n_14483;
assign n_14936 = n_14757 ^ n_14770;
assign n_14937 = n_14771 ^ n_14484;
assign n_14938 = n_14772 ^ n_14485;
assign n_14939 = n_14783 ^ n_14508;
assign n_14940 = n_14566 ^ n_14791;
assign n_14941 = n_14798 ^ n_14603;
assign n_14942 = n_14800 ^ n_14607;
assign n_14943 = n_14802 ^ n_14611;
assign n_14944 = n_14803 ^ n_6646;
assign n_14945 = n_14803 ^ n_6536;
assign n_14946 = ~x0 & ~n_14804;
assign n_14947 = n_14805 ^ x5;
assign n_14948 = n_14806 ^ x8;
assign n_14949 = n_14807 ^ x11;
assign n_14950 = n_14808 ^ x14;
assign n_14951 = n_14809 ^ x17;
assign n_14952 = n_14810 ^ x20;
assign n_14953 = n_14811 ^ x23;
assign n_14954 = n_14812 ^ x26;
assign n_14955 = n_14813 ^ x29;
assign n_14956 = n_14814 ^ x32;
assign n_14957 = n_14815 ^ x35;
assign n_14958 = n_14816 ^ x38;
assign n_14959 = n_14817 ^ x41;
assign n_14960 = n_14818 ^ x44;
assign n_14961 = n_14819 ^ x47;
assign n_14962 = n_14820 ^ x50;
assign n_14963 = n_14821 ^ x53;
assign n_14964 = n_14822 ^ x56;
assign n_14965 = n_14823 ^ x59;
assign n_14966 = n_4982 ^ n_14824;
assign n_14967 = n_14824 ^ x114;
assign n_14968 = ~n_14824 & n_3521;
assign n_14969 = n_14824 ^ x113;
assign n_14970 = n_14825 ^ n_2113;
assign n_14971 = n_14826 ^ x119;
assign n_14972 = n_2174 ^ n_14827;
assign n_14973 = n_774 ^ n_14828;
assign n_14974 = n_2245 ^ n_14829;
assign n_14975 = n_2313 ^ n_14830;
assign n_14976 = n_2380 ^ n_14831;
assign n_14977 = n_2447 ^ n_14832;
assign n_14978 = n_2514 ^ n_14833;
assign n_14979 = n_2580 ^ n_14834;
assign n_14980 = n_2645 ^ n_14835;
assign n_14981 = n_2712 ^ n_14836;
assign n_14982 = n_2780 ^ n_14837;
assign n_14983 = n_2847 ^ n_14838;
assign n_14984 = n_2915 ^ n_14839;
assign n_14985 = n_2981 ^ n_14840;
assign n_14986 = n_3050 ^ n_14841;
assign n_14987 = n_3116 ^ n_14842;
assign n_14988 = n_3185 ^ n_14843;
assign n_14989 = n_3249 ^ n_14844;
assign n_14990 = n_3314 ^ n_14845;
assign n_14991 = n_3379 ^ n_14846;
assign n_14992 = n_1 & ~n_14847;
assign n_14993 = n_14847 ^ x120;
assign n_14994 = n_2173 ^ n_14848;
assign n_14995 = n_773 ^ n_14849;
assign n_14996 = n_2244 ^ n_14850;
assign n_14997 = n_2312 ^ n_14851;
assign n_14998 = n_2379 ^ n_14852;
assign n_14999 = n_2446 ^ n_14853;
assign n_15000 = n_2513 ^ n_14854;
assign n_15001 = n_2579 ^ n_14855;
assign n_15002 = n_2644 ^ n_14856;
assign n_15003 = n_2711 ^ n_14857;
assign n_15004 = n_2779 ^ n_14858;
assign n_15005 = n_2846 ^ n_14859;
assign n_15006 = n_2914 ^ n_14860;
assign n_15007 = n_2980 ^ n_14861;
assign n_15008 = n_3049 ^ n_14862;
assign n_15009 = n_3115 ^ n_14863;
assign n_15010 = n_3184 ^ n_14864;
assign n_15011 = n_3248 ^ n_14865;
assign n_15012 = n_3313 ^ n_14866;
assign n_15013 = n_3378 ^ n_14867;
assign n_15014 = n_14868 ^ x120;
assign n_15015 = ~x120 & ~n_14868;
assign n_15016 = n_14869 ^ n_10375;
assign n_15017 = ~n_13683 & n_14870;
assign n_15018 = n_14872 ^ n_14556;
assign n_15019 = n_14874 ^ n_14557;
assign n_15020 = n_14876 ^ n_14558;
assign n_15021 = n_14878 ^ n_14559;
assign n_15022 = n_14880 ^ n_14560;
assign n_15023 = n_14882 ^ n_14561;
assign n_15024 = n_14883 ^ n_13994;
assign n_15025 = n_14883 ^ n_13873;
assign n_15026 = n_14885 ^ n_14564;
assign n_15027 = n_14887 ^ n_14565;
assign n_15028 = n_14888 ^ n_10374;
assign n_15029 = ~n_13755 & n_14889;
assign y26 = n_14890;
assign n_15030 = ~n_13681 & n_14891;
assign n_15031 = n_14893 ^ n_14570;
assign n_15032 = n_14895 ^ n_14571;
assign n_15033 = n_14897 ^ n_14572;
assign n_15034 = n_14899 ^ n_14573;
assign n_15035 = n_14900 ^ n_13996;
assign n_15036 = n_14900 ^ n_13875;
assign n_15037 = n_14901 ^ n_14449;
assign n_15038 = n_14901 ^ n_14792;
assign n_15039 = n_14902 ^ n_14451;
assign n_15040 = n_14902 ^ n_14793;
assign n_15041 = n_14903 ^ n_14453;
assign n_15042 = n_14903 ^ n_14794;
assign n_15043 = n_14904 ^ n_14455;
assign n_15044 = n_14904 ^ n_14795;
assign n_15045 = n_14905 ^ n_14457;
assign n_15046 = n_14905 ^ n_14796;
assign n_15047 = n_14906 ^ n_14459;
assign n_15048 = n_14906 ^ n_14797;
assign n_15049 = n_14798 ^ n_14908;
assign n_15050 = n_14909 ^ n_14799;
assign n_15051 = n_14909 ^ n_14605;
assign n_15052 = n_14911 ^ n_14800;
assign n_15053 = n_14912 ^ n_14801;
assign n_15054 = n_14912 ^ n_14609;
assign n_15055 = n_3511 & n_14914;
assign n_15056 = n_14486 ^ n_14924;
assign n_15057 = ~n_6415 & ~n_14925;
assign n_15058 = n_14926 ^ n_14774;
assign n_15059 = n_14926 ^ n_14643;
assign n_15060 = n_14927 ^ n_14775;
assign n_15061 = n_14927 ^ n_14644;
assign n_15062 = n_14928 ^ n_14776;
assign n_15063 = n_14928 ^ n_14645;
assign n_15064 = n_14929 ^ n_14777;
assign n_15065 = n_14929 ^ n_14646;
assign n_15066 = n_14930 ^ n_14778;
assign n_15067 = n_14930 ^ n_14584;
assign n_15068 = n_14931 ^ n_14779;
assign n_15069 = n_14931 ^ n_14648;
assign n_15070 = n_14932 ^ n_14907;
assign n_15071 = n_14932 ^ n_14649;
assign n_15072 = n_14934 ^ n_14589;
assign n_15073 = n_14935 ^ n_14651;
assign n_15074 = n_14937 ^ n_14781;
assign n_15075 = n_14937 ^ n_14652;
assign n_15076 = n_14938 ^ n_14653;
assign n_15077 = n_14941 ^ n_14908;
assign n_15078 = n_6646 & n_14945;
assign n_15079 = n_14946 ^ n_14676;
assign n_15080 = n_14915 ^ n_14954;
assign n_15081 = n_14614 ^ n_14954;
assign n_15082 = n_14955 ^ n_14916;
assign n_15083 = n_14955 ^ n_14616;
assign n_15084 = n_14956 ^ n_14917;
assign n_15085 = n_14956 ^ n_14618;
assign n_15086 = n_14957 ^ n_14918;
assign n_15087 = n_14957 ^ n_14620;
assign n_15088 = n_14958 ^ n_14919;
assign n_15089 = n_14958 ^ n_14622;
assign n_15090 = n_14959 ^ n_14920;
assign n_15091 = n_14959 ^ n_14624;
assign n_15092 = n_14960 ^ n_14921;
assign n_15093 = n_14960 ^ n_14626;
assign n_15094 = n_14961 ^ n_14933;
assign n_15095 = n_14961 ^ n_14767;
assign n_15096 = n_14962 ^ n_14629;
assign n_15097 = n_14963 ^ n_14757;
assign n_15098 = n_14964 ^ n_14632;
assign n_15099 = n_14965 ^ n_14486;
assign n_15100 = ~n_265 & ~n_14967;
assign n_15101 = ~n_263 & ~n_14969;
assign n_15102 = ~x0 & n_14970;
assign n_15103 = n_14971 ^ n_2114;
assign n_15104 = n_5047 ^ n_14972;
assign n_15105 = n_5110 ^ n_14973;
assign n_15106 = n_5173 ^ n_14974;
assign n_15107 = n_5234 ^ n_14975;
assign n_15108 = n_5298 ^ n_14976;
assign n_15109 = n_5362 ^ n_14977;
assign n_15110 = n_5426 ^ n_14978;
assign n_15111 = n_5490 ^ n_14979;
assign n_15112 = n_5551 ^ n_14980;
assign n_15113 = n_5614 ^ n_14981;
assign n_15114 = n_5677 ^ n_14982;
assign n_15115 = n_5741 ^ n_14983;
assign n_15116 = n_5807 ^ n_14984;
assign n_15117 = n_5869 ^ n_14985;
assign n_15118 = n_5933 ^ n_14986;
assign n_15119 = n_5996 ^ n_14987;
assign n_15120 = n_6060 ^ n_14988;
assign n_15121 = n_6124 ^ n_14989;
assign n_15122 = n_6186 ^ n_14990;
assign n_15123 = n_6248 ^ n_14991;
assign n_15124 = n_14992 ^ x1;
assign n_15125 = n_655 & n_14993;
assign n_15126 = n_784 & n_14993;
assign n_15127 = ~n_3665 & n_14993;
assign n_15128 = n_854 & n_14993;
assign n_15129 = n_920 & n_14993;
assign n_15130 = n_986 & n_14993;
assign n_15131 = n_1052 & n_14993;
assign n_15132 = n_1117 & n_14993;
assign n_15133 = n_1181 & n_14993;
assign n_15134 = n_1248 & n_14993;
assign n_15135 = n_1314 & n_14993;
assign n_15136 = n_1380 & n_14993;
assign n_15137 = n_1445 & n_14993;
assign n_15138 = n_1510 & n_14993;
assign n_15139 = n_1576 & n_14993;
assign n_15140 = n_1641 & n_14993;
assign n_15141 = n_1706 & n_14993;
assign n_15142 = n_1771 & n_14993;
assign n_15143 = n_14993 & n_1835;
assign n_15144 = n_14993 & n_1899;
assign n_15145 = n_5046 ^ n_14994;
assign n_15146 = n_5109 ^ n_14995;
assign n_15147 = n_5172 ^ n_14996;
assign n_15148 = n_5233 ^ n_14997;
assign n_15149 = n_5297 ^ n_14998;
assign n_15150 = n_5361 ^ n_14999;
assign n_15151 = n_5425 ^ n_15000;
assign n_15152 = n_5489 ^ n_15001;
assign n_15153 = n_5550 ^ n_15002;
assign n_15154 = n_5613 ^ n_15003;
assign n_15155 = n_5676 ^ n_15004;
assign n_15156 = n_5740 ^ n_15005;
assign n_15157 = n_5806 ^ n_15006;
assign n_15158 = n_5868 ^ n_15007;
assign n_15159 = n_5932 ^ n_15008;
assign n_15160 = n_5995 ^ n_15009;
assign n_15161 = n_6059 ^ n_15010;
assign n_15162 = n_6123 ^ n_15011;
assign n_15163 = n_6185 ^ n_15012;
assign n_15164 = n_6247 ^ n_15013;
assign n_15165 = n_1 & ~n_15014;
assign n_15166 = n_15014 ^ x121;
assign n_15167 = x121 & ~n_15015;
assign n_15168 = n_15015 ^ n_15014;
assign n_15169 = n_15017 ^ n_14703;
assign n_15170 = n_15018 ^ n_13983;
assign n_15171 = n_15018 ^ n_13861;
assign n_15172 = n_15019 ^ n_13985;
assign n_15173 = n_15019 ^ n_13863;
assign n_15174 = n_15020 ^ n_13685;
assign n_15175 = n_15020 ^ n_13606;
assign n_15176 = n_15021 ^ n_13989;
assign n_15177 = n_15021 ^ n_13867;
assign n_15178 = n_15022 ^ n_13991;
assign n_15179 = n_15022 ^ n_13869;
assign n_15180 = n_15023 ^ n_13871;
assign n_15181 = n_15023 ^ n_13763;
assign n_15182 = n_15024 ^ n_10385;
assign n_15183 = ~n_13994 & n_15025;
assign n_15184 = n_15026 ^ n_13888;
assign n_15185 = n_15026 ^ n_13775;
assign n_15186 = n_15027 ^ n_14136;
assign n_15187 = n_15027 ^ n_13675;
assign n_15188 = n_15029 ^ n_14722;
assign n_15189 = n_15030 ^ n_14723;
assign n_15190 = n_15031 ^ n_14126;
assign n_15191 = n_15031 ^ n_14000;
assign n_15192 = n_15032 ^ n_14402;
assign n_15193 = n_15032 ^ n_14247;
assign n_15194 = n_15033 ^ n_14010;
assign n_15195 = n_15033 ^ n_13886;
assign n_15196 = n_15034 ^ n_14408;
assign n_15197 = n_15034 ^ n_14253;
assign n_15198 = n_15035 ^ n_13300;
assign n_15199 = n_13996 & ~n_15036;
assign n_15200 = n_15037 ^ n_14792;
assign n_15201 = ~n_15037 & n_15038;
assign n_15202 = n_15039 ^ n_14793;
assign n_15203 = ~n_15039 & n_15040;
assign n_15204 = n_15041 ^ n_14794;
assign n_15205 = n_15041 & n_15042;
assign n_15206 = n_15043 ^ n_14795;
assign n_15207 = ~n_15043 & n_15044;
assign n_15208 = n_15045 ^ n_14796;
assign n_15209 = ~n_15045 & n_15046;
assign n_15210 = n_15047 ^ n_14797;
assign n_15211 = ~n_15047 & n_15048;
assign n_15212 = n_14941 & n_15049;
assign n_15213 = n_15050 ^ n_14605;
assign n_15214 = n_15050 & n_15051;
assign n_15215 = n_15052 ^ n_14607;
assign n_15216 = n_15052 & n_14942;
assign n_15217 = n_15053 ^ n_14609;
assign n_15218 = n_15053 & n_15054;
assign n_15219 = n_15055 ^ n_596;
assign n_15220 = n_15057 ^ n_14782;
assign n_15221 = n_15057 ^ n_14654;
assign n_15222 = ~n_14774 & n_15059;
assign n_15223 = n_14775 & n_15061;
assign n_15224 = n_14776 & n_15063;
assign n_15225 = n_14777 & n_15065;
assign n_15226 = ~n_14778 & n_15067;
assign n_15227 = ~n_14779 & n_15069;
assign n_15228 = n_14907 & ~n_15071;
assign n_15229 = n_15072 ^ n_14650;
assign n_15230 = ~n_15072 & n_14780;
assign n_15231 = n_15073 ^ n_14743;
assign n_15232 = n_15073 & ~n_14910;
assign n_15233 = ~n_14781 & n_15075;
assign n_15234 = n_15078 ^ n_14803;
assign n_15235 = n_14915 & ~n_15081;
assign n_15236 = n_14916 & ~n_15083;
assign n_15237 = ~n_14917 & n_15085;
assign n_15238 = n_14918 & ~n_15087;
assign n_15239 = ~n_14919 & n_15089;
assign n_15240 = n_14920 & n_15091;
assign n_15241 = n_14921 & ~n_15093;
assign n_15242 = n_14933 & ~n_15095;
assign n_15243 = n_15096 ^ n_14756;
assign n_15244 = n_15096 & ~n_14922;
assign n_15245 = n_15097 ^ n_14770;
assign n_15246 = n_15097 & n_14936;
assign n_15247 = n_15098 ^ n_14758;
assign n_15248 = ~n_15098 & n_14923;
assign n_15249 = n_15099 ^ n_14924;
assign n_15250 = n_15099 & n_15056;
assign n_15251 = n_15100 ^ x114;
assign n_15252 = n_15101 ^ x113;
assign n_15253 = n_15102 ^ n_14825;
assign n_15254 = ~x0 & n_15103;
assign n_15255 = n_15104 ^ x5;
assign n_15256 = n_15105 ^ x8;
assign n_15257 = n_15106 ^ x11;
assign n_15258 = n_15107 ^ x14;
assign n_15259 = n_15108 ^ x17;
assign n_15260 = n_15109 ^ x20;
assign n_15261 = n_15110 ^ x23;
assign n_15262 = n_15111 ^ x26;
assign n_15263 = n_15112 ^ x29;
assign n_15264 = n_15113 ^ x32;
assign n_15265 = n_15114 ^ x35;
assign n_15266 = n_15115 ^ x38;
assign n_15267 = n_15116 ^ x41;
assign n_15268 = n_15117 ^ x44;
assign n_15269 = n_15118 ^ x47;
assign n_15270 = n_15119 ^ x50;
assign n_15271 = n_15120 ^ x53;
assign n_15272 = n_15121 ^ x56;
assign n_15273 = n_15122 ^ x59;
assign n_15274 = n_15123 ^ x62;
assign n_15275 = n_15124 ^ x120;
assign n_15276 = n_2175 ^ n_15125;
assign n_15277 = n_775 ^ n_15126;
assign n_15278 = n_2246 ^ n_15127;
assign n_15279 = n_2314 ^ n_15128;
assign n_15280 = n_2381 ^ n_15129;
assign n_15281 = n_2448 ^ n_15130;
assign n_15282 = n_2515 ^ n_15131;
assign n_15283 = n_2581 ^ n_15132;
assign n_15284 = n_2646 ^ n_15133;
assign n_15285 = n_2713 ^ n_15134;
assign n_15286 = n_2781 ^ n_15135;
assign n_15287 = n_2848 ^ n_15136;
assign n_15288 = n_2916 ^ n_15137;
assign n_15289 = n_2982 ^ n_15138;
assign n_15290 = n_3051 ^ n_15139;
assign n_15291 = n_3117 ^ n_15140;
assign n_15292 = n_3186 ^ n_15141;
assign n_15293 = n_3250 ^ n_15142;
assign n_15294 = n_3315 ^ n_15143;
assign n_15295 = n_3380 ^ n_15144;
assign n_15296 = n_15145 ^ x5;
assign n_15297 = n_15146 ^ x8;
assign n_15298 = n_15147 ^ x11;
assign n_15299 = n_15148 ^ x14;
assign n_15300 = n_15149 ^ x17;
assign n_15301 = n_15150 ^ x20;
assign n_15302 = n_15151 ^ x23;
assign n_15303 = n_15152 ^ x26;
assign n_15304 = n_15153 ^ x29;
assign n_15305 = n_15154 ^ x32;
assign n_15306 = n_15155 ^ x35;
assign n_15307 = n_15156 ^ x38;
assign n_15308 = n_15157 ^ x41;
assign n_15309 = n_15158 ^ x44;
assign n_15310 = n_15159 ^ x47;
assign n_15311 = n_15160 ^ x50;
assign n_15312 = n_15161 ^ x53;
assign n_15313 = n_15162 ^ x56;
assign n_15314 = n_15163 ^ x59;
assign n_15315 = n_15164 ^ x62;
assign n_15316 = n_15165 ^ x1;
assign n_15317 = n_655 & n_15166;
assign n_15318 = n_784 & n_15166;
assign n_15319 = ~n_3665 & n_15166;
assign n_15320 = n_854 & n_15166;
assign n_15321 = n_920 & n_15166;
assign n_15322 = n_986 & n_15166;
assign n_15323 = n_1052 & n_15166;
assign n_15324 = n_1117 & n_15166;
assign n_15325 = n_1181 & n_15166;
assign n_15326 = n_1248 & n_15166;
assign n_15327 = n_1314 & n_15166;
assign n_15328 = n_1380 & n_15166;
assign n_15329 = n_1445 & n_15166;
assign n_15330 = n_1510 & n_15166;
assign n_15331 = n_1576 & n_15166;
assign n_15332 = n_1641 & n_15166;
assign n_15333 = n_1706 & n_15166;
assign n_15334 = n_1771 & n_15166;
assign n_15335 = n_1835 & n_15166;
assign n_15336 = n_15166 & n_1899;
assign n_15337 = ~x122 & ~n_15167;
assign n_15338 = ~x121 & n_15168;
assign n_15339 = n_15169 ^ n_14006;
assign n_15340 = n_15169 ^ n_13882;
assign n_15341 = n_15170 ^ n_10377;
assign n_15342 = ~n_13983 & n_15171;
assign n_15343 = n_15172 ^ n_10378;
assign n_15344 = ~n_13985 & n_15173;
assign n_15345 = n_15174 ^ n_10379;
assign n_15346 = n_13685 & ~n_15175;
assign n_15347 = n_15176 ^ n_10382;
assign n_15348 = ~n_13989 & n_15177;
assign n_15349 = n_15178 ^ n_10383;
assign n_15350 = ~n_13991 & n_15179;
assign n_15351 = n_15180 ^ n_10384;
assign n_15352 = ~n_13871 & n_15181;
assign n_15353 = n_15183 ^ n_14883;
assign n_15354 = n_15184 ^ n_12233;
assign n_15355 = ~n_13888 & n_15185;
assign n_15356 = n_15186 ^ n_14474;
assign n_15357 = ~n_14136 & n_15187;
assign n_15358 = n_15188 ^ n_14113;
assign n_15359 = n_15188 ^ n_13979;
assign n_15360 = n_15189 ^ n_14004;
assign n_15361 = n_15189 ^ n_13880;
assign n_15362 = n_15190 ^ n_10753;
assign n_15363 = ~n_14126 & n_15191;
assign n_15364 = n_15192 ^ n_10677;
assign n_15365 = ~n_14402 & n_15193;
assign n_15366 = n_15194 ^ n_10681;
assign n_15367 = ~n_14010 & n_15195;
assign n_15368 = n_15196 ^ n_10682;
assign n_15369 = ~n_14408 & n_15197;
assign n_15370 = n_15199 ^ n_14900;
assign n_15371 = n_15201 ^ n_14792;
assign n_15372 = n_15203 ^ n_14793;
assign n_15373 = n_15205 ^ n_14794;
assign n_15374 = n_15207 ^ n_14795;
assign n_15375 = n_15209 ^ n_14796;
assign n_15376 = n_15211 ^ n_14797;
assign n_15377 = n_15212 ^ n_14908;
assign n_15378 = n_15214 ^ n_14799;
assign n_15379 = n_15216 ^ n_14911;
assign n_15380 = n_15218 ^ n_14801;
assign n_15381 = ~n_14913 & ~n_15219;
assign n_15382 = n_14782 & n_15221;
assign n_15383 = n_15222 ^ n_14926;
assign n_15384 = n_15223 ^ n_14927;
assign n_15385 = n_15224 ^ n_14928;
assign n_15386 = n_15225 ^ n_14929;
assign n_15387 = n_15226 ^ n_14647;
assign n_15388 = n_15227 ^ n_14931;
assign n_15389 = n_15228 ^ n_14740;
assign n_15390 = n_15230 ^ n_14934;
assign n_15391 = n_15232 ^ n_14935;
assign n_15392 = n_15233 ^ n_14937;
assign n_15393 = n_15234 ^ n_14966;
assign n_15394 = n_15235 ^ n_14748;
assign n_15395 = n_15236 ^ n_14955;
assign n_15396 = n_15237 ^ n_14956;
assign n_15397 = n_15238 ^ n_14957;
assign n_15398 = n_15239 ^ n_14958;
assign n_15399 = n_15240 ^ n_14959;
assign n_15400 = n_15241 ^ n_14960;
assign n_15401 = n_15242 ^ n_14961;
assign n_15402 = n_15244 ^ n_14962;
assign n_15403 = n_15246 ^ n_14963;
assign n_15404 = n_15248 ^ n_14964;
assign n_15405 = n_15250 ^ n_14965;
assign n_15406 = n_67 & ~n_15251;
assign n_15407 = n_15252 ^ n_266;
assign n_15408 = n_15254 ^ n_14971;
assign n_15409 = n_15262 ^ n_15200;
assign n_15410 = n_15263 ^ n_15202;
assign n_15411 = n_15204 ^ n_15264;
assign n_15412 = n_15265 ^ n_15206;
assign n_15413 = n_15210 ^ n_15267;
assign n_15414 = n_15077 ^ n_15268;
assign n_15415 = n_15213 ^ n_15269;
assign n_15416 = n_15270 ^ n_15215;
assign n_15417 = n_15271 ^ n_15217;
assign n_15418 = n_15273 ^ n_14944;
assign n_15419 = n_15274 ^ n_6494;
assign n_15420 = n_15275 ^ n_2115;
assign n_15421 = n_5048 ^ n_15276;
assign n_15422 = n_5111 ^ n_15277;
assign n_15423 = n_5174 ^ n_15278;
assign n_15424 = n_5235 ^ n_15279;
assign n_15425 = n_5299 ^ n_15280;
assign n_15426 = n_5363 ^ n_15281;
assign n_15427 = n_5427 ^ n_15282;
assign n_15428 = n_5491 ^ n_15283;
assign n_15429 = n_5552 ^ n_15284;
assign n_15430 = n_5615 ^ n_15285;
assign n_15431 = n_5678 ^ n_15286;
assign n_15432 = n_5742 ^ n_15287;
assign n_15433 = n_5808 ^ n_15288;
assign n_15434 = n_5870 ^ n_15289;
assign n_15435 = n_5934 ^ n_15290;
assign n_15436 = n_5997 ^ n_15291;
assign n_15437 = n_6061 ^ n_15292;
assign n_15438 = n_6125 ^ n_15293;
assign n_15439 = n_6187 ^ n_15294;
assign n_15440 = n_6249 ^ n_15295;
assign n_15441 = n_15303 ^ n_15058;
assign n_15442 = n_15304 ^ n_15060;
assign n_15443 = n_15305 ^ n_15062;
assign n_15444 = n_15306 ^ n_15064;
assign n_15445 = n_15307 ^ n_15066;
assign n_15446 = n_15308 ^ n_15068;
assign n_15447 = n_15070 ^ n_15309;
assign n_15448 = n_15229 ^ n_15310;
assign n_15449 = n_15311 ^ n_15231;
assign n_15450 = n_15312 ^ n_15074;
assign n_15451 = n_15314 ^ n_15220;
assign n_15452 = n_15315 ^ n_6361;
assign n_15453 = n_15316 ^ x121;
assign n_15454 = n_2176 ^ n_15317;
assign n_15455 = n_776 ^ n_15318;
assign n_15456 = n_2247 ^ n_15319;
assign n_15457 = n_2315 ^ n_15320;
assign n_15458 = n_2382 ^ n_15321;
assign n_15459 = n_2449 ^ n_15322;
assign n_15460 = n_2516 ^ n_15323;
assign n_15461 = n_2582 ^ n_15324;
assign n_15462 = n_2647 ^ n_15325;
assign n_15463 = n_2714 ^ n_15326;
assign n_15464 = n_2782 ^ n_15327;
assign n_15465 = n_2849 ^ n_15328;
assign n_15466 = n_2917 ^ n_15329;
assign n_15467 = n_2983 ^ n_15330;
assign n_15468 = n_3052 ^ n_15331;
assign n_15469 = n_3118 ^ n_15332;
assign n_15470 = n_3187 ^ n_15333;
assign n_15471 = n_3251 ^ n_15334;
assign n_15472 = n_3316 ^ n_15335;
assign n_15473 = n_3381 ^ n_15336;
assign n_15474 = ~x124 & n_15337;
assign n_15475 = n_15167 ^ n_15338;
assign n_15476 = x122 & ~n_15338;
assign n_15477 = n_15339 ^ n_10676;
assign n_15478 = ~n_14006 & n_15340;
assign n_15479 = n_15342 ^ n_15018;
assign n_15480 = n_15344 ^ n_15019;
assign n_15481 = n_15346 ^ n_15020;
assign n_15482 = n_15348 ^ n_15021;
assign n_15483 = n_15350 ^ n_15022;
assign n_15484 = n_15352 ^ n_15023;
assign n_15485 = n_15353 ^ n_14415;
assign n_15486 = n_15353 ^ n_14261;
assign n_15487 = n_15355 ^ n_15026;
assign n_15488 = n_15357 ^ n_15027;
assign n_15489 = n_15358 ^ n_10675;
assign n_15490 = ~n_14113 & n_15359;
assign y27 = ~n_15360;
assign n_15491 = n_14004 & ~n_15361;
assign n_15492 = n_15363 ^ n_15031;
assign n_15493 = n_15365 ^ n_15032;
assign n_15494 = n_15367 ^ n_15033;
assign n_15495 = n_15369 ^ n_15034;
assign n_15496 = n_15370 ^ n_14417;
assign n_15497 = n_15370 ^ n_14263;
assign n_15498 = n_15371 ^ n_15082;
assign n_15499 = n_15372 ^ n_15084;
assign n_15500 = n_15373 ^ n_15086;
assign n_15501 = n_15374 ^ n_15088;
assign n_15502 = n_15375 ^ n_15090;
assign n_15503 = n_15376 ^ n_15092;
assign n_15504 = n_15377 ^ n_15094;
assign n_15505 = n_15378 ^ n_15243;
assign n_15506 = n_15247 ^ n_15380;
assign n_15507 = n_15381 ^ n_14312;
assign n_15508 = n_15381 ^ n_14178;
assign n_15509 = n_15382 ^ n_15057;
assign n_15510 = n_15262 ^ n_15383;
assign n_15511 = n_15202 ^ n_15384;
assign n_15512 = n_15385 ^ n_15204;
assign n_15513 = n_15386 ^ n_15265;
assign n_15514 = n_15387 ^ n_15208;
assign n_15515 = n_15387 ^ n_15266;
assign n_15516 = n_15388 ^ n_15210;
assign n_15517 = n_15389 ^ n_15077;
assign n_15518 = n_15390 ^ n_15213;
assign n_15519 = n_15215 ^ n_15391;
assign n_15520 = n_15217 ^ n_15392;
assign n_15521 = n_15394 ^ n_15303;
assign n_15522 = n_15395 ^ n_15304;
assign n_15523 = n_15396 ^ n_15305;
assign n_15524 = n_15397 ^ n_15306;
assign n_15525 = n_15398 ^ n_15066;
assign n_15526 = n_15399 ^ n_15308;
assign n_15527 = n_15400 ^ n_15070;
assign n_15528 = n_15401 ^ n_15310;
assign n_15529 = n_15402 ^ n_15311;
assign n_15530 = n_15403 ^ n_15312;
assign n_15531 = n_15405 ^ n_15314;
assign n_15532 = n_15406 ^ n_14968;
assign n_15533 = x62 & ~n_15407;
assign n_15534 = n_15409 ^ n_15383;
assign n_15535 = n_15410 ^ n_15384;
assign n_15536 = n_15416 ^ n_15391;
assign n_15537 = n_15417 ^ n_15392;
assign n_15538 = n_15419 ^ n_3417;
assign n_15539 = ~n_15419 & ~n_6609;
assign n_15540 = ~x0 & n_15420;
assign n_15541 = n_15421 ^ x5;
assign n_15542 = n_15422 ^ x8;
assign n_15543 = n_15423 ^ x11;
assign n_15544 = n_15424 ^ x14;
assign n_15545 = n_15425 ^ x17;
assign n_15546 = n_15426 ^ x20;
assign n_15547 = n_15427 ^ x23;
assign n_15548 = n_15428 ^ x26;
assign n_15549 = n_15429 ^ x29;
assign n_15550 = n_15430 ^ x32;
assign n_15551 = n_15431 ^ x35;
assign n_15552 = n_15432 ^ x38;
assign n_15553 = n_15433 ^ x41;
assign n_15554 = n_15434 ^ x44;
assign n_15555 = n_15435 ^ x47;
assign n_15556 = n_15436 ^ x50;
assign n_15557 = n_15437 ^ x53;
assign n_15558 = n_15438 ^ x56;
assign n_15559 = n_15439 ^ x59;
assign n_15560 = n_15440 ^ x62;
assign n_15561 = n_15394 ^ n_15441;
assign n_15562 = n_15395 ^ n_15442;
assign n_15563 = n_15396 ^ n_15443;
assign n_15564 = n_15397 ^ n_15444;
assign n_15565 = n_15398 ^ n_15445;
assign n_15566 = n_15399 ^ n_15446;
assign n_15567 = n_15401 ^ n_15448;
assign n_15568 = n_15453 ^ n_2116;
assign n_15569 = n_5049 ^ n_15454;
assign n_15570 = n_5112 ^ n_15455;
assign n_15571 = n_5175 ^ n_15456;
assign n_15572 = n_5236 ^ n_15457;
assign n_15573 = n_5300 ^ n_15458;
assign n_15574 = n_5364 ^ n_15459;
assign n_15575 = n_5428 ^ n_15460;
assign n_15576 = n_5492 ^ n_15461;
assign n_15577 = n_5553 ^ n_15462;
assign n_15578 = n_5616 ^ n_15463;
assign n_15579 = n_5679 ^ n_15464;
assign n_15580 = n_5743 ^ n_15465;
assign n_15581 = n_5809 ^ n_15466;
assign n_15582 = n_5871 ^ n_15467;
assign n_15583 = n_5935 ^ n_15468;
assign n_15584 = n_5998 ^ n_15469;
assign n_15585 = n_6062 ^ n_15470;
assign n_15586 = n_6126 ^ n_15471;
assign n_15587 = n_6188 ^ n_15472;
assign n_15588 = n_6250 ^ n_15473;
assign n_15589 = n_1 & n_15475;
assign n_15590 = n_15475 ^ x122;
assign n_15591 = n_15337 ^ n_15476;
assign n_15592 = x124 & n_15476;
assign n_15593 = n_15478 ^ n_15169;
assign n_15594 = n_15479 ^ n_14404;
assign n_15595 = n_15479 ^ n_14249;
assign n_15596 = n_15480 ^ n_14406;
assign n_15597 = n_15480 ^ n_14251;
assign n_15598 = n_15481 ^ n_14008;
assign n_15599 = n_15481 ^ n_13884;
assign n_15600 = n_15482 ^ n_14410;
assign n_15601 = n_15482 ^ n_14255;
assign n_15602 = n_15483 ^ n_14412;
assign n_15603 = n_15483 ^ n_14257;
assign n_15604 = n_15484 ^ n_14259;
assign n_15605 = n_15484 ^ n_14121;
assign n_15606 = n_15485 ^ n_11135;
assign n_15607 = n_14415 & ~n_15486;
assign n_15608 = n_15487 ^ n_14276;
assign n_15609 = n_15487 ^ n_14133;
assign n_15610 = n_15488 ^ n_14301;
assign n_15611 = n_15488 ^ n_13998;
assign n_15612 = n_15490 ^ n_15188;
assign n_15613 = n_15491 ^ n_15189;
assign n_15614 = n_15492 ^ n_14567;
assign n_15615 = n_15492 ^ n_14420;
assign n_15616 = n_15493 ^ n_14871;
assign n_15617 = n_15493 ^ n_14704;
assign n_15618 = n_15494 ^ n_14430;
assign n_15619 = n_15494 ^ n_14274;
assign n_15620 = n_15495 ^ n_14877;
assign n_15621 = n_15495 ^ n_14710;
assign n_15622 = n_15496 ^ n_13468;
assign n_15623 = ~n_14417 & n_15497;
assign n_15624 = n_15507 ^ n_15076;
assign n_15625 = n_15507 ^ n_14653;
assign n_15626 = n_14312 & n_15508;
assign n_15627 = n_15509 ^ n_15418;
assign n_15628 = n_15509 ^ n_15273;
assign n_15629 = ~n_15409 & n_15510;
assign n_15630 = n_15410 & ~n_15511;
assign n_15631 = n_15512 ^ n_15264;
assign n_15632 = ~n_15512 & n_15411;
assign n_15633 = n_15513 ^ n_15206;
assign n_15634 = n_15513 & ~n_15412;
assign n_15635 = n_15514 ^ n_15266;
assign n_15636 = ~n_15514 & n_15515;
assign n_15637 = n_15516 ^ n_15267;
assign n_15638 = n_15516 & ~n_15413;
assign n_15639 = n_15517 ^ n_15268;
assign n_15640 = ~n_15517 & n_15414;
assign n_15641 = n_15518 ^ n_15269;
assign n_15642 = ~n_15518 & n_15415;
assign n_15643 = ~n_15416 & n_15519;
assign n_15644 = ~n_15417 & n_15520;
assign n_15645 = ~n_15441 & n_15521;
assign n_15646 = n_15442 & n_15522;
assign n_15647 = n_15443 & n_15523;
assign n_15648 = n_15444 & n_15524;
assign n_15649 = ~n_15445 & n_15525;
assign n_15650 = ~n_15446 & n_15526;
assign n_15651 = n_15527 ^ n_15309;
assign n_15652 = n_15527 & ~n_15447;
assign n_15653 = ~n_15448 & ~n_15528;
assign n_15654 = n_15529 ^ n_15231;
assign n_15655 = n_15529 & ~n_15449;
assign n_15656 = n_15530 ^ n_15074;
assign n_15657 = n_15530 & ~n_15450;
assign n_15658 = n_15531 ^ n_15220;
assign n_15659 = n_15531 & n_15451;
assign n_15660 = n_15533 ^ n_266;
assign n_15661 = n_15539 ^ n_15274;
assign n_15662 = n_15540 ^ n_15275;
assign n_15663 = n_15080 ^ n_15547;
assign n_15664 = n_15548 ^ n_15498;
assign n_15665 = n_15548 ^ n_15082;
assign n_15666 = n_15549 ^ n_15499;
assign n_15667 = n_15549 ^ n_15084;
assign n_15668 = n_15550 ^ n_15500;
assign n_15669 = n_15550 ^ n_15373;
assign n_15670 = n_15551 ^ n_15501;
assign n_15671 = n_15551 ^ n_15374;
assign n_15672 = n_15552 ^ n_15502;
assign n_15673 = n_15552 ^ n_15090;
assign n_15674 = n_15553 ^ n_15503;
assign n_15675 = n_15553 ^ n_15092;
assign n_15676 = n_15554 ^ n_15504;
assign n_15677 = n_15554 ^ n_15094;
assign n_15678 = n_15555 ^ n_15505;
assign n_15679 = n_15555 ^ n_15378;
assign n_15680 = n_15556 ^ n_15379;
assign n_15681 = n_15556 ^ n_15245;
assign n_15682 = n_15557 ^ n_15247;
assign n_15683 = n_15558 ^ n_15249;
assign n_15684 = n_15559 ^ n_15393;
assign n_15685 = n_15559 ^ n_15234;
assign n_15686 = ~x0 & n_15568;
assign n_15687 = n_15569 ^ x5;
assign n_15688 = n_15570 ^ x8;
assign n_15689 = n_15571 ^ x11;
assign n_15690 = n_15572 ^ x14;
assign n_15691 = n_15573 ^ x17;
assign n_15692 = n_15574 ^ x20;
assign n_15693 = n_15575 ^ x23;
assign n_15694 = n_15576 ^ x26;
assign n_15695 = n_15577 ^ x29;
assign n_15696 = n_15578 ^ x32;
assign n_15697 = n_15579 ^ x35;
assign n_15698 = n_15580 ^ x38;
assign n_15699 = n_15581 ^ x41;
assign n_15700 = n_15582 ^ x44;
assign n_15701 = n_15583 ^ x47;
assign n_15702 = n_15584 ^ x50;
assign n_15703 = n_15585 ^ x53;
assign n_15704 = n_15586 ^ x56;
assign n_15705 = n_15587 ^ x59;
assign n_15706 = n_15588 ^ x62;
assign n_15707 = n_15589 ^ x1;
assign n_15708 = n_655 & ~n_15590;
assign n_15709 = n_784 & ~n_15590;
assign n_15710 = ~n_3665 & ~n_15590;
assign n_15711 = n_854 & ~n_15590;
assign n_15712 = n_920 & ~n_15590;
assign n_15713 = n_986 & ~n_15590;
assign n_15714 = n_1052 & ~n_15590;
assign n_15715 = n_1117 & ~n_15590;
assign n_15716 = n_1181 & ~n_15590;
assign n_15717 = n_1248 & ~n_15590;
assign n_15718 = n_1314 & ~n_15590;
assign n_15719 = n_1380 & ~n_15590;
assign n_15720 = n_1445 & ~n_15590;
assign n_15721 = n_1510 & ~n_15590;
assign n_15722 = n_1576 & ~n_15590;
assign n_15723 = n_1641 & ~n_15590;
assign n_15724 = n_1706 & ~n_15590;
assign n_15725 = n_1771 & ~n_15590;
assign n_15726 = n_1835 & ~n_15590;
assign n_15727 = ~n_15590 & n_1899;
assign n_15728 = n_1 & n_15591;
assign n_15729 = n_15591 & n_286;
assign n_15730 = n_15591 ^ x123;
assign n_15731 = ~x123 & ~n_15592;
assign n_15732 = n_15593 ^ n_14426;
assign n_15733 = n_15593 ^ n_14270;
assign n_15734 = n_15594 ^ n_10678;
assign n_15735 = n_14404 & ~n_15595;
assign n_15736 = n_15596 ^ n_10679;
assign n_15737 = ~n_14406 & n_15597;
assign n_15738 = n_15598 ^ n_10680;
assign n_15739 = n_14008 & ~n_15599;
assign n_15740 = n_15600 ^ n_10683;
assign n_15741 = n_14410 & ~n_15601;
assign n_15742 = n_15602 ^ n_10684;
assign n_15743 = n_14412 & ~n_15603;
assign n_15744 = n_15604 ^ n_10685;
assign n_15745 = ~n_14259 & n_15605;
assign n_15746 = n_15607 ^ n_15353;
assign n_15747 = n_15608 ^ n_12525;
assign n_15748 = n_14276 & ~n_15609;
assign n_15749 = n_15610 ^ n_14642;
assign n_15750 = ~n_14301 & n_15611;
assign n_15751 = n_15612 ^ n_14554;
assign n_15752 = n_15612 ^ n_14400;
assign n_15753 = n_15613 ^ n_14424;
assign n_15754 = n_15613 ^ n_14268;
assign n_15755 = n_15614 ^ n_10852;
assign n_15756 = ~n_14567 & n_15615;
assign n_15757 = n_15616 ^ n_10780;
assign n_15758 = ~n_14871 & n_15617;
assign n_15759 = n_15618 ^ n_10784;
assign n_15760 = ~n_14430 & n_15619;
assign n_15761 = n_15620 ^ n_10785;
assign n_15762 = ~n_14877 & n_15621;
assign n_15763 = n_15623 ^ n_15370;
assign n_15764 = n_15624 ^ n_15313;
assign n_15765 = n_15624 ^ n_15404;
assign n_15766 = n_15076 & n_15625;
assign n_15767 = n_15626 ^ n_15381;
assign n_15768 = n_15418 & n_15628;
assign n_15769 = n_15629 ^ n_15383;
assign n_15770 = n_15630 ^ n_15263;
assign n_15771 = n_15632 ^ n_15385;
assign n_15772 = n_15634 ^ n_15386;
assign n_15773 = n_15636 ^ n_15266;
assign n_15774 = n_15638 ^ n_15388;
assign n_15775 = n_15640 ^ n_15389;
assign n_15776 = n_15642 ^ n_15390;
assign n_15777 = n_15643 ^ n_15270;
assign n_15778 = n_15644 ^ n_15271;
assign n_15779 = n_15645 ^ n_15394;
assign n_15780 = n_15646 ^ n_15395;
assign n_15781 = n_15647 ^ n_15396;
assign n_15782 = n_15648 ^ n_15397;
assign n_15783 = n_15649 ^ n_15307;
assign n_15784 = n_15650 ^ n_15399;
assign n_15785 = n_15652 ^ n_15400;
assign n_15786 = n_15653 ^ n_15229;
assign n_15787 = n_15655 ^ n_15402;
assign n_15788 = n_15657 ^ n_15403;
assign n_15789 = n_15659 ^ n_15405;
assign n_15790 = x63 & n_15660;
assign n_15791 = n_15661 ^ ~n_6537;
assign n_15792 = ~n_6537 & ~n_15661;
assign n_15793 = n_15498 & ~n_15665;
assign n_15794 = ~n_15499 & n_15667;
assign n_15795 = n_15500 & n_15669;
assign n_15796 = n_15501 & ~n_15671;
assign n_15797 = n_15502 & ~n_15673;
assign n_15798 = n_15503 & ~n_15675;
assign n_15799 = ~n_15504 & n_15677;
assign n_15800 = n_15505 & ~n_15679;
assign n_15801 = n_15680 ^ n_15245;
assign n_15802 = n_15680 & n_15681;
assign n_15803 = n_15682 ^ n_15380;
assign n_15804 = ~n_15682 & n_15506;
assign n_15805 = n_15393 & n_15685;
assign n_15806 = n_15686 ^ n_15453;
assign n_15807 = n_15561 ^ n_15693;
assign n_15808 = n_15562 ^ n_15694;
assign n_15809 = n_15563 ^ n_15695;
assign n_15810 = n_15564 ^ n_15696;
assign n_15811 = n_15565 ^ n_15697;
assign n_15812 = n_15566 ^ n_15698;
assign n_15813 = n_15651 ^ n_15699;
assign n_15814 = n_15700 ^ n_15567;
assign n_15815 = n_15654 ^ n_15701;
assign n_15816 = n_15702 ^ n_15656;
assign n_15817 = n_15658 ^ n_15704;
assign n_15818 = n_15706 ^ n_6419;
assign n_15819 = n_15707 ^ x122;
assign n_15820 = n_2177 ^ n_15708;
assign n_15821 = n_777 ^ n_15709;
assign n_15822 = n_2248 ^ n_15710;
assign n_15823 = n_2316 ^ n_15711;
assign n_15824 = n_2383 ^ n_15712;
assign n_15825 = n_2450 ^ n_15713;
assign n_15826 = n_2517 ^ n_15714;
assign n_15827 = n_2583 ^ n_15715;
assign n_15828 = n_2648 ^ n_15716;
assign n_15829 = n_2715 ^ n_15717;
assign n_15830 = n_2783 ^ n_15718;
assign n_15831 = n_2850 ^ n_15719;
assign n_15832 = n_2918 ^ n_15720;
assign n_15833 = n_2984 ^ n_15721;
assign n_15834 = n_3053 ^ n_15722;
assign n_15835 = n_3119 ^ n_15723;
assign n_15836 = n_3188 ^ n_15724;
assign n_15837 = n_3252 ^ n_15725;
assign n_15838 = n_3317 ^ n_15726;
assign n_15839 = n_3382 ^ n_15727;
assign n_15840 = n_15728 ^ x1;
assign n_15841 = n_1 & ~n_15729;
assign n_15842 = n_15729 ^ x124;
assign n_15843 = n_655 & ~n_15730;
assign n_15844 = n_784 & ~n_15730;
assign n_15845 = ~n_3665 & ~n_15730;
assign n_15846 = n_854 & ~n_15730;
assign n_15847 = n_920 & ~n_15730;
assign n_15848 = n_986 & ~n_15730;
assign n_15849 = n_1052 & ~n_15730;
assign n_15850 = n_1117 & ~n_15730;
assign n_15851 = n_1181 & ~n_15730;
assign n_15852 = n_1248 & ~n_15730;
assign n_15853 = n_1314 & ~n_15730;
assign n_15854 = n_1380 & ~n_15730;
assign n_15855 = n_1445 & ~n_15730;
assign n_15856 = n_1510 & ~n_15730;
assign n_15857 = n_1576 & ~n_15730;
assign n_15858 = n_1641 & ~n_15730;
assign n_15859 = n_1706 & ~n_15730;
assign n_15860 = n_1771 & ~n_15730;
assign n_15861 = n_1835 & ~n_15730;
assign n_15862 = ~n_15730 & n_1899;
assign n_15863 = ~n_15474 & ~n_15731;
assign n_15864 = ~n_15731 & n_616;
assign n_15865 = n_15732 ^ n_10779;
assign n_15866 = ~n_14426 & n_15733;
assign n_15867 = n_15735 ^ n_15479;
assign n_15868 = n_15737 ^ n_15480;
assign n_15869 = n_15739 ^ n_15481;
assign n_15870 = n_15741 ^ n_15482;
assign n_15871 = n_15743 ^ n_15483;
assign n_15872 = n_15745 ^ n_15484;
assign n_15873 = n_15746 ^ n_14884;
assign n_15874 = n_15746 ^ n_14718;
assign n_15875 = n_15748 ^ n_15487;
assign n_15876 = n_15750 ^ n_15488;
assign n_15877 = n_15751 ^ n_10778;
assign n_15878 = ~n_14554 & n_15752;
assign y28 = n_15753;
assign n_15879 = ~n_14424 & n_15754;
assign n_15880 = n_15756 ^ n_15492;
assign n_15881 = n_15758 ^ n_15493;
assign n_15882 = n_15760 ^ n_15494;
assign n_15883 = n_15762 ^ n_15495;
assign n_15884 = n_15763 ^ n_14886;
assign n_15885 = n_15763 ^ n_14720;
assign n_15886 = n_15764 ^ n_15404;
assign n_15887 = n_15764 & ~n_15765;
assign n_15888 = n_15766 ^ n_14938;
assign n_15889 = n_15767 ^ n_14943;
assign n_15890 = n_15767 ^ n_14611;
assign n_15891 = n_15768 ^ n_15509;
assign n_15892 = n_15769 ^ n_15664;
assign n_15893 = n_15770 ^ n_15666;
assign n_15894 = n_15771 ^ n_15668;
assign n_15895 = n_15772 ^ n_15670;
assign n_15896 = n_15773 ^ n_15672;
assign n_15897 = n_15774 ^ n_15674;
assign n_15898 = n_15775 ^ n_15676;
assign n_15899 = n_15776 ^ n_15678;
assign n_15900 = n_15779 ^ n_15534;
assign n_15901 = n_15780 ^ n_15535;
assign n_15902 = n_15781 ^ n_15631;
assign n_15903 = n_15782 ^ n_15633;
assign n_15904 = n_15783 ^ n_15635;
assign n_15905 = n_15784 ^ n_15637;
assign n_15906 = n_15785 ^ n_15639;
assign n_15907 = n_15786 ^ n_15641;
assign n_15908 = n_15536 ^ n_15787;
assign n_15909 = n_15788 ^ n_15537;
assign n_15910 = ~n_15532 & ~n_15790;
assign n_15911 = n_15560 ^ n_15791;
assign n_15912 = n_15792 ^ n_6418;
assign n_15913 = n_15793 ^ n_15548;
assign n_15914 = n_15794 ^ n_15549;
assign n_15915 = n_15795 ^ n_15550;
assign n_15916 = n_15796 ^ n_15088;
assign n_15917 = n_15797 ^ n_15552;
assign n_15918 = n_15798 ^ n_15553;
assign n_15919 = n_15799 ^ n_15377;
assign n_15920 = n_15800 ^ n_15243;
assign n_15921 = n_15801 ^ n_15777;
assign n_15922 = n_15802 ^ n_15379;
assign n_15923 = n_15803 ^ n_15778;
assign n_15924 = n_15804 ^ n_15557;
assign n_15925 = n_15805 ^ n_15559;
assign n_15926 = n_15819 ^ n_2117;
assign n_15927 = n_5050 ^ n_15820;
assign n_15928 = n_5113 ^ n_15821;
assign n_15929 = n_5176 ^ n_15822;
assign n_15930 = n_5237 ^ n_15823;
assign n_15931 = n_5301 ^ n_15824;
assign n_15932 = n_5365 ^ n_15825;
assign n_15933 = n_5429 ^ n_15826;
assign n_15934 = n_5493 ^ n_15827;
assign n_15935 = n_5554 ^ n_15828;
assign n_15936 = n_5617 ^ n_15829;
assign n_15937 = n_5680 ^ n_15830;
assign n_15938 = n_5744 ^ n_15831;
assign n_15939 = n_5810 ^ n_15832;
assign n_15940 = n_5872 ^ n_15833;
assign n_15941 = n_5936 ^ n_15834;
assign n_15942 = n_5999 ^ n_15835;
assign n_15943 = n_6063 ^ n_15836;
assign n_15944 = n_6127 ^ n_15837;
assign n_15945 = n_6189 ^ n_15838;
assign n_15946 = n_6251 ^ n_15839;
assign n_15947 = n_15840 ^ x123;
assign n_15948 = n_15841 ^ x1;
assign n_15949 = n_655 & n_15842;
assign n_15950 = n_784 & n_15842;
assign n_15951 = ~n_3665 & n_15842;
assign n_15952 = n_854 & n_15842;
assign n_15953 = n_920 & n_15842;
assign n_15954 = n_986 & n_15842;
assign n_15955 = n_1052 & n_15842;
assign n_15956 = n_1117 & n_15842;
assign n_15957 = n_1181 & n_15842;
assign n_15958 = n_1248 & n_15842;
assign n_15959 = n_1314 & n_15842;
assign n_15960 = n_1380 & n_15842;
assign n_15961 = n_1445 & n_15842;
assign n_15962 = n_1510 & n_15842;
assign n_15963 = n_1576 & n_15842;
assign n_15964 = n_1641 & n_15842;
assign n_15965 = n_1706 & n_15842;
assign n_15966 = n_1771 & n_15842;
assign n_15967 = n_1835 & n_15842;
assign n_15968 = n_1899 & n_15842;
assign n_15969 = n_2178 ^ n_15843;
assign n_15970 = n_778 ^ n_15844;
assign n_15971 = n_2249 ^ n_15845;
assign n_15972 = n_2317 ^ n_15846;
assign n_15973 = n_2384 ^ n_15847;
assign n_15974 = n_2451 ^ n_15848;
assign n_15975 = n_2518 ^ n_15849;
assign n_15976 = n_2584 ^ n_15850;
assign n_15977 = n_2649 ^ n_15851;
assign n_15978 = n_2716 ^ n_15852;
assign n_15979 = n_2784 ^ n_15853;
assign n_15980 = n_2851 ^ n_15854;
assign n_15981 = n_2919 ^ n_15855;
assign n_15982 = n_2985 ^ n_15856;
assign n_15983 = n_3054 ^ n_15857;
assign n_15984 = n_3120 ^ n_15858;
assign n_15985 = n_3189 ^ n_15859;
assign n_15986 = n_3253 ^ n_15860;
assign n_15987 = n_3318 ^ n_15861;
assign n_15988 = n_3383 ^ n_15862;
assign n_15989 = n_15863 ^ x124;
assign n_15990 = ~n_15863 & n_292;
assign n_15991 = n_293 ^ n_15863;
assign n_15992 = ~n_15864 & n_617;
assign n_15993 = n_15866 ^ n_15593;
assign n_15994 = n_15867 ^ n_14873;
assign n_15995 = n_15867 ^ n_14706;
assign n_15996 = n_15868 ^ n_14875;
assign n_15997 = n_15868 ^ n_14708;
assign n_15998 = n_15869 ^ n_14428;
assign n_15999 = n_15869 ^ n_14272;
assign n_16000 = n_15870 ^ n_14879;
assign n_16001 = n_15870 ^ n_14712;
assign n_16002 = n_15871 ^ n_14881;
assign n_16003 = n_15871 ^ n_14714;
assign n_16004 = n_15872 ^ n_14716;
assign n_16005 = n_15872 ^ n_14562;
assign n_16006 = n_15873 ^ n_11890;
assign n_16007 = n_14884 & ~n_15874;
assign n_16008 = n_15875 ^ n_14732;
assign n_16009 = n_15875 ^ n_14574;
assign n_16010 = n_15876 ^ n_14940;
assign n_16011 = n_15876 ^ n_14566;
assign n_16012 = n_15878 ^ n_15612;
assign n_16013 = n_15879 ^ n_15613;
assign n_16014 = n_15880 ^ n_15028;
assign n_16015 = n_15880 ^ n_14888;
assign n_16016 = n_15881 ^ n_15341;
assign n_16017 = n_15881 ^ n_15170;
assign n_16018 = n_15882 ^ n_14898;
assign n_16019 = n_15882 ^ n_14730;
assign n_16020 = n_15883 ^ n_15347;
assign n_16021 = n_15883 ^ n_15176;
assign n_16022 = n_15884 ^ n_14321;
assign n_16023 = ~n_14886 & n_15885;
assign n_16024 = n_15703 ^ n_15886;
assign n_16025 = n_15887 ^ n_15404;
assign n_16026 = n_15889 ^ n_15272;
assign n_16027 = n_15889 ^ n_15888;
assign n_16028 = n_14943 & ~n_15890;
assign n_16029 = n_15684 ^ n_15891;
assign n_16030 = n_15910 ^ n_15452;
assign n_16031 = n_15910 ^ n_15315;
assign n_16032 = n_15912 ^ n_15818;
assign n_16033 = n_15912 ^ n_15706;
assign n_16034 = n_15913 ^ n_15562;
assign n_16035 = n_15914 ^ n_15563;
assign n_16036 = n_15915 ^ n_15564;
assign n_16037 = n_15916 ^ n_15565;
assign n_16038 = n_15917 ^ n_15566;
assign n_16039 = n_15918 ^ n_15651;
assign n_16040 = n_15919 ^ n_15814;
assign n_16041 = n_15919 ^ n_15700;
assign n_16042 = n_15920 ^ n_15815;
assign n_16043 = n_15920 ^ n_15701;
assign n_16044 = n_15922 ^ n_15702;
assign n_16045 = n_15924 ^ n_15703;
assign n_16046 = n_15925 ^ n_15705;
assign n_16047 = ~x0 & n_15926;
assign n_16048 = n_15927 ^ x5;
assign n_16049 = n_15928 ^ x8;
assign n_16050 = n_15929 ^ x11;
assign n_16051 = n_15930 ^ x14;
assign n_16052 = n_15931 ^ x17;
assign n_16053 = n_15932 ^ x20;
assign n_16054 = n_15933 ^ x23;
assign n_16055 = n_15934 ^ x26;
assign n_16056 = n_15935 ^ x29;
assign n_16057 = n_15936 ^ x32;
assign n_16058 = n_15937 ^ x35;
assign n_16059 = n_15938 ^ x38;
assign n_16060 = n_15939 ^ x41;
assign n_16061 = n_15940 ^ x44;
assign n_16062 = n_15941 ^ x47;
assign n_16063 = n_15942 ^ x50;
assign n_16064 = n_15943 ^ x53;
assign n_16065 = n_15944 ^ x56;
assign n_16066 = n_15945 ^ x59;
assign n_16067 = n_15946 ^ x62;
assign n_16068 = n_15947 ^ n_2118;
assign n_16069 = n_15948 ^ x124;
assign n_16070 = n_2179 ^ n_15949;
assign n_16071 = n_779 ^ n_15950;
assign n_16072 = n_2250 ^ n_15951;
assign n_16073 = n_2318 ^ n_15952;
assign n_16074 = n_2385 ^ n_15953;
assign n_16075 = n_2452 ^ n_15954;
assign n_16076 = n_2519 ^ n_15955;
assign n_16077 = n_2585 ^ n_15956;
assign n_16078 = n_2650 ^ n_15957;
assign n_16079 = n_2717 ^ n_15958;
assign n_16080 = n_2785 ^ n_15959;
assign n_16081 = n_2852 ^ n_15960;
assign n_16082 = n_2920 ^ n_15961;
assign n_16083 = n_2986 ^ n_15962;
assign n_16084 = n_3055 ^ n_15963;
assign n_16085 = n_3121 ^ n_15964;
assign n_16086 = n_3190 ^ n_15965;
assign n_16087 = n_3254 ^ n_15966;
assign n_16088 = n_3319 ^ n_15967;
assign n_16089 = n_3384 ^ n_15968;
assign n_16090 = n_5051 ^ n_15969;
assign n_16091 = n_5114 ^ n_15970;
assign n_16092 = n_5177 ^ n_15971;
assign n_16093 = n_5238 ^ n_15972;
assign n_16094 = n_5302 ^ n_15973;
assign n_16095 = n_5366 ^ n_15974;
assign n_16096 = n_5430 ^ n_15975;
assign n_16097 = n_5494 ^ n_15976;
assign n_16098 = n_5555 ^ n_15977;
assign n_16099 = n_5618 ^ n_15978;
assign n_16100 = n_5681 ^ n_15979;
assign n_16101 = n_5745 ^ n_15980;
assign n_16102 = n_5811 ^ n_15981;
assign n_16103 = n_5873 ^ n_15982;
assign n_16104 = n_5937 ^ n_15983;
assign n_16105 = n_6000 ^ n_15984;
assign n_16106 = n_6064 ^ n_15985;
assign n_16107 = n_6128 ^ n_15986;
assign n_16108 = n_6190 ^ n_15987;
assign n_16109 = n_6252 ^ n_15988;
assign n_16110 = n_1 & ~n_15989;
assign n_16111 = n_15990 ^ n_15864;
assign n_16112 = ~n_15990 & n_296;
assign n_16113 = n_655 & n_15991;
assign n_16114 = n_784 & n_15991;
assign n_16115 = ~n_3665 & n_15991;
assign n_16116 = n_854 & n_15991;
assign n_16117 = n_920 & n_15991;
assign n_16118 = n_986 & n_15991;
assign n_16119 = n_1052 & n_15991;
assign n_16120 = n_1117 & n_15991;
assign n_16121 = n_1181 & n_15991;
assign n_16122 = n_1248 & n_15991;
assign n_16123 = n_1314 & n_15991;
assign n_16124 = n_1380 & n_15991;
assign n_16125 = n_1445 & n_15991;
assign n_16126 = n_1510 & n_15991;
assign n_16127 = n_1576 & n_15991;
assign n_16128 = n_1641 & n_15991;
assign n_16129 = n_1706 & n_15991;
assign n_16130 = n_1771 & n_15991;
assign n_16131 = n_1835 & n_15991;
assign n_16132 = n_1899 & n_15991;
assign n_16133 = ~n_15992 & n_622;
assign n_16134 = n_15993 ^ n_14894;
assign n_16135 = n_15993 ^ n_14726;
assign n_16136 = n_15994 ^ n_10781;
assign n_16137 = ~n_14873 & n_15995;
assign n_16138 = n_15996 ^ n_10782;
assign n_16139 = ~n_14875 & n_15997;
assign n_16140 = n_15998 ^ n_10783;
assign n_16141 = ~n_14428 & n_15999;
assign n_16142 = n_16000 ^ n_10786;
assign n_16143 = ~n_14879 & n_16001;
assign n_16144 = n_16002 ^ n_10787;
assign n_16145 = ~n_14881 & n_16003;
assign n_16146 = n_16004 ^ n_10788;
assign n_16147 = ~n_14716 & n_16005;
assign n_16148 = n_16007 ^ n_15746;
assign n_16149 = n_16008 ^ n_13127;
assign n_16150 = n_14732 & ~n_16009;
assign n_16151 = n_16010 ^ n_15261;
assign n_16152 = n_14940 & ~n_16011;
assign n_16153 = n_16012 ^ n_15016;
assign n_16154 = n_16012 ^ n_14869;
assign n_16155 = n_16013 ^ n_14892;
assign n_16156 = n_16013 ^ n_14724;
assign n_16157 = n_16014 ^ n_10954;
assign n_16158 = ~n_15028 & n_16015;
assign n_16159 = n_16016 ^ n_10856;
assign n_16160 = ~n_15341 & n_16017;
assign n_16161 = n_16018 ^ n_10860;
assign n_16162 = ~n_14898 & n_16019;
assign n_16163 = n_16020 ^ n_10861;
assign n_16164 = ~n_15347 & n_16021;
assign n_16165 = n_16023 ^ n_15763;
assign n_16166 = n_16026 ^ n_15888;
assign n_16167 = n_16026 & ~n_16027;
assign n_16168 = n_16028 ^ n_14802;
assign n_16169 = n_15705 ^ n_16030;
assign n_16170 = n_15452 & n_16031;
assign n_16171 = n_15818 & ~n_16033;
assign n_16172 = n_16034 ^ n_15694;
assign n_16173 = ~n_16034 & n_15808;
assign n_16174 = n_16035 ^ n_15695;
assign n_16175 = ~n_16035 & n_15809;
assign n_16176 = n_16036 ^ n_15696;
assign n_16177 = ~n_16036 & n_15810;
assign n_16178 = n_16037 ^ n_15697;
assign n_16179 = ~n_16037 & n_15811;
assign n_16180 = n_16038 ^ n_15698;
assign n_16181 = n_16038 & ~n_15812;
assign n_16182 = n_16039 ^ n_15699;
assign n_16183 = n_16039 & ~n_15813;
assign n_16184 = n_15814 & n_16041;
assign n_16185 = n_15815 & ~n_16043;
assign n_16186 = n_16044 ^ n_15656;
assign n_16187 = n_16044 & ~n_15816;
assign n_16188 = n_16045 ^ n_15886;
assign n_16189 = n_16045 & n_16024;
assign n_16190 = n_16046 ^ n_16030;
assign n_16191 = n_16047 ^ n_15819;
assign n_16192 = n_16048 ^ n_15256;
assign n_16193 = n_15900 ^ n_16054;
assign n_16194 = n_15534 ^ n_16054;
assign n_16195 = n_15901 ^ n_16055;
assign n_16196 = n_15780 ^ n_16055;
assign n_16197 = n_15902 ^ n_16056;
assign n_16198 = n_15781 ^ n_16056;
assign n_16199 = n_15903 ^ n_16057;
assign n_16200 = n_15782 ^ n_16057;
assign n_16201 = n_15904 ^ n_16058;
assign n_16202 = n_15783 ^ n_16058;
assign n_16203 = n_15905 ^ n_16059;
assign n_16204 = n_15784 ^ n_16059;
assign n_16205 = n_15906 ^ n_16060;
assign n_16206 = n_15785 ^ n_16060;
assign n_16207 = n_15907 ^ n_16061;
assign n_16208 = n_15786 ^ n_16061;
assign n_16209 = n_16062 ^ n_15536;
assign n_16210 = n_15909 ^ n_16063;
assign n_16211 = n_15537 ^ n_16063;
assign n_16212 = n_16065 ^ n_15789;
assign n_16213 = n_16065 ^ n_15627;
assign n_16214 = n_16066 ^ n_15538;
assign n_16215 = n_16067 ^ n_6647;
assign n_16216 = n_16067 ^ n_6538;
assign n_16217 = ~x0 & n_16068;
assign n_16218 = n_16069 ^ n_2119;
assign n_16219 = n_5052 ^ n_16070;
assign n_16220 = n_5115 ^ n_16071;
assign n_16221 = n_5178 ^ n_16072;
assign n_16222 = n_5239 ^ n_16073;
assign n_16223 = n_5303 ^ n_16074;
assign n_16224 = n_5367 ^ n_16075;
assign n_16225 = n_5431 ^ n_16076;
assign n_16226 = n_5495 ^ n_16077;
assign n_16227 = n_5556 ^ n_16078;
assign n_16228 = n_5619 ^ n_16079;
assign n_16229 = n_5682 ^ n_16080;
assign n_16230 = n_5746 ^ n_16081;
assign n_16231 = n_5812 ^ n_16082;
assign n_16232 = n_5874 ^ n_16083;
assign n_16233 = n_5938 ^ n_16084;
assign n_16234 = n_6001 ^ n_16085;
assign n_16235 = n_6065 ^ n_16086;
assign n_16236 = n_6129 ^ n_16087;
assign n_16237 = n_6191 ^ n_16088;
assign n_16238 = n_6253 ^ n_16089;
assign n_16239 = n_16090 ^ x5;
assign n_16240 = n_16091 ^ x8;
assign n_16241 = n_16092 ^ x11;
assign n_16242 = n_16093 ^ x14;
assign n_16243 = n_16094 ^ x17;
assign n_16244 = n_16095 ^ x20;
assign n_16245 = n_16096 ^ x23;
assign n_16246 = n_16097 ^ x26;
assign n_16247 = n_16098 ^ x29;
assign n_16248 = n_16099 ^ x32;
assign n_16249 = n_16100 ^ x35;
assign n_16250 = n_16101 ^ x38;
assign n_16251 = n_16102 ^ x41;
assign n_16252 = n_16103 ^ x44;
assign n_16253 = n_16104 ^ x47;
assign n_16254 = n_16105 ^ x50;
assign n_16255 = n_16106 ^ x53;
assign n_16256 = n_16107 ^ x56;
assign n_16257 = n_16108 ^ x59;
assign n_16258 = n_16109 ^ x62;
assign n_16259 = n_16110 ^ x1;
assign n_16260 = n_1 & ~n_16111;
assign n_16261 = n_16111 ^ x126;
assign n_16262 = n_16112 ^ n_15992;
assign n_16263 = ~n_16112 & n_303;
assign n_16264 = n_2180 ^ n_16113;
assign n_16265 = n_780 ^ n_16114;
assign n_16266 = n_2251 ^ n_16115;
assign n_16267 = n_2319 ^ n_16116;
assign n_16268 = n_2386 ^ n_16117;
assign n_16269 = n_2453 ^ n_16118;
assign n_16270 = n_2520 ^ n_16119;
assign n_16271 = n_2586 ^ n_16120;
assign n_16272 = n_2651 ^ n_16121;
assign n_16273 = n_2718 ^ n_16122;
assign n_16274 = n_2786 ^ n_16123;
assign n_16275 = n_2853 ^ n_16124;
assign n_16276 = n_2921 ^ n_16125;
assign n_16277 = n_2987 ^ n_16126;
assign n_16278 = n_3056 ^ n_16127;
assign n_16279 = n_3122 ^ n_16128;
assign n_16280 = n_3191 ^ n_16129;
assign n_16281 = n_3255 ^ n_16130;
assign n_16282 = n_3320 ^ n_16131;
assign n_16283 = n_3385 ^ n_16132;
assign n_16284 = n_16134 ^ n_10855;
assign n_16285 = ~n_14894 & n_16135;
assign n_16286 = n_16137 ^ n_15867;
assign n_16287 = n_16139 ^ n_15868;
assign n_16288 = n_16141 ^ n_15869;
assign n_16289 = n_16143 ^ n_15870;
assign n_16290 = n_16145 ^ n_15871;
assign n_16291 = n_16147 ^ n_15872;
assign n_16292 = n_16148 ^ n_15354;
assign n_16293 = n_16148 ^ n_15184;
assign n_16294 = n_16150 ^ n_15875;
assign n_16295 = n_16152 ^ n_15876;
assign n_16296 = n_16153 ^ n_10854;
assign n_16297 = ~n_15016 & n_16154;
assign y29 = ~n_16155;
assign n_16298 = n_14892 & ~n_16156;
assign n_16299 = n_16158 ^ n_15880;
assign n_16300 = n_16160 ^ n_15881;
assign n_16301 = n_16162 ^ n_15882;
assign n_16302 = n_16164 ^ n_15883;
assign n_16303 = n_16165 ^ n_15356;
assign n_16304 = n_16165 ^ n_15186;
assign n_16305 = n_16166 ^ n_16064;
assign n_16306 = n_16166 ^ n_16025;
assign n_16307 = n_16167 ^ n_15272;
assign n_16308 = n_16168 ^ n_15558;
assign n_16309 = n_16046 & n_16169;
assign n_16310 = n_16170 ^ n_15910;
assign n_16311 = n_16171 ^ n_15912;
assign n_16312 = n_16173 ^ n_15913;
assign n_16313 = n_16175 ^ n_15914;
assign n_16314 = n_16177 ^ n_15915;
assign n_16315 = n_16179 ^ n_15916;
assign n_16316 = n_16181 ^ n_15917;
assign n_16317 = n_16183 ^ n_15918;
assign n_16318 = n_16184 ^ n_15919;
assign n_16319 = n_16185 ^ n_15654;
assign n_16320 = n_16187 ^ n_15922;
assign n_16321 = n_16189 ^ n_15924;
assign n_16322 = n_16191 ^ n_15255;
assign n_16323 = n_15255 & n_16191;
assign n_16324 = n_15900 & ~n_16194;
assign n_16325 = ~n_15901 & n_16196;
assign n_16326 = n_15902 & n_16198;
assign n_16327 = ~n_15903 & n_16200;
assign n_16328 = ~n_15904 & n_16202;
assign n_16329 = ~n_15905 & n_16204;
assign n_16330 = n_15906 & n_16206;
assign n_16331 = ~n_15907 & ~n_16208;
assign n_16332 = n_16209 ^ n_15787;
assign n_16333 = ~n_16209 & n_15908;
assign n_16334 = ~n_15909 & n_16211;
assign n_16335 = n_16212 ^ n_15627;
assign n_16336 = n_16212 & n_16213;
assign n_16337 = n_6647 & n_16216;
assign n_16338 = n_16217 ^ n_15947;
assign n_16339 = ~x0 & n_16218;
assign n_16340 = n_16219 ^ x5;
assign n_16341 = n_16220 ^ x8;
assign n_16342 = n_16221 ^ x11;
assign n_16343 = n_16222 ^ x14;
assign n_16344 = n_16223 ^ x17;
assign n_16345 = n_16224 ^ x20;
assign n_16346 = n_16225 ^ x23;
assign n_16347 = n_16226 ^ x26;
assign n_16348 = n_16227 ^ x29;
assign n_16349 = n_16228 ^ x32;
assign n_16350 = n_16229 ^ x35;
assign n_16351 = n_16230 ^ x38;
assign n_16352 = n_16231 ^ x41;
assign n_16353 = n_16232 ^ x44;
assign n_16354 = n_16233 ^ x47;
assign n_16355 = n_16234 ^ x50;
assign n_16356 = n_16235 ^ x53;
assign n_16357 = n_16236 ^ x56;
assign n_16358 = n_16237 ^ x59;
assign n_16359 = n_16238 ^ x62;
assign n_16360 = n_16239 ^ n_15542;
assign n_16361 = n_16240 ^ n_15543;
assign n_16362 = n_16245 ^ n_15892;
assign n_16363 = n_16245 ^ n_15769;
assign n_16364 = n_16246 ^ n_15893;
assign n_16365 = n_16246 ^ n_15770;
assign n_16366 = n_16247 ^ n_15894;
assign n_16367 = n_16247 ^ n_15771;
assign n_16368 = n_16248 ^ n_15895;
assign n_16369 = n_16248 ^ n_15772;
assign n_16370 = n_16249 ^ n_15896;
assign n_16371 = n_16249 ^ n_15773;
assign n_16372 = n_16250 ^ n_15897;
assign n_16373 = n_16250 ^ n_15774;
assign n_16374 = n_16251 ^ n_15898;
assign n_16375 = n_16251 ^ n_15775;
assign n_16376 = n_16252 ^ n_15899;
assign n_16377 = n_16252 ^ n_15776;
assign n_16378 = n_15921 ^ n_16253;
assign n_16379 = n_15801 ^ n_16253;
assign n_16380 = n_16254 ^ n_15803;
assign n_16381 = n_16256 ^ n_15684;
assign n_16382 = n_16257 ^ n_15560;
assign n_16383 = n_16258 ^ ~n_6729;
assign n_16384 = ~n_6729 & n_16258;
assign n_16385 = n_16259 ^ x125;
assign n_16386 = n_16260 ^ x1;
assign n_16387 = n_655 & n_16261;
assign n_16388 = n_784 & n_16261;
assign n_16389 = ~n_3665 & n_16261;
assign n_16390 = n_854 & n_16261;
assign n_16391 = n_920 & n_16261;
assign n_16392 = n_986 & n_16261;
assign n_16393 = n_1052 & n_16261;
assign n_16394 = n_1117 & n_16261;
assign n_16395 = n_1181 & n_16261;
assign n_16396 = n_1248 & n_16261;
assign n_16397 = n_1314 & n_16261;
assign n_16398 = n_1380 & n_16261;
assign n_16399 = n_1445 & n_16261;
assign n_16400 = n_1510 & n_16261;
assign n_16401 = n_1576 & n_16261;
assign n_16402 = n_1641 & n_16261;
assign n_16403 = n_1706 & n_16261;
assign n_16404 = n_1771 & n_16261;
assign n_16405 = n_1835 & n_16261;
assign n_16406 = n_1899 & n_16261;
assign n_16407 = n_1 & ~n_16262;
assign n_16408 = n_16262 ^ x127;
assign n_16409 = n_16263 ^ n_16133;
assign n_16410 = n_16263 ^ x2;
assign n_16411 = n_16263 ^ x127;
assign n_16412 = ~n_16263 & ~n_624;
assign n_16413 = ~n_16263 & ~n_625;
assign n_16414 = ~n_16263 & ~n_626;
assign n_16415 = n_5053 ^ n_16264;
assign n_16416 = n_5116 ^ n_16265;
assign n_16417 = n_5179 ^ n_16266;
assign n_16418 = n_5240 ^ n_16267;
assign n_16419 = n_5304 ^ n_16268;
assign n_16420 = n_5368 ^ n_16269;
assign n_16421 = n_5432 ^ n_16270;
assign n_16422 = n_5496 ^ n_16271;
assign n_16423 = n_5557 ^ n_16272;
assign n_16424 = n_5620 ^ n_16273;
assign n_16425 = n_5683 ^ n_16274;
assign n_16426 = n_5747 ^ n_16275;
assign n_16427 = n_5813 ^ n_16276;
assign n_16428 = n_5875 ^ n_16277;
assign n_16429 = n_5939 ^ n_16278;
assign n_16430 = n_6002 ^ n_16279;
assign n_16431 = n_6066 ^ n_16280;
assign n_16432 = n_6130 ^ n_16281;
assign n_16433 = n_6192 ^ n_16282;
assign n_16434 = n_6254 ^ n_16283;
assign n_16435 = n_16285 ^ n_15993;
assign n_16436 = n_16286 ^ n_15343;
assign n_16437 = n_16286 ^ n_15172;
assign n_16438 = n_16287 ^ n_15345;
assign n_16439 = n_16287 ^ n_15174;
assign n_16440 = n_16288 ^ n_14896;
assign n_16441 = n_16288 ^ n_14728;
assign n_16442 = n_16289 ^ n_15349;
assign n_16443 = n_16289 ^ n_15178;
assign n_16444 = n_16290 ^ n_15351;
assign n_16445 = n_16290 ^ n_15180;
assign n_16446 = n_16291 ^ n_15182;
assign n_16447 = n_16291 ^ n_15024;
assign n_16448 = n_16292 ^ n_12807;
assign n_16449 = ~n_15354 & n_16293;
assign n_16450 = n_16294 ^ n_15198;
assign n_16451 = n_16294 ^ n_15035;
assign n_16452 = n_16295 ^ n_15663;
assign n_16453 = n_16295 ^ n_15080;
assign n_16454 = n_16297 ^ n_16012;
assign n_16455 = n_16298 ^ n_16013;
assign n_16456 = n_16299 ^ n_15489;
assign n_16457 = n_16299 ^ n_15358;
assign n_16458 = n_16300 ^ n_15734;
assign n_16459 = n_16300 ^ n_15594;
assign n_16460 = n_16301 ^ n_15368;
assign n_16461 = n_16301 ^ n_15196;
assign n_16462 = n_16302 ^ n_15740;
assign n_16463 = n_16302 ^ n_15600;
assign n_16464 = n_16303 ^ n_14953;
assign n_16465 = ~n_15356 & n_16304;
assign n_16466 = n_16305 ^ n_16025;
assign n_16467 = n_16305 & ~n_16306;
assign n_16468 = n_16308 ^ n_15249;
assign n_16469 = n_16308 & n_15683;
assign n_16470 = n_16309 ^ n_15925;
assign n_16471 = n_16310 ^ n_16214;
assign n_16472 = n_16310 ^ n_15538;
assign n_16473 = n_16312 ^ n_16195;
assign n_16474 = n_16313 ^ n_16197;
assign n_16475 = n_16314 ^ n_16199;
assign n_16476 = n_16315 ^ n_16201;
assign n_16477 = n_16316 ^ n_16203;
assign n_16478 = n_16317 ^ n_16205;
assign n_16479 = n_16318 ^ n_16207;
assign n_16480 = n_16320 ^ n_16210;
assign n_16481 = n_16323 ^ n_16322;
assign n_16482 = n_16324 ^ n_15779;
assign n_16483 = n_16325 ^ n_16055;
assign n_16484 = n_16326 ^ n_16056;
assign n_16485 = n_16327 ^ n_16057;
assign n_16486 = n_16328 ^ n_16058;
assign n_16487 = n_16329 ^ n_16059;
assign n_16488 = n_16330 ^ n_16060;
assign n_16489 = n_16331 ^ n_16061;
assign n_16490 = n_16319 ^ n_16332;
assign n_16491 = n_16333 ^ n_16062;
assign n_16492 = n_16334 ^ n_15788;
assign n_16493 = n_16336 ^ n_15789;
assign n_16494 = n_16337 ^ n_16067;
assign n_16495 = n_16338 ^ n_15541;
assign n_16496 = n_16339 ^ n_16069;
assign n_16497 = n_16340 ^ n_15688;
assign n_16498 = n_16172 ^ n_16346;
assign n_16499 = n_16174 ^ n_16347;
assign n_16500 = n_16176 ^ n_16348;
assign n_16501 = n_16178 ^ n_16349;
assign n_16502 = n_16180 ^ n_16350;
assign n_16503 = n_16182 ^ n_16351;
assign n_16504 = n_16040 ^ n_16352;
assign n_16505 = n_16042 ^ n_16353;
assign n_16506 = n_16186 ^ n_16354;
assign n_16507 = n_16188 ^ n_16355;
assign n_16508 = n_16190 ^ n_16357;
assign n_16509 = n_16358 ^ n_16032;
assign n_16510 = n_16359 ^ n_6496;
assign n_16511 = n_15892 & n_16363;
assign n_16512 = ~n_15893 & n_16365;
assign n_16513 = n_15894 & n_16367;
assign n_16514 = ~n_15895 & n_16369;
assign n_16515 = n_15896 & n_16371;
assign n_16516 = n_15897 & n_16373;
assign n_16517 = n_15898 & n_16375;
assign n_16518 = ~n_15899 & n_16377;
assign n_16519 = ~n_15921 & n_16379;
assign n_16520 = n_16380 ^ n_15778;
assign n_16521 = ~n_16380 & n_15923;
assign n_16522 = n_16381 ^ n_15891;
assign n_16523 = ~n_16381 & n_16029;
assign n_16524 = n_16382 ^ n_15791;
assign n_16525 = n_16382 & ~n_15911;
assign n_16526 = n_16384 ^ n_6500;
assign n_16527 = n_16385 ^ n_2120;
assign n_16528 = n_16386 ^ x126;
assign n_16529 = n_2181 ^ n_16387;
assign n_16530 = n_781 ^ n_16388;
assign n_16531 = n_2252 ^ n_16389;
assign n_16532 = n_2320 ^ n_16390;
assign n_16533 = n_2387 ^ n_16391;
assign n_16534 = n_2454 ^ n_16392;
assign n_16535 = n_2521 ^ n_16393;
assign n_16536 = n_2587 ^ n_16394;
assign n_16537 = n_2652 ^ n_16395;
assign n_16538 = n_2719 ^ n_16396;
assign n_16539 = n_2787 ^ n_16397;
assign n_16540 = n_2854 ^ n_16398;
assign n_16541 = n_2922 ^ n_16399;
assign n_16542 = n_2988 ^ n_16400;
assign n_16543 = n_3057 ^ n_16401;
assign n_16544 = n_3123 ^ n_16402;
assign n_16545 = n_3192 ^ n_16403;
assign n_16546 = n_3256 ^ n_16404;
assign n_16547 = n_3321 ^ n_16405;
assign n_16548 = n_3386 ^ n_16406;
assign n_16549 = n_16407 ^ x1;
assign n_16550 = n_655 & n_16408;
assign n_16551 = n_784 & n_16408;
assign n_16552 = ~n_3665 & n_16408;
assign n_16553 = n_854 & n_16408;
assign n_16554 = n_920 & n_16408;
assign n_16555 = n_986 & n_16408;
assign n_16556 = n_1052 & n_16408;
assign n_16557 = n_1117 & n_16408;
assign n_16558 = n_1181 & n_16408;
assign n_16559 = n_1248 & n_16408;
assign n_16560 = n_1314 & n_16408;
assign n_16561 = n_1380 & n_16408;
assign n_16562 = n_1445 & n_16408;
assign n_16563 = n_1510 & n_16408;
assign n_16564 = n_1576 & n_16408;
assign n_16565 = n_1641 & n_16408;
assign n_16566 = n_1706 & n_16408;
assign n_16567 = n_1771 & n_16408;
assign n_16568 = n_1835 & n_16408;
assign n_16569 = n_1899 & n_16408;
assign n_16570 = n_1 & ~n_16409;
assign n_16571 = n_655 & n_16409;
assign n_16572 = n_784 & n_16409;
assign n_16573 = ~n_3665 & n_16409;
assign n_16574 = n_854 & n_16409;
assign n_16575 = n_920 & n_16409;
assign n_16576 = n_986 & n_16409;
assign n_16577 = n_1052 & n_16409;
assign n_16578 = n_1117 & n_16409;
assign n_16579 = n_1181 & n_16409;
assign n_16580 = n_1248 & n_16409;
assign n_16581 = n_1314 & n_16409;
assign n_16582 = n_1380 & n_16409;
assign n_16583 = n_1445 & n_16409;
assign n_16584 = n_1510 & n_16409;
assign n_16585 = n_1576 & n_16409;
assign n_16586 = n_1641 & n_16409;
assign n_16587 = n_1706 & n_16409;
assign n_16588 = n_1771 & n_16409;
assign n_16589 = n_1835 & n_16409;
assign n_16590 = n_1899 & n_16409;
assign n_16591 = x0 & ~n_16410;
assign n_16592 = n_3 & n_16411;
assign n_16593 = n_15 & n_16411;
assign n_16594 = n_18 & n_16411;
assign n_16595 = n_21 & n_16411;
assign n_16596 = n_24 & n_16411;
assign n_16597 = n_1117 & n_16411;
assign n_16598 = n_30 & n_16411;
assign n_16599 = n_36 & n_16411;
assign n_16600 = n_39 & n_16411;
assign n_16601 = n_1445 & n_16411;
assign n_16602 = n_45 & n_16411;
assign n_16603 = n_48 & n_16411;
assign n_16604 = n_51 & n_16411;
assign n_16605 = n_54 & n_16411;
assign n_16606 = n_1771 & n_16411;
assign n_16607 = n_1835 & n_16411;
assign n_16608 = n_1899 & n_16411;
assign n_16609 = n_16412 ^ x8;
assign n_16610 = n_16413 ^ x11;
assign n_16611 = n_16414 ^ x32;
assign n_16612 = n_16415 ^ x5;
assign n_16613 = n_16416 ^ x8;
assign n_16614 = n_16417 ^ x11;
assign n_16615 = n_16418 ^ x14;
assign n_16616 = n_16419 ^ x17;
assign n_16617 = n_16420 ^ x20;
assign n_16618 = n_16421 ^ x23;
assign n_16619 = n_16422 ^ x26;
assign n_16620 = n_16423 ^ x29;
assign n_16621 = n_16424 ^ x32;
assign n_16622 = n_16425 ^ x35;
assign n_16623 = n_16426 ^ x38;
assign n_16624 = n_16427 ^ x41;
assign n_16625 = n_16428 ^ x44;
assign n_16626 = n_16429 ^ x47;
assign n_16627 = n_16430 ^ x50;
assign n_16628 = n_16431 ^ x53;
assign n_16629 = n_16432 ^ x56;
assign n_16630 = n_16433 ^ x59;
assign n_16631 = n_16434 ^ x62;
assign n_16632 = n_16435 ^ n_15364;
assign n_16633 = n_16435 ^ n_15192;
assign n_16634 = n_16436 ^ n_10857;
assign n_16635 = ~n_15343 & n_16437;
assign n_16636 = n_16438 ^ n_10858;
assign n_16637 = n_15345 & ~n_16439;
assign n_16638 = n_16440 ^ n_10859;
assign n_16639 = ~n_14896 & n_16441;
assign n_16640 = n_16442 ^ n_10862;
assign n_16641 = ~n_15349 & n_16443;
assign n_16642 = n_16444 ^ n_10863;
assign n_16643 = ~n_15351 & n_16445;
assign n_16644 = n_16446 ^ n_10864;
assign n_16645 = ~n_15182 & n_16447;
assign n_16646 = n_16449 ^ n_16148;
assign n_16647 = n_16450 ^ n_14031;
assign n_16648 = n_15198 & ~n_16451;
assign n_16649 = n_16452 ^ n_16244;
assign n_16650 = ~n_15663 & n_16453;
assign n_16651 = n_16454 ^ n_15477;
assign n_16652 = n_16454 ^ n_15339;
assign n_16653 = n_16455 ^ n_15362;
assign n_16654 = n_16455 ^ n_15190;
assign n_16655 = n_16456 ^ n_11220;
assign n_16656 = ~n_15489 & n_16457;
assign n_16657 = n_16458 ^ n_11127;
assign n_16658 = n_15734 & ~n_16459;
assign n_16659 = n_16460 ^ n_11131;
assign n_16660 = ~n_15368 & n_16461;
assign n_16661 = n_16462 ^ n_11132;
assign n_16662 = n_15740 & ~n_16463;
assign n_16663 = n_16465 ^ n_16165;
assign n_16664 = n_16466 ^ n_16321;
assign n_16665 = n_16467 ^ n_16064;
assign n_16666 = n_16468 ^ n_16255;
assign n_16667 = n_16468 ^ n_16307;
assign n_16668 = n_16469 ^ n_16168;
assign n_16669 = n_16470 ^ n_16471;
assign n_16670 = n_16214 & ~n_16472;
assign n_16671 = n_16482 ^ n_16362;
assign n_16672 = n_16483 ^ n_16364;
assign n_16673 = n_16484 ^ n_16366;
assign n_16674 = n_16485 ^ n_16368;
assign n_16675 = n_16486 ^ n_16370;
assign n_16676 = n_16487 ^ n_16372;
assign n_16677 = n_16488 ^ n_16374;
assign n_16678 = n_16489 ^ n_16376;
assign n_16679 = n_16491 ^ n_16378;
assign n_16680 = n_16494 ^ n_16383;
assign n_16681 = n_16496 ^ n_15687;
assign n_16682 = ~n_15687 & ~n_16496;
assign n_16683 = n_16511 ^ n_16245;
assign n_16684 = n_16512 ^ n_16246;
assign n_16685 = n_16513 ^ n_16247;
assign n_16686 = n_16514 ^ n_16248;
assign n_16687 = n_16515 ^ n_16249;
assign n_16688 = n_16516 ^ n_16250;
assign n_16689 = n_16517 ^ n_16251;
assign n_16690 = n_16518 ^ n_16252;
assign n_16691 = n_16519 ^ n_15777;
assign n_16692 = n_16520 ^ n_16492;
assign n_16693 = n_16521 ^ n_16254;
assign n_16694 = n_16493 ^ n_16522;
assign n_16695 = n_16523 ^ n_16256;
assign n_16696 = n_16525 ^ n_16257;
assign n_16697 = n_16526 ^ n_16510;
assign n_16698 = n_16526 ^ n_16359;
assign n_16699 = ~x0 & n_16527;
assign n_16700 = n_16528 ^ n_6501;
assign n_16701 = n_5054 ^ n_16529;
assign n_16702 = n_5117 ^ n_16530;
assign n_16703 = n_5180 ^ n_16531;
assign n_16704 = n_5241 ^ n_16532;
assign n_16705 = n_5305 ^ n_16533;
assign n_16706 = n_5369 ^ n_16534;
assign n_16707 = n_5433 ^ n_16535;
assign n_16708 = n_5497 ^ n_16536;
assign n_16709 = n_5558 ^ n_16537;
assign n_16710 = n_5621 ^ n_16538;
assign n_16711 = n_5684 ^ n_16539;
assign n_16712 = n_5748 ^ n_16540;
assign n_16713 = n_5814 ^ n_16541;
assign n_16714 = n_5876 ^ n_16542;
assign n_16715 = n_5940 ^ n_16543;
assign n_16716 = n_6003 ^ n_16544;
assign n_16717 = n_6067 ^ n_16545;
assign n_16718 = n_6131 ^ n_16546;
assign n_16719 = n_6193 ^ n_16547;
assign n_16720 = n_6255 ^ n_16548;
assign n_16721 = n_16549 ^ x127;
assign n_16722 = n_2182 ^ n_16550;
assign n_16723 = n_782 ^ n_16551;
assign n_16724 = n_2253 ^ n_16552;
assign n_16725 = n_2321 ^ n_16553;
assign n_16726 = n_2388 ^ n_16554;
assign n_16727 = n_2455 ^ n_16555;
assign n_16728 = n_2522 ^ n_16556;
assign n_16729 = n_2588 ^ n_16557;
assign n_16730 = n_2653 ^ n_16558;
assign n_16731 = n_2720 ^ n_16559;
assign n_16732 = n_2788 ^ n_16560;
assign n_16733 = n_2855 ^ n_16561;
assign n_16734 = n_2923 ^ n_16562;
assign n_16735 = n_2989 ^ n_16563;
assign n_16736 = n_3058 ^ n_16564;
assign n_16737 = n_3124 ^ n_16565;
assign n_16738 = n_3193 ^ n_16566;
assign n_16739 = n_3257 ^ n_16567;
assign n_16740 = n_3322 ^ n_16568;
assign n_16741 = n_3387 ^ n_16569;
assign n_16742 = n_16570 ^ x1;
assign n_16743 = n_3597 ^ n_16571;
assign n_16744 = n_3661 ^ n_16572;
assign n_16745 = n_3788 ^ n_16573;
assign n_16746 = n_3851 ^ n_16574;
assign n_16747 = n_3916 ^ n_16575;
assign n_16748 = n_3981 ^ n_16576;
assign n_16749 = n_4046 ^ n_16577;
assign n_16750 = n_4111 ^ n_16578;
assign n_16751 = n_4174 ^ n_16579;
assign n_16752 = n_4238 ^ n_16580;
assign n_16753 = n_4304 ^ n_16581;
assign n_16754 = n_4369 ^ n_16582;
assign n_16755 = n_4436 ^ n_16583;
assign n_16756 = n_4500 ^ n_16584;
assign n_16757 = n_4565 ^ n_16585;
assign n_16758 = n_4629 ^ n_16586;
assign n_16759 = n_4694 ^ n_16587;
assign n_16760 = n_4759 ^ n_16588;
assign n_16761 = n_4823 ^ n_16589;
assign n_16762 = n_4887 ^ n_16590;
assign n_16763 = n_16591 ^ x2;
assign n_16764 = n_16592 ^ n_2185;
assign n_16765 = n_16593 ^ n_2324;
assign n_16766 = n_16594 ^ n_2391;
assign n_16767 = n_16595 ^ n_2458;
assign n_16768 = n_16596 ^ n_2525;
assign n_16769 = n_16597 ^ n_4112;
assign n_16770 = n_16598 ^ n_2656;
assign n_16771 = n_16599 ^ n_2791;
assign n_16772 = n_16600 ^ n_2858;
assign n_16773 = n_4437 ^ n_16601;
assign n_16774 = n_16602 ^ n_2992;
assign n_16775 = n_16603 ^ n_2996;
assign n_16776 = n_16604 ^ n_3127;
assign n_16777 = n_16605 ^ n_3131;
assign n_16778 = n_16606 ^ n_4760;
assign n_16779 = n_16607 ^ n_4824;
assign n_16780 = n_16608 ^ n_4888;
assign n_16781 = n_342 & ~n_16609;
assign n_16782 = n_351 & ~n_16610;
assign n_16783 = n_392 & ~n_16611;
assign n_16784 = n_16612 ^ n_16049;
assign n_16785 = n_16193 ^ n_16617;
assign n_16786 = n_16473 ^ n_16618;
assign n_16787 = n_16195 ^ n_16618;
assign n_16788 = n_16474 ^ n_16619;
assign n_16789 = n_16197 ^ n_16619;
assign n_16790 = n_16475 ^ n_16620;
assign n_16791 = n_16199 ^ n_16620;
assign n_16792 = n_16476 ^ n_16621;
assign n_16793 = n_16201 ^ n_16621;
assign n_16794 = n_16477 ^ n_16622;
assign n_16795 = n_16316 ^ n_16622;
assign n_16796 = n_16478 ^ n_16623;
assign n_16797 = n_16205 ^ n_16623;
assign n_16798 = n_16479 ^ n_16624;
assign n_16799 = n_16318 ^ n_16624;
assign n_16800 = n_16625 ^ n_16332;
assign n_16801 = n_16320 ^ n_16626;
assign n_16802 = n_16466 ^ n_16627;
assign n_16803 = n_16470 ^ n_16629;
assign n_16804 = n_16311 ^ n_16630;
assign n_16805 = n_16630 ^ n_16215;
assign n_16806 = n_16631 ^ n_6728;
assign n_16807 = n_16632 ^ n_11126;
assign n_16808 = ~n_15364 & n_16633;
assign n_16809 = n_16635 ^ n_16286;
assign n_16810 = n_16637 ^ n_16287;
assign n_16811 = n_16639 ^ n_16288;
assign n_16812 = n_16641 ^ n_16289;
assign n_16813 = n_16643 ^ n_16290;
assign n_16814 = n_16645 ^ n_16291;
assign n_16815 = n_16646 ^ n_15747;
assign n_16816 = n_16646 ^ n_15608;
assign n_16817 = n_16648 ^ n_16294;
assign n_16818 = n_16650 ^ n_16295;
assign n_16819 = n_16651 ^ n_11125;
assign n_16820 = ~n_15477 & n_16652;
assign y30 = n_16653;
assign n_16821 = ~n_15362 & n_16654;
assign n_16822 = n_16656 ^ n_16299;
assign n_16823 = n_16658 ^ n_16300;
assign n_16824 = n_16660 ^ n_16301;
assign n_16825 = n_16662 ^ n_16302;
assign n_16826 = n_16663 ^ n_15749;
assign n_16827 = n_16663 ^ n_15610;
assign n_16828 = n_16666 ^ n_16307;
assign n_16829 = ~n_16666 & n_16667;
assign n_16830 = n_16668 ^ n_15817;
assign n_16831 = n_16668 ^ n_15704;
assign n_16832 = n_16670 ^ n_16066;
assign n_16833 = n_16682 ^ n_16681;
assign n_16834 = n_16498 ^ n_16683;
assign n_16835 = n_16346 ^ n_16683;
assign n_16836 = n_16499 ^ n_16684;
assign n_16837 = n_16347 ^ n_16684;
assign n_16838 = n_16500 ^ n_16685;
assign n_16839 = n_16348 ^ n_16685;
assign n_16840 = n_16501 ^ n_16686;
assign n_16841 = n_16349 ^ n_16686;
assign n_16842 = n_16502 ^ n_16687;
assign n_16843 = n_16350 ^ n_16687;
assign n_16844 = n_16503 ^ n_16688;
assign n_16845 = n_16351 ^ n_16688;
assign n_16846 = n_16689 ^ n_16504;
assign n_16847 = n_16689 ^ n_16352;
assign n_16848 = n_16690 ^ n_16042;
assign n_16849 = n_16506 ^ n_16691;
assign n_16850 = n_16354 ^ n_16691;
assign n_16851 = n_16507 ^ n_16693;
assign n_16852 = n_16355 ^ n_16693;
assign n_16853 = n_16508 ^ n_16695;
assign n_16854 = n_16357 ^ n_16695;
assign n_16855 = n_16696 ^ n_16358;
assign n_16856 = n_16510 & n_16698;
assign n_16857 = n_16699 ^ n_16385;
assign n_16858 = ~x0 & ~n_16700;
assign n_16859 = n_16701 ^ x5;
assign n_16860 = n_16702 ^ x8;
assign n_16861 = n_16703 ^ x11;
assign n_16862 = n_16704 ^ x14;
assign n_16863 = n_16705 ^ x17;
assign n_16864 = n_16706 ^ x20;
assign n_16865 = n_16707 ^ x23;
assign n_16866 = n_16708 ^ x26;
assign n_16867 = n_16709 ^ x29;
assign n_16868 = n_16710 ^ x32;
assign n_16869 = n_16711 ^ x35;
assign n_16870 = n_16712 ^ x38;
assign n_16871 = n_16713 ^ x41;
assign n_16872 = n_16714 ^ x44;
assign n_16873 = n_16715 ^ x47;
assign n_16874 = n_16716 ^ x50;
assign n_16875 = n_16717 ^ x53;
assign n_16876 = n_16718 ^ x56;
assign n_16877 = n_16719 ^ x59;
assign n_16878 = n_16720 ^ x62;
assign n_16879 = n_16721 ^ n_3531;
assign n_16880 = n_5055 ^ n_16722;
assign n_16881 = n_5118 ^ n_16723;
assign n_16882 = n_5181 ^ n_16724;
assign n_16883 = n_5242 ^ n_16725;
assign n_16884 = n_5306 ^ n_16726;
assign n_16885 = n_5370 ^ n_16727;
assign n_16886 = n_5434 ^ n_16728;
assign n_16887 = n_5498 ^ n_16729;
assign n_16888 = n_5559 ^ n_16730;
assign n_16889 = n_5622 ^ n_16731;
assign n_16890 = n_5685 ^ n_16732;
assign n_16891 = n_5749 ^ n_16733;
assign n_16892 = n_5815 ^ n_16734;
assign n_16893 = n_5877 ^ n_16735;
assign n_16894 = n_5941 ^ n_16736;
assign n_16895 = n_6004 ^ n_16737;
assign n_16896 = n_6068 ^ n_16738;
assign n_16897 = n_6132 ^ n_16739;
assign n_16898 = n_6194 ^ n_16740;
assign n_16899 = n_6256 ^ n_16741;
assign n_16900 = n_16742 ^ n_3533;
assign n_16901 = n_2183 ^ n_16743;
assign n_16902 = n_783 ^ n_16744;
assign n_16903 = n_2254 ^ n_16745;
assign n_16904 = n_2322 ^ n_16746;
assign n_16905 = n_2389 ^ n_16747;
assign n_16906 = n_2456 ^ n_16748;
assign n_16907 = n_2523 ^ n_16749;
assign n_16908 = n_2589 ^ n_16750;
assign n_16909 = n_2654 ^ n_16751;
assign n_16910 = n_2721 ^ n_16752;
assign n_16911 = n_2789 ^ n_16753;
assign n_16912 = n_2856 ^ n_16754;
assign n_16913 = n_2924 ^ n_16755;
assign n_16914 = n_2990 ^ n_16756;
assign n_16915 = n_3059 ^ n_16757;
assign n_16916 = n_3125 ^ n_16758;
assign n_16917 = n_3194 ^ n_16759;
assign n_16918 = n_3258 ^ n_16760;
assign n_16919 = n_3323 ^ n_16761;
assign n_16920 = n_3388 ^ n_16762;
assign n_16921 = n_16763 ^ n_1;
assign n_16922 = ~n_5056 & ~n_16764;
assign n_16923 = ~n_5243 & ~n_16765;
assign n_16924 = ~n_5307 & ~n_16766;
assign n_16925 = ~n_5371 & ~n_16767;
assign n_16926 = ~n_5435 & ~n_16768;
assign n_16927 = n_16769 ^ x26;
assign n_16928 = ~n_5560 & ~n_16770;
assign n_16929 = ~n_5686 & ~n_16771;
assign n_16930 = ~n_5750 & ~n_16772;
assign n_16931 = n_16773 ^ x41;
assign n_16932 = ~n_5878 & ~n_16774;
assign n_16933 = ~n_5942 & ~n_16775;
assign n_16934 = ~n_6005 & ~n_16776;
assign n_16935 = ~n_6069 & ~n_16777;
assign n_16936 = n_16778 ^ x56;
assign n_16937 = n_16779 ^ x59;
assign n_16938 = n_16780 ^ n_3530;
assign n_16939 = n_16780 ^ x125;
assign n_16940 = n_16780 ^ x126;
assign n_16941 = n_3663 & ~n_16781;
assign n_16942 = n_3789 & ~n_16782;
assign n_16943 = n_4240 & ~n_16783;
assign n_16944 = ~n_16473 & n_16787;
assign n_16945 = n_16474 & ~n_16789;
assign n_16946 = ~n_16475 & n_16791;
assign n_16947 = ~n_16476 & n_16793;
assign n_16948 = ~n_16477 & n_16795;
assign n_16949 = n_16478 & ~n_16797;
assign n_16950 = ~n_16479 & n_16799;
assign n_16951 = n_16319 ^ n_16800;
assign n_16952 = ~n_16800 & n_16490;
assign n_16953 = n_16801 ^ n_16210;
assign n_16954 = n_16801 & n_16480;
assign n_16955 = n_16802 ^ n_16321;
assign n_16956 = n_16802 & ~n_16664;
assign n_16957 = n_16803 ^ n_16471;
assign n_16958 = n_16803 & ~n_16669;
assign n_16959 = n_16804 ^ n_16215;
assign n_16960 = ~n_16804 & n_16805;
assign n_16961 = n_16806 ^ n_3420;
assign n_16962 = ~n_16806 & ~n_6850;
assign n_16963 = n_16808 ^ n_16435;
assign n_16964 = n_16809 ^ n_15736;
assign n_16965 = n_16809 ^ n_15596;
assign n_16966 = n_16810 ^ n_15738;
assign n_16967 = n_16810 ^ n_15598;
assign n_16968 = n_16811 ^ n_15366;
assign n_16969 = n_16811 ^ n_15194;
assign n_16970 = n_16812 ^ n_15742;
assign n_16971 = n_16812 ^ n_15602;
assign n_16972 = n_16813 ^ n_15744;
assign n_16973 = n_16813 ^ n_15604;
assign n_16974 = n_16814 ^ n_15606;
assign n_16975 = n_16814 ^ n_15485;
assign n_16976 = n_16815 ^ n_12965;
assign n_16977 = n_15747 & ~n_16816;
assign n_16978 = n_16817 ^ n_15622;
assign n_16979 = n_16817 ^ n_15496;
assign n_16980 = n_16818 ^ n_15807;
assign n_16981 = n_16818 ^ n_15561;
assign n_16982 = n_16820 ^ n_16454;
assign n_16983 = n_16821 ^ n_16455;
assign n_16984 = n_16822 ^ n_15877;
assign n_16985 = n_16822 ^ n_15751;
assign n_16986 = n_16823 ^ n_16136;
assign n_16987 = n_16823 ^ n_15994;
assign n_16988 = n_16824 ^ n_15761;
assign n_16989 = n_16824 ^ n_15620;
assign n_16990 = n_16825 ^ n_16142;
assign n_16991 = n_16825 ^ n_10786;
assign n_16992 = n_16826 ^ n_15302;
assign n_16993 = ~n_15749 & n_16827;
assign n_16994 = n_16828 ^ n_16665;
assign n_16995 = n_16829 ^ n_16255;
assign n_16996 = n_16830 ^ n_16356;
assign n_16997 = ~n_15817 & ~n_16831;
assign n_16998 = n_16832 ^ n_16524;
assign n_16999 = n_16498 & n_16835;
assign n_17000 = n_16499 & n_16837;
assign n_17001 = n_16500 & n_16839;
assign n_17002 = n_16501 & n_16841;
assign n_17003 = ~n_16502 & n_16843;
assign n_17004 = ~n_16503 & n_16845;
assign n_17005 = n_16504 & n_16847;
assign n_17006 = n_16848 ^ n_16353;
assign n_17007 = n_16848 & ~n_16505;
assign n_17008 = ~n_16506 & n_16850;
assign n_17009 = n_16507 & n_16852;
assign n_17010 = n_16508 & n_16854;
assign n_17011 = n_16855 ^ n_16032;
assign n_17012 = n_16855 & ~n_16509;
assign n_17013 = n_16856 ^ n_16526;
assign n_17014 = n_16857 ^ n_16192;
assign n_17015 = n_16857 ^ n_16048;
assign n_17016 = n_16858 ^ n_16528;
assign n_17017 = n_16671 ^ n_16864;
assign n_17018 = n_16482 ^ n_16864;
assign n_17019 = n_16865 ^ n_16672;
assign n_17020 = n_16865 ^ n_16364;
assign n_17021 = n_16866 ^ n_16673;
assign n_17022 = n_16866 ^ n_16366;
assign n_17023 = n_16867 ^ n_16674;
assign n_17024 = n_16867 ^ n_16485;
assign n_17025 = n_16868 ^ n_16675;
assign n_17026 = n_16868 ^ n_16370;
assign n_17027 = n_16869 ^ n_16676;
assign n_17028 = n_16869 ^ n_16372;
assign n_17029 = n_16870 ^ n_16677;
assign n_17030 = n_16870 ^ n_16374;
assign n_17031 = n_16871 ^ n_16678;
assign n_17032 = n_16871 ^ n_16489;
assign n_17033 = n_16872 ^ n_16679;
assign n_17034 = n_16872 ^ n_16491;
assign n_17035 = n_16873 ^ n_16520;
assign n_17036 = n_16828 ^ n_16874;
assign n_17037 = n_16875 ^ n_16493;
assign n_17038 = n_16832 ^ n_16876;
assign n_17039 = n_16877 ^ n_16680;
assign n_17040 = n_16877 ^ n_16494;
assign n_17041 = ~x0 & n_16879;
assign n_17042 = n_16880 ^ x5;
assign n_17043 = n_16881 ^ x8;
assign n_17044 = n_16882 ^ x11;
assign n_17045 = n_16883 ^ x14;
assign n_17046 = n_16884 ^ x17;
assign n_17047 = n_16885 ^ x20;
assign n_17048 = n_16886 ^ x23;
assign n_17049 = n_16887 ^ x26;
assign n_17050 = n_16888 ^ x29;
assign n_17051 = n_16889 ^ x32;
assign n_17052 = n_16890 ^ x35;
assign n_17053 = n_16891 ^ x38;
assign n_17054 = n_16892 ^ x41;
assign n_17055 = n_16893 ^ x44;
assign n_17056 = n_16894 ^ x47;
assign n_17057 = n_16895 ^ x50;
assign n_17058 = n_16896 ^ x53;
assign n_17059 = n_16897 ^ x56;
assign n_17060 = n_16898 ^ x59;
assign n_17061 = n_16899 ^ x62;
assign n_17062 = ~x0 & n_16900;
assign n_17063 = n_16901 ^ x5;
assign n_17064 = n_16902 ^ x8;
assign n_17065 = n_16903 ^ x11;
assign n_17066 = n_16904 ^ x14;
assign n_17067 = n_16905 ^ x17;
assign n_17068 = n_16906 ^ x20;
assign n_17069 = n_16907 ^ x23;
assign n_17070 = n_16908 ^ x26;
assign n_17071 = n_16909 ^ x29;
assign n_17072 = n_16910 ^ x32;
assign n_17073 = n_16911 ^ x35;
assign n_17074 = n_16912 ^ x38;
assign n_17075 = n_16913 ^ x41;
assign n_17076 = n_16914 ^ x44;
assign n_17077 = n_16915 ^ x47;
assign n_17078 = n_16916 ^ x50;
assign n_17079 = n_16917 ^ x53;
assign n_17080 = n_16918 ^ x56;
assign n_17081 = n_16919 ^ x59;
assign n_17082 = n_16920 ^ x62;
assign n_17083 = n_311 & n_16921;
assign n_17084 = n_16922 ^ x4;
assign n_17085 = n_16923 ^ x13;
assign n_17086 = n_16924 ^ x16;
assign n_17087 = n_16925 ^ x19;
assign n_17088 = n_16926 ^ x22;
assign n_17089 = n_16928 ^ x28;
assign n_17090 = n_16929 ^ x34;
assign n_17091 = n_16930 ^ x37;
assign n_17092 = n_16932 ^ x43;
assign n_17093 = n_16933 ^ x46;
assign n_17094 = n_16934 ^ x49;
assign n_17095 = n_16935 ^ x52;
assign n_17096 = ~n_293 & ~n_16939;
assign n_17097 = ~n_297 & ~n_16940;
assign n_17098 = n_16944 ^ n_16618;
assign n_17099 = n_16945 ^ n_16619;
assign n_17100 = n_16946 ^ n_16620;
assign n_17101 = n_16947 ^ n_16621;
assign n_17102 = n_16948 ^ n_16622;
assign n_17103 = n_16949 ^ n_16623;
assign n_17104 = n_16950 ^ n_16624;
assign n_17105 = n_16952 ^ n_16625;
assign n_17106 = n_16954 ^ n_16626;
assign n_17107 = n_16956 ^ n_16627;
assign n_17108 = n_16958 ^ n_16629;
assign n_17109 = n_16960 ^ n_16311;
assign n_17110 = n_16962 ^ n_16631;
assign n_17111 = n_16963 ^ n_15757;
assign n_17112 = n_16963 ^ n_15616;
assign n_17113 = n_16964 ^ n_11128;
assign n_17114 = ~n_15736 & n_16965;
assign n_17115 = n_16966 ^ n_11129;
assign n_17116 = n_15738 & ~n_16967;
assign n_17117 = n_16968 ^ n_11130;
assign n_17118 = ~n_15366 & n_16969;
assign n_17119 = n_16970 ^ n_11133;
assign n_17120 = n_15742 & ~n_16971;
assign n_17121 = n_16972 ^ n_11134;
assign n_17122 = ~n_15744 & n_16973;
assign n_17123 = n_16974 ^ n_11728;
assign n_17124 = n_15606 & ~n_16975;
assign n_17125 = n_16977 ^ n_16646;
assign n_17126 = n_16978 ^ n_14166;
assign n_17127 = ~n_15622 & n_16979;
assign n_17128 = n_16980 ^ n_16345;
assign n_17129 = ~n_15807 & n_16981;
assign n_17130 = n_16982 ^ n_15865;
assign n_17131 = n_16982 ^ n_15732;
assign n_17132 = n_16983 ^ n_15755;
assign n_17133 = n_16983 ^ n_15614;
assign n_17134 = n_16984 ^ n_11586;
assign n_17135 = ~n_15877 & n_16985;
assign n_17136 = n_16986 ^ n_11440;
assign n_17137 = ~n_16136 & n_16987;
assign n_17138 = n_16988 ^ n_11444;
assign n_17139 = ~n_15761 & n_16989;
assign n_17140 = n_16990 ^ n_11445;
assign n_17141 = n_16142 & ~n_16991;
assign n_17142 = n_16993 ^ n_16663;
assign n_17143 = n_16356 ^ n_16995;
assign n_17144 = n_16996 ^ n_16995;
assign n_17145 = n_16997 ^ n_15658;
assign n_17146 = n_16998 ^ n_16876;
assign n_17147 = n_16999 ^ n_16683;
assign n_17148 = n_17000 ^ n_16684;
assign n_17149 = n_17001 ^ n_16685;
assign n_17150 = n_17002 ^ n_16686;
assign n_17151 = n_17003 ^ n_16687;
assign n_17152 = n_17004 ^ n_16688;
assign n_17153 = n_17005 ^ n_16689;
assign n_17154 = n_17007 ^ n_16690;
assign n_17155 = n_17008 ^ n_16691;
assign n_17156 = n_17009 ^ n_16693;
assign n_17157 = n_17010 ^ n_16695;
assign n_17158 = n_17012 ^ n_16696;
assign n_17159 = n_17013 ^ n_16961;
assign n_17160 = n_16671 & n_17018;
assign n_17161 = ~n_16672 & n_17020;
assign n_17162 = n_16673 & ~n_17022;
assign n_17163 = n_16927 ^ n_17023;
assign n_17164 = ~n_17023 & ~n_16927;
assign n_17165 = ~n_16674 & n_17024;
assign n_17166 = n_16675 & ~n_17026;
assign n_17167 = n_16943 ^ n_17027;
assign n_17168 = n_16676 & ~n_17028;
assign n_17169 = n_16677 & ~n_17030;
assign n_17170 = ~n_16678 & n_17032;
assign n_17171 = n_17033 & ~n_16931;
assign n_17172 = n_16931 ^ n_17033;
assign n_17173 = n_16679 & n_17034;
assign n_17174 = n_17035 ^ n_16492;
assign n_17175 = ~n_17035 & n_16692;
assign n_17176 = n_17036 ^ n_16665;
assign n_17177 = ~n_17036 & n_16994;
assign n_17178 = n_17037 ^ n_16522;
assign n_17179 = n_17037 & n_16694;
assign n_17180 = ~n_16998 & n_17038;
assign n_17181 = ~n_16680 & n_17040;
assign n_17182 = n_17041 ^ n_16721;
assign n_17183 = n_17047 ^ n_16834;
assign n_17184 = ~n_16834 & n_17047;
assign n_17185 = n_17048 ^ n_16836;
assign n_17186 = n_17049 ^ n_16838;
assign n_17187 = n_17050 ^ n_16840;
assign n_17188 = n_17051 ^ n_16842;
assign n_17189 = ~n_16842 & ~n_17051;
assign n_17190 = n_17052 ^ n_16844;
assign n_17191 = n_17053 ^ n_16846;
assign n_17192 = n_17055 ^ n_16849;
assign n_17193 = n_17056 ^ n_16851;
assign n_17194 = n_17058 ^ n_16853;
assign n_17195 = n_17011 ^ n_17059;
assign n_17196 = n_17059 & n_17011;
assign n_17197 = n_17060 ^ n_16697;
assign n_17198 = n_17061 ^ n_6422;
assign n_17199 = n_17062 ^ n_16742;
assign n_17200 = n_16786 ^ n_17068;
assign n_17201 = n_16788 ^ n_17069;
assign n_17202 = n_16790 ^ n_17070;
assign n_17203 = n_16792 ^ n_17071;
assign n_17204 = n_16794 ^ n_17072;
assign n_17205 = n_16796 ^ n_17073;
assign n_17206 = n_17073 & ~n_16796;
assign n_17207 = n_16798 ^ n_17074;
assign n_17208 = n_16951 ^ n_17075;
assign n_17209 = n_16953 ^ n_17076;
assign n_17210 = n_16955 ^ n_17077;
assign n_17211 = n_17077 & n_16955;
assign n_17212 = n_16957 ^ n_17079;
assign n_17213 = n_16959 ^ n_17080;
assign n_17214 = n_17013 ^ n_17081;
assign n_17215 = n_17082 ^ n_6540;
assign n_17216 = n_17083 ^ n_16591;
assign n_17217 = n_17086 ^ n_17017;
assign n_17218 = n_17088 ^ n_17021;
assign n_17219 = n_17089 ^ n_17025;
assign n_17220 = n_17090 ^ n_17029;
assign n_17221 = n_17091 ^ n_17031;
assign n_17222 = n_17096 ^ x125;
assign n_17223 = n_17097 ^ x126;
assign n_17224 = n_16939 ^ n_17097;
assign n_17225 = n_17087 ^ n_17098;
assign n_17226 = ~n_17098 & ~n_17087;
assign n_17227 = n_17099 ^ n_17021;
assign n_17228 = n_17101 ^ n_17025;
assign n_17229 = n_17027 ^ n_17102;
assign n_17230 = n_17103 ^ n_17029;
assign n_17231 = n_17104 ^ n_17031;
assign n_17232 = n_17105 ^ n_16931;
assign n_17233 = n_17092 ^ n_17106;
assign n_17234 = n_17109 ^ n_16936;
assign n_17235 = n_16936 & ~n_17109;
assign n_17236 = n_17110 ^ ~n_6539;
assign n_17237 = ~n_6539 & ~n_17110;
assign n_17238 = n_17111 ^ n_11439;
assign n_17239 = ~n_15757 & n_17112;
assign n_17240 = n_17114 ^ n_16809;
assign n_17241 = n_17116 ^ n_16810;
assign n_17242 = n_17118 ^ n_16811;
assign n_17243 = n_17120 ^ n_16812;
assign n_17244 = n_17122 ^ n_16813;
assign n_17245 = n_17124 ^ n_16814;
assign n_17246 = n_17125 ^ n_16149;
assign n_17247 = n_17125 ^ n_16008;
assign n_17248 = n_17127 ^ n_16817;
assign n_17249 = n_17129 ^ n_16818;
assign n_17250 = n_17130 ^ n_11438;
assign n_17251 = ~n_15865 & n_17131;
assign y31 = n_17132;
assign n_17252 = ~n_15755 & n_17133;
assign n_17253 = n_17135 ^ n_16822;
assign n_17254 = n_17137 ^ n_16823;
assign n_17255 = n_17139 ^ n_16824;
assign n_17256 = n_17141 ^ n_16000;
assign n_17257 = n_17142 ^ n_16151;
assign n_17258 = n_17142 ^ n_16010;
assign n_17259 = n_16996 & n_17143;
assign n_17260 = n_17144 ^ n_17057;
assign n_17261 = ~n_17057 & n_17144;
assign n_17262 = n_17145 ^ n_16628;
assign n_17263 = n_17145 ^ n_16335;
assign n_17264 = n_17095 ^ n_17146;
assign n_17265 = n_17146 ^ n_17108;
assign n_17266 = n_17147 ^ n_16786;
assign n_17267 = n_17148 ^ n_16788;
assign n_17268 = n_17149 ^ n_16790;
assign n_17269 = n_17150 ^ n_16792;
assign n_17270 = n_17151 ^ n_16794;
assign n_17271 = n_17153 ^ n_16798;
assign n_17272 = n_17154 ^ n_16951;
assign n_17273 = n_17155 ^ n_16953;
assign n_17274 = n_17157 ^ n_16957;
assign n_17275 = n_17158 ^ n_16959;
assign n_17276 = n_17159 ^ n_17081;
assign n_17277 = n_17160 ^ n_16864;
assign n_17278 = n_17161 ^ n_16865;
assign n_17279 = n_17162 ^ n_16866;
assign n_17280 = n_17100 ^ n_17163;
assign n_17281 = n_17164 ^ n_17163;
assign n_17282 = n_17165 ^ n_16867;
assign n_17283 = n_17166 ^ n_16868;
assign n_17284 = n_17167 ^ n_17102;
assign n_17285 = n_17168 ^ n_16869;
assign n_17286 = n_17169 ^ n_16870;
assign n_17287 = n_17170 ^ n_16871;
assign n_17288 = ~n_17105 & n_17171;
assign n_17289 = n_17171 ^ n_17172;
assign n_17290 = n_17173 ^ n_16872;
assign n_17291 = ~n_17174 & n_17092;
assign n_17292 = n_17092 ^ n_17174;
assign n_17293 = n_17175 ^ n_16873;
assign n_17294 = n_17093 ^ n_17176;
assign n_17295 = n_17176 ^ n_17107;
assign n_17296 = n_17177 ^ n_16874;
assign n_17297 = n_17179 ^ n_16875;
assign n_17298 = n_17180 ^ n_16876;
assign n_17299 = n_17181 ^ n_16877;
assign n_17300 = n_17184 ^ n_17183;
assign n_17301 = n_17189 ^ n_17188;
assign n_17302 = n_17196 ^ n_17195;
assign n_17303 = ~n_621 & ~n_17199;
assign n_17304 = n_17205 ^ n_17152;
assign n_17305 = n_17206 ^ n_17205;
assign n_17306 = n_17210 ^ n_17156;
assign n_17307 = n_17211 ^ n_17210;
assign n_17308 = ~n_17159 & n_17214;
assign n_17309 = n_17215 ^ n_3423;
assign n_17310 = n_17215 & n_6648;
assign n_17311 = n_17216 ^ x2;
assign n_17312 = n_17222 ^ n_17223;
assign n_17313 = x63 & ~n_17224;
assign n_17314 = n_17226 ^ n_17225;
assign n_17315 = n_17088 ^ n_17227;
assign n_17316 = n_17227 & ~n_17218;
assign n_17317 = n_17089 ^ n_17228;
assign n_17318 = n_17228 & ~n_17219;
assign n_17319 = ~n_17167 & n_17229;
assign n_17320 = n_17090 ^ n_17230;
assign n_17321 = n_17230 & ~n_17220;
assign n_17322 = n_17091 ^ n_17231;
assign n_17323 = ~n_17231 & n_17221;
assign n_17324 = n_17232 ^ n_17033;
assign n_17325 = n_17233 ^ n_17174;
assign n_17326 = n_17235 ^ n_17234;
assign n_17327 = n_17236 ^ n_16878;
assign n_17328 = ~n_16878 & ~n_17236;
assign n_17329 = n_17237 ^ n_6421;
assign n_17330 = n_17239 ^ n_16963;
assign n_17331 = n_17240 ^ n_16138;
assign n_17332 = n_17240 ^ n_15996;
assign n_17333 = n_17241 ^ n_16140;
assign n_17334 = n_17241 ^ n_15998;
assign n_17335 = n_17242 ^ n_15759;
assign n_17336 = n_17242 ^ n_15618;
assign n_17337 = n_17243 ^ n_16144;
assign n_17338 = n_17243 ^ n_16002;
assign n_17339 = n_17244 ^ n_16146;
assign n_17340 = n_17244 ^ n_16004;
assign n_17341 = n_17245 ^ n_16006;
assign n_17342 = n_17245 ^ n_15873;
assign n_17343 = n_17246 ^ n_13642;
assign n_17344 = n_16149 & ~n_17247;
assign n_17345 = n_17248 ^ n_16022;
assign n_17346 = n_17248 ^ n_15884;
assign n_17347 = n_17249 ^ n_16193;
assign n_17348 = n_17251 ^ n_16982;
assign n_17349 = n_17252 ^ n_16983;
assign n_17350 = n_17253 ^ n_16296;
assign n_17351 = n_17253 ^ n_16153;
assign n_17352 = n_17254 ^ n_16634;
assign n_17353 = n_17254 ^ n_16436;
assign n_17354 = n_17255 ^ n_16163;
assign n_17355 = n_17255 ^ n_16020;
assign n_17356 = n_17256 ^ n_16640;
assign n_17357 = n_17256 ^ n_10862;
assign n_17358 = n_17257 ^ n_16053;
assign n_17359 = n_16151 & ~n_17258;
assign n_17360 = n_17259 ^ n_16995;
assign n_17361 = n_17261 ^ n_17260;
assign n_17362 = n_17262 ^ n_16335;
assign n_17363 = ~n_17262 & ~n_17263;
assign n_17364 = n_17264 ^ n_17108;
assign n_17365 = n_17264 & ~n_17265;
assign n_17366 = n_17266 ^ n_17068;
assign n_17367 = n_17266 & ~n_17200;
assign n_17368 = n_17267 ^ n_17069;
assign n_17369 = ~n_17267 & n_17201;
assign n_17370 = n_17268 ^ n_17070;
assign n_17371 = n_17268 & ~n_17202;
assign n_17372 = n_17269 ^ n_17071;
assign n_17373 = n_17269 & ~n_17203;
assign n_17374 = n_17270 ^ n_17072;
assign n_17375 = n_17270 & ~n_17204;
assign n_17376 = n_17271 ^ n_17074;
assign n_17377 = n_17271 & ~n_17207;
assign n_17378 = n_17272 ^ n_17075;
assign n_17379 = ~n_17272 & n_17208;
assign n_17380 = n_17273 ^ n_17076;
assign n_17381 = ~n_17273 & n_17209;
assign n_17382 = n_17274 ^ n_17079;
assign n_17383 = n_17274 & ~n_17212;
assign n_17384 = n_17275 ^ n_17080;
assign n_17385 = n_17275 & ~n_17213;
assign n_17386 = n_17277 ^ n_17183;
assign n_17387 = n_17278 ^ n_17185;
assign n_17388 = n_17278 ^ n_16836;
assign n_17389 = n_17279 ^ n_17186;
assign n_17390 = n_17279 ^ n_17049;
assign n_17391 = n_17049 & n_17279;
assign n_17392 = n_17282 ^ n_17187;
assign n_17393 = n_17282 ^ n_17050;
assign n_17394 = n_17189 ^ n_17283;
assign n_17395 = n_17285 ^ n_17190;
assign n_17396 = n_17285 ^ n_16844;
assign n_17397 = n_17286 ^ n_17191;
assign n_17398 = n_17286 ^ n_17053;
assign n_17399 = n_17287 ^ n_17054;
assign n_17400 = ~n_17054 & ~n_17287;
assign n_17401 = n_17105 & n_17289;
assign n_17402 = n_17290 ^ n_17192;
assign n_17403 = n_17290 ^ n_17055;
assign n_17404 = n_17291 ^ n_17292;
assign n_17405 = n_17293 ^ n_17193;
assign n_17406 = n_17293 ^ n_17056;
assign n_17407 = n_17294 ^ n_17107;
assign n_17408 = ~n_17294 & n_17295;
assign n_17409 = n_17261 ^ n_17296;
assign n_17410 = n_17297 ^ n_17194;
assign n_17411 = n_17297 ^ n_17058;
assign n_17412 = n_17299 ^ n_17060;
assign n_17413 = n_17308 ^ n_17081;
assign n_17414 = n_17310 ^ n_17082;
assign n_17415 = n_17311 ^ x127;
assign n_17416 = ~x63 & n_17312;
assign n_17417 = n_17313 ^ n_16780;
assign n_17418 = n_17314 ^ n_17019;
assign n_17419 = n_17316 ^ n_17088;
assign n_17420 = n_17318 ^ n_17089;
assign n_17421 = n_17319 ^ n_16943;
assign n_17422 = ~n_17305 & ~n_17320;
assign n_17423 = n_17321 ^ n_17090;
assign n_17424 = n_17323 ^ n_17091;
assign n_17425 = n_17326 ^ n_17039;
assign n_17426 = n_17328 ^ n_17327;
assign n_17427 = n_17329 ^ n_17198;
assign n_17428 = n_17329 ^ n_17061;
assign n_17429 = n_17330 ^ n_16159;
assign n_17430 = n_17330 ^ n_16016;
assign n_17431 = n_17331 ^ n_11441;
assign n_17432 = ~n_16138 & n_17332;
assign n_17433 = n_17333 ^ n_11442;
assign n_17434 = ~n_16140 & n_17334;
assign n_17435 = n_17335 ^ n_11443;
assign n_17436 = ~n_15759 & n_17336;
assign n_17437 = n_17337 ^ n_11446;
assign n_17438 = ~n_16144 & n_17338;
assign n_17439 = n_17339 ^ n_11447;
assign n_17440 = ~n_16146 & n_17340;
assign n_17441 = n_17341 ^ n_12665;
assign n_17442 = n_16006 & ~n_17342;
assign n_17443 = n_17344 ^ n_17125;
assign n_17444 = n_17345 ^ n_14790;
assign n_17445 = ~n_16022 & n_17346;
assign n_17446 = n_17347 ^ n_16617;
assign n_17447 = n_17347 & ~n_16785;
assign n_17448 = n_17348 ^ n_16284;
assign n_17449 = n_17348 ^ n_16134;
assign n_17450 = n_17349 ^ n_16157;
assign n_17451 = n_17349 ^ n_16014;
assign n_17452 = n_17350 ^ n_11696;
assign n_17453 = ~n_16296 & n_17351;
assign n_17454 = n_17352 ^ n_11632;
assign n_17455 = ~n_16634 & n_17353;
assign n_17456 = n_17354 ^ n_11636;
assign n_17457 = ~n_16163 & n_17355;
assign n_17458 = n_17356 ^ n_11637;
assign n_17459 = n_16640 & ~n_17357;
assign n_17460 = n_17359 ^ n_17142;
assign n_17461 = n_17362 ^ n_17360;
assign n_17462 = n_17362 ^ n_17078;
assign n_17463 = n_17363 ^ n_16628;
assign n_17464 = n_17365 ^ n_17095;
assign n_17465 = n_17300 ^ n_17366;
assign n_17466 = n_17367 ^ n_17147;
assign n_17467 = n_17369 ^ n_17148;
assign n_17468 = n_17371 ^ n_17149;
assign n_17469 = n_17373 ^ n_17150;
assign n_17470 = n_17374 ^ n_17301;
assign n_17471 = n_17301 ^ ~n_17374;
assign n_17472 = n_17375 ^ n_17151;
assign n_17473 = n_17377 ^ n_17153;
assign n_17474 = n_17379 ^ n_17154;
assign n_17475 = n_17381 ^ n_17155;
assign n_17476 = n_17383 ^ n_17157;
assign n_17477 = n_17384 ^ n_17196;
assign n_17478 = n_17385 ^ n_17158;
assign n_17479 = n_17387 ^ n_17226;
assign n_17480 = ~n_17185 & n_17388;
assign n_17481 = n_17391 ^ n_17390;
assign n_17482 = n_17391 ^ n_17370;
assign n_17483 = n_17392 ^ n_17281;
assign n_17484 = n_17187 & n_17393;
assign n_17485 = n_17190 & ~n_17396;
assign n_17486 = n_17191 & n_17398;
assign n_17487 = n_17400 ^ n_17006;
assign n_17488 = n_17400 ^ n_17399;
assign n_17489 = n_17288 ^ n_17401;
assign n_17490 = ~n_17192 & n_17403;
assign n_17491 = n_17405 ^ n_17404;
assign n_17492 = n_17193 & n_17406;
assign n_17493 = n_17307 & ~n_17407;
assign n_17494 = n_17408 ^ n_17093;
assign n_17495 = n_17194 & n_17411;
assign n_17496 = n_17412 ^ n_16697;
assign n_17497 = n_17412 & n_17197;
assign n_17498 = n_17413 ^ n_16937;
assign n_17499 = ~n_16937 & ~n_17413;
assign n_17500 = n_17414 ^ n_16938;
assign n_17501 = n_1 & n_17415;
assign n_17502 = n_17416 ^ n_17222;
assign n_17503 = n_17419 ^ n_17389;
assign n_17504 = ~n_17049 & ~n_17419;
assign n_17505 = n_17419 ^ n_16838;
assign n_17506 = ~n_16838 & n_17419;
assign n_17507 = n_17420 ^ n_17283;
assign n_17508 = ~n_17283 & ~n_17420;
assign n_17509 = n_17421 ^ n_17395;
assign n_17510 = n_17423 ^ n_17397;
assign n_17511 = n_17424 ^ n_17006;
assign n_17512 = n_17006 & n_17424;
assign n_17513 = n_17198 & ~n_17428;
assign n_17514 = n_17429 ^ n_11631;
assign n_17515 = ~n_16159 & n_17430;
assign n_17516 = n_17432 ^ n_17240;
assign n_17517 = n_17434 ^ n_17241;
assign n_17518 = n_17436 ^ n_17242;
assign n_17519 = n_17438 ^ n_17243;
assign n_17520 = n_17440 ^ n_17244;
assign n_17521 = n_17442 ^ n_17245;
assign n_17522 = n_17443 ^ n_16647;
assign n_17523 = n_17443 ^ n_16450;
assign n_17524 = n_17445 ^ n_17248;
assign n_17525 = n_17067 & n_17446;
assign n_17526 = n_17446 ^ n_17067;
assign n_17527 = n_17447 ^ n_17249;
assign n_17528 = n_17448 ^ n_11630;
assign n_17529 = ~n_16284 & n_17449;
assign y32 = n_17450;
assign n_17530 = ~n_16157 & n_17451;
assign n_17531 = n_17453 ^ n_17253;
assign n_17532 = n_17455 ^ n_17254;
assign n_17533 = n_17457 ^ n_17255;
assign n_17534 = n_17459 ^ n_16442;
assign n_17535 = n_17460 ^ n_16452;
assign n_17536 = n_17461 ^ n_17078;
assign n_17537 = n_17461 & ~n_17462;
assign n_17538 = n_17094 ^ n_17463;
assign n_17539 = n_17463 & n_17094;
assign n_17540 = n_17464 ^ n_17298;
assign n_17541 = ~n_17298 & ~n_17464;
assign n_17542 = n_17466 ^ n_17019;
assign n_17543 = n_17019 & n_17466;
assign n_17544 = n_17315 ^ n_17467;
assign n_17545 = n_17468 ^ n_17280;
assign n_17546 = n_17100 & n_17468;
assign n_17547 = n_17468 ^ n_17100;
assign n_17548 = n_17317 ^ n_17469;
assign n_17549 = n_17472 ^ n_17284;
assign n_17550 = n_17322 ^ n_17473;
assign n_17551 = n_17474 ^ n_17324;
assign n_17552 = n_17474 & n_17401;
assign n_17553 = n_17325 ^ n_17475;
assign n_17554 = n_17475 & n_17106;
assign n_17555 = n_17106 ^ n_17475;
assign n_17556 = n_17364 ^ n_17476;
assign n_17557 = n_17478 ^ n_17039;
assign n_17558 = ~n_17039 & ~n_17478;
assign n_17559 = n_17480 ^ n_17048;
assign n_17560 = n_17484 ^ n_17282;
assign n_17561 = n_17485 ^ n_17052;
assign n_17562 = n_17486 ^ n_17286;
assign n_17563 = n_17378 ^ n_17488;
assign n_17564 = n_17489 ^ n_17324;
assign n_17565 = n_17490 ^ n_17290;
assign n_17566 = n_17492 ^ n_17293;
assign n_17567 = n_17494 ^ n_17296;
assign n_17568 = n_17296 & n_17494;
assign n_17569 = n_17495 ^ n_17297;
assign n_17570 = ~n_17235 ^ n_17496;
assign n_17571 = n_17497 ^ n_17299;
assign n_17572 = n_17498 ^ n_17327;
assign n_17573 = n_17499 ^ n_17498;
assign n_17574 = n_17499 & n_17328;
assign n_17575 = n_17426 ^ n_17499;
assign n_17576 = ~n_17499 & n_17427;
assign n_17577 = ~n_17499 & ~n_17426;
assign n_17578 = n_17501 ^ n_1;
assign n_17579 = n_17502 ^ n_17417;
assign n_17580 = n_17503 ^ n_17279;
assign n_17581 = n_17503 ^ n_16838;
assign n_17582 = n_17505 ^ n_17506;
assign n_17583 = n_17506 ^ n_17370;
assign n_17584 = n_17507 ^ n_17188;
assign n_17585 = n_17189 ^ n_17507;
assign n_17586 = ~n_17507 & ~n_17301;
assign n_17587 = n_17507 & ~n_17394;
assign n_17588 = n_17508 ^ n_17507;
assign n_17589 = ~n_17508 & n_17471;
assign n_17590 = n_17511 ^ n_17399;
assign n_17591 = n_17511 & n_17487;
assign n_17592 = n_17488 ^ n_17511;
assign n_17593 = n_17512 ^ n_17511;
assign n_17594 = n_17378 ^ n_17512;
assign n_17595 = n_17513 ^ n_17329;
assign n_17596 = n_17515 ^ n_17330;
assign n_17597 = n_17516 ^ n_16636;
assign n_17598 = n_17516 ^ n_16438;
assign n_17599 = n_17517 ^ n_16638;
assign n_17600 = n_17517 ^ n_16440;
assign n_17601 = n_17518 ^ n_16161;
assign n_17602 = n_17518 ^ n_16018;
assign n_17603 = n_17519 ^ n_16642;
assign n_17604 = n_17519 ^ n_16444;
assign n_17605 = n_17520 ^ n_16644;
assign n_17606 = n_17520 ^ n_16446;
assign n_17607 = n_17521 ^ n_16448;
assign n_17608 = n_17521 ^ n_16292;
assign n_17609 = n_17522 ^ n_14473;
assign n_17610 = n_16647 & ~n_17523;
assign n_17611 = n_17524 ^ n_16464;
assign n_17612 = n_17524 ^ n_16303;
assign n_17613 = n_17525 ^ n_17526;
assign n_17614 = n_17217 ^ n_17527;
assign n_17615 = n_17086 ^ n_17527;
assign n_17616 = n_17529 ^ n_17348;
assign n_17617 = n_17530 ^ n_17349;
assign n_17618 = n_17531 ^ n_16819;
assign n_17619 = n_17531 ^ n_16651;
assign n_17620 = n_17532 ^ n_17113;
assign n_17621 = n_17532 ^ n_16964;
assign n_17622 = n_17533 ^ n_16661;
assign n_17623 = n_17533 ^ n_16462;
assign n_17624 = n_17534 ^ n_17119;
assign n_17625 = n_17534 ^ n_11133;
assign n_17626 = n_17535 ^ n_16244;
assign n_17627 = n_17535 & ~n_16649;
assign n_17628 = ~n_17361 ^ ~n_17536;
assign n_17629 = n_17537 ^ n_17360;
assign n_17630 = n_17539 ^ n_17178;
assign n_17631 = n_17539 ^ n_17538;
assign n_17632 = n_17540 ^ n_17195;
assign n_17633 = n_17540 & n_17196;
assign n_17634 = n_17541 ^ n_17540;
assign n_17635 = ~n_17541 & n_17477;
assign n_17636 = n_17225 ^ n_17542;
assign n_17637 = n_17542 & n_17418;
assign n_17638 = n_17543 ^ n_17542;
assign n_17639 = ~n_17543 & n_17479;
assign n_17640 = ~n_17546 & n_17281;
assign n_17641 = ~n_17546 & n_17164;
assign n_17642 = ~n_17546 ^ n_17392;
assign n_17643 = n_17546 ^ n_17547;
assign n_17644 = n_17554 ^ n_17174;
assign n_17645 = n_17554 ^ n_17555;
assign n_17646 = n_17291 & n_17555;
assign n_17647 = n_17555 ^ n_17404;
assign n_17648 = n_17557 ^ n_17234;
assign n_17649 = n_17557 & n_17235;
assign n_17650 = n_17326 ^ n_17557;
assign n_17651 = n_17557 & n_17425;
assign n_17652 = n_17558 ^ n_17557;
assign n_17653 = n_17559 ^ n_17368;
assign n_17654 = n_17560 ^ n_17372;
assign n_17655 = n_17561 ^ n_17304;
assign n_17656 = ~n_17152 & ~n_17561;
assign n_17657 = n_17561 ^ n_17152;
assign n_17658 = n_17562 ^ n_17376;
assign n_17659 = ~n_17474 & ~n_17564;
assign n_17660 = n_17565 ^ n_17380;
assign n_17661 = n_17566 ^ n_17306;
assign n_17662 = n_17156 & n_17566;
assign n_17663 = n_17566 ^ n_17156;
assign n_17664 = n_17567 ^ n_17260;
assign n_17665 = n_17567 & n_17409;
assign n_17666 = n_17260 & ~n_17568;
assign n_17667 = n_17568 ^ n_17567;
assign n_17668 = n_17536 ^ n_17568;
assign n_17669 = n_17569 ^ n_17382;
assign n_17670 = ~n_17558 & n_17570;
assign n_17671 = n_17571 ^ n_17276;
assign n_17672 = n_17328 ^ n_17573;
assign n_17673 = ~n_17573 & ~n_17426;
assign n_17674 = n_17573 & n_17328;
assign n_17675 = n_17573 & ~n_17427;
assign n_17676 = n_17577 ^ n_17576;
assign n_17677 = n_17578 ^ x2;
assign n_17678 = x62 & n_17579;
assign n_17679 = ~n_17580 & n_17581;
assign n_17680 = n_17582 ^ n_17279;
assign n_17681 = n_17583 & n_17481;
assign n_17682 = n_17587 ^ n_17283;
assign n_17683 = n_17588 ^ n_17374;
assign n_17684 = n_17591 ^ n_17424;
assign n_17685 = n_17593 & n_17563;
assign n_17686 = n_17595 ^ n_17309;
assign n_17687 = n_17596 ^ n_16657;
assign n_17688 = n_17596 ^ n_16458;
assign n_17689 = n_17597 ^ n_11633;
assign n_17690 = n_16636 & ~n_17598;
assign n_17691 = n_17599 ^ n_11634;
assign n_17692 = ~n_16638 & n_17600;
assign n_17693 = n_17601 ^ n_11635;
assign n_17694 = ~n_16161 & n_17602;
assign n_17695 = n_17603 ^ n_11638;
assign n_17696 = ~n_16642 & n_17604;
assign n_17697 = n_17605 ^ n_11639;
assign n_17698 = ~n_16644 & n_17606;
assign n_17699 = n_17607 ^ n_13299;
assign n_17700 = ~n_16448 & n_17608;
assign n_17701 = n_17610 ^ n_17443;
assign n_17702 = n_17611 ^ n_15546;
assign n_17703 = ~n_16464 & n_17612;
assign n_17704 = n_17614 ^ n_17525;
assign n_17705 = n_17217 & n_17615;
assign n_17706 = n_17616 ^ n_16807;
assign n_17707 = n_17616 ^ n_16632;
assign n_17708 = n_17617 ^ n_16655;
assign n_17709 = n_17617 ^ n_16456;
assign n_17710 = n_17618 ^ n_11797;
assign n_17711 = ~n_16819 & n_17619;
assign n_17712 = n_17620 ^ n_11721;
assign n_17713 = ~n_17113 & n_17621;
assign n_17714 = n_17622 ^ n_11725;
assign n_17715 = n_16661 & ~n_17623;
assign n_17716 = n_17624 ^ n_11726;
assign n_17717 = ~n_17119 & ~n_17625;
assign n_17718 = n_17626 ^ n_16863;
assign n_17719 = n_17627 ^ n_17460;
assign n_17720 = n_17629 ^ n_17178;
assign n_17721 = n_17178 & ~n_17629;
assign n_17722 = n_17631 ^ ~n_17410;
assign n_17723 = ~n_17302 & n_17634;
assign n_17724 = n_17634 & ~n_17384;
assign n_17725 = n_17637 ^ n_17466;
assign n_17726 = n_17314 ^ n_17638;
assign n_17727 = n_17638 & ~n_17387;
assign n_17728 = n_17640 ^ n_17641;
assign n_17729 = ~n_17164 & n_17642;
assign n_17730 = n_17643 ^ n_16927;
assign n_17731 = ~n_17643 ^ n_17281;
assign n_17732 = n_17643 & n_17483;
assign n_17733 = ~n_17292 & n_17644;
assign n_17734 = n_17405 ^ n_17645;
assign n_17735 = n_17651 ^ n_17478;
assign n_17736 = n_17652 ^ n_17496;
assign n_17737 = n_17656 ^ n_17206;
assign n_17738 = n_17320 ^ n_17656;
assign n_17739 = n_17656 ^ n_17657;
assign n_17740 = n_17659 ^ n_17288;
assign n_17741 = ~n_17288 & ~n_17659;
assign n_17742 = ~n_17210 & n_17662;
assign n_17743 = n_17662 & n_17307;
assign n_17744 = n_17662 ^ n_17663;
assign n_17745 = n_17665 ^ n_17494;
assign n_17746 = n_17260 & n_17667;
assign n_17747 = n_17667 & n_17628;
assign n_17748 = ~n_17261 & n_17668;
assign n_17749 = ~n_17674 & n_17576;
assign n_17750 = ~n_17426 & ~n_17675;
assign n_17751 = ~n_17328 & ~n_17675;
assign n_17752 = n_17678 ^ n_17417;
assign n_17753 = n_17390 & ~n_17680;
assign n_17754 = n_17588 ^ n_17682;
assign n_17755 = ~n_17189 & ~n_17683;
assign n_17756 = n_17593 ^ n_17684;
assign n_17757 = n_17684 & ~n_17378;
assign n_17758 = n_17687 ^ n_11720;
assign n_17759 = n_16657 & ~n_17688;
assign n_17760 = n_17690 ^ n_17516;
assign n_17761 = n_17692 ^ n_17517;
assign n_17762 = n_17694 ^ n_17518;
assign n_17763 = n_17696 ^ n_17519;
assign n_17764 = n_17698 ^ n_17520;
assign n_17765 = n_17700 ^ n_17521;
assign n_17766 = n_17701 ^ n_17126;
assign n_17767 = n_17701 ^ n_16978;
assign n_17768 = n_17703 ^ n_17524;
assign n_17769 = n_17705 ^ n_17527;
assign n_17770 = n_17706 ^ n_11719;
assign n_17771 = ~n_16807 & n_17707;
assign y33 = n_17708;
assign n_17772 = ~n_16655 & n_17709;
assign n_17773 = n_17711 ^ n_17531;
assign n_17774 = n_17713 ^ n_17532;
assign n_17775 = n_17715 ^ n_17533;
assign n_17776 = n_17717 ^ n_16970;
assign n_17777 = n_17719 ^ n_17128;
assign n_17778 = n_17719 ^ n_16980;
assign n_17779 = n_17720 ^ n_17538;
assign n_17780 = ~n_17720 & n_17630;
assign n_17781 = ~n_17538 & ~n_17721;
assign n_17782 = n_17721 ^ n_17720;
assign n_17783 = n_17410 ^ n_17721;
assign n_17784 = ~n_17541 & ~n_17723;
assign n_17785 = n_17387 & ~n_17725;
assign n_17786 = n_17314 & ~n_17727;
assign n_17787 = n_17163 & ~n_17730;
assign n_17788 = n_17733 ^ n_17092;
assign n_17789 = ~n_17291 & ~n_17734;
assign n_17790 = ~n_17496 & n_17735;
assign n_17791 = ~n_17326 & n_17736;
assign n_17792 = ~n_17206 & n_17738;
assign n_17793 = n_17739 ^ n_17305;
assign n_17794 = n_17739 ^ n_16796;
assign n_17795 = n_17739 & ~n_17422;
assign n_17796 = n_17740 ^ n_17741;
assign n_17797 = n_17402 & n_17741;
assign n_17798 = n_17743 ^ n_17407;
assign n_17799 = n_17744 ^ n_17210;
assign n_17800 = n_17407 ^ n_17744;
assign n_17801 = n_17745 & n_17536;
assign n_17802 = ~n_17749 & ~n_17750;
assign n_17803 = n_17751 ^ n_17676;
assign n_17804 = n_17752 ^ n_6503;
assign n_17805 = n_17753 ^ n_17279;
assign n_17806 = n_17374 & n_17754;
assign n_17807 = ~n_17589 ^ ~n_17755;
assign n_17808 = n_17759 ^ n_17596;
assign n_17809 = n_17760 ^ n_17115;
assign n_17810 = n_17760 ^ n_16966;
assign n_17811 = n_17761 ^ n_17117;
assign n_17812 = n_17761 ^ n_16968;
assign n_17813 = n_17762 ^ n_16659;
assign n_17814 = n_17762 ^ n_16460;
assign n_17815 = n_17763 ^ n_17121;
assign n_17816 = n_17763 ^ n_16972;
assign n_17817 = n_17764 ^ n_17123;
assign n_17818 = n_17764 ^ n_16974;
assign n_17819 = n_17765 ^ n_16976;
assign n_17820 = n_17765 ^ n_16815;
assign n_17821 = n_17766 ^ n_14641;
assign n_17822 = ~n_17126 & n_17767;
assign n_17823 = n_17768 ^ n_16992;
assign n_17824 = n_17768 ^ n_16826;
assign n_17825 = n_17769 ^ n_17386;
assign n_17826 = n_17277 & n_17769;
assign n_17827 = n_17769 ^ n_17277;
assign n_17828 = n_17771 ^ n_17616;
assign n_17829 = n_17772 ^ n_17617;
assign n_17830 = n_17773 ^ n_17250;
assign n_17831 = n_17773 ^ n_17130;
assign n_17832 = n_17774 ^ n_17431;
assign n_17833 = n_17774 ^ n_17331;
assign n_17834 = n_17775 ^ n_17140;
assign n_17835 = n_17775 ^ n_16990;
assign n_17836 = n_17776 ^ n_17437;
assign n_17837 = n_17776 ^ n_11446;
assign n_17838 = n_17777 ^ n_17046;
assign n_17839 = ~n_17128 & n_17778;
assign n_17840 = n_17780 ^ n_17629;
assign n_17841 = ~n_17538 & ~n_17782;
assign n_17842 = ~n_17782 & n_17722;
assign n_17843 = ~n_17539 & n_17783;
assign n_17844 = n_17784 ^ n_17541;
assign n_17845 = n_17784 & n_17384;
assign n_17846 = n_17226 & n_17786;
assign n_17847 = ~n_17786 ^ ~n_17639;
assign n_17848 = n_17787 ^ n_17023;
assign n_17849 = n_17405 & ~n_17788;
assign n_17850 = ~n_17205 & ~n_17794;
assign n_17851 = n_17656 & n_17795;
assign n_17852 = ~n_17795 ^ ~n_17792;
assign n_17853 = n_17796 ^ n_17552;
assign n_17854 = ~n_17552 & ~n_17797;
assign n_17855 = ~n_17211 & ~n_17800;
assign n_17856 = n_17370 & n_17805;
assign n_17857 = n_17806 ^ n_17588;
assign n_17858 = n_17808 ^ n_17136;
assign n_17859 = n_17808 ^ n_16986;
assign n_17860 = n_17809 ^ n_11722;
assign n_17861 = n_17115 & ~n_17810;
assign n_17862 = n_17811 ^ n_11723;
assign n_17863 = ~n_17117 & n_17812;
assign n_17864 = n_17813 ^ n_11724;
assign n_17865 = ~n_16659 & n_17814;
assign n_17866 = n_17815 ^ n_11727;
assign n_17867 = ~n_17121 & n_17816;
assign n_17868 = n_17817 ^ n_12524;
assign n_17869 = n_17123 & ~n_17818;
assign n_17870 = n_17819 ^ n_13467;
assign n_17871 = n_16976 & ~n_17820;
assign n_17872 = n_17822 ^ n_17701;
assign n_17873 = n_17823 ^ n_15692;
assign n_17874 = ~n_16992 & n_17824;
assign n_17875 = n_17047 & n_17826;
assign n_17876 = ~n_17826 & ~n_17465;
assign n_17877 = n_17826 ^ n_17827;
assign n_17878 = n_17828 ^ n_17238;
assign n_17879 = n_17828 ^ n_17111;
assign n_17880 = n_17829 ^ n_17134;
assign n_17881 = n_17829 ^ n_16984;
assign n_17882 = n_17830 ^ n_11941;
assign n_17883 = ~n_17250 & n_17831;
assign n_17884 = n_17832 ^ n_11883;
assign n_17885 = ~n_17431 & n_17833;
assign n_17886 = n_17834 ^ n_11887;
assign n_17887 = ~n_17140 & n_17835;
assign n_17888 = n_17836 ^ n_11888;
assign n_17889 = n_17437 & n_17837;
assign n_17890 = n_17839 ^ n_17719;
assign n_17891 = ~n_17840 & n_17410;
assign n_17892 = n_17844 ^ n_17633;
assign n_17893 = ~n_17846 & ~n_17785;
assign n_17894 = n_17848 ^ ~n_17731;
assign n_17895 = n_17848 & ~n_17392;
assign n_17896 = n_17850 ^ n_17073;
assign n_17897 = n_17853 ^ n_17551;
assign n_17898 = ~n_17470 & n_17857;
assign n_17899 = n_17858 ^ n_11882;
assign n_17900 = ~n_17136 & n_17859;
assign n_17901 = n_17861 ^ n_17760;
assign n_17902 = n_17863 ^ n_17761;
assign n_17903 = n_17865 ^ n_17762;
assign n_17904 = n_17867 ^ n_17763;
assign n_17905 = n_17869 ^ n_17764;
assign n_17906 = n_17871 ^ n_17765;
assign n_17907 = n_17872 ^ n_17444;
assign n_17908 = n_17872 ^ n_17345;
assign n_17909 = n_17874 ^ n_17768;
assign n_17910 = n_17877 ^ n_16834;
assign n_17911 = n_17877 ^ n_17825;
assign n_17912 = n_17877 & n_17184;
assign n_17913 = n_17877 & n_17366;
assign n_17914 = n_17878 ^ n_11881;
assign n_17915 = ~n_17238 & n_17879;
assign y34 = n_17880;
assign n_17916 = ~n_17134 & n_17881;
assign n_17917 = n_17883 ^ n_17773;
assign n_17918 = n_17885 ^ n_17774;
assign n_17919 = n_17887 ^ n_17775;
assign n_17920 = n_17889 ^ n_17337;
assign n_17921 = n_17890 ^ n_17446;
assign n_17922 = n_17320 & ~n_17896;
assign n_17923 = n_17897 ^ n_17741;
assign n_17924 = n_17898 ^ n_17301;
assign n_17925 = n_17900 ^ n_17808;
assign n_17926 = n_17901 ^ n_17433;
assign n_17927 = n_17901 ^ n_17333;
assign n_17928 = n_17902 ^ n_17435;
assign n_17929 = n_17902 ^ n_17335;
assign n_17930 = n_17903 ^ n_17138;
assign n_17931 = n_17903 ^ n_16988;
assign n_17932 = n_17904 ^ n_17439;
assign n_17933 = n_17904 ^ n_17339;
assign n_17934 = n_17905 ^ n_17441;
assign n_17935 = n_17905 ^ n_17341;
assign n_17936 = n_17906 ^ n_17343;
assign n_17937 = n_17906 ^ n_17246;
assign n_17938 = n_17907 ^ n_15260;
assign n_17939 = ~n_17444 & n_17908;
assign n_17940 = n_17909 ^ n_17358;
assign n_17941 = n_17909 ^ n_17257;
assign n_17942 = n_17910 & n_17911;
assign n_17943 = n_17912 ^ n_17366;
assign n_17944 = n_17915 ^ n_17828;
assign n_17945 = n_17916 ^ n_17829;
assign n_17946 = n_17917 ^ n_17528;
assign n_17947 = n_17917 ^ n_17448;
assign n_17948 = n_17918 ^ n_17689;
assign n_17949 = n_17918 ^ n_17597;
assign n_17950 = n_17919 ^ n_17458;
assign n_17951 = n_17919 ^ n_17356;
assign n_17952 = n_17920 ^ n_17695;
assign n_17953 = n_17920 ^ n_11638;
assign n_17954 = n_17921 ^ n_17067;
assign n_17955 = ~n_17922 & ~n_17851;
assign n_17956 = ~n_17402 ^ n_17923;
assign n_17957 = n_17925 ^ n_17454;
assign n_17958 = n_17925 ^ n_17352;
assign n_17959 = n_17926 ^ n_11884;
assign n_17960 = ~n_17433 & n_17927;
assign n_17961 = n_17928 ^ n_11885;
assign n_17962 = ~n_17435 & n_17929;
assign n_17963 = n_17930 ^ n_11886;
assign n_17964 = ~n_17138 & n_17931;
assign n_17965 = n_17932 ^ n_11889;
assign n_17966 = ~n_17439 & n_17933;
assign n_17967 = n_17934 ^ n_13126;
assign n_17968 = n_17441 & ~n_17935;
assign n_17969 = n_17936 ^ n_14320;
assign n_17970 = n_17343 & ~n_17937;
assign n_17971 = n_17939 ^ n_17872;
assign n_17972 = n_17940 ^ n_16616;
assign n_17973 = n_17358 & ~n_17941;
assign n_17974 = n_17944 ^ n_17514;
assign n_17975 = n_17944 ^ n_17429;
assign n_17976 = n_17945 ^ n_17452;
assign n_17977 = n_17945 ^ n_17350;
assign n_17978 = n_17946 ^ n_12305;
assign n_17979 = ~n_17528 & n_17947;
assign n_17980 = n_17948 ^ n_12226;
assign n_17981 = n_17689 & ~n_17949;
assign n_17982 = n_17950 ^ n_12230;
assign n_17983 = ~n_17458 & n_17951;
assign n_17984 = n_17952 ^ n_12231;
assign n_17985 = n_17695 & ~n_17953;
assign n_17986 = n_17796 & n_17956;
assign n_17987 = n_17957 ^ n_12225;
assign n_17988 = ~n_17454 & n_17958;
assign n_17989 = n_17960 ^ n_17901;
assign n_17990 = n_17962 ^ n_17902;
assign n_17991 = n_17964 ^ n_17903;
assign n_17992 = n_17966 ^ n_17904;
assign n_17993 = n_17968 ^ n_17905;
assign n_17994 = n_17970 ^ n_17906;
assign n_17995 = n_17971 ^ n_17702;
assign n_17996 = n_17971 ^ n_17611;
assign n_17997 = n_17973 ^ n_17909;
assign n_17998 = n_17974 ^ n_12224;
assign n_17999 = ~n_17514 & n_17975;
assign y35 = n_17976;
assign n_18000 = ~n_17452 & n_17977;
assign n_18001 = n_17979 ^ n_17917;
assign n_18002 = n_17981 ^ n_17918;
assign n_18003 = n_17983 ^ n_17919;
assign n_18004 = n_17985 ^ n_17603;
assign n_18005 = n_17988 ^ n_17925;
assign n_18006 = n_17989 ^ n_17691;
assign n_18007 = n_17989 ^ n_17599;
assign n_18008 = n_17990 ^ n_17693;
assign n_18009 = n_17990 ^ n_17601;
assign n_18010 = n_17991 ^ n_17456;
assign n_18011 = n_17991 ^ n_17354;
assign n_18012 = n_17992 ^ n_17697;
assign n_18013 = n_17992 ^ n_17605;
assign n_18014 = n_17993 ^ n_17699;
assign n_18015 = n_17993 ^ n_17607;
assign n_18016 = n_17994 ^ n_17609;
assign n_18017 = n_17994 ^ n_17522;
assign n_18018 = n_17995 ^ n_16243;
assign n_18019 = ~n_17702 & n_17996;
assign n_18020 = n_17997 ^ n_17626;
assign n_18021 = n_17999 ^ n_17944;
assign n_18022 = n_18000 ^ n_17945;
assign n_18023 = n_18001 ^ n_17770;
assign n_18024 = n_18001 ^ n_17706;
assign n_18025 = n_18002 ^ n_17860;
assign n_18026 = n_18002 ^ n_17809;
assign n_18027 = n_18003 ^ n_17716;
assign n_18028 = n_18003 ^ n_17624;
assign n_18029 = n_18004 ^ n_17866;
assign n_18030 = n_18004 ^ n_17815;
assign n_18031 = n_18005 ^ n_17712;
assign n_18032 = n_18005 ^ n_17620;
assign n_18033 = n_18006 ^ n_12227;
assign n_18034 = ~n_17691 & n_18007;
assign n_18035 = n_18008 ^ n_12228;
assign n_18036 = ~n_17693 & n_18009;
assign n_18037 = n_18010 ^ n_12229;
assign n_18038 = ~n_17456 & n_18011;
assign n_18039 = n_18012 ^ n_12232;
assign n_18040 = ~n_17697 & n_18013;
assign n_18041 = n_18014 ^ n_14030;
assign n_18042 = ~n_17699 & n_18015;
assign n_18043 = n_18016 ^ n_14952;
assign n_18044 = n_17609 & ~n_18017;
assign n_18045 = n_18019 ^ n_17971;
assign n_18046 = n_18020 ^ n_16863;
assign n_18047 = n_18020 & ~n_17718;
assign n_18048 = n_18021 ^ n_17758;
assign n_18049 = n_18021 ^ n_17687;
assign n_18050 = n_18022 ^ n_17710;
assign n_18051 = n_18022 ^ n_17618;
assign n_18052 = n_18023 ^ n_12641;
assign n_18053 = ~n_17770 & n_18024;
assign n_18054 = n_18025 ^ n_12518;
assign n_18055 = n_17860 & ~n_18026;
assign n_18056 = n_18027 ^ n_12522;
assign n_18057 = n_17716 & ~n_18028;
assign n_18058 = n_18029 ^ n_12523;
assign n_18059 = ~n_17866 & n_18030;
assign n_18060 = n_18031 ^ n_12517;
assign n_18061 = ~n_17712 & n_18032;
assign n_18062 = n_18034 ^ n_17989;
assign n_18063 = n_18036 ^ n_17990;
assign n_18064 = n_18038 ^ n_17991;
assign n_18065 = n_18040 ^ n_17992;
assign n_18066 = n_18042 ^ n_17993;
assign n_18067 = n_18044 ^ n_17994;
assign n_18068 = n_18045 ^ n_17873;
assign n_18069 = n_18045 ^ n_17823;
assign n_18070 = n_18046 ^ n_17085;
assign n_18071 = n_17085 & n_18046;
assign n_18072 = n_18047 ^ n_17997;
assign n_18073 = n_18048 ^ n_12516;
assign n_18074 = n_17758 & ~n_18049;
assign y36 = n_18050;
assign n_18075 = ~n_17710 & n_18051;
assign n_18076 = n_18053 ^ n_18001;
assign n_18077 = n_18055 ^ n_18002;
assign n_18078 = n_18057 ^ n_18003;
assign n_18079 = n_18059 ^ n_18004;
assign n_18080 = n_18061 ^ n_18005;
assign n_18081 = n_18062 ^ n_17862;
assign n_18082 = n_18062 ^ n_17811;
assign n_18083 = n_18063 ^ n_17864;
assign n_18084 = n_18063 ^ n_17813;
assign n_18085 = n_18064 ^ n_17714;
assign n_18086 = n_18064 ^ n_17622;
assign n_18087 = n_18065 ^ n_17868;
assign n_18088 = n_18065 ^ n_17817;
assign n_18089 = n_18066 ^ n_17870;
assign n_18090 = n_18066 ^ n_17819;
assign n_18091 = n_18067 ^ n_17821;
assign n_18092 = n_18067 ^ n_17766;
assign n_18093 = n_18068 ^ n_16344;
assign n_18094 = ~n_17873 & n_18069;
assign n_18095 = n_18071 ^ n_18070;
assign n_18096 = n_18072 ^ n_17838;
assign n_18097 = n_18072 ^ n_17777;
assign n_18098 = n_18074 ^ n_18021;
assign n_18099 = n_18075 ^ n_18022;
assign n_18100 = n_18076 ^ n_17914;
assign n_18101 = n_18076 ^ n_17878;
assign n_18102 = n_18077 ^ n_17959;
assign n_18103 = n_18077 ^ n_17926;
assign n_18104 = n_18078 ^ n_17888;
assign n_18105 = n_18078 ^ n_17836;
assign n_18106 = n_18079 ^ n_17965;
assign n_18107 = n_18079 ^ n_17932;
assign n_18108 = n_18080 ^ n_17884;
assign n_18109 = n_18080 ^ n_17832;
assign n_18110 = n_18081 ^ n_12519;
assign n_18111 = ~n_17862 & n_18082;
assign n_18112 = n_18083 ^ n_12520;
assign n_18113 = ~n_17864 & n_18084;
assign n_18114 = n_18085 ^ n_12521;
assign n_18115 = n_17714 & ~n_18086;
assign n_18116 = n_18087 ^ n_12964;
assign n_18117 = n_17868 & ~n_18088;
assign n_18118 = n_18089 ^ n_14165;
assign n_18119 = n_17870 & ~n_18090;
assign n_18120 = n_18091 ^ n_15301;
assign n_18121 = ~n_17821 & n_18092;
assign n_18122 = n_18094 ^ n_18045;
assign n_18123 = n_18095 & n_18096;
assign n_18124 = ~n_17838 & n_18097;
assign n_18125 = n_18098 ^ n_17899;
assign n_18126 = n_18098 ^ n_17858;
assign n_18127 = n_18099 ^ n_17882;
assign n_18128 = n_18099 ^ n_17830;
assign n_18129 = n_18100 ^ n_12783;
assign n_18130 = ~n_17914 & n_18101;
assign n_18131 = n_18102 ^ n_12659;
assign n_18132 = ~n_17959 & n_18103;
assign n_18133 = n_18104 ^ n_12663;
assign n_18134 = n_17888 & ~n_18105;
assign n_18135 = n_18106 ^ n_12664;
assign n_18136 = ~n_17965 & n_18107;
assign n_18137 = n_18108 ^ n_12658;
assign n_18138 = ~n_17884 & n_18109;
assign n_18139 = n_18111 ^ n_18062;
assign n_18140 = n_18113 ^ n_18063;
assign n_18141 = n_18115 ^ n_18064;
assign n_18142 = n_18117 ^ n_18065;
assign n_18143 = n_18119 ^ n_18066;
assign n_18144 = n_18121 ^ n_18067;
assign n_18145 = n_18122 ^ n_17972;
assign n_18146 = n_18122 ^ n_17940;
assign n_18147 = n_18124 ^ n_18072;
assign n_18148 = n_18125 ^ n_12657;
assign n_18149 = ~n_17899 & n_18126;
assign y37 = n_18127;
assign n_18150 = ~n_17882 & n_18128;
assign n_18151 = n_18130 ^ n_18076;
assign n_18152 = n_18132 ^ n_18077;
assign n_18153 = n_18134 ^ n_18078;
assign n_18154 = n_18136 ^ n_18079;
assign n_18155 = n_18138 ^ n_18080;
assign n_18156 = n_18139 ^ n_17961;
assign n_18157 = n_18139 ^ n_17928;
assign n_18158 = n_18140 ^ n_17963;
assign n_18159 = n_18140 ^ n_17930;
assign n_18160 = n_18141 ^ n_17886;
assign n_18161 = n_18141 ^ n_17834;
assign n_18162 = n_18142 ^ n_17967;
assign n_18163 = n_18142 ^ n_17934;
assign n_18164 = n_18143 ^ n_17969;
assign n_18165 = n_18143 ^ n_17936;
assign n_18166 = n_18144 ^ n_17938;
assign n_18167 = n_18144 ^ n_17907;
assign n_18168 = n_18145 ^ n_17066;
assign n_18169 = n_17972 & ~n_18146;
assign n_18170 = n_18147 ^ n_17954;
assign n_18171 = ~n_17890 & ~n_18147;
assign n_18172 = n_18147 ^ n_17890;
assign n_18173 = n_18149 ^ n_18098;
assign n_18174 = n_18150 ^ n_18099;
assign n_18175 = n_18151 ^ n_17998;
assign n_18176 = n_18151 ^ n_17974;
assign n_18177 = n_18152 ^ n_18033;
assign n_18178 = n_18152 ^ n_18006;
assign n_18179 = n_18153 ^ n_17984;
assign n_18180 = n_18153 ^ n_17952;
assign n_18181 = n_18154 ^ n_18039;
assign n_18182 = n_18154 ^ n_18012;
assign n_18183 = n_18155 ^ n_17980;
assign n_18184 = n_18155 ^ n_17948;
assign n_18185 = n_18156 ^ n_12660;
assign n_18186 = ~n_17961 & n_18157;
assign n_18187 = n_18158 ^ n_12661;
assign n_18188 = ~n_17963 & n_18159;
assign n_18189 = n_18160 ^ n_12662;
assign n_18190 = ~n_17886 & n_18161;
assign n_18191 = n_18162 ^ n_13641;
assign n_18192 = n_17967 & ~n_18163;
assign n_18193 = n_18164 ^ n_14789;
assign n_18194 = n_17969 & ~n_18165;
assign n_18195 = n_18166 ^ n_16052;
assign n_18196 = ~n_17938 & n_18167;
assign n_18197 = n_18169 ^ n_18122;
assign n_18198 = n_17525 ^ n_18171;
assign n_18199 = n_18171 & ~n_17613;
assign n_18200 = ~n_18171 & ~n_17704;
assign n_18201 = n_18171 ^ n_18172;
assign n_18202 = n_18173 ^ n_17987;
assign n_18203 = n_18173 ^ n_17957;
assign n_18204 = n_18174 ^ n_17978;
assign n_18205 = n_18174 ^ n_17946;
assign n_18206 = n_18175 ^ n_12919;
assign n_18207 = ~n_17998 & n_18176;
assign n_18208 = n_18177 ^ n_12801;
assign n_18209 = ~n_18033 & n_18178;
assign n_18210 = n_18179 ^ n_12805;
assign n_18211 = ~n_17984 & n_18180;
assign n_18212 = n_18181 ^ n_12806;
assign n_18213 = ~n_18039 & n_18182;
assign n_18214 = n_18183 ^ n_12800;
assign n_18215 = n_17980 & ~n_18184;
assign n_18216 = n_18186 ^ n_18139;
assign n_18217 = n_18188 ^ n_18140;
assign n_18218 = n_18190 ^ n_18141;
assign n_18219 = n_18192 ^ n_18142;
assign n_18220 = n_18194 ^ n_18143;
assign n_18221 = n_18196 ^ n_18144;
assign n_18222 = n_18197 ^ n_18070;
assign n_18223 = ~n_18201 & n_17525;
assign n_18224 = n_17613 ^ n_18201;
assign n_18225 = n_18201 & ~n_17613;
assign n_18226 = n_18201 & n_17614;
assign n_18227 = n_18202 ^ n_12799;
assign n_18228 = ~n_17987 & n_18203;
assign y38 = n_18204;
assign n_18229 = ~n_17978 & n_18205;
assign n_18230 = n_18207 ^ n_18151;
assign n_18231 = n_18209 ^ n_18152;
assign n_18232 = n_18211 ^ n_18153;
assign n_18233 = n_18213 ^ n_18154;
assign n_18234 = n_18215 ^ n_18155;
assign n_18235 = n_18216 ^ n_18035;
assign n_18236 = n_18216 ^ n_18008;
assign n_18237 = n_18217 ^ n_18037;
assign n_18238 = n_18217 ^ n_18010;
assign n_18239 = n_18218 ^ n_17982;
assign n_18240 = n_18218 ^ n_17950;
assign n_18241 = n_18219 ^ n_18041;
assign n_18242 = n_18219 ^ n_18014;
assign n_18243 = n_18220 ^ n_18043;
assign n_18244 = n_18220 ^ n_18016;
assign n_18245 = n_18221 ^ n_18018;
assign n_18246 = n_18221 ^ n_17995;
assign n_18247 = n_18225 ^ n_17614;
assign n_18248 = n_18228 ^ n_18173;
assign n_18249 = n_18229 ^ n_18174;
assign n_18250 = n_18230 ^ n_18073;
assign n_18251 = n_18230 ^ n_18048;
assign n_18252 = n_18231 ^ n_18110;
assign n_18253 = n_18231 ^ n_18081;
assign n_18254 = n_18232 ^ n_18058;
assign n_18255 = n_18232 ^ n_18029;
assign n_18256 = n_18233 ^ n_18116;
assign n_18257 = n_18233 ^ n_18087;
assign n_18258 = n_18234 ^ n_18054;
assign n_18259 = n_18234 ^ n_18025;
assign n_18260 = n_18235 ^ n_12802;
assign n_18261 = ~n_18035 & n_18236;
assign n_18262 = n_18237 ^ n_12803;
assign n_18263 = ~n_18037 & n_18238;
assign n_18264 = n_18239 ^ n_12804;
assign n_18265 = ~n_17982 & n_18240;
assign n_18266 = n_18241 ^ n_14472;
assign n_18267 = ~n_18041 & n_18242;
assign n_18268 = n_18243 ^ n_15545;
assign n_18269 = n_18043 & ~n_18244;
assign n_18270 = n_18245 ^ n_16862;
assign n_18271 = ~n_18018 & n_18246;
assign n_18272 = n_18248 ^ n_18060;
assign n_18273 = n_18248 ^ n_18031;
assign n_18274 = n_18249 ^ n_18052;
assign n_18275 = n_18249 ^ n_18023;
assign n_18276 = n_18250 ^ n_13064;
assign n_18277 = n_18073 & ~n_18251;
assign n_18278 = n_18252 ^ n_12959;
assign n_18279 = ~n_18110 & n_18253;
assign n_18280 = n_18254 ^ n_12963;
assign n_18281 = ~n_18058 & n_18255;
assign n_18282 = n_18256 ^ n_13466;
assign n_18283 = n_18116 & ~n_18257;
assign n_18284 = n_18258 ^ n_12958;
assign n_18285 = n_18054 & ~n_18259;
assign n_18286 = n_18261 ^ n_18216;
assign n_18287 = n_18263 ^ n_18217;
assign n_18288 = n_18265 ^ n_18218;
assign n_18289 = n_18267 ^ n_18219;
assign n_18290 = n_18269 ^ n_18220;
assign n_18291 = n_18271 ^ n_18221;
assign n_18292 = n_18272 ^ n_12957;
assign n_18293 = ~n_18060 & n_18273;
assign y39 = n_18274;
assign n_18294 = ~n_18052 & n_18275;
assign n_18295 = n_18277 ^ n_18230;
assign n_18296 = n_18279 ^ n_18231;
assign n_18297 = n_18281 ^ n_18232;
assign n_18298 = n_18283 ^ n_18233;
assign n_18299 = n_18285 ^ n_18234;
assign n_18300 = n_18286 ^ n_18112;
assign n_18301 = n_18286 ^ n_18083;
assign n_18302 = n_18287 ^ n_18114;
assign n_18303 = n_18287 ^ n_18085;
assign n_18304 = n_18288 ^ n_18056;
assign n_18305 = n_18288 ^ n_18027;
assign n_18306 = n_18289 ^ n_18118;
assign n_18307 = n_18289 ^ n_18089;
assign n_18308 = n_18290 ^ n_18120;
assign n_18309 = n_18290 ^ n_18091;
assign n_18310 = n_18291 ^ n_18093;
assign n_18311 = n_18291 ^ n_18068;
assign n_18312 = n_18293 ^ n_18248;
assign n_18313 = n_18294 ^ n_18249;
assign n_18314 = n_18295 ^ n_18148;
assign n_18315 = n_18295 ^ n_18125;
assign n_18316 = n_18296 ^ n_18185;
assign n_18317 = n_18296 ^ n_18156;
assign n_18318 = n_18297 ^ n_18135;
assign n_18319 = n_18297 ^ n_18106;
assign n_18320 = n_18298 ^ n_18191;
assign n_18321 = n_18298 ^ n_18162;
assign n_18322 = n_18299 ^ n_18131;
assign n_18323 = n_18299 ^ n_18102;
assign n_18324 = n_18300 ^ n_12960;
assign n_18325 = ~n_18112 & n_18301;
assign n_18326 = n_18302 ^ n_12961;
assign n_18327 = n_18114 & ~n_18303;
assign n_18328 = n_18304 ^ n_12962;
assign n_18329 = n_18056 & ~n_18305;
assign n_18330 = n_18306 ^ n_14640;
assign n_18331 = n_18118 & ~n_18307;
assign n_18332 = n_18308 ^ n_15691;
assign n_18333 = ~n_18120 & n_18309;
assign n_18334 = n_18310 ^ n_17045;
assign n_18335 = ~n_18093 & n_18311;
assign n_18336 = n_18312 ^ n_18137;
assign n_18337 = n_18312 ^ n_18108;
assign n_18338 = n_18313 ^ n_18129;
assign n_18339 = n_18313 ^ n_18100;
assign n_18340 = n_18314 ^ n_13200;
assign n_18341 = ~n_18148 & n_18315;
assign n_18342 = n_18316 ^ n_13121;
assign n_18343 = ~n_18185 & n_18317;
assign n_18344 = n_18318 ^ n_13125;
assign n_18345 = ~n_18135 & n_18319;
assign n_18346 = n_18320 ^ n_14319;
assign n_18347 = n_18191 & ~n_18321;
assign n_18348 = n_18322 ^ n_13120;
assign n_18349 = ~n_18131 & n_18323;
assign n_18350 = n_18325 ^ n_18286;
assign n_18351 = n_18327 ^ n_18287;
assign n_18352 = n_18329 ^ n_18288;
assign n_18353 = n_18331 ^ n_18289;
assign n_18354 = n_18333 ^ n_18290;
assign n_18355 = n_18335 ^ n_18291;
assign n_18356 = n_18336 ^ n_13119;
assign n_18357 = ~n_18137 & n_18337;
assign y40 = n_18338;
assign n_18358 = ~n_18129 & n_18339;
assign n_18359 = n_18341 ^ n_18295;
assign n_18360 = n_18343 ^ n_18296;
assign n_18361 = n_18345 ^ n_18297;
assign n_18362 = n_18347 ^ n_18298;
assign n_18363 = n_18349 ^ n_18299;
assign n_18364 = n_18350 ^ n_18187;
assign n_18365 = n_18350 ^ n_18158;
assign n_18366 = n_18351 ^ n_18189;
assign n_18367 = n_18351 ^ n_18160;
assign n_18368 = n_18352 ^ n_18133;
assign n_18369 = n_18352 ^ n_18104;
assign n_18370 = n_18353 ^ n_18193;
assign n_18371 = n_18353 ^ n_18164;
assign n_18372 = n_18354 ^ n_18195;
assign n_18373 = n_18354 ^ n_18166;
assign n_18374 = n_18355 ^ n_18168;
assign n_18375 = n_18355 ^ n_18145;
assign n_18376 = n_18357 ^ n_18312;
assign n_18377 = n_18358 ^ n_18313;
assign n_18378 = n_18359 ^ n_18227;
assign n_18379 = n_18359 ^ n_18202;
assign n_18380 = n_18360 ^ n_18260;
assign n_18381 = n_18360 ^ n_18235;
assign n_18382 = n_18361 ^ n_18212;
assign n_18383 = n_18361 ^ n_18181;
assign n_18384 = n_18362 ^ n_18266;
assign n_18385 = n_18362 ^ n_18241;
assign n_18386 = n_18363 ^ n_18208;
assign n_18387 = n_18363 ^ n_18177;
assign n_18388 = n_18364 ^ n_13122;
assign n_18389 = ~n_18187 & n_18365;
assign n_18390 = n_18366 ^ n_13123;
assign n_18391 = ~n_18189 & n_18367;
assign n_18392 = n_18368 ^ n_13124;
assign n_18393 = n_18133 & ~n_18369;
assign n_18394 = n_18370 ^ n_15259;
assign n_18395 = n_18193 & ~n_18371;
assign n_18396 = n_18372 ^ n_16615;
assign n_18397 = ~n_18195 & n_18373;
assign n_18398 = n_18168 & ~n_18375;
assign n_18399 = n_18376 ^ n_18214;
assign n_18400 = n_18376 ^ n_18183;
assign n_18401 = n_18377 ^ n_18206;
assign n_18402 = n_18377 ^ n_18175;
assign n_18403 = n_18378 ^ n_13419;
assign n_18404 = ~n_18227 & n_18379;
assign n_18405 = n_18380 ^ n_13294;
assign n_18406 = ~n_18260 & n_18381;
assign n_18407 = n_18382 ^ n_13298;
assign n_18408 = ~n_18212 & n_18383;
assign n_18409 = n_18384 ^ n_14951;
assign n_18410 = ~n_18266 & n_18385;
assign n_18411 = n_18386 ^ n_13293;
assign n_18412 = ~n_18208 & n_18387;
assign n_18413 = n_18389 ^ n_18350;
assign n_18414 = n_18391 ^ n_18351;
assign n_18415 = n_18393 ^ n_18352;
assign n_18416 = n_18395 ^ n_18353;
assign n_18417 = n_18397 ^ n_18354;
assign n_18418 = n_18398 ^ n_18355;
assign n_18419 = n_18399 ^ n_13292;
assign n_18420 = n_18214 & ~n_18400;
assign y41 = n_18401;
assign n_18421 = ~n_18206 & n_18402;
assign n_18422 = n_18404 ^ n_18359;
assign n_18423 = n_18406 ^ n_18360;
assign n_18424 = n_18408 ^ n_18361;
assign n_18425 = n_18410 ^ n_18362;
assign n_18426 = n_18412 ^ n_18363;
assign n_18427 = n_18413 ^ n_18262;
assign n_18428 = n_18413 ^ n_18237;
assign n_18429 = n_18414 ^ n_18264;
assign n_18430 = n_18414 ^ n_18239;
assign n_18431 = n_18415 ^ n_18210;
assign n_18432 = n_18415 ^ n_18179;
assign n_18433 = n_18416 ^ n_18268;
assign n_18434 = n_18416 ^ n_18243;
assign n_18435 = n_18417 ^ n_18270;
assign n_18436 = n_18417 ^ n_18245;
assign n_18437 = n_18418 ^ n_18222;
assign n_18438 = n_18418 ^ n_18197;
assign n_18439 = n_18197 & n_18418;
assign n_18440 = n_18420 ^ n_18376;
assign n_18441 = n_18421 ^ n_18377;
assign n_18442 = n_18422 ^ n_18292;
assign n_18443 = n_18422 ^ n_18272;
assign n_18444 = n_18423 ^ n_18324;
assign n_18445 = n_18423 ^ n_18300;
assign n_18446 = n_18424 ^ n_18282;
assign n_18447 = n_18424 ^ n_18256;
assign n_18448 = n_18425 ^ n_18330;
assign n_18449 = n_18425 ^ n_18306;
assign n_18450 = n_18426 ^ n_18278;
assign n_18451 = n_18426 ^ n_18252;
assign n_18452 = n_18427 ^ n_13295;
assign n_18453 = ~n_18262 & n_18428;
assign n_18454 = n_18429 ^ n_13296;
assign n_18455 = ~n_18264 & n_18430;
assign n_18456 = n_18431 ^ n_13297;
assign n_18457 = ~n_18210 & n_18432;
assign n_18458 = n_18433 ^ n_16242;
assign n_18459 = n_18268 & ~n_18434;
assign n_18460 = n_18435 ^ n_16942;
assign n_18461 = ~n_18270 & n_18436;
assign n_18462 = n_18437 ^ n_18197;
assign n_18463 = n_18439 ^ n_18438;
assign n_18464 = n_18095 & n_18439;
assign n_18465 = n_18440 ^ n_18284;
assign n_18466 = n_18440 ^ n_18258;
assign n_18467 = n_18441 ^ n_18276;
assign n_18468 = n_18441 ^ n_18250;
assign n_18469 = n_18442 ^ n_13538;
assign n_18470 = ~n_18292 & n_18443;
assign n_18471 = n_18444 ^ n_13462;
assign n_18472 = ~n_18324 & n_18445;
assign n_18473 = n_18446 ^ n_14164;
assign n_18474 = n_18282 & ~n_18447;
assign n_18475 = n_18448 ^ n_15300;
assign n_18476 = n_18330 & ~n_18449;
assign n_18477 = n_18450 ^ n_13461;
assign n_18478 = ~n_18278 & n_18451;
assign n_18479 = n_18453 ^ n_18413;
assign n_18480 = n_18455 ^ n_18414;
assign n_18481 = n_18457 ^ n_18415;
assign n_18482 = n_18459 ^ n_18416;
assign n_18483 = n_18461 ^ n_18417;
assign n_18484 = n_18462 & ~n_18438;
assign n_18485 = n_18463 ^ n_18096;
assign n_18486 = n_18464 ^ n_18096;
assign n_18487 = n_18465 ^ n_13460;
assign n_18488 = n_18284 & ~n_18466;
assign y42 = ~n_18467;
assign n_18489 = n_18276 & ~n_18468;
assign n_18490 = n_18470 ^ n_18422;
assign n_18491 = n_18472 ^ n_18423;
assign n_18492 = n_18474 ^ n_18424;
assign n_18493 = n_18476 ^ n_18425;
assign n_18494 = n_18478 ^ n_18426;
assign n_18495 = n_18479 ^ n_18326;
assign n_18496 = n_18479 ^ n_18302;
assign n_18497 = n_18480 ^ n_18328;
assign n_18498 = n_18480 ^ n_18304;
assign n_18499 = n_18481 ^ n_18280;
assign n_18500 = n_18481 ^ n_18254;
assign n_18501 = n_18482 ^ n_18332;
assign n_18502 = n_18482 ^ n_18308;
assign n_18503 = n_18483 ^ n_18334;
assign n_18504 = n_18483 ^ n_18310;
assign n_18505 = ~n_18071 & n_18485;
assign n_18506 = n_18488 ^ n_18440;
assign n_18507 = n_18489 ^ n_18441;
assign n_18508 = n_18490 ^ n_18356;
assign n_18509 = n_18490 ^ n_18336;
assign n_18510 = n_18491 ^ n_18388;
assign n_18511 = n_18491 ^ n_18364;
assign n_18512 = n_18492 ^ n_18346;
assign n_18513 = n_18492 ^ n_18320;
assign n_18514 = n_18493 ^ n_18394;
assign n_18515 = n_18493 ^ n_18370;
assign n_18516 = n_18494 ^ n_18342;
assign n_18517 = n_18494 ^ n_18316;
assign n_18518 = n_18495 ^ n_13463;
assign n_18519 = n_18326 & ~n_18496;
assign n_18520 = n_18497 ^ n_13464;
assign n_18521 = n_18328 & ~n_18498;
assign n_18522 = n_18499 ^ n_13465;
assign n_18523 = ~n_18280 & n_18500;
assign n_18524 = n_18501 ^ n_16343;
assign n_18525 = ~n_18332 & n_18502;
assign n_18526 = ~n_18334 & n_18504;
assign n_18527 = n_18506 ^ n_18348;
assign n_18528 = n_18506 ^ n_18322;
assign n_18529 = n_18507 ^ n_18340;
assign n_18530 = n_18507 ^ n_18314;
assign n_18531 = n_18508 ^ n_13790;
assign n_18532 = ~n_18356 & n_18509;
assign n_18533 = n_18510 ^ n_13637;
assign n_18534 = ~n_18388 & n_18511;
assign n_18535 = n_18512 ^ n_14788;
assign n_18536 = n_18346 & ~n_18513;
assign n_18537 = n_18514 ^ n_16051;
assign n_18538 = n_18394 & ~n_18515;
assign n_18539 = n_18516 ^ n_13636;
assign n_18540 = ~n_18342 & n_18517;
assign n_18541 = n_18519 ^ n_18479;
assign n_18542 = n_18521 ^ n_18480;
assign n_18543 = n_18523 ^ n_18481;
assign n_18544 = n_18525 ^ n_18482;
assign n_18545 = n_18526 ^ n_18483;
assign n_18546 = n_18527 ^ n_13635;
assign n_18547 = ~n_18348 & n_18528;
assign y43 = n_18529;
assign n_18548 = ~n_18340 & n_18530;
assign n_18549 = n_18532 ^ n_18490;
assign n_18550 = n_18534 ^ n_18491;
assign n_18551 = n_18536 ^ n_18492;
assign n_18552 = n_18538 ^ n_18493;
assign n_18553 = n_18540 ^ n_18494;
assign n_18554 = n_18541 ^ n_18390;
assign n_18555 = n_18541 ^ n_18366;
assign n_18556 = n_18542 ^ n_18392;
assign n_18557 = n_18542 ^ n_18368;
assign n_18558 = n_18543 ^ n_18344;
assign n_18559 = n_18543 ^ n_18318;
assign n_18560 = n_18544 ^ n_18396;
assign n_18561 = n_18544 ^ n_18372;
assign n_18562 = n_18545 ^ n_18374;
assign n_18563 = n_18547 ^ n_18506;
assign n_18564 = n_18548 ^ n_18507;
assign n_18565 = n_18549 ^ n_18419;
assign n_18566 = n_18549 ^ n_18399;
assign n_18567 = n_18550 ^ n_18452;
assign n_18568 = n_18550 ^ n_18427;
assign n_18569 = n_18551 ^ n_18409;
assign n_18570 = n_18551 ^ n_18384;
assign n_18571 = n_18552 ^ n_18458;
assign n_18572 = n_18552 ^ n_18433;
assign n_18573 = n_18553 ^ n_18405;
assign n_18574 = n_18553 ^ n_18380;
assign n_18575 = n_18554 ^ n_13638;
assign n_18576 = ~n_18390 & n_18555;
assign n_18577 = n_18556 ^ n_13639;
assign n_18578 = n_18392 & ~n_18557;
assign n_18579 = n_18558 ^ n_13640;
assign n_18580 = ~n_18344 & n_18559;
assign n_18581 = n_18560 ^ n_17065;
assign n_18582 = ~n_18396 & n_18561;
assign n_18583 = n_18563 ^ n_18411;
assign n_18584 = n_18563 ^ n_18386;
assign n_18585 = n_18564 ^ n_18403;
assign n_18586 = n_18564 ^ n_18378;
assign n_18587 = n_18565 ^ n_14135;
assign n_18588 = n_18419 & ~n_18566;
assign n_18589 = n_18567 ^ n_14026;
assign n_18590 = ~n_18452 & n_18568;
assign n_18591 = n_18569 ^ n_15544;
assign n_18592 = ~n_18409 & n_18570;
assign n_18593 = n_18571 ^ n_16861;
assign n_18594 = n_18458 & ~n_18572;
assign n_18595 = n_18573 ^ n_14025;
assign n_18596 = ~n_18405 & n_18574;
assign n_18597 = n_18576 ^ n_18541;
assign n_18598 = n_18578 ^ n_18542;
assign n_18599 = n_18580 ^ n_18543;
assign n_18600 = n_18582 ^ n_18544;
assign n_18601 = n_18583 ^ n_14024;
assign n_18602 = ~n_18411 & n_18584;
assign y44 = n_18585;
assign n_18603 = ~n_18403 & n_18586;
assign n_18604 = n_18588 ^ n_18549;
assign n_18605 = n_18590 ^ n_18550;
assign n_18606 = n_18592 ^ n_18551;
assign n_18607 = n_18594 ^ n_18552;
assign n_18608 = n_18596 ^ n_18553;
assign n_18609 = n_18597 ^ n_18454;
assign n_18610 = n_18597 ^ n_18429;
assign n_18611 = n_18598 ^ n_18456;
assign n_18612 = n_18598 ^ n_18431;
assign n_18613 = n_18599 ^ n_18407;
assign n_18614 = n_18599 ^ n_18382;
assign n_18615 = n_18600 ^ n_18460;
assign n_18616 = n_18600 ^ n_18435;
assign n_18617 = n_18602 ^ n_18563;
assign n_18618 = n_18603 ^ n_18564;
assign n_18619 = n_18604 ^ n_18487;
assign n_18620 = n_18604 ^ n_18465;
assign n_18621 = n_18605 ^ n_18518;
assign n_18622 = n_18605 ^ n_18495;
assign n_18623 = n_18606 ^ n_18475;
assign n_18624 = n_18606 ^ n_18448;
assign n_18625 = n_18607 ^ n_18524;
assign n_18626 = n_18607 ^ n_18501;
assign n_18627 = n_18471 ^ n_18608;
assign n_18628 = n_13462 ^ n_18608;
assign n_18629 = n_18609 ^ n_14027;
assign n_18630 = ~n_18454 & n_18610;
assign n_18631 = n_18611 ^ n_14028;
assign n_18632 = ~n_18456 & n_18612;
assign n_18633 = n_18613 ^ n_14029;
assign n_18634 = ~n_18407 & n_18614;
assign n_18635 = ~n_18460 & n_18616;
assign n_18636 = n_18617 ^ n_18477;
assign n_18637 = n_18617 ^ n_18450;
assign n_18638 = n_18618 ^ n_18469;
assign n_18639 = n_18618 ^ n_18442;
assign n_18640 = n_18619 ^ n_14300;
assign n_18641 = n_18487 & ~n_18620;
assign n_18642 = n_18621 ^ n_14161;
assign n_18643 = n_18518 & ~n_18622;
assign n_18644 = n_18623 ^ n_15690;
assign n_18645 = n_18475 & ~n_18624;
assign n_18646 = n_18625 ^ n_17044;
assign n_18647 = ~n_18524 & n_18626;
assign n_18648 = n_18627 ^ n_14160;
assign n_18649 = ~n_18471 & n_18628;
assign n_18650 = n_18630 ^ n_18597;
assign n_18651 = n_18632 ^ n_18598;
assign n_18652 = n_18634 ^ n_18599;
assign n_18653 = n_18635 ^ n_18600;
assign n_18654 = n_18636 ^ n_14159;
assign n_18655 = ~n_18477 & n_18637;
assign y45 = n_18638;
assign n_18656 = ~n_18469 & n_18639;
assign n_18657 = n_18641 ^ n_18604;
assign n_18658 = n_18643 ^ n_18605;
assign n_18659 = n_18645 ^ n_18606;
assign n_18660 = n_18647 ^ n_18607;
assign n_18661 = n_18649 ^ n_18608;
assign n_18662 = n_18650 ^ n_18520;
assign n_18663 = n_18650 ^ n_18497;
assign n_18664 = n_18651 ^ n_18522;
assign n_18665 = n_18651 ^ n_18499;
assign n_18666 = n_18652 ^ n_18473;
assign n_18667 = n_18652 ^ n_18446;
assign n_18668 = n_18653 ^ n_18503;
assign n_18669 = n_18655 ^ n_18617;
assign n_18670 = n_18656 ^ n_18618;
assign n_18671 = n_18657 ^ n_18546;
assign n_18672 = n_18657 ^ n_18527;
assign n_18673 = n_18658 ^ n_18575;
assign n_18674 = n_18658 ^ n_18554;
assign n_18675 = n_18659 ^ n_18537;
assign n_18676 = n_18659 ^ n_16051;
assign n_18677 = n_18660 ^ n_18581;
assign n_18678 = n_18660 ^ n_18560;
assign n_18679 = n_18661 ^ n_18533;
assign n_18680 = n_18661 ^ n_18510;
assign n_18681 = n_18662 ^ n_14162;
assign n_18682 = n_18520 & ~n_18663;
assign n_18683 = n_18664 ^ n_14163;
assign n_18684 = ~n_18522 & n_18665;
assign n_18685 = n_18666 ^ n_14639;
assign n_18686 = n_18473 & ~n_18667;
assign n_18687 = n_18669 ^ n_18539;
assign n_18688 = n_18669 ^ n_18516;
assign n_18689 = n_18670 ^ n_18531;
assign n_18690 = n_18670 ^ n_18508;
assign n_18691 = n_18671 ^ n_14447;
assign n_18692 = ~n_18546 & n_18672;
assign n_18693 = n_18673 ^ n_14316;
assign n_18694 = ~n_18575 & n_18674;
assign n_18695 = n_18675 ^ n_16614;
assign n_18696 = ~n_18537 & ~n_18676;
assign n_18697 = ~n_18581 & n_18678;
assign n_18698 = n_18679 ^ n_14315;
assign n_18699 = ~n_18533 & n_18680;
assign n_18700 = n_18682 ^ n_18650;
assign n_18701 = n_18684 ^ n_18651;
assign n_18702 = n_18686 ^ n_18652;
assign n_18703 = n_18687 ^ n_14314;
assign n_18704 = ~n_18539 & n_18688;
assign y46 = n_18689;
assign n_18705 = ~n_18531 & n_18690;
assign n_18706 = n_18692 ^ n_18657;
assign n_18707 = n_18694 ^ n_18658;
assign n_18708 = n_18696 ^ n_18514;
assign n_18709 = n_18697 ^ n_18660;
assign n_18710 = n_18699 ^ n_18661;
assign n_18711 = n_18700 ^ n_18577;
assign n_18712 = n_18700 ^ n_18556;
assign n_18713 = n_18701 ^ n_18579;
assign n_18714 = n_18701 ^ n_18558;
assign n_18715 = n_18702 ^ n_18535;
assign n_18716 = n_18702 ^ n_18512;
assign n_18717 = n_18704 ^ n_18669;
assign n_18718 = n_18705 ^ n_18670;
assign n_18719 = n_18706 ^ n_18601;
assign n_18720 = n_18706 ^ n_18583;
assign n_18721 = n_18707 ^ n_18629;
assign n_18722 = n_18707 ^ n_18609;
assign n_18723 = n_18708 ^ n_18593;
assign n_18724 = n_18708 ^ n_18571;
assign n_18725 = n_18709 ^ n_18615;
assign n_18726 = n_18710 ^ n_18589;
assign n_18727 = n_18710 ^ n_18567;
assign n_18728 = n_18711 ^ n_14317;
assign n_18729 = n_18577 & ~n_18712;
assign n_18730 = n_18713 ^ n_14318;
assign n_18731 = ~n_18579 & n_18714;
assign n_18732 = n_18715 ^ n_15258;
assign n_18733 = n_18535 & ~n_18716;
assign n_18734 = n_18717 ^ n_18595;
assign n_18735 = n_18717 ^ n_18573;
assign n_18736 = n_18718 ^ n_18587;
assign n_18737 = n_18718 ^ n_18565;
assign n_18738 = n_18719 ^ n_14613;
assign n_18739 = ~n_18601 & n_18720;
assign n_18740 = n_18721 ^ n_14469;
assign n_18741 = ~n_18629 & n_18722;
assign n_18742 = n_18723 ^ n_16941;
assign n_18743 = n_16941 & n_18723;
assign n_18744 = n_18593 & n_18724;
assign n_18745 = n_18726 ^ n_14468;
assign n_18746 = ~n_18589 & n_18727;
assign n_18747 = n_18729 ^ n_18700;
assign n_18748 = n_18731 ^ n_18701;
assign n_18749 = n_18733 ^ n_18702;
assign n_18750 = n_18734 ^ n_14467;
assign n_18751 = ~n_18595 & n_18735;
assign y47 = ~n_18736;
assign n_18752 = n_18587 & ~n_18737;
assign n_18753 = n_18739 ^ n_18706;
assign n_18754 = n_18741 ^ n_18707;
assign n_18755 = n_18743 ^ n_18742;
assign n_18756 = n_18744 ^ n_18708;
assign n_18757 = n_18746 ^ n_18710;
assign n_18758 = n_18747 ^ n_18631;
assign n_18759 = n_18747 ^ n_18611;
assign n_18760 = n_18748 ^ n_18633;
assign n_18761 = n_18748 ^ n_18613;
assign n_18762 = n_18749 ^ n_18591;
assign n_18763 = n_18749 ^ n_18569;
assign n_18764 = n_18751 ^ n_18717;
assign n_18765 = n_18752 ^ n_18718;
assign n_18766 = n_18753 ^ n_18654;
assign n_18767 = n_18753 ^ n_18636;
assign n_18768 = n_18754 ^ n_18681;
assign n_18769 = n_18754 ^ n_18662;
assign n_18770 = n_18756 ^ n_18646;
assign n_18771 = n_18756 ^ n_17044;
assign n_18772 = n_18757 ^ n_18642;
assign n_18773 = n_18757 ^ n_18621;
assign n_18774 = n_18758 ^ n_14470;
assign n_18775 = ~n_18631 & n_18759;
assign n_18776 = n_18760 ^ n_14471;
assign n_18777 = ~n_18633 & n_18761;
assign n_18778 = n_18762 ^ n_16241;
assign n_18779 = ~n_18591 & n_18763;
assign n_18780 = n_18764 ^ n_18648;
assign n_18781 = n_18764 ^ n_18627;
assign n_18782 = n_18765 ^ n_18640;
assign n_18783 = n_18765 ^ n_18619;
assign n_18784 = n_18766 ^ n_14773;
assign n_18785 = ~n_18654 & n_18767;
assign n_18786 = n_18768 ^ n_14637;
assign n_18787 = n_18681 & ~n_18769;
assign n_18788 = n_18646 & n_18771;
assign n_18789 = n_18772 ^ n_14636;
assign n_18790 = n_18642 & ~n_18773;
assign n_18791 = n_18775 ^ n_18747;
assign n_18792 = n_18777 ^ n_18748;
assign n_18793 = n_18779 ^ n_18749;
assign n_18794 = n_18780 ^ n_14635;
assign n_18795 = ~n_18648 & n_18781;
assign y48 = ~n_18782;
assign n_18796 = n_18640 & ~n_18783;
assign n_18797 = n_18785 ^ n_18753;
assign n_18798 = n_18787 ^ n_18754;
assign n_18799 = n_18788 ^ n_18625;
assign n_18800 = n_18790 ^ n_18757;
assign n_18801 = n_18791 ^ n_18683;
assign n_18802 = n_18791 ^ n_18664;
assign n_18803 = n_18792 ^ n_18685;
assign n_18804 = n_18792 ^ n_18666;
assign n_18805 = n_18793 ^ n_18644;
assign n_18806 = n_18793 ^ n_18623;
assign n_18807 = n_18795 ^ n_18764;
assign n_18808 = n_18796 ^ n_18765;
assign n_18809 = n_18797 ^ n_18703;
assign n_18810 = n_18797 ^ n_18687;
assign n_18811 = n_18798 ^ n_18728;
assign n_18812 = n_18798 ^ n_18711;
assign n_18813 = n_18799 ^ n_18677;
assign n_18814 = n_18800 ^ n_18693;
assign n_18815 = n_18800 ^ n_18673;
assign n_18816 = n_18801 ^ n_14638;
assign n_18817 = ~n_18683 & n_18802;
assign n_18818 = n_18803 ^ n_15299;
assign n_18819 = n_18685 & ~n_18804;
assign n_18820 = n_18805 ^ n_16342;
assign n_18821 = n_18644 & ~n_18806;
assign n_18822 = n_18807 ^ n_18698;
assign n_18823 = n_18807 ^ n_18679;
assign n_18824 = n_18808 ^ n_18691;
assign n_18825 = n_18808 ^ n_18671;
assign n_18826 = n_18809 ^ n_14939;
assign n_18827 = ~n_18703 & n_18810;
assign n_18828 = n_18811 ^ n_14786;
assign n_18829 = n_18728 & ~n_18812;
assign n_18830 = n_18814 ^ n_14785;
assign n_18831 = ~n_18693 & n_18815;
assign n_18832 = n_18817 ^ n_18791;
assign n_18833 = n_18819 ^ n_18792;
assign n_18834 = n_18821 ^ n_18793;
assign n_18835 = n_18822 ^ n_14784;
assign n_18836 = ~n_18698 & n_18823;
assign y49 = n_18824;
assign n_18837 = ~n_18691 & n_18825;
assign n_18838 = n_18827 ^ n_18797;
assign n_18839 = n_18829 ^ n_18798;
assign n_18840 = n_18831 ^ n_18800;
assign n_18841 = n_18832 ^ n_18730;
assign n_18842 = n_18832 ^ n_18713;
assign n_18843 = n_18833 ^ n_18732;
assign n_18844 = n_18833 ^ n_18715;
assign n_18845 = n_18834 ^ n_18695;
assign n_18846 = n_18834 ^ n_18675;
assign n_18847 = n_18836 ^ n_18807;
assign n_18848 = n_18837 ^ n_18808;
assign n_18849 = n_18838 ^ n_18750;
assign n_18850 = n_18838 ^ n_18734;
assign n_18851 = n_18839 ^ n_18774;
assign n_18852 = n_18839 ^ n_18758;
assign n_18853 = n_18840 ^ n_18740;
assign n_18854 = n_18840 ^ n_18721;
assign n_18855 = n_18841 ^ n_14787;
assign n_18856 = ~n_18730 & n_18842;
assign n_18857 = n_18843 ^ n_16050;
assign n_18858 = n_18732 & ~n_18844;
assign n_18859 = n_18845 ^ n_17064;
assign n_18860 = n_18695 & ~n_18846;
assign n_18861 = n_18847 ^ n_18745;
assign n_18862 = n_18847 ^ n_18726;
assign n_18863 = n_18848 ^ n_18738;
assign n_18864 = n_18848 ^ n_18719;
assign n_18865 = n_18849 ^ n_15079;
assign n_18866 = ~n_18750 & n_18850;
assign n_18867 = n_18851 ^ n_14949;
assign n_18868 = ~n_18774 & n_18852;
assign n_18869 = n_18853 ^ n_14948;
assign n_18870 = ~n_18740 & n_18854;
assign n_18871 = n_18856 ^ n_18832;
assign n_18872 = n_18858 ^ n_18833;
assign n_18873 = n_18860 ^ n_18834;
assign n_18874 = n_18861 ^ n_14947;
assign n_18875 = ~n_18745 & n_18862;
assign y50 = n_18863;
assign n_18876 = ~n_18738 & n_18864;
assign n_18877 = n_18866 ^ n_18838;
assign n_18878 = n_18868 ^ n_18839;
assign n_18879 = n_18870 ^ n_18840;
assign n_18880 = n_18871 ^ n_18776;
assign n_18881 = n_18871 ^ n_18760;
assign n_18882 = n_18872 ^ n_18778;
assign n_18883 = n_18872 ^ n_18762;
assign n_18884 = n_18873 ^ n_18742;
assign n_18885 = n_18873 & n_18743;
assign n_18886 = ~n_18873 & ~n_18755;
assign n_18887 = n_18875 ^ n_18847;
assign n_18888 = n_18876 ^ n_18848;
assign n_18889 = n_18877 ^ n_18794;
assign n_18890 = n_18877 ^ n_18780;
assign n_18891 = n_18878 ^ n_18816;
assign n_18892 = n_18878 ^ n_18801;
assign n_18893 = n_18879 ^ n_18786;
assign n_18894 = n_18879 ^ n_18768;
assign n_18895 = n_18880 ^ n_14950;
assign n_18896 = ~n_18776 & n_18881;
assign n_18897 = n_18882 ^ n_16860;
assign n_18898 = ~n_18778 & n_18883;
assign n_18899 = n_18770 & ~n_18885;
assign n_18900 = n_18885 ^ n_18886;
assign n_18901 = n_18887 ^ n_18789;
assign n_18902 = n_18887 ^ n_18772;
assign n_18903 = n_18888 ^ n_18784;
assign n_18904 = n_18888 ^ n_18766;
assign n_18905 = n_18889 ^ n_15253;
assign n_18906 = ~n_18794 & n_18890;
assign n_18907 = n_18891 ^ n_15298;
assign n_18908 = ~n_18816 & n_18892;
assign n_18909 = n_18893 ^ n_15297;
assign n_18910 = n_18786 & ~n_18894;
assign n_18911 = n_18896 ^ n_18871;
assign n_18912 = n_18898 ^ n_18872;
assign n_18913 = ~n_18886 & ~n_18899;
assign n_18914 = n_18900 ^ n_18742;
assign n_18915 = n_18901 ^ n_15296;
assign n_18916 = n_18789 & ~n_18902;
assign y51 = n_18903;
assign n_18917 = ~n_18784 & n_18904;
assign n_18918 = n_18906 ^ n_18877;
assign n_18919 = n_18908 ^ n_18878;
assign n_18920 = n_18910 ^ n_18879;
assign n_18921 = n_18911 ^ n_18818;
assign n_18922 = n_18911 ^ n_18803;
assign n_18923 = n_18912 ^ n_18820;
assign n_18924 = n_18912 ^ n_18805;
assign n_18925 = n_18914 ^ n_18873;
assign n_18926 = n_18916 ^ n_18887;
assign n_18927 = n_18917 ^ n_18888;
assign n_18928 = n_18918 ^ n_18835;
assign n_18929 = n_18918 ^ n_18822;
assign n_18930 = n_18919 ^ n_18855;
assign n_18931 = n_18919 ^ n_18841;
assign n_18932 = n_18920 ^ n_18828;
assign n_18933 = n_18920 ^ n_18811;
assign n_18934 = n_18921 ^ n_15689;
assign n_18935 = n_18818 & ~n_18922;
assign n_18936 = n_18923 ^ n_17043;
assign n_18937 = n_18820 & ~n_18924;
assign n_18938 = n_18925 ^ n_18770;
assign n_18939 = n_18770 & n_18925;
assign n_18940 = n_18926 ^ n_18830;
assign n_18941 = n_18926 ^ n_18814;
assign n_18942 = n_18927 ^ n_18826;
assign n_18943 = n_18927 ^ n_18809;
assign n_18944 = n_18928 ^ n_15408;
assign n_18945 = ~n_18835 & n_18929;
assign n_18946 = n_18930 ^ n_15257;
assign n_18947 = ~n_18855 & n_18931;
assign n_18948 = n_18932 ^ n_17014;
assign n_18949 = n_18932 ^ n_15256;
assign n_18950 = n_18828 & ~n_18933;
assign n_18951 = n_18935 ^ n_18911;
assign n_18952 = n_18937 ^ n_18912;
assign n_18953 = n_18938 ^ n_18939;
assign n_18954 = n_18940 ^ n_16322;
assign n_18955 = n_18940 & n_16323;
assign n_18956 = ~n_18940 & ~n_16481;
assign n_18957 = ~n_18830 & n_18941;
assign y52 = n_18942;
assign n_18958 = ~n_18826 & n_18943;
assign n_18959 = n_18945 ^ n_18918;
assign n_18960 = n_18947 ^ n_18919;
assign n_18961 = n_18950 ^ n_18920;
assign n_18962 = n_18951 ^ n_18857;
assign n_18963 = n_18951 ^ n_18843;
assign n_18964 = n_18952 ^ n_18859;
assign n_18965 = n_18952 ^ n_18845;
assign n_18966 = n_18955 ^ n_16322;
assign n_18967 = n_18957 ^ n_18926;
assign n_18968 = n_18958 ^ n_18927;
assign n_18969 = n_18959 ^ n_18874;
assign n_18970 = n_18959 ^ n_18861;
assign n_18971 = n_18960 ^ n_18895;
assign n_18972 = n_18960 ^ n_18880;
assign n_18973 = n_18961 ^ n_18867;
assign n_18974 = n_18961 ^ n_18851;
assign n_18975 = n_18962 ^ n_16613;
assign n_18976 = n_18857 & ~n_18963;
assign n_18977 = n_18859 & ~n_18965;
assign n_18978 = n_18966 ^ n_18956;
assign n_18979 = n_18967 ^ n_18869;
assign n_18980 = n_18967 ^ n_18853;
assign n_18981 = n_18968 ^ n_18865;
assign n_18982 = n_18968 ^ n_18849;
assign n_18983 = n_18969 ^ n_15662;
assign n_18984 = ~n_18874 & n_18970;
assign n_18985 = n_18971 ^ n_16361;
assign n_18986 = n_18971 ^ n_16240;
assign n_18987 = ~n_18895 & n_18972;
assign n_18988 = n_18973 ^ n_16360;
assign n_18989 = n_18973 ^ n_16239;
assign n_18990 = ~n_18867 & n_18974;
assign n_18991 = n_18976 ^ n_18951;
assign n_18992 = n_18977 ^ n_18952;
assign n_18993 = n_18978 ^ n_18940;
assign n_18994 = n_18979 ^ n_16495;
assign n_18995 = n_18979 ^ n_16338;
assign n_18996 = ~n_18869 & n_18980;
assign y53 = n_18981;
assign n_18997 = ~n_18865 & n_18982;
assign n_18998 = n_18984 ^ n_18959;
assign n_18999 = n_18985 ^ n_16859;
assign n_19000 = ~n_16361 & n_18986;
assign n_19001 = n_18987 ^ n_18960;
assign n_19002 = n_18988 ^ n_17016;
assign n_19003 = ~n_16360 & n_18989;
assign n_19004 = n_18990 ^ n_18961;
assign n_19005 = n_18991 ^ n_18897;
assign n_19006 = n_18991 ^ n_18882;
assign n_19007 = n_18992 ^ n_18884;
assign n_19008 = ~n_18992 & n_18900;
assign n_19009 = n_18992 & ~n_18925;
assign n_19010 = n_18913 ^ n_18992;
assign n_19011 = ~n_18992 & ~n_18913;
assign n_19012 = ~n_16495 & n_18995;
assign n_19013 = n_18996 ^ n_18967;
assign n_19014 = n_18997 ^ n_18968;
assign n_19015 = n_18998 ^ n_18915;
assign n_19016 = n_18998 ^ n_18901;
assign n_19017 = n_19000 ^ n_18971;
assign n_19018 = n_19001 ^ n_18934;
assign n_19019 = n_19001 ^ n_18921;
assign n_19020 = n_19003 ^ n_18973;
assign n_19021 = n_19004 ^ n_18907;
assign n_19022 = n_19004 ^ n_18891;
assign n_19023 = n_19005 ^ n_17084;
assign n_19024 = ~n_18897 & n_19006;
assign n_19025 = n_19008 ^ n_18885;
assign n_19026 = n_19009 ^ n_18885;
assign n_19027 = n_19010 ^ n_19011;
assign n_19028 = ~n_18939 & ~n_19011;
assign n_19029 = n_19012 ^ n_18979;
assign n_19030 = n_19013 ^ n_18909;
assign n_19031 = n_19013 ^ n_18893;
assign n_19032 = n_19014 ^ n_18905;
assign n_19033 = n_19014 ^ n_18889;
assign n_19034 = n_19015 ^ n_15806;
assign n_19035 = n_18915 & ~n_19016;
assign n_19036 = n_19018 ^ n_19017;
assign n_19037 = n_19018 ^ n_16341;
assign n_19038 = n_18934 & ~n_19019;
assign n_19039 = n_17182 ^ n_19020;
assign n_19040 = n_19021 ^ n_16497;
assign n_19041 = n_19021 ^ n_16340;
assign n_19042 = ~n_18907 & n_19022;
assign n_19043 = n_19024 ^ n_18991;
assign n_19044 = n_18953 & n_19027;
assign n_19045 = n_19029 ^ n_15687;
assign n_19046 = n_16682 ^ n_19029;
assign n_19047 = n_19030 ^ n_19029;
assign n_19048 = ~n_19029 & n_19030;
assign n_19049 = n_18909 & ~n_19031;
assign y54 = n_19032;
assign n_19050 = ~n_18905 & n_19033;
assign n_19051 = n_19035 ^ n_18998;
assign n_19052 = n_19036 ^ n_16341;
assign n_19053 = ~n_19036 & n_19037;
assign n_19054 = n_19038 ^ n_19001;
assign n_19055 = n_19040 ^ n_17182;
assign n_19056 = ~n_16497 & n_19041;
assign n_19057 = n_19042 ^ n_19004;
assign n_19058 = n_19043 ^ n_18936;
assign n_19059 = n_19043 ^ n_18923;
assign n_19060 = n_19045 ^ n_19030;
assign n_19061 = n_19047 ^ n_16681;
assign n_19062 = ~n_19047 & ~n_19046;
assign n_19063 = n_16682 & n_19048;
assign n_19064 = n_19048 ^ n_19047;
assign n_19065 = n_19049 ^ n_19013;
assign n_19066 = n_19050 ^ n_19014;
assign n_19067 = n_19051 ^ n_18954;
assign n_19068 = n_18955 ^ n_19051;
assign n_19069 = n_19051 & n_18955;
assign n_19070 = ~n_19051 & n_18993;
assign n_19071 = ~n_19051 & n_18956;
assign n_19072 = n_19052 ^ n_17042;
assign n_19073 = n_19053 ^ n_19017;
assign n_19074 = n_19054 ^ n_18975;
assign n_19075 = n_19054 ^ n_18962;
assign n_19076 = n_19055 ^ n_19020;
assign n_19077 = n_19055 & ~n_19039;
assign n_19078 = n_19056 ^ n_19021;
assign n_19079 = n_19057 ^ n_18946;
assign n_19080 = n_19057 ^ n_18930;
assign n_19081 = n_18936 & ~n_19059;
assign n_19082 = n_19048 & n_19060;
assign n_19083 = n_19062 ^ n_19029;
assign n_19084 = ~n_16833 & n_19064;
assign n_19085 = n_19064 ^ n_16496;
assign n_19086 = n_19065 ^ n_18948;
assign n_19087 = n_19065 ^ n_18932;
assign n_19088 = n_18949 ^ n_19065;
assign n_19089 = n_19066 ^ n_18944;
assign n_19090 = n_19066 ^ n_18928;
assign n_19091 = n_19068 ^ n_19069;
assign n_19092 = ~n_18956 & ~n_19070;
assign n_19093 = n_19071 ^ n_19069;
assign n_19094 = n_18994 & ~n_19071;
assign n_19095 = n_19074 ^ n_17063;
assign n_19096 = n_19074 ^ n_19073;
assign n_19097 = n_18975 & ~n_19075;
assign n_19098 = n_19077 ^ n_19040;
assign n_19099 = n_17303 ^ n_19078;
assign n_19100 = n_19079 ^ n_16784;
assign n_19101 = n_19079 ^ n_16612;
assign n_19102 = ~n_18946 & n_19080;
assign n_19103 = n_19081 ^ n_19043;
assign n_19104 = n_19082 ^ n_19060;
assign n_19105 = n_19063 ^ n_19084;
assign n_19106 = ~n_19086 & n_19083;
assign n_19107 = ~n_19086 & ~n_19063;
assign n_19108 = n_19064 ^ n_19086;
assign n_19109 = n_18949 & ~n_19087;
assign n_19110 = n_19088 ^ n_16048;
assign y55 = n_19089;
assign n_19111 = ~n_18944 & n_19090;
assign n_19112 = ~n_18993 & n_19091;
assign n_19113 = n_18994 & n_19092;
assign n_19114 = n_19095 ^ n_19073;
assign n_19115 = n_19095 & ~n_19096;
assign n_19116 = n_19097 ^ n_19054;
assign n_19117 = n_19100 ^ n_17303;
assign n_19118 = ~n_16784 & n_19101;
assign n_19119 = n_19102 ^ n_19057;
assign n_19120 = n_19103 ^ n_18964;
assign n_19121 = n_19085 & ~n_19104;
assign n_19122 = n_19105 ^ n_19061;
assign n_19123 = ~n_16833 ^ ~n_19108;
assign n_19124 = n_19109 ^ n_19065;
assign n_19125 = n_17015 & n_19110;
assign n_19126 = n_19111 ^ n_19066;
assign n_19127 = n_19112 ^ n_19092;
assign n_19128 = n_19094 ^ n_19112;
assign n_19129 = ~n_19069 & ~n_19113;
assign n_19130 = n_19115 ^ n_19073;
assign n_19131 = n_19116 ^ n_19023;
assign n_19132 = n_17084 & n_19116;
assign n_19133 = n_19116 ^ n_17084;
assign n_19134 = n_19117 ^ n_19078;
assign n_19135 = ~n_19117 & n_19099;
assign n_19136 = n_19118 ^ n_19079;
assign n_19137 = n_19119 ^ n_18999;
assign n_19138 = n_19119 ^ n_18985;
assign n_19139 = n_19121 ^ n_16496;
assign n_19140 = n_19124 ^ n_19002;
assign n_19141 = n_19124 ^ n_18988;
assign n_19142 = n_19125 ^ n_16857;
assign n_19143 = n_19126 ^ n_18983;
assign n_19144 = n_19126 ^ n_18969;
assign n_19145 = ~n_19130 & ~n_19005;
assign n_19146 = n_19005 ^ n_19130;
assign n_19147 = n_19131 ^ n_19130;
assign n_19148 = n_19132 & ~n_19058;
assign n_19149 = n_19132 ^ n_19133;
assign n_19150 = n_19134 ^ n_19098;
assign n_19151 = n_19135 ^ n_19100;
assign n_19152 = n_19136 ^ n_17677;
assign n_19153 = n_17677 ^ n_19137;
assign n_19154 = ~n_18999 & n_19138;
assign n_19155 = n_19139 ^ n_19122;
assign n_19156 = ~n_19139 ^ ~n_19107;
assign n_19157 = ~n_19002 & n_19141;
assign n_19158 = n_19140 ^ n_19142;
assign y56 = n_19143;
assign n_19159 = ~n_18983 & n_19144;
assign n_19160 = n_19132 ^ n_19145;
assign n_19161 = ~n_19145 & ~n_19058;
assign n_19162 = ~n_19145 & n_19132;
assign n_19163 = n_19145 ^ n_19146;
assign n_19164 = n_19152 ^ n_19137;
assign n_19165 = n_19152 & ~n_19153;
assign n_19166 = n_19154 ^ n_19119;
assign n_19167 = n_19157 ^ n_19124;
assign n_19168 = n_19159 ^ n_19126;
assign n_19169 = n_19161 ^ n_19162;
assign n_19170 = n_19149 ^ n_19163;
assign n_19171 = n_19058 ^ n_19163;
assign n_19172 = n_19164 ^ n_19151;
assign n_19173 = n_19165 ^ n_19136;
assign n_19174 = n_19166 ^ n_19052;
assign n_19175 = n_19167 ^ n_19076;
assign n_19176 = n_19168 ^ n_19034;
assign n_19177 = n_19168 ^ n_19015;
assign n_19178 = n_19149 & n_19171;
assign n_19179 = n_19174 ^ n_17042;
assign n_19180 = ~n_19174 & n_19072;
assign y57 = ~n_19176;
assign n_19181 = n_19034 & ~n_19177;
assign n_19182 = n_19179 ^ n_19173;
assign n_19183 = n_19180 ^ n_19166;
assign n_19184 = n_19181 ^ n_19168;
assign n_19185 = n_19183 ^ n_19114;
assign n_19186 = n_19184 ^ n_19067;
assign n_19187 = n_19184 & ~n_19127;
assign n_19188 = n_19184 & n_19128;
assign y58 = n_19186;
assign n_19189 = n_19187 ^ n_19092;
assign n_19190 = n_19129 & ~n_19188;
assign n_19191 = n_19189 & ~n_19093;
assign n_19192 = n_19190 ^ n_19061;
assign n_19193 = ~n_19190 & ~n_19122;
assign n_19194 = n_19190 & n_19123;
assign n_19195 = n_19191 ^ n_18994;
assign y60 = n_19192;
assign n_19196 = n_19155 ^ n_19193;
assign n_19197 = n_19156 & ~n_19194;
assign y59 = n_19195;
assign n_19198 = ~n_19105 & n_19196;
assign n_19199 = ~n_19106 & ~n_19197;
assign n_19200 = n_19198 ^ n_19086;
assign n_19201 = n_19199 ^ n_19158;
assign n_19202 = n_19199 ^ n_19140;
assign y61 = ~n_19200;
assign y62 = ~n_19201;
assign n_19203 = ~n_19158 & ~n_19202;
assign n_19204 = n_19203 ^ n_19199;
assign n_19205 = n_19204 ^ n_19175;
assign n_19206 = n_19204 ^ n_19167;
assign y63 = ~n_19205;
assign n_19207 = ~n_19175 & ~n_19206;
assign n_19208 = n_19207 ^ n_19204;
assign n_19209 = n_19208 ^ n_19150;
assign n_19210 = n_19208 ^ n_19134;
assign y64 = n_19209;
assign n_19211 = n_19150 & n_19210;
assign n_19212 = n_19211 ^ n_19208;
assign n_19213 = n_19212 ^ n_19172;
assign n_19214 = n_19212 ^ n_19164;
assign y65 = ~n_19213;
assign n_19215 = ~n_19172 & ~n_19214;
assign n_19216 = n_19215 ^ n_19212;
assign n_19217 = n_19216 ^ n_19182;
assign n_19218 = n_19216 ^ n_19179;
assign y66 = n_19217;
assign n_19219 = n_19182 & n_19218;
assign n_19220 = n_19219 ^ n_19216;
assign n_19221 = n_19220 ^ n_19185;
assign n_19222 = n_19220 ^ n_19183;
assign y67 = n_19221;
assign n_19223 = n_19185 & ~n_19222;
assign n_19224 = n_19223 ^ n_19220;
assign n_19225 = n_19224 ^ n_19147;
assign n_19226 = n_19224 ^ n_19130;
assign n_19227 = n_19224 & n_19163;
assign n_19228 = n_19161 ^ n_19224;
assign y68 = ~n_19225;
assign n_19229 = n_19226 ^ n_19005;
assign n_19230 = n_19169 & ~n_19227;
assign n_19231 = n_19178 & ~n_19228;
assign n_19232 = n_19229 & n_19160;
assign n_19233 = ~n_19229 & n_19170;
assign n_19234 = ~n_19148 & ~n_19231;
assign n_19235 = n_19232 ^ n_19233;
assign n_19236 = ~n_19230 & n_19234;
assign n_19237 = n_19058 ^ n_19235;
assign n_19238 = n_19236 ^ n_19120;
assign n_19239 = n_19236 ^ n_19103;
assign y69 = n_19237;
assign y70 = n_19238;
assign n_19240 = n_19120 & ~n_19239;
assign n_19241 = n_19240 ^ n_19236;
assign n_19242 = n_19241 ^ n_19007;
assign n_19243 = n_19007 & n_19241;
assign n_19244 = ~n_19241 & n_19028;
assign y71 = ~n_19242;
assign n_19245 = n_19243 ^ n_19026;
assign n_19246 = n_19044 & ~n_19244;
assign n_19247 = ~n_19025 ^ ~n_19245;
assign n_19248 = n_19246 ^ n_18813;
assign n_19249 = n_19246 ^ n_18799;
assign n_19250 = ~n_19247 ^ n_18770;
assign y73 = ~n_19248;
assign n_19251 = ~n_18813 & ~n_19249;
assign y72 = ~n_19250;
assign n_19252 = n_19251 ^ n_19246;
assign n_19253 = n_19252 ^ n_18725;
assign n_19254 = n_19252 ^ n_18709;
assign y74 = ~n_19253;
assign n_19255 = ~n_18725 & ~n_19254;
assign n_19256 = n_19255 ^ n_19252;
assign n_19257 = n_19256 ^ n_18668;
assign n_19258 = n_19256 ^ n_18653;
assign y75 = ~n_19257;
assign n_19259 = ~n_18668 & ~n_19258;
assign n_19260 = n_19259 ^ n_19256;
assign n_19261 = n_19260 ^ n_18562;
assign n_19262 = n_19260 ^ n_18545;
assign y76 = n_19261;
assign n_19263 = n_18562 & ~n_19262;
assign n_19264 = n_19263 ^ n_19260;
assign n_19265 = n_19264 ^ n_18437;
assign n_19266 = n_18437 & ~n_19264;
assign n_19267 = ~n_19264 & n_18486;
assign n_19268 = n_19264 ^ n_18418;
assign y77 = ~n_19265;
assign n_19269 = n_19266 ^ n_18484;
assign n_19270 = n_18505 & ~n_19267;
assign n_19271 = n_18438 & ~n_19268;
assign n_19272 = n_18095 ^ n_19269;
assign n_19273 = n_19271 ^ n_18418;
assign n_19274 = n_18096 ^ n_19272;
assign n_19275 = ~n_18123 & ~n_19273;
assign y78 = n_19274;
assign n_19276 = ~n_19270 & ~n_19275;
assign n_19277 = n_19276 ^ n_18170;
assign n_19278 = n_18171 ^ n_19276;
assign n_19279 = n_18201 ^ n_19276;
assign n_19280 = ~n_19276 & n_18247;
assign n_19281 = n_19276 ^ n_17446;
assign y79 = n_19277;
assign n_19282 = n_19278 & n_18198;
assign n_19283 = n_19279 & n_18224;
assign n_19284 = n_18200 & ~n_19280;
assign n_19285 = n_17526 & n_19281;
assign n_19286 = n_19282 ^ n_18223;
assign n_19287 = n_18199 ^ n_19283;
assign n_19288 = n_19285 ^ n_17446;
assign n_19289 = n_19286 ^ n_19287;
assign n_19290 = ~n_18226 & n_19288;
assign n_19291 = n_17614 ^ n_19289;
assign n_19292 = ~n_19284 & ~n_19290;
assign y80 = n_19291;
assign n_19293 = n_19292 ^ n_17825;
assign n_19294 = ~n_17825 & n_19292;
assign n_19295 = ~n_19292 & n_17943;
assign n_19296 = n_19292 ^ n_17047;
assign y81 = n_19293;
assign n_19297 = n_19294 ^ n_17942;
assign n_19298 = n_17876 & ~n_19295;
assign n_19299 = ~n_17183 & ~n_19296;
assign n_19300 = n_17875 ^ n_19297;
assign n_19301 = n_19299 ^ n_17047;
assign n_19302 = n_17366 ^ n_19300;
assign n_19303 = ~n_17913 & ~n_19301;
assign y82 = ~n_19302;
assign n_19304 = ~n_19298 & ~n_19303;
assign n_19305 = n_19304 ^ n_17636;
assign n_19306 = n_19304 ^ n_17542;
assign n_19307 = ~n_19304 & n_17847;
assign y83 = n_19305;
assign n_19308 = n_17636 & n_19306;
assign n_19309 = n_17893 & ~n_19307;
assign n_19310 = n_19308 ^ n_17726;
assign n_19311 = n_19309 ^ n_17653;
assign n_19312 = n_19309 ^ n_17559;
assign n_19313 = n_17387 ^ n_19310;
assign y85 = ~n_19311;
assign n_19314 = n_17653 & n_19312;
assign y84 = n_19313;
assign n_19315 = n_19314 ^ n_19309;
assign n_19316 = n_19315 ^ n_17544;
assign n_19317 = n_19315 ^ n_17467;
assign y86 = ~n_19316;
assign n_19318 = n_17544 & n_19317;
assign n_19319 = n_19318 ^ n_19315;
assign n_19320 = n_19319 ^ n_17503;
assign n_19321 = ~n_17503 & n_19319;
assign n_19322 = n_19319 & n_17681;
assign n_19323 = n_19319 ^ n_16838;
assign y87 = ~n_19320;
assign n_19324 = n_19321 ^ n_17679;
assign n_19325 = ~n_17856 & ~n_19322;
assign n_19326 = ~n_17505 & n_19323;
assign n_19327 = n_19324 ^ n_17504;
assign n_19328 = n_19326 ^ n_17419;
assign n_19329 = n_17370 ^ n_19327;
assign n_19330 = n_17482 & n_19328;
assign y88 = ~n_19329;
assign n_19331 = n_19325 & ~n_19330;
assign n_19332 = n_19331 ^ n_17545;
assign n_19333 = n_17163 & n_19331;
assign n_19334 = n_19331 & ~n_17546;
assign n_19335 = ~n_19331 & n_17729;
assign y89 = ~n_19332;
assign n_19336 = n_17643 & ~n_19334;
assign n_19337 = ~n_19334 & n_17732;
assign n_19338 = ~n_17895 & ~n_19335;
assign n_19339 = n_17894 ^ n_19336;
assign n_19340 = ~n_19337 & n_19338;
assign n_19341 = n_19339 ^ ~n_17731;
assign n_19342 = n_19340 ^ n_17654;
assign n_19343 = n_19340 ^ n_17560;
assign n_19344 = n_17728 ^ n_19341;
assign y91 = ~n_19342;
assign n_19345 = ~n_17654 & ~n_19343;
assign n_19346 = n_19333 ^ n_19344;
assign n_19347 = n_19345 ^ n_19340;
assign n_19348 = n_17392 ^ n_19346;
assign n_19349 = n_19347 ^ n_17548;
assign n_19350 = n_19347 ^ n_17469;
assign y90 = ~n_19348;
assign y92 = n_19349;
assign n_19351 = n_17548 & ~n_19350;
assign n_19352 = n_19351 ^ n_19347;
assign n_19353 = n_19352 ^ n_17584;
assign n_19354 = n_17189 ^ n_19352;
assign n_19355 = ~n_19352 & ~n_17301;
assign n_19356 = ~n_19352 & n_17807;
assign y93 = ~n_19353;
assign n_19357 = ~n_19354 & ~n_17585;
assign n_19358 = n_19355 ^ n_17586;
assign n_19359 = n_17924 & ~n_19356;
assign n_19360 = n_19357 ^ n_19358;
assign n_19361 = n_19359 ^ n_17549;
assign n_19362 = n_19359 ^ n_17472;
assign n_19363 = n_17508 ^ n_19360;
assign y95 = n_19361;
assign n_19364 = n_17549 & ~n_19362;
assign n_19365 = n_17374 ^ n_19363;
assign n_19366 = n_19364 ^ n_19359;
assign y94 = ~n_19365;
assign n_19367 = n_19366 ^ n_17509;
assign n_19368 = n_19366 ^ n_17421;
assign y96 = ~n_19367;
assign n_19369 = ~n_17509 & ~n_19368;
assign n_19370 = n_19369 ^ n_19366;
assign n_19371 = n_19370 ^ n_17655;
assign n_19372 = n_19370 ^ n_17152;
assign n_19373 = n_19370 & n_17852;
assign y97 = n_19371;
assign n_19374 = n_19372 ^ n_17561;
assign n_19375 = n_17955 & ~n_19373;
assign n_19376 = n_19374 & n_17737;
assign n_19377 = ~n_19374 & ~n_17793;
assign n_19378 = n_19375 ^ n_17510;
assign n_19379 = n_19375 ^ n_17423;
assign n_19380 = n_19376 ^ n_19377;
assign y99 = ~n_19378;
assign n_19381 = n_17510 & n_19379;
assign n_19382 = n_17320 ^ n_19380;
assign n_19383 = n_19381 ^ n_19375;
assign y98 = n_19382;
assign n_19384 = n_19383 ^ n_17658;
assign n_19385 = n_19383 ^ n_17562;
assign y100 = n_19384;
assign n_19386 = ~n_17658 & n_19385;
assign n_19387 = n_19386 ^ n_19383;
assign n_19388 = n_19387 ^ n_17550;
assign n_19389 = n_19387 ^ n_17473;
assign y101 = n_19388;
assign n_19390 = ~n_17550 & n_19389;
assign n_19391 = n_19390 ^ n_19387;
assign n_19392 = n_19391 ^ n_17590;
assign n_19393 = n_19391 & n_17400;
assign n_19394 = n_17488 ^ n_19391;
assign n_19395 = n_19391 & n_17685;
assign n_19396 = n_19391 ^ n_17054;
assign y102 = n_19392;
assign n_19397 = n_17756 ^ n_19393;
assign n_19398 = n_19394 & n_17592;
assign n_19399 = ~n_17757 & ~n_19395;
assign n_19400 = n_17399 & ~n_19396;
assign n_19401 = n_19397 ^ n_19398;
assign n_19402 = n_19400 ^ n_17287;
assign n_19403 = n_19401 ^ n_17512;
assign n_19404 = ~n_17594 & n_19402;
assign n_19405 = n_17378 ^ n_19403;
assign n_19406 = n_19399 & ~n_19404;
assign y103 = n_19405;
assign n_19407 = n_19406 ^ n_17551;
assign n_19408 = ~n_19406 & n_17897;
assign n_19409 = ~n_19406 & n_17986;
assign y104 = n_19407;
assign n_19410 = n_19408 ^ n_17741;
assign n_19411 = n_17854 & ~n_19409;
assign n_19412 = n_17853 & n_19410;
assign n_19413 = n_19411 ^ n_17660;
assign n_19414 = n_19411 ^ n_17380;
assign n_19415 = n_19412 ^ n_17402;
assign y106 = n_19413;
assign n_19416 = ~n_17660 & ~n_19414;
assign y105 = n_19415;
assign n_19417 = n_19416 ^ n_17565;
assign n_19418 = n_19417 ^ n_17553;
assign n_19419 = ~n_19417 & n_17291;
assign n_19420 = n_17404 ^ n_19417;
assign n_19421 = ~n_19417 & n_17789;
assign n_19422 = n_19417 ^ n_17475;
assign y107 = ~n_19418;
assign n_19423 = n_19419 ^ n_17646;
assign n_19424 = n_19420 & ~n_17647;
assign n_19425 = ~n_17849 & ~n_19421;
assign n_19426 = n_17555 & n_19422;
assign n_19427 = n_19423 ^ n_19424;
assign n_19428 = n_19426 ^ n_17475;
assign n_19429 = n_17645 ^ n_19427;
assign n_19430 = n_17491 & ~n_19428;
assign n_19431 = n_17405 ^ n_19429;
assign n_19432 = n_19425 & ~n_19430;
assign y108 = ~n_19431;
assign n_19433 = n_19432 ^ n_17661;
assign n_19434 = n_19432 & n_17662;
assign n_19435 = n_17744 ^ n_19432;
assign n_19436 = n_19432 & ~n_17798;
assign n_19437 = n_19432 ^ n_17566;
assign y109 = n_19433;
assign n_19438 = n_17742 ^ n_19434;
assign n_19439 = ~n_19435 & n_17799;
assign n_19440 = n_17855 & ~n_19436;
assign n_19441 = n_17663 & n_19437;
assign n_19442 = n_19438 ^ n_19439;
assign n_19443 = n_19441 ^ n_17566;
assign n_19444 = n_17307 ^ n_19442;
assign n_19445 = ~n_17493 & ~n_19443;
assign n_19446 = n_17407 ^ n_19444;
assign n_19447 = ~n_19440 & ~n_19445;
assign y110 = ~n_19446;
assign n_19448 = n_19447 ^ n_17664;
assign n_19449 = ~n_19447 & n_17745;
assign n_19450 = ~n_19447 & n_17568;
assign n_19451 = ~n_19447 & ~n_17361;
assign n_19452 = n_19447 & n_17747;
assign y111 = ~n_19448;
assign n_19453 = n_19449 ^ n_19450;
assign n_19454 = n_17568 ^ n_19451;
assign n_19455 = ~n_19451 & n_17746;
assign n_19456 = ~n_19451 & n_17748;
assign n_19457 = ~n_17801 & ~n_19452;
assign n_19458 = ~n_17666 & ~n_19454;
assign n_19459 = ~n_19456 & n_19457;
assign n_19460 = n_19458 ^ n_19455;
assign n_19461 = n_19459 ^ n_17779;
assign n_19462 = ~n_19459 & ~n_17840;
assign n_19463 = ~n_19459 & n_17721;
assign n_19464 = ~n_19459 & n_17631;
assign n_19465 = n_19459 & n_17842;
assign n_19466 = n_19453 ^ n_19460;
assign y113 = n_19461;
assign n_19467 = n_19462 ^ n_19463;
assign n_19468 = n_17721 ^ n_19464;
assign n_19469 = ~n_19464 & n_17841;
assign n_19470 = ~n_19464 & n_17843;
assign n_19471 = ~n_17891 & ~n_19465;
assign n_19472 = n_19466 ^ n_17361;
assign n_19473 = ~n_17781 & ~n_19468;
assign n_19474 = ~n_19470 & n_19471;
assign n_19475 = n_17536 ^ n_19472;
assign n_19476 = n_19473 ^ n_19469;
assign n_19477 = n_19474 ^ n_17669;
assign n_19478 = n_19474 ^ n_17382;
assign y112 = n_19475;
assign n_19479 = n_19467 ^ n_19476;
assign y115 = n_19477;
assign n_19480 = n_17669 & ~n_19478;
assign n_19481 = n_19479 ^ n_17631;
assign n_19482 = n_19480 ^ n_17569;
assign n_19483 = n_17410 ^ n_19481;
assign n_19484 = n_19482 ^ n_17556;
assign n_19485 = n_19482 ^ n_17364;
assign y114 = n_19483;
assign y116 = n_19484;
assign n_19486 = n_17556 & ~n_19485;
assign n_19487 = n_19486 ^ n_17476;
assign n_19488 = n_19487 ^ n_17632;
assign n_19489 = n_19487 & ~n_17634;
assign n_19490 = ~n_19487 & ~n_17541;
assign n_19491 = ~n_19487 & ~n_17196;
assign n_19492 = n_19487 & n_17635;
assign y117 = n_19488;
assign n_19493 = n_19489 ^ n_19490;
assign n_19494 = n_17302 & ~n_19491;
assign n_19495 = ~n_17845 & ~n_19492;
assign n_19496 = n_17892 ^ n_19494;
assign n_19497 = n_19494 & ~n_17724;
assign n_19498 = n_19493 ^ n_19496;
assign n_19499 = n_19495 & ~n_19497;
assign n_19500 = n_17384 ^ n_19498;
assign n_19501 = n_19499 ^ n_17648;
assign n_19502 = n_19499 & ~n_17235;
assign n_19503 = n_17326 ^ n_19499;
assign n_19504 = ~n_19499 & n_17670;
assign y118 = ~n_19500;
assign y119 = n_19501;
assign n_19505 = n_19502 ^ n_19499;
assign n_19506 = ~n_19502 & n_17791;
assign n_19507 = ~n_19503 & ~n_17650;
assign n_19508 = ~n_17790 & ~n_19504;
assign n_19509 = n_19505 ^ n_17649;
assign n_19510 = ~n_19506 & n_19508;
assign n_19511 = n_19509 ^ n_19507;
assign n_19512 = n_19510 ^ n_17671;
assign n_19513 = n_19510 ^ n_17571;
assign n_19514 = n_17558 ^ n_19511;
assign y121 = ~n_19512;
assign n_19515 = ~n_17671 & ~n_19513;
assign n_19516 = n_17496 ^ n_19514;
assign n_19517 = n_19515 ^ n_19510;
assign y120 = n_19516;
assign n_19518 = n_19517 ^ n_17572;
assign n_19519 = n_17573 ^ n_19517;
assign n_19520 = n_17499 ^ n_19517;
assign n_19521 = ~n_19517 & n_17803;
assign y122 = ~n_19518;
assign n_19522 = ~n_19519 & ~n_17672;
assign n_19523 = ~n_19520 & ~n_17575;
assign n_19524 = n_17802 & ~n_19521;
assign n_19525 = n_19522 ^ n_17574;
assign n_19526 = n_19523 ^ n_17673;
assign n_19527 = n_19524 ^ n_17686;
assign n_19528 = n_19524 ^ n_17309;
assign n_19529 = n_19525 ^ n_19526;
assign y124 = ~n_19527;
assign n_19530 = n_17686 & ~n_19528;
assign n_19531 = n_17427 ^ n_19529;
assign n_19532 = n_19530 ^ n_17595;
assign y123 = ~n_19531;
assign n_19533 = n_19532 ^ n_17500;
assign n_19534 = n_19532 ^ n_17414;
assign y125 = n_19533;
assign n_19535 = n_17500 & ~n_19534;
assign n_19536 = n_19535 ^ n_19532;
assign n_19537 = n_19536 ^ n_17804;
assign n_19538 = n_19536 ^ n_17752;
assign y126 = n_19537;
assign n_19539 = n_17804 & ~n_19538;
assign n_19540 = n_19539 ^ n_19536;
assign n_19541 = n_19540 ^ n_6612;
assign y127 = n_19541;
endmodule