module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n307 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n617 , n618 , n619 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n758 , n759 , n760 , n766 , n767 , n768 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n781 , n784 , n785 , n786 , n787 , n788 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n927 , n930 , n931 , n932 , n933 , n934 , n935 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1020 , n1021 , n1022 , n1023 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1072 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1143 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1278 , n1279 , n1280 , n1281 , n1282 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1297 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1567 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1706 , n1707 , n1708 , n1709 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1763 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1882 , n1883 , n1884 , n1885 , n1886 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1906 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1938 , n1939 , n1940 , n1941 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1956 , n1957 , n1958 , n1959 , n1962 , n1963 , n1964 , n1966 , n1967 , n1968 , n1972 , n1973 , n1974 , n1975 , n1977 , n1978 , n1979 , n1986 , n1987 , n1988 , n1990 , n1991 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2018 , n2019 , n2020 , n2021 , n2022 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2883 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3170 , n3171 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3387 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4114 , n4115 , n4116 , n4117 , n4118 , n4121 , n4122 , n4123 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4351 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5312 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5823 , n5824 , n5825 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6356 , n6357 , n6358 , n6359 , n6360 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6519 , n6520 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7156 , n7157 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7996 , n7997 , n7998 , n7999 , n8000 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8185 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8197 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9534 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9824 , n9825 , n9826 , n9827 , n9828 , n9830 , n9832 , n9833 , n9834 , n9835 , n9838 , n9839 , n9840 , n9841 , n9845 , n9846 , n9847 , n9849 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9873 , n9874 , n9875 , n9877 , n9879 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9897 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9931 , n9934 , n9936 , n9937 , n9938 , n9942 , n9943 , n9944 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9954 , n9955 , n9956 , n9959 , n9960 , n9961 , n9962 , n9963 , n9968 , n9969 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10008 , n10009 , n10011 , n10012 , n10013 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10039 , n10040 , n10041 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10052 , n10053 , n10054 , n10055 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10069 , n10070 , n10071 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10566 , n10567 , n10568 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10849 , n10850 , n10851 , n10852 , n10853 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10979 , n10980 , n10981 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11336 , n11337 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11548 , n11549 , n11550 , n11551 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14230 , n14231 , n14232 , n14234 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 ;
  assign n136 = x125 & ~x126 ;
  assign n129 = x124 & ~x125 ;
  assign n135 = ~x126 & ~n129 ;
  assign n137 = n136 ^ n135 ;
  assign n134 = x126 & ~x127 ;
  assign n138 = n137 ^ n134 ;
  assign n183 = n134 ^ x127 ;
  assign n2950 = ~x74 & ~x75 ;
  assign n2951 = ~x76 & n2950 ;
  assign n130 = n129 ^ x125 ;
  assign n1003 = ~n130 & ~n183 ;
  assign n837 = ~x100 & ~x101 ;
  assign n838 = ~x102 & n837 ;
  assign n352 = x112 & ~x113 ;
  assign n146 = x122 & ~x123 ;
  assign n147 = n146 ^ x123 ;
  assign n166 = n147 ^ x124 ;
  assign n148 = ~x124 & ~n147 ;
  assign n167 = n166 ^ n148 ;
  assign n168 = x125 & ~n167 ;
  assign n141 = x127 ^ x126 ;
  assign n142 = n141 ^ n137 ;
  assign n143 = n142 ^ x125 ;
  assign n144 = n143 ^ x127 ;
  assign n145 = n144 ^ n137 ;
  assign n149 = n148 ^ n145 ;
  assign n150 = n148 ^ x127 ;
  assign n151 = n150 ^ x127 ;
  assign n154 = x126 & n151 ;
  assign n155 = n154 ^ x127 ;
  assign n156 = ~n149 & ~n155 ;
  assign n157 = n156 ^ n142 ;
  assign n160 = ~n146 & ~n157 ;
  assign n132 = ~x120 & ~x121 ;
  assign n133 = ~x122 & n132 ;
  assign n139 = n138 ^ n133 ;
  assign n140 = n138 ^ x123 ;
  assign n158 = n157 ^ n140 ;
  assign n159 = n139 & ~n158 ;
  assign n161 = n160 ^ n159 ;
  assign n162 = n161 ^ x123 ;
  assign n169 = n162 ^ x126 ;
  assign n170 = n168 & ~n169 ;
  assign n131 = n130 ^ x127 ;
  assign n163 = ~x125 & n162 ;
  assign n164 = n163 ^ n148 ;
  assign n165 = n131 & n164 ;
  assign n171 = n170 ^ n165 ;
  assign n172 = n137 ^ x125 ;
  assign n173 = n147 ^ x126 ;
  assign n174 = ~x125 & x127 ;
  assign n175 = ~x124 & n174 ;
  assign n176 = n173 & n175 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n177 ^ x127 ;
  assign n179 = n178 ^ n162 ;
  assign n180 = ~x124 & x127 ;
  assign n181 = ~n136 & n147 ;
  assign n182 = n180 & ~n181 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = n179 & ~n184 ;
  assign n186 = n172 & n185 ;
  assign n187 = n186 ^ n178 ;
  assign n188 = ~n171 & ~n187 ;
  assign n247 = n188 ^ x119 ;
  assign n203 = n188 ^ n157 ;
  assign n201 = n188 ^ x121 ;
  assign n202 = n201 ^ x120 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = n204 ^ n203 ;
  assign n206 = n205 ^ n201 ;
  assign n211 = ~n201 & n203 ;
  assign n207 = ~x118 & ~x119 ;
  assign n208 = n207 ^ n201 ;
  assign n209 = n201 ^ n157 ;
  assign n210 = ~n208 & ~n209 ;
  assign n212 = n211 ^ n210 ;
  assign n213 = ~n206 & n212 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ n157 ;
  assign n216 = n215 ^ n138 ;
  assign n218 = n132 ^ x122 ;
  assign n190 = n157 ^ n132 ;
  assign n217 = n188 & ~n190 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = n219 ^ n215 ;
  assign n221 = n216 & ~n220 ;
  assign n222 = n221 ^ n138 ;
  assign n198 = n139 ^ x123 ;
  assign n199 = n198 ^ n157 ;
  assign n189 = n138 ^ n132 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = n191 ^ n189 ;
  assign n193 = n189 ^ x122 ;
  assign n194 = n193 ^ n189 ;
  assign n195 = ~n192 & n194 ;
  assign n196 = n195 ^ n189 ;
  assign n197 = n188 & ~n196 ;
  assign n200 = n199 ^ n197 ;
  assign n223 = n222 ^ n200 ;
  assign n238 = n163 & n178 ;
  assign n232 = x127 ^ x124 ;
  assign n233 = x125 & ~n147 ;
  assign n234 = ~n232 & n233 ;
  assign n235 = n234 ^ n182 ;
  assign n236 = n162 & n235 ;
  assign n237 = n236 ^ n182 ;
  assign n239 = n238 ^ n237 ;
  assign n226 = n167 ^ x127 ;
  assign n227 = ~n162 & n226 ;
  assign n228 = n227 ^ n167 ;
  assign n229 = n129 & ~n228 ;
  assign n230 = n229 ^ n167 ;
  assign n231 = n169 & ~n230 ;
  assign n240 = n239 ^ n231 ;
  assign n241 = n240 ^ n183 ;
  assign n242 = n241 ^ n200 ;
  assign n243 = n242 ^ n240 ;
  assign n244 = ~n223 & ~n243 ;
  assign n245 = n244 ^ n241 ;
  assign n248 = n247 ^ n245 ;
  assign n250 = n188 ^ x118 ;
  assign n249 = ~x116 & ~x117 ;
  assign n251 = n250 ^ n249 ;
  assign n252 = ~n248 & ~n251 ;
  assign n260 = n252 ^ n203 ;
  assign n246 = n245 ^ n188 ;
  assign n257 = n246 & n247 ;
  assign n258 = n257 ^ n252 ;
  assign n259 = x118 & n258 ;
  assign n261 = n260 ^ n259 ;
  assign n273 = n207 ^ n188 ;
  assign n274 = ~n245 & ~n273 ;
  assign n275 = n274 ^ n188 ;
  assign n276 = n275 ^ x120 ;
  assign n277 = n276 ^ n157 ;
  assign n278 = ~n261 & ~n277 ;
  assign n279 = n278 ^ n276 ;
  assign n280 = n279 ^ n138 ;
  assign n284 = x120 & ~n275 ;
  assign n281 = n207 ^ n157 ;
  assign n282 = ~n245 & ~n281 ;
  assign n283 = n282 ^ n201 ;
  assign n285 = n284 ^ n283 ;
  assign n286 = n285 ^ n279 ;
  assign n287 = ~n280 & ~n286 ;
  assign n288 = n287 ^ n138 ;
  assign n262 = n216 & ~n245 ;
  assign n263 = n262 ^ n219 ;
  assign n289 = n183 & ~n263 ;
  assign n290 = n288 & ~n289 ;
  assign n265 = n263 ^ n200 ;
  assign n264 = n263 ^ n240 ;
  assign n266 = n265 ^ n264 ;
  assign n269 = n222 & n266 ;
  assign n270 = n269 ^ n265 ;
  assign n271 = n183 & n270 ;
  assign n272 = n271 ^ n263 ;
  assign n291 = n290 ^ n272 ;
  assign n298 = n249 ^ n245 ;
  assign n299 = ~n291 & ~n298 ;
  assign n300 = n299 ^ n249 ;
  assign n303 = n300 ^ x118 ;
  assign n304 = n303 ^ n188 ;
  assign n305 = n291 ^ x117 ;
  assign n307 = n291 ^ n245 ;
  assign n315 = n305 & ~n307 ;
  assign n311 = ~x114 & ~x115 ;
  assign n312 = n311 ^ n305 ;
  assign n313 = n305 ^ n245 ;
  assign n314 = n312 & n313 ;
  assign n316 = n315 ^ n314 ;
  assign n317 = ~x116 & n316 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n318 ^ n245 ;
  assign n320 = n319 ^ n303 ;
  assign n321 = n304 & ~n320 ;
  assign n322 = n321 ^ n188 ;
  assign n301 = x118 & n300 ;
  assign n295 = n249 ^ n188 ;
  assign n296 = n291 & ~n295 ;
  assign n294 = n245 ^ x119 ;
  assign n297 = n296 ^ n294 ;
  assign n302 = n301 ^ n297 ;
  assign n323 = n322 ^ n302 ;
  assign n324 = n302 ^ n157 ;
  assign n325 = ~n323 & n324 ;
  assign n326 = n325 ^ n322 ;
  assign n292 = n261 & n291 ;
  assign n293 = n292 ^ n276 ;
  assign n327 = n326 ^ n293 ;
  assign n332 = n293 ^ n138 ;
  assign n333 = n327 & ~n332 ;
  assign n328 = ~n280 & n291 ;
  assign n329 = n328 ^ n285 ;
  assign n330 = n329 ^ n138 ;
  assign n334 = n333 ^ n330 ;
  assign n339 = n329 ^ n183 ;
  assign n340 = n334 & n339 ;
  assign n335 = n289 ^ n183 ;
  assign n336 = n335 ^ n272 ;
  assign n337 = n288 & n336 ;
  assign n338 = n337 ^ n289 ;
  assign n341 = n340 ^ n338 ;
  assign n342 = n326 ^ n138 ;
  assign n343 = ~n341 & n342 ;
  assign n344 = n343 ^ n293 ;
  assign n388 = n322 ^ n157 ;
  assign n389 = ~n341 & n388 ;
  assign n390 = n389 ^ n302 ;
  assign n350 = n291 ^ x115 ;
  assign n351 = n350 ^ n341 ;
  assign n354 = n291 ^ x114 ;
  assign n353 = n352 ^ x113 ;
  assign n355 = n354 ^ n353 ;
  assign n356 = n351 & ~n355 ;
  assign n364 = n356 ^ n307 ;
  assign n349 = n341 ^ n291 ;
  assign n361 = ~n349 & ~n350 ;
  assign n362 = n361 ^ n356 ;
  assign n363 = x114 & n362 ;
  assign n365 = n364 ^ n363 ;
  assign n366 = n311 ^ n291 ;
  assign n367 = ~n341 & n366 ;
  assign n368 = n367 ^ n291 ;
  assign n369 = n368 ^ x116 ;
  assign n370 = n369 ^ n245 ;
  assign n371 = n365 & n370 ;
  assign n372 = n371 ^ n369 ;
  assign n373 = n372 ^ n188 ;
  assign n377 = x116 & n368 ;
  assign n374 = n311 ^ n245 ;
  assign n375 = ~n341 & ~n374 ;
  assign n376 = n375 ^ n305 ;
  assign n378 = n377 ^ n376 ;
  assign n379 = n378 ^ n372 ;
  assign n380 = n373 & ~n379 ;
  assign n381 = n380 ^ n203 ;
  assign n382 = n319 ^ n188 ;
  assign n383 = ~n341 & n382 ;
  assign n384 = n383 ^ n303 ;
  assign n385 = n384 ^ n157 ;
  assign n386 = ~n381 & n385 ;
  assign n387 = n386 ^ n384 ;
  assign n391 = n390 ^ n387 ;
  assign n392 = n390 ^ n138 ;
  assign n393 = n391 & ~n392 ;
  assign n394 = n393 ^ n138 ;
  assign n400 = n344 & ~n394 ;
  assign n346 = n329 & n341 ;
  assign n347 = ~n334 & n346 ;
  assign n345 = n344 ^ n334 ;
  assign n348 = n347 ^ n345 ;
  assign n398 = n394 ^ n348 ;
  assign n399 = n183 & n398 ;
  assign n401 = n400 ^ n399 ;
  assign n431 = ~n352 & ~n401 ;
  assign n422 = ~x110 & ~x111 ;
  assign n423 = ~x112 & n422 ;
  assign n424 = n423 ^ n341 ;
  assign n427 = n401 ^ x113 ;
  assign n428 = n427 ^ n423 ;
  assign n429 = n424 & n428 ;
  assign n425 = n291 ^ x113 ;
  assign n430 = n429 ^ n425 ;
  assign n432 = n431 ^ n430 ;
  assign n397 = n387 ^ n138 ;
  assign n402 = n397 & ~n401 ;
  assign n403 = n402 ^ n390 ;
  assign n405 = n403 ^ n183 ;
  assign n406 = n381 & ~n401 ;
  assign n407 = n406 ^ n384 ;
  assign n408 = n407 ^ n138 ;
  assign n442 = n373 & ~n401 ;
  assign n443 = n442 ^ n378 ;
  assign n409 = ~n365 & ~n401 ;
  assign n410 = n409 ^ n369 ;
  assign n411 = n410 ^ n188 ;
  assign n416 = n353 ^ n341 ;
  assign n417 = ~n401 & n416 ;
  assign n418 = n417 ^ n341 ;
  assign n419 = x114 & ~n418 ;
  assign n413 = n353 ^ n291 ;
  assign n414 = ~n401 & ~n413 ;
  assign n412 = n341 ^ x115 ;
  assign n415 = n414 ^ n412 ;
  assign n420 = n419 ^ n415 ;
  assign n421 = n420 ^ n245 ;
  assign n433 = n418 ^ x114 ;
  assign n434 = n433 ^ n291 ;
  assign n435 = ~n432 & n434 ;
  assign n436 = n435 ^ n307 ;
  assign n437 = ~n421 & n436 ;
  assign n438 = n437 ^ n420 ;
  assign n439 = n438 ^ n410 ;
  assign n440 = n411 & n439 ;
  assign n441 = n440 ^ n188 ;
  assign n444 = n443 ^ n441 ;
  assign n445 = n441 ^ n157 ;
  assign n446 = n444 & ~n445 ;
  assign n447 = n446 ^ n443 ;
  assign n448 = n447 ^ n407 ;
  assign n449 = n408 & ~n448 ;
  assign n450 = n449 ^ n138 ;
  assign n451 = n450 ^ n403 ;
  assign n395 = n348 & n394 ;
  assign n396 = n395 ^ n344 ;
  assign n452 = n451 ^ n396 ;
  assign n453 = n405 & n452 ;
  assign n404 = n403 ^ n396 ;
  assign n454 = n453 ^ n404 ;
  assign n455 = ~n396 & ~n453 ;
  assign n456 = ~n454 & n455 ;
  assign n457 = n456 ^ n454 ;
  assign n458 = ~n432 & n457 ;
  assign n459 = n458 ^ n433 ;
  assign n460 = n459 ^ n245 ;
  assign n461 = n457 ^ n401 ;
  assign n463 = n401 ^ x111 ;
  assign n476 = ~n461 & n463 ;
  assign n464 = n463 ^ n457 ;
  assign n467 = n401 ^ x110 ;
  assign n465 = x108 & ~x109 ;
  assign n466 = n465 ^ x109 ;
  assign n468 = n467 ^ n466 ;
  assign n469 = n464 & n468 ;
  assign n477 = n476 ^ n469 ;
  assign n478 = x110 & n477 ;
  assign n462 = n401 ^ n341 ;
  assign n470 = n469 ^ n462 ;
  assign n479 = n478 ^ n470 ;
  assign n481 = n422 ^ n401 ;
  assign n482 = n457 & ~n481 ;
  assign n480 = n401 ^ x112 ;
  assign n483 = n482 ^ n480 ;
  assign n484 = n483 ^ n341 ;
  assign n485 = n479 & ~n484 ;
  assign n486 = n485 ^ n349 ;
  assign n487 = n423 ^ n401 ;
  assign n488 = n487 ^ n341 ;
  assign n496 = n488 ^ x113 ;
  assign n493 = ~x112 & ~n401 ;
  assign n494 = n493 ^ n488 ;
  assign n495 = ~n457 & n494 ;
  assign n497 = n496 ^ n495 ;
  assign n498 = n497 ^ n291 ;
  assign n499 = ~n486 & ~n498 ;
  assign n500 = n499 ^ n307 ;
  assign n501 = ~n460 & n500 ;
  assign n502 = n501 ^ n459 ;
  assign n503 = n502 ^ n188 ;
  assign n504 = ~n436 & n457 ;
  assign n505 = n504 ^ n420 ;
  assign n506 = n505 ^ n502 ;
  assign n507 = ~n503 & ~n506 ;
  assign n508 = n507 ^ n203 ;
  assign n511 = n447 ^ n138 ;
  assign n512 = n457 & n511 ;
  assign n513 = n512 ^ n407 ;
  assign n514 = n513 ^ n183 ;
  assign n516 = n438 ^ n188 ;
  assign n517 = n457 & ~n516 ;
  assign n518 = n517 ^ n410 ;
  assign n519 = n518 ^ n157 ;
  assign n520 = ~n508 & n519 ;
  assign n521 = n520 ^ n518 ;
  assign n522 = n521 ^ n138 ;
  assign n523 = n445 & n457 ;
  assign n524 = n523 ^ n443 ;
  assign n525 = n524 ^ n521 ;
  assign n526 = n522 & ~n525 ;
  assign n527 = n526 ^ n138 ;
  assign n509 = n404 & n450 ;
  assign n510 = n509 ^ n403 ;
  assign n515 = n513 ^ n510 ;
  assign n528 = n527 ^ n515 ;
  assign n529 = ~n514 & ~n528 ;
  assign n530 = n529 ^ n513 ;
  assign n531 = n530 ^ n510 ;
  assign n532 = ~n510 & n531 ;
  assign n533 = ~n529 & n532 ;
  assign n534 = n533 ^ n531 ;
  assign n535 = n508 & ~n534 ;
  assign n536 = n535 ^ n518 ;
  assign n537 = n536 ^ n138 ;
  assign n584 = ~n503 & ~n534 ;
  assign n585 = n584 ^ n505 ;
  assign n538 = ~n486 & ~n534 ;
  assign n539 = n538 ^ n497 ;
  assign n540 = n539 ^ n245 ;
  assign n550 = n534 ^ x109 ;
  assign n551 = n550 ^ n457 ;
  assign n555 = x106 & ~x107 ;
  assign n556 = n555 ^ x107 ;
  assign n557 = ~x108 & ~n556 ;
  assign n558 = n557 ^ n457 ;
  assign n559 = n551 & ~n558 ;
  assign n554 = ~n465 & ~n534 ;
  assign n560 = n559 ^ n554 ;
  assign n561 = n560 ^ x109 ;
  assign n562 = n561 ^ n401 ;
  assign n545 = n466 ^ n457 ;
  assign n546 = n534 & ~n545 ;
  assign n547 = n546 ^ n466 ;
  assign n563 = n547 ^ x110 ;
  assign n564 = n563 ^ n561 ;
  assign n565 = n562 & n564 ;
  assign n566 = n565 ^ n401 ;
  assign n548 = x110 & ~n547 ;
  assign n542 = n466 ^ n401 ;
  assign n543 = ~n534 & n542 ;
  assign n541 = n457 ^ x111 ;
  assign n544 = n543 ^ n541 ;
  assign n549 = n548 ^ n544 ;
  assign n567 = n566 ^ n549 ;
  assign n568 = n566 ^ n341 ;
  assign n569 = ~n567 & n568 ;
  assign n570 = n569 ^ n349 ;
  assign n571 = n479 & ~n534 ;
  assign n572 = n571 ^ n483 ;
  assign n573 = n572 ^ n291 ;
  assign n574 = ~n570 & n573 ;
  assign n575 = n574 ^ n307 ;
  assign n576 = n540 & n575 ;
  assign n577 = n576 ^ n539 ;
  assign n578 = n577 ^ n188 ;
  assign n579 = ~n500 & ~n534 ;
  assign n580 = n579 ^ n459 ;
  assign n581 = n580 ^ n577 ;
  assign n582 = n578 & n581 ;
  assign n583 = n582 ^ n188 ;
  assign n586 = n585 ^ n583 ;
  assign n587 = n583 ^ n157 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = n588 ^ n585 ;
  assign n590 = n589 ^ n536 ;
  assign n591 = n537 & n590 ;
  assign n592 = n591 ^ n138 ;
  assign n600 = ~n183 & n510 ;
  assign n601 = n600 ^ n515 ;
  assign n602 = n527 & ~n601 ;
  assign n593 = n522 & ~n534 ;
  assign n594 = n593 ^ n524 ;
  assign n595 = n594 ^ n513 ;
  assign n603 = n602 ^ n595 ;
  assign n617 = n592 & n603 ;
  assign n618 = n617 ^ n594 ;
  assign n619 = n183 & n618 ;
  assign n604 = n183 & ~n603 ;
  assign n605 = n594 ^ n183 ;
  assign n606 = n605 ^ n604 ;
  assign n607 = ~n604 & ~n606 ;
  assign n608 = n592 & n607 ;
  assign n609 = n608 ^ n606 ;
  assign n610 = n589 ^ n138 ;
  assign n611 = n609 & ~n610 ;
  assign n612 = n611 ^ n536 ;
  assign n692 = n612 ^ n183 ;
  assign n622 = n578 & n609 ;
  assign n623 = n622 ^ n580 ;
  assign n624 = n623 ^ n157 ;
  assign n625 = ~n575 & n609 ;
  assign n626 = n625 ^ n539 ;
  assign n627 = n626 ^ n188 ;
  assign n628 = n568 & n609 ;
  assign n629 = n628 ^ n549 ;
  assign n630 = n629 ^ n291 ;
  assign n631 = n562 & n609 ;
  assign n632 = n631 ^ n563 ;
  assign n633 = n632 ^ n341 ;
  assign n660 = n558 ^ n550 ;
  assign n657 = x108 & ~n534 ;
  assign n658 = n657 ^ n558 ;
  assign n659 = ~n609 & n658 ;
  assign n661 = n660 ^ n659 ;
  assign n635 = n556 ^ n534 ;
  assign n636 = n609 & n635 ;
  assign n634 = n534 ^ x108 ;
  assign n637 = n636 ^ n634 ;
  assign n638 = n637 ^ n457 ;
  assign n649 = ~n555 & n609 ;
  assign n639 = x104 & ~x105 ;
  assign n640 = n639 ^ x105 ;
  assign n641 = ~x106 & ~n640 ;
  assign n642 = n641 ^ n534 ;
  assign n643 = n457 ^ x107 ;
  assign n644 = n643 ^ n534 ;
  assign n645 = n644 ^ n457 ;
  assign n646 = n645 ^ n609 ;
  assign n647 = n642 & n646 ;
  assign n648 = n647 ^ n643 ;
  assign n650 = n649 ^ n648 ;
  assign n651 = n638 & n650 ;
  assign n652 = n651 ^ n637 ;
  assign n662 = n661 ^ n652 ;
  assign n663 = n661 ^ n401 ;
  assign n664 = ~n662 & ~n663 ;
  assign n665 = n664 ^ n462 ;
  assign n666 = ~n633 & n665 ;
  assign n667 = n666 ^ n349 ;
  assign n668 = ~n630 & ~n667 ;
  assign n669 = n668 ^ n307 ;
  assign n670 = ~n570 & n609 ;
  assign n671 = n670 ^ n572 ;
  assign n672 = n671 ^ n245 ;
  assign n673 = n669 & ~n672 ;
  assign n674 = n673 ^ n671 ;
  assign n675 = n674 ^ n626 ;
  assign n676 = n627 & n675 ;
  assign n677 = n676 ^ n203 ;
  assign n678 = ~n624 & ~n677 ;
  assign n679 = n678 ^ n623 ;
  assign n680 = n679 ^ n138 ;
  assign n681 = n587 & n609 ;
  assign n682 = n681 ^ n585 ;
  assign n683 = n682 ^ n679 ;
  assign n684 = ~n680 & ~n683 ;
  assign n685 = n684 ^ n138 ;
  assign n693 = n685 ^ n612 ;
  assign n694 = ~n692 & n693 ;
  assign n695 = n694 ^ n612 ;
  assign n696 = ~n619 & ~n695 ;
  assign n839 = n838 ^ n696 ;
  assign n688 = ~n619 & n685 ;
  assign n689 = n688 ^ n183 ;
  assign n690 = ~n612 & n689 ;
  assign n686 = n685 ^ n183 ;
  assign n691 = n690 ^ n686 ;
  assign n697 = ~n680 & ~n696 ;
  assign n698 = n697 ^ n682 ;
  assign n699 = n698 ^ n183 ;
  assign n4971 = n137 ^ x127 ;
  assign n702 = n674 ^ n188 ;
  assign n703 = ~n696 & ~n702 ;
  assign n704 = n703 ^ n626 ;
  assign n705 = n704 ^ n157 ;
  assign n706 = ~n669 & ~n696 ;
  assign n707 = n706 ^ n671 ;
  assign n708 = n707 ^ n188 ;
  assign n715 = n665 & ~n696 ;
  assign n716 = n715 ^ n632 ;
  assign n717 = n716 ^ n291 ;
  assign n758 = n652 ^ n401 ;
  assign n759 = ~n696 & ~n758 ;
  assign n760 = n759 ^ n661 ;
  assign n807 = n760 ^ n349 ;
  assign n719 = ~n650 & ~n696 ;
  assign n720 = n719 ^ n637 ;
  assign n721 = n720 ^ n401 ;
  assign n729 = n642 ^ x107 ;
  assign n730 = n729 ^ n609 ;
  assign n726 = x106 & n609 ;
  assign n727 = n726 ^ n642 ;
  assign n728 = n696 & ~n727 ;
  assign n731 = n730 ^ n728 ;
  assign n732 = n731 ^ n457 ;
  assign n750 = n534 ^ n457 ;
  assign n735 = n640 ^ x106 ;
  assign n733 = n640 ^ n609 ;
  assign n734 = n696 & ~n733 ;
  assign n736 = n735 ^ n734 ;
  assign n737 = n736 ^ n534 ;
  assign n747 = ~n639 & ~n696 ;
  assign n738 = ~x102 & ~x103 ;
  assign n739 = ~x104 & n738 ;
  assign n740 = n739 ^ n609 ;
  assign n743 = n609 ^ x105 ;
  assign n744 = n743 ^ n696 ;
  assign n745 = ~n740 & n744 ;
  assign n741 = n534 ^ x105 ;
  assign n746 = n745 ^ n741 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = ~n737 & n748 ;
  assign n751 = n750 ^ n749 ;
  assign n752 = n732 & n751 ;
  assign n753 = n752 ^ n731 ;
  assign n754 = n753 ^ n720 ;
  assign n755 = ~n721 & ~n754 ;
  assign n756 = n755 ^ n401 ;
  assign n808 = n807 ^ n756 ;
  assign n809 = n808 ^ n349 ;
  assign n810 = n756 ^ n341 ;
  assign n813 = n809 & n810 ;
  assign n718 = n716 ^ n341 ;
  assign n766 = n813 ^ n718 ;
  assign n767 = n717 & n766 ;
  assign n768 = n767 ^ n307 ;
  assign n709 = ~n667 & ~n696 ;
  assign n710 = n709 ^ n629 ;
  assign n798 = n710 ^ n188 ;
  assign n799 = n798 ^ n246 ;
  assign n802 = n768 & n799 ;
  assign n711 = n710 ^ n707 ;
  assign n772 = n802 ^ n711 ;
  assign n773 = ~n708 & n772 ;
  assign n774 = n773 ^ n203 ;
  assign n775 = n705 & ~n774 ;
  assign n776 = n775 ^ n704 ;
  assign n700 = n677 & ~n696 ;
  assign n701 = n700 ^ n623 ;
  assign n777 = n776 ^ n701 ;
  assign n778 = n776 ^ n138 ;
  assign n779 = n777 & n778 ;
  assign n781 = n4971 ^ n779 ;
  assign n784 = n699 & n781 ;
  assign n785 = n784 ^ n698 ;
  assign n786 = ~n691 & n785 ;
  assign n842 = n786 ^ n696 ;
  assign n843 = ~n839 & n842 ;
  assign n836 = x102 & ~n786 ;
  assign n840 = n839 ^ n836 ;
  assign n841 = ~x103 & ~n840 ;
  assign n844 = n843 ^ n841 ;
  assign n835 = n696 ^ n609 ;
  assign n845 = n844 ^ n835 ;
  assign n847 = n738 ^ n696 ;
  assign n848 = n786 & ~n847 ;
  assign n846 = n738 ^ x104 ;
  assign n849 = n848 ^ n846 ;
  assign n850 = n849 ^ n609 ;
  assign n851 = ~n845 & ~n850 ;
  assign n834 = n609 ^ n534 ;
  assign n852 = n851 ^ n834 ;
  assign n788 = n781 ^ n183 ;
  assign n791 = ~n691 & n788 ;
  assign n792 = n791 ^ n183 ;
  assign n793 = n698 & n792 ;
  assign n794 = n793 ^ n781 ;
  assign n795 = n774 & ~n786 ;
  assign n796 = n795 ^ n704 ;
  assign n797 = n796 ^ n138 ;
  assign n803 = n802 ^ n798 ;
  assign n804 = ~n786 & n803 ;
  assign n805 = n804 ^ n707 ;
  assign n806 = n805 ^ n157 ;
  assign n875 = ~n768 & ~n786 ;
  assign n876 = n875 ^ n710 ;
  assign n814 = n813 ^ n349 ;
  assign n815 = ~n786 & ~n814 ;
  assign n816 = n815 ^ n716 ;
  assign n817 = n816 ^ n245 ;
  assign n818 = ~n786 & n810 ;
  assign n819 = n818 ^ n760 ;
  assign n820 = n819 ^ n291 ;
  assign n830 = n740 ^ x105 ;
  assign n831 = n830 ^ n696 ;
  assign n827 = x104 & ~n696 ;
  assign n828 = n827 ^ n740 ;
  assign n829 = n786 & n828 ;
  assign n832 = n831 ^ n829 ;
  assign n833 = n832 ^ n534 ;
  assign n853 = ~n833 & ~n852 ;
  assign n854 = n853 ^ n750 ;
  assign n855 = n748 & ~n786 ;
  assign n856 = n855 ^ n736 ;
  assign n857 = n856 ^ n457 ;
  assign n858 = n854 & n857 ;
  assign n859 = n858 ^ n856 ;
  assign n821 = ~n751 & ~n786 ;
  assign n822 = n821 ^ n731 ;
  assign n860 = n859 ^ n822 ;
  assign n861 = n859 ^ n401 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = n862 ^ n401 ;
  assign n864 = n863 ^ n341 ;
  assign n865 = n753 ^ n401 ;
  assign n866 = ~n786 & ~n865 ;
  assign n867 = n866 ^ n720 ;
  assign n868 = n867 ^ n863 ;
  assign n869 = n864 & n868 ;
  assign n870 = n869 ^ n349 ;
  assign n871 = n820 & ~n870 ;
  assign n872 = n871 ^ n307 ;
  assign n873 = ~n817 & n872 ;
  assign n874 = n873 ^ n816 ;
  assign n877 = n876 ^ n874 ;
  assign n878 = n876 ^ n188 ;
  assign n879 = n877 & n878 ;
  assign n880 = n879 ^ n203 ;
  assign n881 = ~n806 & ~n880 ;
  assign n882 = n881 ^ n805 ;
  assign n883 = n882 ^ n796 ;
  assign n884 = n797 & n883 ;
  assign n885 = n884 ^ n138 ;
  assign n886 = n885 ^ n183 ;
  assign n887 = n778 & ~n786 ;
  assign n888 = n887 ^ n701 ;
  assign n889 = n888 ^ n885 ;
  assign n890 = ~n886 & ~n889 ;
  assign n891 = n890 ^ n885 ;
  assign n892 = ~n794 & ~n891 ;
  assign n903 = ~n852 & ~n892 ;
  assign n904 = n903 ^ n832 ;
  assign n905 = n904 ^ n457 ;
  assign n908 = ~x101 & n836 ;
  assign n909 = ~x102 & n696 ;
  assign n910 = n786 ^ x100 ;
  assign n913 = ~x101 & ~n910 ;
  assign n914 = n913 ^ n786 ;
  assign n915 = ~n892 & ~n914 ;
  assign n916 = n909 & n915 ;
  assign n917 = n916 ^ n696 ;
  assign n918 = n892 & n917 ;
  assign n919 = n908 & n918 ;
  assign n920 = n919 ^ n917 ;
  assign n921 = ~x98 & ~x99 ;
  assign n922 = ~x100 & n921 ;
  assign n923 = n920 & n922 ;
  assign n927 = n892 ^ n786 ;
  assign n930 = x101 & ~n927 ;
  assign n924 = n786 ^ x102 ;
  assign n931 = n930 ^ n924 ;
  assign n932 = n923 & n931 ;
  assign n933 = n932 ^ n920 ;
  assign n943 = n922 ^ n892 ;
  assign n944 = n922 ^ x101 ;
  assign n945 = ~n943 & ~n944 ;
  assign n946 = n945 ^ n922 ;
  assign n947 = n786 & ~n946 ;
  assign n934 = n892 ^ x101 ;
  assign n940 = ~n910 & n943 ;
  assign n935 = n892 ^ x100 ;
  assign n941 = n940 ^ n935 ;
  assign n942 = ~n934 & ~n941 ;
  assign n948 = n947 ^ n942 ;
  assign n953 = x102 & n948 ;
  assign n954 = n953 ^ n942 ;
  assign n955 = ~n933 & ~n954 ;
  assign n956 = n955 ^ n609 ;
  assign n958 = n839 ^ x103 ;
  assign n959 = n958 ^ n786 ;
  assign n957 = ~n840 & n892 ;
  assign n960 = n959 ^ n957 ;
  assign n961 = n960 ^ n955 ;
  assign n962 = n956 & n961 ;
  assign n963 = n962 ^ n609 ;
  assign n906 = ~n845 & ~n892 ;
  assign n907 = n906 ^ n849 ;
  assign n964 = n963 ^ n907 ;
  assign n965 = n963 ^ n534 ;
  assign n966 = n964 & ~n965 ;
  assign n967 = n966 ^ n750 ;
  assign n968 = n905 & n967 ;
  assign n969 = n968 ^ n904 ;
  assign n970 = n969 ^ n401 ;
  assign n971 = ~n854 & ~n892 ;
  assign n972 = n971 ^ n856 ;
  assign n973 = n972 ^ n969 ;
  assign n974 = ~n970 & ~n973 ;
  assign n975 = n974 ^ n462 ;
  assign n976 = ~n861 & ~n892 ;
  assign n977 = n976 ^ n822 ;
  assign n978 = n977 ^ n341 ;
  assign n979 = n975 & ~n978 ;
  assign n980 = n979 ^ n349 ;
  assign n1012 = ~n886 & ~n892 ;
  assign n1013 = n1012 ^ n888 ;
  assign n893 = n882 ^ n138 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = n894 ^ n796 ;
  assign n1014 = n895 ^ n183 ;
  assign n896 = n874 ^ n188 ;
  assign n897 = ~n892 & ~n896 ;
  assign n898 = n897 ^ n876 ;
  assign n899 = n898 ^ n157 ;
  assign n988 = ~n872 & ~n892 ;
  assign n989 = n988 ^ n816 ;
  assign n900 = n864 & ~n892 ;
  assign n901 = n900 ^ n867 ;
  assign n902 = n901 ^ n291 ;
  assign n981 = n902 & ~n980 ;
  assign n982 = n981 ^ n307 ;
  assign n983 = ~n870 & ~n892 ;
  assign n984 = n983 ^ n819 ;
  assign n985 = n984 ^ n245 ;
  assign n986 = n982 & ~n985 ;
  assign n987 = n986 ^ n984 ;
  assign n990 = n989 ^ n987 ;
  assign n991 = n989 ^ n188 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = n992 ^ n203 ;
  assign n994 = n899 & ~n993 ;
  assign n995 = n994 ^ n898 ;
  assign n996 = n995 ^ n138 ;
  assign n997 = n880 & ~n892 ;
  assign n998 = n997 ^ n805 ;
  assign n999 = n998 ^ n995 ;
  assign n1000 = n996 & n999 ;
  assign n1001 = n1000 ^ n138 ;
  assign n1031 = n1001 ^ n895 ;
  assign n1032 = ~n1014 & n1031 ;
  assign n1033 = n1032 ^ n895 ;
  assign n1034 = n1013 & ~n1033 ;
  assign n1044 = ~n980 & ~n1034 ;
  assign n1045 = n1044 ^ n901 ;
  assign n1046 = n1045 ^ n245 ;
  assign n1047 = ~n967 & ~n1034 ;
  assign n1048 = n1047 ^ n904 ;
  assign n1049 = n1048 ^ n401 ;
  assign n1050 = ~n965 & ~n1034 ;
  assign n1051 = n1050 ^ n907 ;
  assign n1052 = n1051 ^ n457 ;
  assign n1054 = ~x100 & ~n892 ;
  assign n1057 = n1054 ^ x101 ;
  assign n1053 = n927 ^ n922 ;
  assign n1055 = n1054 ^ n1053 ;
  assign n1056 = ~n1034 & n1055 ;
  assign n1058 = n1057 ^ n1056 ;
  assign n1059 = n1058 ^ n696 ;
  assign n1072 = n1034 ^ n892 ;
  assign n1160 = n1034 ^ x99 ;
  assign n1075 = ~n1072 & n1160 ;
  assign n1060 = n892 ^ x99 ;
  assign n1061 = n1060 ^ n1034 ;
  assign n1062 = ~x96 & ~x97 ;
  assign n1063 = n1062 ^ x98 ;
  assign n1064 = n1063 ^ n892 ;
  assign n1065 = ~n1061 & ~n1064 ;
  assign n1066 = n1065 ^ n927 ;
  assign n1067 = n1066 ^ x99 ;
  assign n1068 = n1067 ^ n786 ;
  assign n1076 = n1075 ^ n1068 ;
  assign n1077 = x98 & n1076 ;
  assign n1078 = n1077 ^ n1066 ;
  assign n1081 = n921 ^ x100 ;
  assign n1079 = n921 ^ n892 ;
  assign n1080 = n1034 & ~n1079 ;
  assign n1082 = n1081 ^ n1080 ;
  assign n1085 = n1082 ^ n786 ;
  assign n1086 = ~n1078 & n1085 ;
  assign n1083 = n1082 ^ n696 ;
  assign n1087 = n1086 ^ n1083 ;
  assign n1088 = n1059 & n1087 ;
  assign n1089 = n1088 ^ n835 ;
  assign n1093 = n948 ^ n696 ;
  assign n1094 = ~n1034 & n1093 ;
  assign n1090 = n837 ^ n786 ;
  assign n1091 = ~n892 & ~n1090 ;
  assign n1092 = n1091 ^ n924 ;
  assign n1095 = n1094 ^ n1092 ;
  assign n1096 = n1095 ^ n609 ;
  assign n1097 = ~n1089 & n1096 ;
  assign n1098 = n1097 ^ n834 ;
  assign n1099 = n956 & ~n1034 ;
  assign n1100 = n1099 ^ n960 ;
  assign n1101 = n1100 ^ n534 ;
  assign n1102 = ~n1098 & n1101 ;
  assign n1103 = n1102 ^ n750 ;
  assign n1104 = ~n1052 & n1103 ;
  assign n1105 = n1104 ^ n1051 ;
  assign n1106 = n1105 ^ n1048 ;
  assign n1107 = ~n1049 & n1106 ;
  assign n1108 = n1107 ^ n401 ;
  assign n1109 = n1108 ^ n341 ;
  assign n1110 = ~n970 & ~n1034 ;
  assign n1111 = n1110 ^ n972 ;
  assign n1112 = n1111 ^ n1108 ;
  assign n1113 = n1109 & n1112 ;
  assign n1114 = n1113 ^ n349 ;
  assign n1115 = n975 & ~n1034 ;
  assign n1116 = n1115 ^ n977 ;
  assign n1117 = n1116 ^ n291 ;
  assign n1118 = ~n1114 & n1117 ;
  assign n1119 = n1118 ^ n307 ;
  assign n1120 = ~n1046 & n1119 ;
  assign n1121 = n1120 ^ n1045 ;
  assign n1042 = ~n982 & ~n1034 ;
  assign n1043 = n1042 ^ n984 ;
  assign n1122 = n1121 ^ n1043 ;
  assign n1123 = n1121 ^ n188 ;
  assign n1124 = ~n1122 & ~n1123 ;
  assign n1125 = n1124 ^ n203 ;
  assign n1025 = n995 & n1003 ;
  assign n1026 = n1013 & n1025 ;
  assign n1015 = n1014 ^ n1013 ;
  assign n1020 = n998 & n1013 ;
  assign n1021 = n1020 ^ n1001 ;
  assign n1022 = n1015 & ~n1021 ;
  assign n1023 = n1022 ^ n1013 ;
  assign n1027 = n1026 ^ n1023 ;
  assign n1002 = n1001 ^ n183 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1355 = n1003 ^ n183 ;
  assign n4969 = n1355 ^ n137 ;
  assign n4970 = n4969 ^ x127 ;
  assign n1008 = n4970 ^ n1002 ;
  assign n1009 = ~n999 & ~n1008 ;
  assign n1010 = n1009 ^ n1002 ;
  assign n1011 = ~n1004 & ~n1010 ;
  assign n1028 = n1027 ^ n1011 ;
  assign n1029 = n895 & n1028 ;
  assign n1030 = n1029 ^ n1027 ;
  assign n1035 = n993 & ~n1034 ;
  assign n1036 = n1035 ^ n898 ;
  assign n1037 = n1036 ^ n138 ;
  assign n1038 = n987 ^ n188 ;
  assign n1039 = ~n1034 & ~n1038 ;
  assign n1040 = n1039 ^ n989 ;
  assign n1041 = n1040 ^ n157 ;
  assign n1126 = ~n1041 & ~n1125 ;
  assign n1127 = n1126 ^ n1040 ;
  assign n1128 = n1127 ^ n1036 ;
  assign n1129 = n1037 & n1128 ;
  assign n1130 = n1129 ^ n138 ;
  assign n1131 = n1030 & n1130 ;
  assign n1132 = n996 & ~n1034 ;
  assign n1133 = n1132 ^ n998 ;
  assign n1134 = n1133 ^ n183 ;
  assign n1135 = n1131 & n1134 ;
  assign n1136 = n1135 ^ n1030 ;
  assign n1170 = n1125 & ~n1136 ;
  assign n1171 = n1170 ^ n1040 ;
  assign n1172 = n138 & ~n1171 ;
  assign n1222 = ~n1123 & ~n1136 ;
  assign n1223 = n1222 ^ n1043 ;
  assign n1173 = n1109 & ~n1136 ;
  assign n1174 = n1173 ^ n1111 ;
  assign n1175 = n1174 ^ n291 ;
  assign n1202 = n1105 ^ n401 ;
  assign n1203 = ~n1136 & n1202 ;
  assign n1204 = n1203 ^ n1048 ;
  assign n1176 = ~n1103 & ~n1136 ;
  assign n1177 = n1176 ^ n1051 ;
  assign n1178 = n1177 ^ n401 ;
  assign n1179 = ~n1089 & ~n1136 ;
  assign n1180 = n1179 ^ n1095 ;
  assign n1181 = n1180 ^ n534 ;
  assign n1137 = n1136 ^ x97 ;
  assign n787 = ~x94 & ~x95 ;
  assign n1138 = n1137 ^ n787 ;
  assign n1139 = n1034 ^ n787 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1149 = n1140 ^ n1072 ;
  assign n1143 = n1136 ^ n1034 ;
  assign n1146 = ~n1137 & n1143 ;
  assign n1147 = n1146 ^ n1140 ;
  assign n1148 = x96 & n1147 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1151 = n1062 ^ n1034 ;
  assign n1152 = n1136 & ~n1151 ;
  assign n1153 = n1152 ^ n1062 ;
  assign n1154 = n1153 ^ x98 ;
  assign n1157 = n1154 ^ n892 ;
  assign n1158 = ~n1150 & n1157 ;
  assign n1155 = n1154 ^ n786 ;
  assign n1159 = n1158 ^ n1155 ;
  assign n1164 = x98 & n1153 ;
  assign n1161 = n1062 ^ n892 ;
  assign n1162 = ~n1136 & ~n1161 ;
  assign n1163 = n1162 ^ n1160 ;
  assign n1165 = n1164 ^ n1163 ;
  assign n1166 = n1165 ^ n696 ;
  assign n1167 = n1166 ^ n842 ;
  assign n1168 = ~n1159 & ~n1167 ;
  assign n1169 = n1168 ^ n1166 ;
  assign n1182 = n1078 & ~n1136 ;
  assign n1183 = n1182 ^ n1082 ;
  assign n1184 = n1183 ^ n696 ;
  assign n1185 = ~n1169 & n1184 ;
  assign n1186 = n1185 ^ n835 ;
  assign n1187 = n1087 & ~n1136 ;
  assign n1188 = n1187 ^ n1058 ;
  assign n1189 = n1188 ^ n609 ;
  assign n1190 = ~n1186 & ~n1189 ;
  assign n1191 = n1190 ^ n834 ;
  assign n1192 = ~n1181 & ~n1191 ;
  assign n1193 = n1192 ^ n750 ;
  assign n1194 = ~n1098 & ~n1136 ;
  assign n1195 = n1194 ^ n1100 ;
  assign n1196 = n1195 ^ n457 ;
  assign n1197 = ~n1193 & ~n1196 ;
  assign n1198 = n1197 ^ n457 ;
  assign n1199 = n1198 ^ n1177 ;
  assign n1200 = n1178 & n1199 ;
  assign n1201 = n1200 ^ n401 ;
  assign n1205 = n1204 ^ n1201 ;
  assign n1206 = n1204 ^ n341 ;
  assign n1207 = n1205 & ~n1206 ;
  assign n1208 = n1207 ^ n349 ;
  assign n1209 = n1175 & ~n1208 ;
  assign n1210 = n1209 ^ n307 ;
  assign n1211 = ~n1114 & ~n1136 ;
  assign n1212 = n1211 ^ n1116 ;
  assign n1213 = n1212 ^ n245 ;
  assign n1214 = n1210 & ~n1213 ;
  assign n1215 = n1214 ^ n1212 ;
  assign n1216 = n1215 ^ n188 ;
  assign n1217 = ~n1119 & ~n1136 ;
  assign n1218 = n1217 ^ n1045 ;
  assign n1219 = n1218 ^ n1215 ;
  assign n1220 = ~n1216 & ~n1219 ;
  assign n1221 = n1220 ^ n188 ;
  assign n1224 = n1223 ^ n1221 ;
  assign n1225 = n1221 ^ n157 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1227 = n1226 ^ n1223 ;
  assign n1229 = n1171 & n1227 ;
  assign n1228 = n1227 ^ n1171 ;
  assign n1230 = n1229 ^ n1228 ;
  assign n1231 = n138 & ~n1227 ;
  assign n1243 = n1040 ^ n1036 ;
  assign n1245 = n138 & ~n1243 ;
  assign n1246 = n1245 ^ n1036 ;
  assign n1247 = n1127 & ~n1246 ;
  assign n1248 = n1247 ^ n138 ;
  assign n1256 = n1030 & ~n1036 ;
  assign n1232 = ~n1030 & n1133 ;
  assign n1249 = ~n138 & ~n1232 ;
  assign n1257 = n1256 ^ n1249 ;
  assign n1258 = ~n1248 & n1257 ;
  assign n1233 = n1232 ^ n1133 ;
  assign n1234 = n1130 & ~n1233 ;
  assign n1235 = n1234 ^ n1133 ;
  assign n1250 = n1249 ^ n1235 ;
  assign n1259 = n1258 ^ n1250 ;
  assign n1236 = n1136 ^ n1127 ;
  assign n1237 = n1036 & n1236 ;
  assign n1238 = n1237 ^ n1127 ;
  assign n1239 = n1127 ^ n1037 ;
  assign n1240 = ~n1238 & n1239 ;
  assign n1241 = n1133 & ~n1172 ;
  assign n1242 = n1240 & n1241 ;
  assign n1260 = n1259 ^ n1242 ;
  assign n1261 = ~n183 & n1260 ;
  assign n1262 = n1261 ^ n1235 ;
  assign n1263 = n183 & n1235 ;
  assign n1264 = ~n1240 & n1263 ;
  assign n1266 = ~n1036 & n1127 ;
  assign n1265 = n1238 ^ n1136 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1268 = n1264 & ~n1267 ;
  assign n1269 = n1268 ^ n1263 ;
  assign n1270 = n1262 & ~n1269 ;
  assign n1271 = n1231 & n1270 ;
  assign n1272 = n1271 ^ n1262 ;
  assign n1273 = ~n1230 & n1272 ;
  assign n1278 = n1263 & n1266 ;
  assign n1279 = n1278 ^ n1269 ;
  assign n1280 = n1273 & ~n1279 ;
  assign n1281 = n1280 ^ n1272 ;
  assign n1282 = n1172 & n1281 ;
  assign n1287 = n1127 & n1136 ;
  assign n1288 = n1287 ^ n1128 ;
  assign n1289 = n1282 & n1288 ;
  assign n1290 = n1289 ^ n1281 ;
  assign n1351 = n1227 ^ n138 ;
  assign n1352 = ~n1290 & ~n1351 ;
  assign n1353 = n1352 ^ n1171 ;
  assign n1354 = n1353 ^ n183 ;
  assign n1365 = n138 & ~n1229 ;
  assign n1366 = n1365 ^ n1230 ;
  assign n1374 = n1290 & ~n1365 ;
  assign n1371 = n1365 ^ n183 ;
  assign n1357 = n1127 ^ n138 ;
  assign n1358 = ~n1136 & ~n1357 ;
  assign n1359 = n1358 ^ n1036 ;
  assign n1367 = n1359 ^ n1230 ;
  assign n1368 = ~n183 & n1367 ;
  assign n1372 = n1371 ^ n1368 ;
  assign n1369 = n1171 & n1368 ;
  assign n1370 = n1272 & n1369 ;
  assign n1373 = n1372 ^ n1370 ;
  assign n1375 = n1374 ^ n1373 ;
  assign n1376 = n1366 & n1375 ;
  assign n1362 = n1290 ^ n183 ;
  assign n1363 = n1362 ^ n1359 ;
  assign n1356 = n1229 & ~n1355 ;
  assign n1360 = ~n1262 & n1359 ;
  assign n1361 = n1356 & n1360 ;
  assign n1364 = n1363 ^ n1361 ;
  assign n1377 = n1376 ^ n1364 ;
  assign n1378 = n1225 & ~n1290 ;
  assign n1379 = n1378 ^ n1223 ;
  assign n1380 = n1379 ^ n138 ;
  assign n1383 = ~n1210 & ~n1290 ;
  assign n1384 = n1383 ^ n1212 ;
  assign n1385 = n1384 ^ n188 ;
  assign n1386 = n1201 ^ n341 ;
  assign n1387 = ~n1290 & n1386 ;
  assign n1388 = n1387 ^ n1204 ;
  assign n1389 = n1388 ^ n291 ;
  assign n1291 = ~n1169 & ~n1290 ;
  assign n1292 = n1291 ^ n1183 ;
  assign n1293 = n1292 ^ n609 ;
  assign n1297 = n1136 ^ n787 ;
  assign n1300 = ~x96 & ~n1297 ;
  assign n1301 = n1300 ^ n1143 ;
  assign n1302 = ~n1290 & n1301 ;
  assign n1303 = n1302 ^ x97 ;
  assign n1294 = ~x96 & ~n1136 ;
  assign n1304 = n1303 ^ n1294 ;
  assign n1305 = n1304 ^ n892 ;
  assign n1306 = ~x92 & ~x93 ;
  assign n1307 = n1306 ^ x94 ;
  assign n1308 = n1307 ^ n1136 ;
  assign n1309 = n1307 ^ x95 ;
  assign n1310 = n1309 ^ n1290 ;
  assign n1311 = ~n1308 & ~n1310 ;
  assign n1321 = n1311 ^ n1143 ;
  assign n1312 = n1311 ^ n1290 ;
  assign n1313 = n1312 ^ x95 ;
  assign n1314 = n1313 ^ n1311 ;
  assign n1315 = n1311 ^ n1136 ;
  assign n1316 = n1315 ^ n1290 ;
  assign n1317 = n1316 ^ n1311 ;
  assign n1318 = ~n1314 & n1317 ;
  assign n1319 = n1318 ^ n1311 ;
  assign n1320 = x94 & n1319 ;
  assign n1322 = n1321 ^ n1320 ;
  assign n1324 = n1136 ^ x96 ;
  assign n1323 = ~n1290 & ~n1297 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1326 = n1325 ^ n1034 ;
  assign n1327 = n1322 & ~n1326 ;
  assign n1328 = n1327 ^ n1072 ;
  assign n1329 = n1305 & n1328 ;
  assign n1330 = n1329 ^ n927 ;
  assign n1331 = n1150 & ~n1290 ;
  assign n1332 = n1331 ^ n1154 ;
  assign n1335 = n1332 ^ n786 ;
  assign n1336 = ~n1330 & n1335 ;
  assign n1333 = n1332 ^ n696 ;
  assign n1337 = n1336 ^ n1333 ;
  assign n1338 = n1159 & ~n1290 ;
  assign n1339 = n1338 ^ n1165 ;
  assign n1340 = n1339 ^ n609 ;
  assign n1341 = n1340 ^ n835 ;
  assign n1342 = ~n1337 & ~n1341 ;
  assign n1343 = n1342 ^ n1340 ;
  assign n1344 = ~n1293 & n1343 ;
  assign n1345 = n1344 ^ n834 ;
  assign n1346 = ~n1186 & ~n1290 ;
  assign n1347 = n1346 ^ n1188 ;
  assign n1348 = n1347 ^ n534 ;
  assign n1349 = ~n1345 & n1348 ;
  assign n1350 = n1349 ^ n750 ;
  assign n1393 = ~n1191 & ~n1290 ;
  assign n1394 = n1393 ^ n1180 ;
  assign n1395 = n1394 ^ n457 ;
  assign n1396 = n1350 & n1395 ;
  assign n1397 = n1396 ^ n1394 ;
  assign n1398 = n1397 ^ n401 ;
  assign n1399 = ~n1193 & ~n1290 ;
  assign n1400 = n1399 ^ n1195 ;
  assign n1401 = n1400 ^ n1397 ;
  assign n1402 = ~n1398 & n1401 ;
  assign n1403 = n1402 ^ n401 ;
  assign n1390 = n1198 ^ n401 ;
  assign n1391 = ~n1290 & ~n1390 ;
  assign n1392 = n1391 ^ n1177 ;
  assign n1404 = n1403 ^ n1392 ;
  assign n1405 = n1403 ^ n341 ;
  assign n1406 = ~n1404 & n1405 ;
  assign n1407 = n1406 ^ n349 ;
  assign n1408 = n1389 & ~n1407 ;
  assign n1409 = n1408 ^ n307 ;
  assign n1410 = ~n1208 & ~n1290 ;
  assign n1411 = n1410 ^ n1174 ;
  assign n1412 = n1411 ^ n245 ;
  assign n1413 = n1409 & ~n1412 ;
  assign n1414 = n1413 ^ n1411 ;
  assign n1415 = n1414 ^ n1384 ;
  assign n1416 = ~n1385 & ~n1415 ;
  assign n1417 = n1416 ^ n188 ;
  assign n1381 = ~n1216 & ~n1290 ;
  assign n1382 = n1381 ^ n1218 ;
  assign n1418 = n1417 ^ n1382 ;
  assign n1419 = n1382 ^ n157 ;
  assign n1420 = ~n1418 & n1419 ;
  assign n1421 = n1420 ^ n1417 ;
  assign n1422 = n1421 ^ n1379 ;
  assign n1423 = ~n1380 & n1422 ;
  assign n1424 = n1423 ^ n138 ;
  assign n1425 = ~n1377 & n1424 ;
  assign n1426 = n1354 & n1425 ;
  assign n1427 = n1426 ^ n1377 ;
  assign n1509 = n1417 ^ n157 ;
  assign n1510 = n1427 & n1509 ;
  assign n1511 = n1510 ^ n1382 ;
  assign n1512 = n1003 & ~n1511 ;
  assign n1521 = n138 & n1421 ;
  assign n1520 = n1421 ^ n138 ;
  assign n1522 = n1521 ^ n1520 ;
  assign n1523 = n1522 ^ n1353 ;
  assign n1524 = n1427 & ~n1521 ;
  assign n1525 = n1524 ^ n1521 ;
  assign n1526 = n1522 & n1524 ;
  assign n1527 = n1526 ^ n1379 ;
  assign n1528 = ~n183 & n1527 ;
  assign n1529 = n1525 & n1528 ;
  assign n1530 = n1523 & n1529 ;
  assign n1531 = n1530 ^ n1528 ;
  assign n1532 = n1531 ^ n183 ;
  assign n1535 = n1512 & n1532 ;
  assign n1513 = n1424 ^ n1353 ;
  assign n1514 = n1424 ^ n183 ;
  assign n1517 = ~n1377 & ~n1514 ;
  assign n1518 = n1517 ^ n183 ;
  assign n1519 = ~n1513 & n1518 ;
  assign n1533 = n1532 ^ n1519 ;
  assign n1536 = n1535 ^ n1533 ;
  assign n1537 = n1414 ^ n188 ;
  assign n1538 = n1427 & ~n1537 ;
  assign n1539 = n1538 ^ n1384 ;
  assign n1540 = n1539 ^ n157 ;
  assign n1541 = ~n1407 & n1427 ;
  assign n1542 = n1541 ^ n1388 ;
  assign n1543 = n1542 ^ n245 ;
  assign n1428 = ~n1350 & n1427 ;
  assign n1429 = n1428 ^ n1394 ;
  assign n1430 = n1429 ^ n401 ;
  assign n1431 = ~n1345 & n1427 ;
  assign n1432 = n1431 ^ n1347 ;
  assign n1433 = n1432 ^ n457 ;
  assign n1434 = n1343 & n1427 ;
  assign n1435 = n1434 ^ n1292 ;
  assign n1436 = n1435 ^ n534 ;
  assign n1437 = n1337 & n1427 ;
  assign n1438 = n1437 ^ n1339 ;
  assign n1439 = n1438 ^ n609 ;
  assign n1440 = n1306 ^ n1290 ;
  assign n1441 = ~n1427 & ~n1440 ;
  assign n1442 = n1441 ^ n1307 ;
  assign n1443 = n1442 ^ n1136 ;
  assign n1445 = n1427 ^ x93 ;
  assign n1450 = n1427 ^ n1290 ;
  assign n1451 = n1445 & ~n1450 ;
  assign n1452 = n1451 ^ n1136 ;
  assign n1453 = n1452 ^ n1290 ;
  assign n1449 = n1445 ^ n1136 ;
  assign n1454 = n1453 ^ n1449 ;
  assign n1444 = ~x90 & ~x91 ;
  assign n1446 = n1445 ^ n1444 ;
  assign n1447 = n1444 ^ n1290 ;
  assign n1448 = ~n1446 & n1447 ;
  assign n1455 = n1454 ^ n1448 ;
  assign n1456 = ~x92 & n1455 ;
  assign n1457 = n1456 ^ n1453 ;
  assign n1458 = n1443 & n1457 ;
  assign n1459 = n1458 ^ n1143 ;
  assign n1461 = n1290 ^ n1136 ;
  assign n1462 = n1461 ^ n1440 ;
  assign n1463 = n1462 ^ n1461 ;
  assign n1464 = n1461 ^ x94 ;
  assign n1465 = n1464 ^ n1461 ;
  assign n1466 = ~n1463 & ~n1465 ;
  assign n1467 = n1466 ^ n1461 ;
  assign n1468 = n1427 & n1467 ;
  assign n1469 = n1468 ^ x95 ;
  assign n1460 = ~x94 & ~n1290 ;
  assign n1470 = n1469 ^ n1460 ;
  assign n1473 = n1470 ^ n1034 ;
  assign n1474 = ~n1459 & n1473 ;
  assign n1471 = n1470 ^ n892 ;
  assign n1475 = n1474 ^ n1471 ;
  assign n1476 = n1322 & n1427 ;
  assign n1477 = n1476 ^ n1325 ;
  assign n1478 = n1477 ^ n892 ;
  assign n1479 = n1475 & ~n1478 ;
  assign n1480 = n1479 ^ n927 ;
  assign n1481 = n1328 & n1427 ;
  assign n1482 = n1481 ^ n1304 ;
  assign n1485 = n1482 ^ n786 ;
  assign n1486 = ~n1480 & n1485 ;
  assign n1483 = n1482 ^ n696 ;
  assign n1487 = n1486 ^ n1483 ;
  assign n1488 = n1330 & n1427 ;
  assign n1489 = n1488 ^ n1332 ;
  assign n1490 = n1489 ^ n609 ;
  assign n1491 = n1490 ^ n835 ;
  assign n1492 = ~n1487 & n1491 ;
  assign n1493 = n1492 ^ n1490 ;
  assign n1494 = n1439 & ~n1493 ;
  assign n1495 = n1494 ^ n834 ;
  assign n1496 = n1436 & ~n1495 ;
  assign n1497 = n1496 ^ n750 ;
  assign n1498 = ~n1433 & n1497 ;
  assign n1499 = n1498 ^ n1432 ;
  assign n1500 = n1499 ^ n1429 ;
  assign n1501 = ~n1430 & n1500 ;
  assign n1502 = n1501 ^ n401 ;
  assign n1503 = n1502 ^ n341 ;
  assign n1504 = ~n1398 & n1427 ;
  assign n1505 = n1504 ^ n1400 ;
  assign n1506 = n1505 ^ n1502 ;
  assign n1507 = n1503 & ~n1506 ;
  assign n1508 = n1507 ^ n349 ;
  assign n1544 = n1405 & n1427 ;
  assign n1545 = n1544 ^ n1392 ;
  assign n1546 = n1545 ^ n291 ;
  assign n1547 = ~n1508 & ~n1546 ;
  assign n1548 = n1547 ^ n307 ;
  assign n1549 = ~n1543 & n1548 ;
  assign n1550 = n1549 ^ n1542 ;
  assign n1551 = n1550 ^ n188 ;
  assign n1552 = ~n1409 & n1427 ;
  assign n1553 = n1552 ^ n1411 ;
  assign n1554 = n1553 ^ n1550 ;
  assign n1555 = ~n1551 & ~n1554 ;
  assign n1556 = n1555 ^ n203 ;
  assign n1557 = ~n1540 & ~n1556 ;
  assign n1558 = n1557 ^ n1539 ;
  assign n1559 = n1511 & n1558 ;
  assign n1560 = n1558 ^ n1511 ;
  assign n1561 = n1560 ^ n1559 ;
  assign n1562 = ~n138 & n1561 ;
  assign n1563 = ~n1559 & ~n1562 ;
  assign n1564 = n1536 & n1563 ;
  assign n1569 = ~n183 & ~n1558 ;
  assign n1570 = n1569 ^ n1527 ;
  assign n1571 = n1564 & ~n1570 ;
  assign n1572 = n1571 ^ n1536 ;
  assign n1716 = n1558 ^ n138 ;
  assign n1717 = ~n1572 & ~n1716 ;
  assign n1718 = n1717 ^ n1511 ;
  assign n1719 = n1718 ^ n183 ;
  assign n1565 = n1527 ^ n183 ;
  assign n1696 = n1565 ^ n1563 ;
  assign n1567 = n1558 ^ n1527 ;
  assign n1675 = n1567 ^ n1511 ;
  assign n1676 = n1675 ^ n1558 ;
  assign n1677 = n1558 ^ n1536 ;
  assign n1678 = ~n1511 & n1677 ;
  assign n1679 = n1678 ^ n1558 ;
  assign n1680 = n1676 & ~n1679 ;
  assign n1681 = n1680 ^ n1558 ;
  assign n1682 = n1003 & ~n1681 ;
  assign n1683 = n1682 ^ n1003 ;
  assign n1684 = n1536 ^ n183 ;
  assign n1685 = n1684 ^ n1527 ;
  assign n1686 = n1685 ^ n183 ;
  assign n1689 = n1559 & ~n1686 ;
  assign n1690 = n1689 ^ n183 ;
  assign n1691 = ~n1683 & ~n1690 ;
  assign n1693 = n1527 & ~n1562 ;
  assign n1694 = n1691 & n1693 ;
  assign n1692 = n1691 ^ n1683 ;
  assign n1695 = n1694 ^ n1692 ;
  assign n1697 = n1696 ^ n1695 ;
  assign n1700 = n1697 ^ n1536 ;
  assign n1706 = n1700 ^ n1697 ;
  assign n1707 = ~n1527 & n1706 ;
  assign n1698 = n1697 ^ n1696 ;
  assign n1699 = n1698 ^ n1536 ;
  assign n1708 = n1707 ^ n1699 ;
  assign n1709 = n1697 ^ n1511 ;
  assign n1712 = ~n1698 & n1709 ;
  assign n1713 = n1712 ^ n1511 ;
  assign n1714 = ~n1708 & n1713 ;
  assign n1715 = n1714 ^ n1698 ;
  assign n1720 = n1556 & ~n1572 ;
  assign n1721 = n1720 ^ n1539 ;
  assign n1722 = n1721 ^ n138 ;
  assign n1723 = ~n1551 & ~n1572 ;
  assign n1724 = n1723 ^ n1553 ;
  assign n1725 = n1724 ^ n157 ;
  assign n1573 = ~n1508 & ~n1572 ;
  assign n1574 = n1573 ^ n1545 ;
  assign n1575 = n1574 ^ n245 ;
  assign n1576 = n1499 ^ n401 ;
  assign n1577 = ~n1572 & n1576 ;
  assign n1578 = n1577 ^ n1429 ;
  assign n1579 = n1578 ^ n341 ;
  assign n1580 = ~n1497 & ~n1572 ;
  assign n1581 = n1580 ^ n1432 ;
  assign n1582 = n1581 ^ n401 ;
  assign n1583 = ~n1495 & ~n1572 ;
  assign n1584 = n1583 ^ n1435 ;
  assign n1585 = n1584 ^ n457 ;
  assign n1586 = n1487 & ~n1572 ;
  assign n1587 = n1586 ^ n1489 ;
  assign n1588 = n1587 ^ n609 ;
  assign n1598 = ~x92 & n1427 ;
  assign n1589 = n1450 ^ x92 ;
  assign n1590 = n1589 ^ n1450 ;
  assign n1591 = n1444 ^ n1427 ;
  assign n1594 = ~n1590 & n1591 ;
  assign n1595 = n1594 ^ n1450 ;
  assign n1596 = ~n1572 & ~n1595 ;
  assign n1597 = n1596 ^ x93 ;
  assign n1599 = n1598 ^ n1597 ;
  assign n1600 = n1599 ^ n1136 ;
  assign n1620 = n1427 ^ x92 ;
  assign n1619 = ~n1572 & n1591 ;
  assign n1621 = n1620 ^ n1619 ;
  assign n1624 = n1621 ^ n1136 ;
  assign n1603 = ~x88 & ~x89 ;
  assign n1602 = n1427 ^ x90 ;
  assign n1604 = n1603 ^ n1602 ;
  assign n1605 = n1572 ^ n1427 ;
  assign n1606 = n1605 ^ x91 ;
  assign n1607 = n1604 & n1606 ;
  assign n1608 = n1607 ^ n1450 ;
  assign n1601 = n1290 ^ x91 ;
  assign n1609 = n1608 ^ n1601 ;
  assign n1610 = n1609 ^ n1572 ;
  assign n1611 = n1610 ^ x91 ;
  assign n1612 = n1611 ^ n1609 ;
  assign n1613 = n1609 ^ n1605 ;
  assign n1614 = n1613 ^ n1609 ;
  assign n1615 = n1612 & n1614 ;
  assign n1616 = n1615 ^ n1609 ;
  assign n1617 = x90 & ~n1616 ;
  assign n1618 = n1617 ^ n1608 ;
  assign n1622 = n1621 ^ n1290 ;
  assign n1623 = n1618 & n1622 ;
  assign n1625 = n1624 ^ n1623 ;
  assign n1626 = n1600 & n1625 ;
  assign n1627 = n1626 ^ n1143 ;
  assign n1628 = n1457 & ~n1572 ;
  assign n1629 = n1628 ^ n1442 ;
  assign n1632 = n1629 ^ n1034 ;
  assign n1633 = ~n1627 & n1632 ;
  assign n1630 = n1629 ^ n892 ;
  assign n1634 = n1633 ^ n1630 ;
  assign n1635 = n1459 & ~n1572 ;
  assign n1636 = n1635 ^ n1470 ;
  assign n1637 = n1636 ^ n786 ;
  assign n1638 = n1637 ^ n927 ;
  assign n1639 = ~n1634 & n1638 ;
  assign n1640 = n1639 ^ n1637 ;
  assign n1641 = n1475 & ~n1572 ;
  assign n1642 = n1641 ^ n1477 ;
  assign n1643 = n1642 ^ n786 ;
  assign n1644 = n1640 & ~n1643 ;
  assign n1645 = n1644 ^ n842 ;
  assign n1646 = n1480 & ~n1572 ;
  assign n1647 = n1646 ^ n1482 ;
  assign n1650 = n1647 ^ n696 ;
  assign n1651 = ~n1645 & n1650 ;
  assign n1648 = n1647 ^ n609 ;
  assign n1652 = n1651 ^ n1648 ;
  assign n1653 = ~n1588 & ~n1652 ;
  assign n1654 = n1653 ^ n834 ;
  assign n1655 = ~n1493 & ~n1572 ;
  assign n1656 = n1655 ^ n1438 ;
  assign n1657 = n1656 ^ n534 ;
  assign n1658 = ~n1654 & ~n1657 ;
  assign n1659 = n1658 ^ n750 ;
  assign n1660 = ~n1585 & n1659 ;
  assign n1661 = n1660 ^ n1584 ;
  assign n1662 = n1661 ^ n1581 ;
  assign n1663 = n1582 & ~n1662 ;
  assign n1664 = n1663 ^ n462 ;
  assign n1665 = ~n1579 & n1664 ;
  assign n1666 = n1665 ^ n349 ;
  assign n1667 = n1503 & ~n1572 ;
  assign n1668 = n1667 ^ n1505 ;
  assign n1669 = n1668 ^ n291 ;
  assign n1670 = ~n1666 & ~n1669 ;
  assign n1671 = n1670 ^ n307 ;
  assign n1672 = n1575 & n1671 ;
  assign n1673 = n1672 ^ n1574 ;
  assign n1674 = n1673 ^ n188 ;
  assign n1726 = ~n1548 & ~n1572 ;
  assign n1727 = n1726 ^ n1542 ;
  assign n1728 = n1727 ^ n1673 ;
  assign n1729 = n1674 & n1728 ;
  assign n1730 = n1729 ^ n188 ;
  assign n1731 = n1730 ^ n1724 ;
  assign n1732 = n1725 & ~n1731 ;
  assign n1733 = n1732 ^ n1730 ;
  assign n1734 = n1733 ^ n1721 ;
  assign n1735 = ~n1722 & n1734 ;
  assign n1736 = n1735 ^ n138 ;
  assign n1737 = ~n1715 & n1736 ;
  assign n1738 = n1719 & n1737 ;
  assign n1739 = n1738 ^ n1715 ;
  assign n1745 = n1661 ^ n401 ;
  assign n1746 = n1739 & n1745 ;
  assign n1747 = n1746 ^ n1581 ;
  assign n1748 = n1747 ^ n341 ;
  assign n1829 = ~n1659 & n1739 ;
  assign n1830 = n1829 ^ n1584 ;
  assign n1749 = ~n1654 & n1739 ;
  assign n1750 = n1749 ^ n1656 ;
  assign n1751 = n1750 ^ n457 ;
  assign n1752 = ~n1652 & n1739 ;
  assign n1753 = n1752 ^ n1587 ;
  assign n1754 = n1753 ^ n534 ;
  assign n1756 = ~x86 & ~x87 ;
  assign n1757 = n1756 ^ x88 ;
  assign n1755 = n1739 ^ x89 ;
  assign n1758 = n1757 ^ n1755 ;
  assign n1759 = n1755 ^ n1572 ;
  assign n1760 = n1758 & n1759 ;
  assign n1769 = n1760 ^ n1605 ;
  assign n1763 = n1739 ^ n1572 ;
  assign n1766 = n1755 & ~n1763 ;
  assign n1767 = n1766 ^ n1760 ;
  assign n1768 = x88 & n1767 ;
  assign n1770 = n1769 ^ n1768 ;
  assign n1772 = n1603 ^ n1572 ;
  assign n1773 = ~n1739 & ~n1772 ;
  assign n1771 = n1603 ^ x90 ;
  assign n1774 = n1773 ^ n1771 ;
  assign n1775 = n1774 ^ n1427 ;
  assign n1776 = ~n1770 & ~n1775 ;
  assign n1777 = n1776 ^ n1450 ;
  assign n1786 = ~x90 & ~n1572 ;
  assign n1780 = n1605 ^ x90 ;
  assign n1781 = n1780 ^ n1605 ;
  assign n1782 = ~n1772 & ~n1781 ;
  assign n1783 = n1782 ^ n1605 ;
  assign n1784 = n1739 & ~n1783 ;
  assign n1785 = n1784 ^ x91 ;
  assign n1787 = n1786 ^ n1785 ;
  assign n1788 = n1787 ^ n1290 ;
  assign n1789 = ~n1777 & n1788 ;
  assign n1790 = n1789 ^ n1461 ;
  assign n1791 = ~n1618 & n1739 ;
  assign n1792 = n1791 ^ n1621 ;
  assign n1793 = n1792 ^ n1136 ;
  assign n1794 = n1790 & n1793 ;
  assign n1795 = n1794 ^ n1143 ;
  assign n1796 = n1625 & n1739 ;
  assign n1797 = n1796 ^ n1599 ;
  assign n1800 = n1797 ^ n1034 ;
  assign n1801 = ~n1795 & n1800 ;
  assign n1798 = n1797 ^ n892 ;
  assign n1802 = n1801 ^ n1798 ;
  assign n1803 = n1627 & n1739 ;
  assign n1804 = n1803 ^ n1629 ;
  assign n1805 = n1804 ^ n786 ;
  assign n1806 = n1805 ^ n927 ;
  assign n1807 = ~n1802 & n1806 ;
  assign n1808 = n1807 ^ n1805 ;
  assign n1809 = n1634 & n1739 ;
  assign n1810 = n1809 ^ n1636 ;
  assign n1811 = n1810 ^ n696 ;
  assign n1812 = n1811 ^ n842 ;
  assign n1813 = ~n1808 & n1812 ;
  assign n1814 = n1813 ^ n1811 ;
  assign n1815 = n1640 & n1739 ;
  assign n1816 = n1815 ^ n1642 ;
  assign n1817 = n1816 ^ n696 ;
  assign n1818 = n1814 & ~n1817 ;
  assign n1819 = n1818 ^ n835 ;
  assign n1820 = n1645 & n1739 ;
  assign n1821 = n1820 ^ n1647 ;
  assign n1822 = n1821 ^ n609 ;
  assign n1823 = ~n1819 & ~n1822 ;
  assign n1824 = n1823 ^ n834 ;
  assign n1825 = n1754 & ~n1824 ;
  assign n1826 = n1825 ^ n750 ;
  assign n1827 = n1751 & n1826 ;
  assign n1828 = n1827 ^ n1750 ;
  assign n1831 = n1830 ^ n1828 ;
  assign n1832 = n1830 ^ n401 ;
  assign n1833 = n1831 & n1832 ;
  assign n1834 = n1833 ^ n462 ;
  assign n1835 = n1748 & n1834 ;
  assign n1836 = n1835 ^ n349 ;
  assign n1860 = n1733 ^ n138 ;
  assign n1861 = n1739 & n1860 ;
  assign n1862 = n1861 ^ n1721 ;
  assign n1854 = n1736 ^ n1718 ;
  assign n1855 = n183 & ~n1854 ;
  assign n1856 = ~n1715 & n1855 ;
  assign n1857 = n1736 & n1856 ;
  assign n1858 = n1857 ^ n1855 ;
  assign n1859 = n1858 ^ n183 ;
  assign n1863 = n1862 ^ n1859 ;
  assign n1864 = n1730 ^ n157 ;
  assign n1865 = n1739 & n1864 ;
  assign n1866 = n1865 ^ n1724 ;
  assign n1867 = ~n138 & n1866 ;
  assign n1868 = n1866 ^ n138 ;
  assign n1869 = n1868 ^ n1867 ;
  assign n1870 = ~n1862 & n1869 ;
  assign n1873 = n138 & n1730 ;
  assign n1874 = n157 & n1873 ;
  assign n1875 = n1874 ^ n1739 ;
  assign n1876 = n1733 ^ n1722 ;
  assign n1877 = n1864 ^ n1724 ;
  assign n1878 = n1877 ^ n1864 ;
  assign n1879 = ~n1721 & ~n1878 ;
  assign n1880 = n1879 ^ n1864 ;
  assign n1882 = n138 & n1880 ;
  assign n1883 = n1882 ^ n1721 ;
  assign n1884 = n1876 & ~n1883 ;
  assign n1885 = n1884 ^ n1721 ;
  assign n1886 = n1885 ^ n1884 ;
  assign n1891 = n138 & ~n1724 ;
  assign n1892 = n1886 & n1891 ;
  assign n1893 = n1892 ^ n1886 ;
  assign n1894 = n1893 ^ n1884 ;
  assign n1895 = ~n1875 & n1894 ;
  assign n1896 = n1895 ^ n1884 ;
  assign n1871 = ~n138 & n1721 ;
  assign n1923 = n1896 ^ n1871 ;
  assign n1921 = n1896 ^ n1715 ;
  assign n1920 = n1718 ^ n1715 ;
  assign n1922 = n1921 ^ n1920 ;
  assign n1924 = n1923 ^ n1922 ;
  assign n1927 = n1924 ^ n1920 ;
  assign n1925 = n1924 ^ n1733 ;
  assign n1926 = n1925 ^ n1922 ;
  assign n1986 = n1927 ^ n1926 ;
  assign n1987 = n1986 ^ n1923 ;
  assign n1988 = n1987 ^ n1896 ;
  assign n1990 = n1988 ^ n1986 ;
  assign n1900 = n1733 ^ n1715 ;
  assign n1897 = n1896 ^ n1718 ;
  assign n1872 = n1871 ^ n1715 ;
  assign n1898 = n1897 ^ n1872 ;
  assign n1973 = n1900 ^ n1898 ;
  assign n1903 = n1897 ^ n1715 ;
  assign n1974 = n1973 ^ n1903 ;
  assign n1975 = n1974 ^ n1896 ;
  assign n1977 = n1975 ^ n1973 ;
  assign n1938 = n1898 ^ n1715 ;
  assign n1939 = n1938 ^ n1733 ;
  assign n1940 = n1939 ^ n1896 ;
  assign n1941 = n1940 ^ n1897 ;
  assign n1959 = n1941 ^ n1871 ;
  assign n1901 = n1900 ^ n1897 ;
  assign n1956 = n1941 ^ n1901 ;
  assign n1957 = n1956 ^ n1941 ;
  assign n1958 = n1957 ^ n1897 ;
  assign n1962 = n1959 ^ n1958 ;
  assign n1963 = n1962 ^ n1940 ;
  assign n1964 = n1963 ^ n1718 ;
  assign n1966 = n1964 ^ n1962 ;
  assign n1947 = ~n1733 & n1871 ;
  assign n1948 = n1718 & ~n1896 ;
  assign n1949 = n1948 ^ n1920 ;
  assign n1950 = n1949 ^ n1715 ;
  assign n1951 = n1949 ^ n1948 ;
  assign n1952 = ~n1950 & n1951 ;
  assign n1953 = n1947 & n1952 ;
  assign n1954 = n1953 ^ n1949 ;
  assign n1967 = n1966 ^ n1954 ;
  assign n1968 = n1967 ^ n1956 ;
  assign n1972 = n1968 ^ n1938 ;
  assign n1978 = n1977 ^ n1972 ;
  assign n1979 = n1978 ^ n1871 ;
  assign n1991 = n1990 ^ n1979 ;
  assign n1997 = n1991 ^ n1718 ;
  assign n1899 = n1898 ^ n1897 ;
  assign n1902 = n1901 ^ n1899 ;
  assign n1904 = n1903 ^ n1902 ;
  assign n1906 = n1904 ^ n1896 ;
  assign n1998 = n1997 ^ n1906 ;
  assign n1999 = ~n183 & n1998 ;
  assign n2000 = n1999 ^ n1859 ;
  assign n2001 = n1870 & n2000 ;
  assign n2002 = n2001 ^ n2000 ;
  assign n1740 = n1674 & n1739 ;
  assign n1741 = n1740 ^ n1727 ;
  assign n1742 = n1741 ^ n157 ;
  assign n1837 = n1664 & n1739 ;
  assign n1838 = n1837 ^ n1578 ;
  assign n1839 = n1838 ^ n291 ;
  assign n1840 = ~n1836 & n1839 ;
  assign n1841 = n1840 ^ n307 ;
  assign n1842 = ~n1666 & n1739 ;
  assign n1843 = n1842 ^ n1668 ;
  assign n1844 = n1843 ^ n245 ;
  assign n1845 = ~n1841 & n1844 ;
  assign n1846 = n1845 ^ n245 ;
  assign n1743 = ~n1671 & n1739 ;
  assign n1744 = n1743 ^ n1574 ;
  assign n1847 = n1846 ^ n1744 ;
  assign n1848 = n1846 ^ n188 ;
  assign n1849 = ~n1847 & n1848 ;
  assign n1850 = n1849 ^ n203 ;
  assign n1851 = ~n1742 & ~n1850 ;
  assign n1852 = n1851 ^ n1741 ;
  assign n2003 = n1852 & n2002 ;
  assign n2004 = n2002 & ~n2003 ;
  assign n2005 = ~n1867 & n2004 ;
  assign n2006 = n1863 & n2005 ;
  assign n2007 = n2006 ^ n2004 ;
  assign n2008 = n2007 ^ n2003 ;
  assign n2045 = ~n1836 & ~n2008 ;
  assign n2046 = n2045 ^ n1838 ;
  assign n2047 = n2046 ^ n245 ;
  assign n2048 = n1828 ^ n401 ;
  assign n2049 = ~n2008 & ~n2048 ;
  assign n2050 = n2049 ^ n1830 ;
  assign n2051 = n2050 ^ n341 ;
  assign n2139 = ~n1826 & ~n2008 ;
  assign n2140 = n2139 ^ n1750 ;
  assign n2052 = ~n1824 & ~n2008 ;
  assign n2053 = n2052 ^ n1753 ;
  assign n2054 = n2053 ^ n457 ;
  assign n2055 = ~n1777 & ~n2008 ;
  assign n2056 = n2055 ^ n1787 ;
  assign n2057 = n2056 ^ n1136 ;
  assign n2094 = ~n1770 & ~n2008 ;
  assign n2095 = n2094 ^ n1774 ;
  assign n2098 = n2095 ^ n1136 ;
  assign n2074 = n1756 ^ n1739 ;
  assign n2075 = n2008 & n2074 ;
  assign n2076 = n2075 ^ n1757 ;
  assign n2079 = n2076 ^ n1427 ;
  assign n2058 = n1739 ^ x87 ;
  assign n2059 = n2058 ^ n2008 ;
  assign n2061 = ~x84 & ~x85 ;
  assign n2060 = n1739 ^ x86 ;
  assign n2062 = n2061 ^ n2060 ;
  assign n2063 = n2059 & n2062 ;
  assign n2072 = n2063 ^ n1763 ;
  assign n2064 = n2008 ^ n1739 ;
  assign n2065 = n2064 ^ n2063 ;
  assign n2066 = n2065 ^ n2063 ;
  assign n2069 = ~n2058 & ~n2066 ;
  assign n2070 = n2069 ^ n2063 ;
  assign n2071 = x86 & n2070 ;
  assign n2073 = n2072 ^ n2071 ;
  assign n2077 = n2076 ^ n1572 ;
  assign n2078 = n2073 & n2077 ;
  assign n2080 = n2079 ^ n2078 ;
  assign n2084 = n1763 ^ x88 ;
  assign n2085 = n2084 ^ n1763 ;
  assign n2086 = n2074 & ~n2085 ;
  assign n2087 = n2086 ^ n1763 ;
  assign n2088 = ~n2008 & ~n2087 ;
  assign n2089 = n2088 ^ x89 ;
  assign n2081 = ~x88 & n1739 ;
  assign n2090 = n2089 ^ n2081 ;
  assign n2091 = n2090 ^ n1427 ;
  assign n2092 = ~n2080 & ~n2091 ;
  assign n2093 = n2092 ^ n1450 ;
  assign n2096 = n2095 ^ n1290 ;
  assign n2097 = n2093 & n2096 ;
  assign n2099 = n2098 ^ n2097 ;
  assign n2100 = n2057 & n2099 ;
  assign n2101 = n2100 ^ n1143 ;
  assign n2102 = n1790 & ~n2008 ;
  assign n2103 = n2102 ^ n1792 ;
  assign n2106 = n2103 ^ n1034 ;
  assign n2107 = ~n2101 & n2106 ;
  assign n2104 = n2103 ^ n892 ;
  assign n2108 = n2107 ^ n2104 ;
  assign n2109 = n1795 & ~n2008 ;
  assign n2110 = n2109 ^ n1797 ;
  assign n2111 = n2110 ^ n786 ;
  assign n2112 = n2111 ^ n927 ;
  assign n2113 = ~n2108 & n2112 ;
  assign n2114 = n2113 ^ n2111 ;
  assign n2115 = n1802 & ~n2008 ;
  assign n2116 = n2115 ^ n1804 ;
  assign n2117 = n2116 ^ n696 ;
  assign n2118 = n2117 ^ n842 ;
  assign n2119 = ~n2114 & n2118 ;
  assign n2120 = n2119 ^ n2117 ;
  assign n2121 = n1808 & ~n2008 ;
  assign n2122 = n2121 ^ n1810 ;
  assign n2123 = n2122 ^ n609 ;
  assign n2124 = n2123 ^ n835 ;
  assign n2125 = ~n2120 & n2124 ;
  assign n2126 = n2125 ^ n2123 ;
  assign n2127 = n1814 & ~n2008 ;
  assign n2128 = n2127 ^ n1816 ;
  assign n2129 = n2128 ^ n609 ;
  assign n2130 = ~n2126 & n2129 ;
  assign n2131 = n2130 ^ n834 ;
  assign n2132 = ~n1819 & ~n2008 ;
  assign n2133 = n2132 ^ n1821 ;
  assign n2134 = n2133 ^ n534 ;
  assign n2135 = ~n2131 & n2134 ;
  assign n2136 = n2135 ^ n750 ;
  assign n2137 = ~n2054 & n2136 ;
  assign n2138 = n2137 ^ n2053 ;
  assign n2141 = n2140 ^ n2138 ;
  assign n2142 = n2140 ^ n401 ;
  assign n2143 = n2141 & ~n2142 ;
  assign n2144 = n2143 ^ n462 ;
  assign n2145 = n2051 & n2144 ;
  assign n2146 = n2145 ^ n349 ;
  assign n2147 = n1834 & ~n2008 ;
  assign n2148 = n2147 ^ n1747 ;
  assign n2149 = n2148 ^ n291 ;
  assign n2150 = ~n2146 & ~n2149 ;
  assign n2151 = n2150 ^ n307 ;
  assign n2152 = ~n2047 & n2151 ;
  assign n2153 = n2152 ^ n2046 ;
  assign n2154 = n2153 ^ n188 ;
  assign n2155 = ~n1841 & ~n2008 ;
  assign n2156 = n2155 ^ n1843 ;
  assign n2157 = n2156 ^ n2153 ;
  assign n2158 = ~n2154 & n2157 ;
  assign n2159 = n2158 ^ n188 ;
  assign n2163 = n2159 ^ n157 ;
  assign n2012 = ~n183 & ~n1866 ;
  assign n1853 = n1852 ^ n138 ;
  assign n2038 = n2003 ^ n1852 ;
  assign n2039 = n2038 ^ n2008 ;
  assign n2040 = n1853 & ~n2039 ;
  assign n2043 = n2012 & n2040 ;
  assign n2021 = n1866 ^ n1853 ;
  assign n2030 = n183 & n1862 ;
  assign n2018 = n1862 ^ n183 ;
  assign n2019 = n2018 ^ n2008 ;
  assign n2020 = n2019 ^ n1853 ;
  assign n2031 = n2030 ^ n2020 ;
  assign n2032 = n2021 & n2031 ;
  assign n2022 = n2021 ^ n2020 ;
  assign n2035 = n2032 ^ n2022 ;
  assign n2013 = n1853 ^ n183 ;
  assign n2014 = n2008 ^ n1866 ;
  assign n2015 = ~n2013 & ~n2014 ;
  assign n2033 = n2032 ^ n1866 ;
  assign n2034 = n2015 & n2033 ;
  assign n2036 = n2035 ^ n2034 ;
  assign n2037 = n2036 ^ n2021 ;
  assign n2041 = n2040 ^ n2037 ;
  assign n2044 = n2043 ^ n2041 ;
  assign n2160 = n1848 & ~n2008 ;
  assign n2161 = n2160 ^ n1744 ;
  assign n2162 = n2161 ^ n2159 ;
  assign n2164 = n2162 & ~n2163 ;
  assign n2165 = n2164 ^ n2161 ;
  assign n2166 = n2165 ^ n138 ;
  assign n2167 = n1850 & ~n2008 ;
  assign n2168 = n2167 ^ n1741 ;
  assign n2169 = n2168 ^ n138 ;
  assign n2170 = n2166 & ~n2169 ;
  assign n2171 = n2170 ^ n138 ;
  assign n2172 = n2044 & n2171 ;
  assign n2174 = n2172 ^ n2044 ;
  assign n2009 = ~n1853 & ~n2008 ;
  assign n2010 = n2009 ^ n1866 ;
  assign n2011 = n183 & n2010 ;
  assign n2173 = n2011 & n2172 ;
  assign n2175 = n2174 ^ n2173 ;
  assign n2176 = n2163 & ~n2175 ;
  assign n2177 = n2176 ^ n2161 ;
  assign n2178 = n138 & n2165 ;
  assign n2179 = n2178 ^ n2166 ;
  assign n2180 = ~n2175 & ~n2178 ;
  assign n2181 = n2179 & n2180 ;
  assign n2182 = n2181 ^ n2168 ;
  assign n2183 = ~n2177 & n2182 ;
  assign n2295 = ~n2151 & ~n2175 ;
  assign n2296 = n2295 ^ n2046 ;
  assign n2184 = n2138 ^ n401 ;
  assign n2185 = ~n2175 & n2184 ;
  assign n2186 = n2185 ^ n2140 ;
  assign n2187 = n2186 ^ n341 ;
  assign n2277 = ~n2136 & ~n2175 ;
  assign n2278 = n2277 ^ n2053 ;
  assign n2188 = ~n2131 & ~n2175 ;
  assign n2189 = n2188 ^ n2133 ;
  assign n2190 = n2189 ^ n457 ;
  assign n2191 = n2120 & ~n2175 ;
  assign n2192 = n2191 ^ n2122 ;
  assign n2193 = n2192 ^ n609 ;
  assign n2237 = ~n2093 & ~n2175 ;
  assign n2238 = n2237 ^ n2095 ;
  assign n2226 = ~n2073 & ~n2175 ;
  assign n2227 = n2226 ^ n2076 ;
  assign n2198 = n2061 ^ n2008 ;
  assign n2199 = ~n2175 & ~n2198 ;
  assign n2200 = n2199 ^ n2008 ;
  assign n2201 = x86 & ~n2200 ;
  assign n2196 = n2008 ^ x87 ;
  assign n2194 = n2061 ^ n1739 ;
  assign n2195 = ~n2175 & n2194 ;
  assign n2197 = n2196 ^ n2195 ;
  assign n2202 = n2201 ^ n2197 ;
  assign n2203 = n2202 ^ n1572 ;
  assign n2205 = n2008 ^ x85 ;
  assign n2206 = n2205 ^ n2175 ;
  assign n2207 = ~x82 & ~x83 ;
  assign n2208 = n2207 ^ n2008 ;
  assign n2209 = n2208 ^ x84 ;
  assign n2210 = ~n2206 & ~n2209 ;
  assign n2218 = n2210 ^ n2064 ;
  assign n2204 = n2175 ^ n2008 ;
  assign n2211 = n2210 ^ n2204 ;
  assign n2212 = n2211 ^ n2210 ;
  assign n2215 = n2205 & n2212 ;
  assign n2216 = n2215 ^ n2210 ;
  assign n2217 = x84 & n2216 ;
  assign n2219 = n2218 ^ n2217 ;
  assign n2220 = n2200 ^ x86 ;
  assign n2221 = n2220 ^ n1739 ;
  assign n2222 = ~n2219 & n2221 ;
  assign n2223 = n2222 ^ n1763 ;
  assign n2224 = ~n2203 & n2223 ;
  assign n2225 = n2224 ^ n2202 ;
  assign n2228 = n2227 ^ n2225 ;
  assign n2229 = n2227 ^ n1427 ;
  assign n2230 = n2228 & ~n2229 ;
  assign n2231 = n2230 ^ n1450 ;
  assign n2232 = ~n2080 & ~n2175 ;
  assign n2233 = n2232 ^ n2090 ;
  assign n2234 = n2233 ^ n1290 ;
  assign n2235 = n2231 & n2234 ;
  assign n2236 = n2235 ^ n2233 ;
  assign n2239 = n2238 ^ n2236 ;
  assign n2240 = n2238 ^ n1136 ;
  assign n2241 = ~n2239 & n2240 ;
  assign n2242 = n2241 ^ n1143 ;
  assign n2243 = n2099 & ~n2175 ;
  assign n2244 = n2243 ^ n2056 ;
  assign n2247 = n2244 ^ n1034 ;
  assign n2248 = ~n2242 & n2247 ;
  assign n2245 = n2244 ^ n892 ;
  assign n2249 = n2248 ^ n2245 ;
  assign n2250 = n2101 & ~n2175 ;
  assign n2251 = n2250 ^ n2103 ;
  assign n2252 = n2251 ^ n786 ;
  assign n2253 = n2252 ^ n927 ;
  assign n2254 = ~n2249 & n2253 ;
  assign n2255 = n2254 ^ n2252 ;
  assign n2256 = n2108 & ~n2175 ;
  assign n2257 = n2256 ^ n2110 ;
  assign n2258 = n2257 ^ n696 ;
  assign n2259 = n2258 ^ n842 ;
  assign n2260 = ~n2255 & n2259 ;
  assign n2261 = n2260 ^ n2258 ;
  assign n2262 = n2114 & ~n2175 ;
  assign n2263 = n2262 ^ n2116 ;
  assign n2264 = n2263 ^ n609 ;
  assign n2265 = n2264 ^ n835 ;
  assign n2266 = ~n2261 & n2265 ;
  assign n2267 = n2266 ^ n2264 ;
  assign n2268 = ~n2193 & ~n2267 ;
  assign n2269 = n2268 ^ n834 ;
  assign n2270 = ~n2126 & ~n2175 ;
  assign n2271 = n2270 ^ n2128 ;
  assign n2272 = n2271 ^ n534 ;
  assign n2273 = ~n2269 & ~n2272 ;
  assign n2274 = n2273 ^ n750 ;
  assign n2275 = ~n2190 & n2274 ;
  assign n2276 = n2275 ^ n2189 ;
  assign n2279 = n2278 ^ n2276 ;
  assign n2280 = n2278 ^ n401 ;
  assign n2281 = ~n2279 & n2280 ;
  assign n2282 = n2281 ^ n462 ;
  assign n2283 = ~n2187 & n2282 ;
  assign n2284 = n2283 ^ n349 ;
  assign n2285 = n2144 & ~n2175 ;
  assign n2286 = n2285 ^ n2050 ;
  assign n2287 = n2286 ^ n291 ;
  assign n2288 = ~n2284 & ~n2287 ;
  assign n2289 = n2288 ^ n307 ;
  assign n2290 = ~n2146 & ~n2175 ;
  assign n2291 = n2290 ^ n2148 ;
  assign n2292 = n2291 ^ n245 ;
  assign n2293 = n2289 & n2292 ;
  assign n2294 = n2293 ^ n2291 ;
  assign n2297 = n2296 ^ n2294 ;
  assign n2298 = n2296 ^ n188 ;
  assign n2299 = n2297 & ~n2298 ;
  assign n2300 = n2299 ^ n203 ;
  assign n2301 = ~n2154 & ~n2175 ;
  assign n2302 = n2301 ^ n2156 ;
  assign n2303 = n2302 ^ n157 ;
  assign n2304 = n2300 & n2303 ;
  assign n2305 = n2304 ^ n157 ;
  assign n2340 = n2305 ^ n138 ;
  assign n2341 = n2182 & n2340 ;
  assign n2307 = n138 & n2177 ;
  assign n2306 = n2177 ^ n138 ;
  assign n2308 = n2307 ^ n2306 ;
  assign n2338 = n2308 ^ n2305 ;
  assign n2309 = n2305 & n2308 ;
  assign n2339 = n2338 ^ n2309 ;
  assign n2342 = n2341 ^ n2339 ;
  assign n2310 = n2180 ^ n2010 ;
  assign n2311 = n2310 ^ n2168 ;
  assign n2318 = n2168 & ~n2178 ;
  assign n2319 = n2044 & n2318 ;
  assign n2320 = n2319 ^ n2318 ;
  assign n2321 = n2320 ^ n2168 ;
  assign n2322 = ~n2311 & ~n2321 ;
  assign n2323 = ~n2179 & n2322 ;
  assign n2312 = n2311 ^ n2175 ;
  assign n2313 = n2175 ^ n2010 ;
  assign n2314 = n2313 ^ n2175 ;
  assign n2315 = ~n2312 & n2314 ;
  assign n2316 = n2315 ^ n2175 ;
  assign n2317 = ~n2307 & n2316 ;
  assign n2324 = n2323 ^ n2317 ;
  assign n2325 = ~n2309 & n2324 ;
  assign n2343 = ~n183 & ~n2325 ;
  assign n2344 = ~n2342 & n2343 ;
  assign n2326 = n2319 ^ n2010 ;
  assign n2327 = n2044 ^ n2010 ;
  assign n2328 = n2326 & ~n2327 ;
  assign n2329 = n2328 ^ n2318 ;
  assign n2330 = n2179 & ~n2329 ;
  assign n2331 = n2330 ^ n2010 ;
  assign n2332 = n2331 ^ n2325 ;
  assign n2333 = ~n183 & n2332 ;
  assign n2334 = n2333 ^ n2331 ;
  assign n2345 = n2344 ^ n2334 ;
  assign n2346 = n2345 ^ n2305 ;
  assign n2347 = n2346 ^ n2345 ;
  assign n2350 = n1003 & n2347 ;
  assign n2351 = n2350 ^ n2345 ;
  assign n2352 = n2183 & n2351 ;
  assign n2353 = n2352 ^ n2344 ;
  assign n2354 = ~n183 & ~n2353 ;
  assign n2355 = ~n2307 & ~n2309 ;
  assign n2356 = n2355 ^ n2182 ;
  assign n2357 = n2356 ^ n2183 ;
  assign n2358 = n2334 & ~n2355 ;
  assign n2361 = n2357 & ~n2358 ;
  assign n2362 = n2361 ^ n2183 ;
  assign n2363 = ~n2353 & n2362 ;
  assign n2364 = ~n2354 & ~n2363 ;
  assign n2365 = ~n2182 & n2358 ;
  assign n2366 = n2365 ^ n2334 ;
  assign n2367 = n2340 & ~n2366 ;
  assign n2368 = n2367 ^ n2177 ;
  assign n2369 = n183 & ~n2368 ;
  assign n2373 = ~n2289 & ~n2366 ;
  assign n2374 = n2373 ^ n2291 ;
  assign n2375 = n2374 ^ n188 ;
  assign n2376 = n2276 ^ n401 ;
  assign n2377 = ~n2366 & n2376 ;
  assign n2378 = n2377 ^ n2278 ;
  assign n2379 = n2378 ^ n341 ;
  assign n2479 = ~n2274 & ~n2366 ;
  assign n2480 = n2479 ^ n2189 ;
  assign n2380 = ~n2267 & ~n2366 ;
  assign n2381 = n2380 ^ n2192 ;
  assign n2382 = n2381 ^ n534 ;
  assign n2383 = n2261 & ~n2366 ;
  assign n2384 = n2383 ^ n2263 ;
  assign n2385 = n2384 ^ n609 ;
  assign n2386 = ~n2231 & ~n2366 ;
  assign n2387 = n2386 ^ n2233 ;
  assign n2388 = n2387 ^ n1136 ;
  assign n2435 = n2225 ^ n1427 ;
  assign n2436 = ~n2366 & n2435 ;
  assign n2437 = n2436 ^ n2227 ;
  assign n2440 = n2437 ^ n1136 ;
  assign n2429 = ~n2223 & ~n2366 ;
  assign n2430 = n2429 ^ n2202 ;
  assign n2389 = ~n2219 & ~n2366 ;
  assign n2390 = n2389 ^ n2220 ;
  assign n2391 = n2390 ^ n1572 ;
  assign n2393 = n2207 ^ n2175 ;
  assign n2394 = ~n2366 & ~n2393 ;
  assign n2392 = n2175 ^ x84 ;
  assign n2395 = n2394 ^ n2392 ;
  assign n2396 = n2395 ^ n2008 ;
  assign n2399 = n2366 ^ n2175 ;
  assign n2397 = n2175 ^ x83 ;
  assign n2398 = n2397 ^ x82 ;
  assign n2400 = n2399 ^ n2398 ;
  assign n2401 = n2400 ^ n2399 ;
  assign n2402 = n2401 ^ n2397 ;
  assign n2404 = n2397 ^ n2366 ;
  assign n2405 = ~x80 & ~x81 ;
  assign n2406 = n2405 ^ n2400 ;
  assign n2407 = ~n2404 & ~n2406 ;
  assign n2403 = n2397 & n2399 ;
  assign n2408 = n2407 ^ n2403 ;
  assign n2409 = ~n2402 & n2408 ;
  assign n2410 = n2409 ^ n2403 ;
  assign n2411 = n2410 ^ n2175 ;
  assign n2412 = n2411 ^ n2395 ;
  assign n2413 = ~n2396 & n2412 ;
  assign n2414 = n2413 ^ n2064 ;
  assign n2422 = ~x84 & ~n2175 ;
  assign n2415 = n2393 ^ n2208 ;
  assign n2416 = n2415 ^ n2208 ;
  assign n2417 = n2209 ^ n2208 ;
  assign n2418 = ~n2416 & n2417 ;
  assign n2419 = n2418 ^ n2208 ;
  assign n2420 = ~n2366 & ~n2419 ;
  assign n2421 = n2420 ^ x85 ;
  assign n2423 = n2422 ^ n2421 ;
  assign n2424 = n2423 ^ n1739 ;
  assign n2425 = ~n2414 & ~n2424 ;
  assign n2426 = n2425 ^ n1763 ;
  assign n2427 = ~n2391 & n2426 ;
  assign n2428 = n2427 ^ n2390 ;
  assign n2431 = n2430 ^ n2428 ;
  assign n2432 = n2430 ^ n1427 ;
  assign n2433 = ~n2431 & n2432 ;
  assign n2434 = n2433 ^ n1450 ;
  assign n2438 = n2437 ^ n1290 ;
  assign n2439 = n2434 & n2438 ;
  assign n2441 = n2440 ^ n2439 ;
  assign n2442 = n2388 & n2441 ;
  assign n2443 = n2442 ^ n1143 ;
  assign n2444 = n2236 ^ n1136 ;
  assign n2445 = ~n2366 & n2444 ;
  assign n2446 = n2445 ^ n2238 ;
  assign n2449 = n2446 ^ n1034 ;
  assign n2450 = ~n2443 & n2449 ;
  assign n2447 = n2446 ^ n892 ;
  assign n2451 = n2450 ^ n2447 ;
  assign n2452 = n2242 & ~n2366 ;
  assign n2453 = n2452 ^ n2244 ;
  assign n2454 = n2453 ^ n786 ;
  assign n2455 = n2454 ^ n927 ;
  assign n2456 = ~n2451 & n2455 ;
  assign n2457 = n2456 ^ n2454 ;
  assign n2458 = n2249 & ~n2366 ;
  assign n2459 = n2458 ^ n2251 ;
  assign n2460 = n2459 ^ n696 ;
  assign n2461 = n2460 ^ n842 ;
  assign n2462 = ~n2457 & n2461 ;
  assign n2463 = n2462 ^ n2460 ;
  assign n2464 = n2255 & ~n2366 ;
  assign n2465 = n2464 ^ n2257 ;
  assign n2466 = n2465 ^ n609 ;
  assign n2467 = n2466 ^ n835 ;
  assign n2468 = ~n2463 & n2467 ;
  assign n2469 = n2468 ^ n2466 ;
  assign n2470 = ~n2385 & ~n2469 ;
  assign n2471 = n2470 ^ n834 ;
  assign n2472 = n2382 & ~n2471 ;
  assign n2473 = n2472 ^ n750 ;
  assign n2474 = ~n2269 & ~n2366 ;
  assign n2475 = n2474 ^ n2271 ;
  assign n2476 = n2475 ^ n457 ;
  assign n2477 = ~n2473 & n2476 ;
  assign n2478 = n2477 ^ n457 ;
  assign n2481 = n2480 ^ n2478 ;
  assign n2482 = n2480 ^ n401 ;
  assign n2483 = n2481 & n2482 ;
  assign n2484 = n2483 ^ n462 ;
  assign n2485 = n2379 & n2484 ;
  assign n2486 = n2485 ^ n349 ;
  assign n2487 = n2282 & ~n2366 ;
  assign n2488 = n2487 ^ n2186 ;
  assign n2489 = n2488 ^ n291 ;
  assign n2490 = ~n2486 & n2489 ;
  assign n2491 = n2490 ^ n307 ;
  assign n2492 = ~n2284 & ~n2366 ;
  assign n2493 = n2492 ^ n2286 ;
  assign n2494 = n2493 ^ n245 ;
  assign n2495 = n2491 & n2494 ;
  assign n2496 = n2495 ^ n2493 ;
  assign n2497 = n2496 ^ n2374 ;
  assign n2498 = n2375 & ~n2497 ;
  assign n2499 = n2498 ^ n188 ;
  assign n2370 = n2294 ^ n188 ;
  assign n2371 = ~n2366 & n2370 ;
  assign n2372 = n2371 ^ n2296 ;
  assign n2500 = n2499 ^ n2372 ;
  assign n2501 = n2372 ^ n157 ;
  assign n2502 = ~n2500 & n2501 ;
  assign n2503 = n2502 ^ n2499 ;
  assign n2504 = n2503 ^ n138 ;
  assign n2505 = n2300 & ~n2366 ;
  assign n2506 = n2505 ^ n2302 ;
  assign n2507 = n2506 ^ n2503 ;
  assign n2508 = n2504 & ~n2507 ;
  assign n2509 = n2508 ^ n138 ;
  assign n2510 = ~n2369 & n2509 ;
  assign n2511 = n2364 & ~n2510 ;
  assign n2610 = n2499 ^ n157 ;
  assign n2611 = ~n2511 & n2610 ;
  assign n2612 = n2611 ^ n2372 ;
  assign n2613 = n2612 ^ n138 ;
  assign n2647 = n2496 ^ n188 ;
  assign n2648 = ~n2511 & n2647 ;
  assign n2649 = n2648 ^ n2374 ;
  assign n2614 = n2478 ^ n401 ;
  assign n2615 = ~n2511 & ~n2614 ;
  assign n2616 = n2615 ^ n2480 ;
  assign n2617 = n2616 ^ n341 ;
  assign n2512 = ~n2469 & ~n2511 ;
  assign n2513 = n2512 ^ n2384 ;
  assign n2514 = n2513 ^ n534 ;
  assign n2515 = n2463 & ~n2511 ;
  assign n2516 = n2515 ^ n2465 ;
  assign n2606 = n2516 ^ n534 ;
  assign n2517 = n2516 ^ n609 ;
  assign n2574 = ~n2434 & ~n2511 ;
  assign n2575 = n2574 ^ n2437 ;
  assign n2557 = ~n2414 & ~n2511 ;
  assign n2558 = n2557 ^ n2423 ;
  assign n2561 = n2558 ^ n1427 ;
  assign n2522 = n2405 ^ n2366 ;
  assign n2523 = ~n2511 & ~n2522 ;
  assign n2524 = n2523 ^ n2366 ;
  assign n2525 = x82 & ~n2524 ;
  assign n2519 = n2405 ^ n2175 ;
  assign n2520 = ~n2511 & ~n2519 ;
  assign n2518 = n2366 ^ x83 ;
  assign n2521 = n2520 ^ n2518 ;
  assign n2526 = n2525 ^ n2521 ;
  assign n2527 = n2526 ^ n2008 ;
  assign n2528 = n2524 ^ x82 ;
  assign n2529 = n2528 ^ n2175 ;
  assign n2530 = n2511 ^ n2366 ;
  assign n2531 = n2175 ^ x81 ;
  assign n2532 = n2531 ^ n2175 ;
  assign n2533 = n2532 ^ n2511 ;
  assign n2534 = ~n2530 & n2533 ;
  assign n2535 = n2534 ^ n2531 ;
  assign n2541 = n2535 ^ n2399 ;
  assign n2537 = ~x78 & ~x79 ;
  assign n2536 = n2511 ^ x81 ;
  assign n2538 = n2537 ^ n2536 ;
  assign n2539 = n2537 ^ n2366 ;
  assign n2540 = ~n2538 & ~n2539 ;
  assign n2542 = n2541 ^ n2540 ;
  assign n2543 = ~x80 & n2542 ;
  assign n2544 = n2543 ^ n2535 ;
  assign n2545 = ~n2529 & n2544 ;
  assign n2546 = n2545 ^ n2175 ;
  assign n2547 = n2546 ^ n2526 ;
  assign n2548 = ~n2527 & n2547 ;
  assign n2549 = n2548 ^ n2008 ;
  assign n2550 = n2549 ^ n1739 ;
  assign n2551 = n2411 ^ n2008 ;
  assign n2552 = ~n2511 & n2551 ;
  assign n2553 = n2552 ^ n2395 ;
  assign n2554 = n2553 ^ n2549 ;
  assign n2555 = ~n2550 & n2554 ;
  assign n2556 = n2555 ^ n1763 ;
  assign n2559 = n2558 ^ n1572 ;
  assign n2560 = n2556 & n2559 ;
  assign n2562 = n2561 ^ n2560 ;
  assign n2563 = ~n2426 & ~n2511 ;
  assign n2564 = n2563 ^ n2390 ;
  assign n2565 = n2564 ^ n1427 ;
  assign n2566 = ~n2562 & n2565 ;
  assign n2567 = n2566 ^ n1450 ;
  assign n2568 = n2428 ^ n1427 ;
  assign n2569 = ~n2511 & n2568 ;
  assign n2570 = n2569 ^ n2430 ;
  assign n2571 = n2570 ^ n1290 ;
  assign n2572 = n2567 & ~n2571 ;
  assign n2573 = n2572 ^ n2570 ;
  assign n2576 = n2575 ^ n2573 ;
  assign n2577 = n2575 ^ n1136 ;
  assign n2578 = n2576 & n2577 ;
  assign n2579 = n2578 ^ n1143 ;
  assign n2580 = n2441 & ~n2511 ;
  assign n2581 = n2580 ^ n2387 ;
  assign n2584 = n2581 ^ n1034 ;
  assign n2585 = ~n2579 & n2584 ;
  assign n2582 = n2581 ^ n892 ;
  assign n2586 = n2585 ^ n2582 ;
  assign n2587 = n2443 & ~n2511 ;
  assign n2588 = n2587 ^ n2446 ;
  assign n2589 = n2588 ^ n786 ;
  assign n2590 = n2589 ^ n927 ;
  assign n2591 = ~n2586 & n2590 ;
  assign n2592 = n2591 ^ n2589 ;
  assign n2593 = n2451 & ~n2511 ;
  assign n2594 = n2593 ^ n2453 ;
  assign n2595 = n2594 ^ n696 ;
  assign n2596 = n2595 ^ n842 ;
  assign n2597 = ~n2592 & n2596 ;
  assign n2598 = n2597 ^ n2595 ;
  assign n2599 = n2457 & ~n2511 ;
  assign n2600 = n2599 ^ n2459 ;
  assign n2601 = n2600 ^ n609 ;
  assign n2602 = n2601 ^ n835 ;
  assign n2603 = ~n2598 & n2602 ;
  assign n2604 = n2603 ^ n2601 ;
  assign n2605 = ~n2517 & n2604 ;
  assign n2607 = n2606 ^ n2605 ;
  assign n2608 = n2514 & n2607 ;
  assign n2609 = n2608 ^ n750 ;
  assign n2618 = ~n2471 & ~n2511 ;
  assign n2619 = n2618 ^ n2381 ;
  assign n2620 = n2619 ^ n457 ;
  assign n2621 = n2609 & ~n2620 ;
  assign n2622 = n2621 ^ n2619 ;
  assign n2623 = n2622 ^ n401 ;
  assign n2624 = ~n2473 & ~n2511 ;
  assign n2625 = n2624 ^ n2475 ;
  assign n2626 = n2625 ^ n2622 ;
  assign n2627 = n2623 & n2626 ;
  assign n2628 = n2627 ^ n462 ;
  assign n2629 = n2617 & n2628 ;
  assign n2630 = n2629 ^ n349 ;
  assign n2631 = n2484 & ~n2511 ;
  assign n2632 = n2631 ^ n2378 ;
  assign n2633 = n2632 ^ n291 ;
  assign n2634 = ~n2630 & ~n2633 ;
  assign n2635 = n2634 ^ n307 ;
  assign n2636 = ~n2486 & ~n2511 ;
  assign n2637 = n2636 ^ n2488 ;
  assign n2638 = n2637 ^ n245 ;
  assign n2639 = n2635 & ~n2638 ;
  assign n2640 = n2639 ^ n2637 ;
  assign n2641 = n2640 ^ n188 ;
  assign n2642 = ~n2491 & ~n2511 ;
  assign n2643 = n2642 ^ n2493 ;
  assign n2644 = n2643 ^ n2640 ;
  assign n2645 = ~n2641 & n2644 ;
  assign n2646 = n2645 ^ n188 ;
  assign n2650 = n2649 ^ n2646 ;
  assign n2651 = n2646 ^ n157 ;
  assign n2652 = n2650 & ~n2651 ;
  assign n2653 = n2652 ^ n2649 ;
  assign n2654 = n2653 ^ n2612 ;
  assign n2655 = ~n2613 & n2654 ;
  assign n2656 = n2655 ^ n138 ;
  assign n2667 = n138 & ~n2612 ;
  assign n2668 = n2612 & ~n2653 ;
  assign n2669 = n2668 ^ n2654 ;
  assign n2670 = ~n2667 & ~n2669 ;
  assign n2671 = ~n2653 & n2670 ;
  assign n2672 = n2511 ^ n2503 ;
  assign n2676 = n2511 ^ n138 ;
  assign n2677 = n2676 ^ n2368 ;
  assign n2678 = n2677 ^ n2676 ;
  assign n2673 = n2672 ^ n2506 ;
  assign n2679 = n2673 ^ n2511 ;
  assign n2680 = n2679 ^ n2676 ;
  assign n2681 = n2680 ^ n2511 ;
  assign n2682 = n2678 & ~n2681 ;
  assign n2683 = n2682 ^ n2681 ;
  assign n2684 = ~n2672 & ~n2683 ;
  assign n2685 = n2684 ^ n2511 ;
  assign n2686 = n2682 ^ n138 ;
  assign n2687 = n2686 ^ n2684 ;
  assign n2688 = ~n2685 & ~n2687 ;
  assign n2689 = n2688 ^ n2673 ;
  assign n2690 = n2671 & n2689 ;
  assign n2691 = n2690 ^ n2670 ;
  assign n2692 = ~n138 & n2691 ;
  assign n2693 = n2503 ^ n2368 ;
  assign n2694 = ~n2507 & ~n2693 ;
  assign n2695 = n2694 ^ n2503 ;
  assign n2696 = ~n2511 & n2695 ;
  assign n2697 = n2696 ^ n2506 ;
  assign n2698 = n2692 & ~n2697 ;
  assign n2700 = n2698 ^ n2690 ;
  assign n2701 = ~n183 & ~n2700 ;
  assign n2657 = ~n2354 & n2368 ;
  assign n2659 = n2657 ^ n183 ;
  assign n2660 = n2657 ^ n2363 ;
  assign n2661 = n2660 ^ n2657 ;
  assign n2662 = n2659 & n2661 ;
  assign n2663 = n2662 ^ n2657 ;
  assign n2664 = n2509 & n2663 ;
  assign n2665 = n2664 ^ n2657 ;
  assign n2702 = n2701 ^ n2665 ;
  assign n2703 = n2656 & ~n2702 ;
  assign n2704 = n2504 & ~n2511 ;
  assign n2705 = n2704 ^ n2506 ;
  assign n2706 = n2703 & n2705 ;
  assign n2707 = n2706 ^ n2702 ;
  assign n2830 = n2653 ^ n138 ;
  assign n2831 = n2707 & n2830 ;
  assign n2832 = n2831 ^ n2612 ;
  assign n2833 = n2832 ^ n183 ;
  assign n2856 = n2651 & n2707 ;
  assign n2857 = n2856 ^ n2649 ;
  assign n2860 = n2857 ^ n138 ;
  assign n2834 = ~n2641 & n2707 ;
  assign n2835 = n2834 ^ n2643 ;
  assign n2836 = n2835 ^ n157 ;
  assign n2847 = ~n2635 & n2707 ;
  assign n2848 = n2847 ^ n2637 ;
  assign n2708 = ~n2609 & n2707 ;
  assign n2709 = n2708 ^ n2619 ;
  assign n2710 = n2709 ^ n401 ;
  assign n2711 = n2607 & n2707 ;
  assign n2712 = n2711 ^ n2513 ;
  assign n2713 = n2712 ^ n457 ;
  assign n2714 = ~n2604 & n2707 ;
  assign n2715 = n2714 ^ n2516 ;
  assign n2716 = n2715 ^ n534 ;
  assign n2719 = n2592 & n2707 ;
  assign n2720 = n2719 ^ n2594 ;
  assign n2721 = n2720 ^ n696 ;
  assign n2784 = ~n2567 & n2707 ;
  assign n2785 = n2784 ^ n2570 ;
  assign n2722 = n2544 & n2707 ;
  assign n2723 = n2722 ^ n2528 ;
  assign n2724 = n2723 ^ n2008 ;
  assign n2734 = ~x80 & ~n2511 ;
  assign n2725 = n2537 ^ n2511 ;
  assign n2726 = n2725 ^ n2530 ;
  assign n2727 = n2726 ^ n2530 ;
  assign n2728 = n2530 ^ x80 ;
  assign n2729 = n2728 ^ n2530 ;
  assign n2730 = ~n2727 & ~n2729 ;
  assign n2731 = n2730 ^ n2530 ;
  assign n2732 = n2707 & n2731 ;
  assign n2733 = n2732 ^ x81 ;
  assign n2735 = n2734 ^ n2733 ;
  assign n2736 = n2735 ^ n2175 ;
  assign n2738 = n2511 ^ x79 ;
  assign n2739 = n2738 ^ n2707 ;
  assign n2741 = n2511 ^ x78 ;
  assign n2740 = ~x76 & ~x77 ;
  assign n2742 = n2741 ^ n2740 ;
  assign n2743 = n2739 & ~n2742 ;
  assign n2751 = n2743 ^ n2530 ;
  assign n2737 = n2707 ^ n2511 ;
  assign n2744 = n2743 ^ n2737 ;
  assign n2745 = n2744 ^ n2743 ;
  assign n2748 = n2738 & ~n2745 ;
  assign n2749 = n2748 ^ n2743 ;
  assign n2750 = x78 & n2749 ;
  assign n2752 = n2751 ^ n2750 ;
  assign n2754 = n2707 & ~n2725 ;
  assign n2753 = n2511 ^ x80 ;
  assign n2755 = n2754 ^ n2753 ;
  assign n2756 = n2755 ^ n2366 ;
  assign n2757 = n2752 & ~n2756 ;
  assign n2758 = n2757 ^ n2399 ;
  assign n2759 = n2736 & n2758 ;
  assign n2760 = n2759 ^ n2204 ;
  assign n2761 = ~n2724 & n2760 ;
  assign n2762 = n2761 ^ n2064 ;
  assign n2763 = n2546 ^ n2008 ;
  assign n2764 = n2707 & n2763 ;
  assign n2765 = n2764 ^ n2526 ;
  assign n2766 = n2765 ^ n1739 ;
  assign n2767 = ~n2762 & n2766 ;
  assign n2768 = n2767 ^ n1763 ;
  assign n2769 = ~n2550 & n2707 ;
  assign n2770 = n2769 ^ n2553 ;
  assign n2771 = n2770 ^ n1572 ;
  assign n2772 = ~n2768 & ~n2771 ;
  assign n2773 = n2772 ^ n1605 ;
  assign n2774 = ~n2556 & n2707 ;
  assign n2775 = n2774 ^ n2558 ;
  assign n2776 = n2775 ^ n1427 ;
  assign n2777 = ~n2773 & ~n2776 ;
  assign n2778 = n2777 ^ n1450 ;
  assign n2779 = ~n2562 & n2707 ;
  assign n2780 = n2779 ^ n2564 ;
  assign n2781 = n2780 ^ n1290 ;
  assign n2782 = n2778 & ~n2781 ;
  assign n2783 = n2782 ^ n2780 ;
  assign n2786 = n2785 ^ n2783 ;
  assign n2787 = n2785 ^ n1136 ;
  assign n2788 = ~n2786 & ~n2787 ;
  assign n2789 = n2788 ^ n1136 ;
  assign n2790 = n2789 ^ n1034 ;
  assign n2791 = n2573 ^ n1136 ;
  assign n2792 = n2707 & ~n2791 ;
  assign n2793 = n2792 ^ n2575 ;
  assign n2796 = n2793 ^ n2789 ;
  assign n2797 = ~n2790 & n2796 ;
  assign n2794 = n2793 ^ n892 ;
  assign n2798 = n2797 ^ n2794 ;
  assign n2799 = n2579 & n2707 ;
  assign n2800 = n2799 ^ n2581 ;
  assign n2801 = n2800 ^ n786 ;
  assign n2802 = n2801 ^ n927 ;
  assign n2803 = ~n2798 & n2802 ;
  assign n2804 = n2803 ^ n2801 ;
  assign n2805 = n2586 & n2707 ;
  assign n2806 = n2805 ^ n2588 ;
  assign n2807 = n2806 ^ n696 ;
  assign n2808 = n2807 ^ n842 ;
  assign n2809 = ~n2804 & n2808 ;
  assign n2810 = n2809 ^ n2807 ;
  assign n2811 = n2721 & ~n2810 ;
  assign n2812 = n2811 ^ n2720 ;
  assign n2717 = n2598 & n2707 ;
  assign n2718 = n2717 ^ n2600 ;
  assign n2813 = n2812 ^ n2718 ;
  assign n2814 = n2718 ^ n609 ;
  assign n2815 = ~n2813 & ~n2814 ;
  assign n2816 = n2815 ^ n834 ;
  assign n2817 = n2716 & ~n2816 ;
  assign n2818 = n2817 ^ n750 ;
  assign n2819 = ~n2713 & n2818 ;
  assign n2820 = n2819 ^ n2712 ;
  assign n2821 = n2820 ^ n2709 ;
  assign n2822 = n2710 & ~n2821 ;
  assign n2823 = n2822 ^ n401 ;
  assign n2824 = n2823 ^ n341 ;
  assign n2825 = n2623 & n2707 ;
  assign n2826 = n2825 ^ n2625 ;
  assign n2827 = n2826 ^ n2823 ;
  assign n2828 = n2824 & n2827 ;
  assign n2829 = n2828 ^ n349 ;
  assign n2837 = n2628 & n2707 ;
  assign n2838 = n2837 ^ n2616 ;
  assign n2839 = n2838 ^ n291 ;
  assign n2840 = ~n2829 & ~n2839 ;
  assign n2841 = n2840 ^ n307 ;
  assign n2842 = ~n2630 & n2707 ;
  assign n2843 = n2842 ^ n2632 ;
  assign n2844 = n2843 ^ n245 ;
  assign n2845 = n2841 & n2844 ;
  assign n2846 = n2845 ^ n2843 ;
  assign n2849 = n2848 ^ n2846 ;
  assign n2850 = n2848 ^ n188 ;
  assign n2851 = n2849 & ~n2850 ;
  assign n2852 = n2851 ^ n203 ;
  assign n2853 = n2836 & ~n2852 ;
  assign n2854 = n2853 ^ n2835 ;
  assign n2855 = n2854 ^ n138 ;
  assign n2858 = n2857 ^ n2854 ;
  assign n2859 = ~n2855 & ~n2858 ;
  assign n2861 = n2860 ^ n2859 ;
  assign n2862 = n2861 ^ n2854 ;
  assign n2875 = n130 & n2668 ;
  assign n2876 = n2875 ^ n2656 ;
  assign n2877 = ~n183 & n2876 ;
  assign n2878 = n2877 ^ n2656 ;
  assign n2865 = n2705 ^ n2665 ;
  assign n2863 = n2669 ^ n2667 ;
  assign n2864 = n2863 ^ n2670 ;
  assign n2866 = n2865 ^ n2864 ;
  assign n2867 = ~n183 & n2866 ;
  assign n2868 = n2867 ^ n2865 ;
  assign n2869 = n2656 & n2868 ;
  assign n2870 = n2869 ^ n183 ;
  assign n2879 = n2878 ^ n2870 ;
  assign n2880 = n2879 ^ n2707 ;
  assign n2881 = n2880 ^ n2879 ;
  assign n2883 = n2879 ^ n2878 ;
  assign n2886 = n2612 & ~n2883 ;
  assign n2887 = ~n2881 & n2886 ;
  assign n2888 = n2887 ^ n2881 ;
  assign n2889 = n2888 ^ n2880 ;
  assign n2890 = ~n2705 & n2889 ;
  assign n2891 = n2890 ^ n2878 ;
  assign n2892 = ~n2862 & n2891 ;
  assign n2893 = n2833 & n2892 ;
  assign n2894 = n2893 ^ n2891 ;
  assign n3051 = ~n2855 & n2894 ;
  assign n3052 = n2858 & n3051 ;
  assign n3054 = n2854 ^ n183 ;
  assign n3053 = n2861 ^ n2832 ;
  assign n3055 = n3054 ^ n3053 ;
  assign n3058 = n2859 ^ n2832 ;
  assign n3059 = n2857 ^ n2855 ;
  assign n3060 = ~n3058 & n3059 ;
  assign n3061 = n3055 & n3060 ;
  assign n3056 = n3055 ^ n3052 ;
  assign n3062 = n3061 ^ n3056 ;
  assign n3063 = n3062 ^ n2854 ;
  assign n3064 = n3063 ^ n2857 ;
  assign n3065 = n3064 ^ n183 ;
  assign n3066 = n3065 ^ n3062 ;
  assign n3067 = ~n3052 & n3066 ;
  assign n3068 = n3067 ^ n3063 ;
  assign n3069 = n2832 & ~n3068 ;
  assign n3070 = n3069 ^ n3062 ;
  assign n3071 = n2894 & n3070 ;
  assign n3072 = n3071 ^ n3062 ;
  assign n3079 = n2852 & ~n2894 ;
  assign n3080 = n3079 ^ n2835 ;
  assign n3045 = ~n2841 & ~n2894 ;
  assign n3046 = n3045 ^ n2843 ;
  assign n2895 = ~n2829 & ~n2894 ;
  assign n2896 = n2895 ^ n2838 ;
  assign n2897 = n2896 ^ n245 ;
  assign n2898 = n2820 ^ n401 ;
  assign n2899 = ~n2894 & n2898 ;
  assign n2900 = n2899 ^ n2709 ;
  assign n2901 = n2900 ^ n341 ;
  assign n3030 = ~n2818 & ~n2894 ;
  assign n3031 = n3030 ^ n2712 ;
  assign n2902 = ~n2816 & ~n2894 ;
  assign n2903 = n2902 ^ n2715 ;
  assign n2904 = n2903 ^ n457 ;
  assign n2905 = n2812 ^ n609 ;
  assign n2906 = ~n2894 & ~n2905 ;
  assign n2907 = n2906 ^ n2718 ;
  assign n2908 = n2907 ^ n534 ;
  assign n2909 = n2810 & ~n2894 ;
  assign n2910 = n2909 ^ n2720 ;
  assign n3024 = n2910 ^ n534 ;
  assign n2911 = n2910 ^ n609 ;
  assign n2912 = ~n2778 & ~n2894 ;
  assign n2913 = n2912 ^ n2780 ;
  assign n2914 = n2913 ^ n1136 ;
  assign n2989 = ~n2773 & ~n2894 ;
  assign n2990 = n2989 ^ n2775 ;
  assign n2993 = n2990 ^ n1136 ;
  assign n2915 = ~n2768 & ~n2894 ;
  assign n2916 = n2915 ^ n2770 ;
  assign n2917 = n2916 ^ n1427 ;
  assign n2920 = n2752 & ~n2894 ;
  assign n2921 = n2920 ^ n2755 ;
  assign n2922 = n2921 ^ n2175 ;
  assign n2924 = n2740 ^ n2707 ;
  assign n2925 = ~n2894 & n2924 ;
  assign n2926 = n2925 ^ n2707 ;
  assign n2927 = ~x78 & n2926 ;
  assign n2923 = ~n2737 & ~n2894 ;
  assign n2928 = n2927 ^ n2923 ;
  assign n2929 = n2928 ^ x79 ;
  assign n2930 = n2929 ^ n2366 ;
  assign n2966 = ~n2511 & ~n2707 ;
  assign n2967 = n2894 & n2966 ;
  assign n2956 = n2511 & ~n2707 ;
  assign n2963 = n2956 ^ n2366 ;
  assign n2953 = n2951 ^ x78 ;
  assign n2954 = n2953 ^ n2511 ;
  assign n2952 = n2951 ^ n2707 ;
  assign n2955 = n2954 ^ n2952 ;
  assign n2957 = n2956 ^ n2952 ;
  assign n2934 = n2894 ^ x77 ;
  assign n2958 = n2951 ^ n2934 ;
  assign n2959 = n2958 ^ n2952 ;
  assign n2960 = n2957 & ~n2959 ;
  assign n2961 = n2960 ^ n2952 ;
  assign n2962 = n2955 & n2961 ;
  assign n2964 = n2963 ^ n2962 ;
  assign n2936 = n2934 ^ n2707 ;
  assign n2935 = n2934 ^ n2511 ;
  assign n2937 = n2936 ^ n2935 ;
  assign n2931 = ~x76 & ~n2894 ;
  assign n2932 = n2931 ^ n2894 ;
  assign n2933 = ~x77 & ~n2932 ;
  assign n2938 = n2937 ^ n2933 ;
  assign n2939 = n2938 ^ n2933 ;
  assign n2940 = ~n2934 & ~n2936 ;
  assign n2941 = n2939 & n2940 ;
  assign n2942 = n2941 ^ n2938 ;
  assign n2943 = x78 ^ x77 ;
  assign n2944 = n2943 ^ x78 ;
  assign n2945 = n2894 ^ x78 ;
  assign n2946 = n2945 ^ x78 ;
  assign n2947 = n2944 & ~n2946 ;
  assign n2948 = n2947 ^ x78 ;
  assign n2949 = ~n2942 & ~n2948 ;
  assign n2965 = n2964 ^ n2949 ;
  assign n2968 = n2967 ^ n2965 ;
  assign n2969 = n2930 & n2968 ;
  assign n2970 = n2969 ^ n2399 ;
  assign n2971 = ~n2922 & n2970 ;
  assign n2972 = n2971 ^ n2204 ;
  assign n2973 = n2758 & ~n2894 ;
  assign n2974 = n2973 ^ n2735 ;
  assign n2975 = n2974 ^ n2008 ;
  assign n2976 = n2972 & n2975 ;
  assign n2977 = n2976 ^ n2064 ;
  assign n2978 = n2760 & ~n2894 ;
  assign n2979 = n2978 ^ n2723 ;
  assign n2980 = n2979 ^ n1739 ;
  assign n2981 = ~n2977 & n2980 ;
  assign n2982 = n2981 ^ n1739 ;
  assign n2918 = ~n2762 & ~n2894 ;
  assign n2919 = n2918 ^ n2765 ;
  assign n2983 = n2982 ^ n2919 ;
  assign n2984 = n2919 ^ n1572 ;
  assign n2985 = ~n2983 & ~n2984 ;
  assign n2986 = n2985 ^ n1605 ;
  assign n2987 = n2917 & ~n2986 ;
  assign n2988 = n2987 ^ n1450 ;
  assign n2991 = n2990 ^ n1290 ;
  assign n2992 = n2988 & n2991 ;
  assign n2994 = n2993 ^ n2992 ;
  assign n2995 = ~n2914 & n2994 ;
  assign n2996 = n2995 ^ n1143 ;
  assign n2997 = n2783 ^ n1136 ;
  assign n2998 = ~n2894 & ~n2997 ;
  assign n2999 = n2998 ^ n2785 ;
  assign n3000 = n2999 ^ n892 ;
  assign n3001 = n3000 ^ n892 ;
  assign n3002 = n3001 ^ n1034 ;
  assign n3003 = ~n2996 & ~n3002 ;
  assign n3004 = n3003 ^ n3000 ;
  assign n3005 = n2790 & ~n2894 ;
  assign n3006 = n3005 ^ n2793 ;
  assign n3007 = n3006 ^ n786 ;
  assign n3008 = n3007 ^ n927 ;
  assign n3009 = n3004 & n3008 ;
  assign n3010 = n3009 ^ n3007 ;
  assign n3011 = n2798 & ~n2894 ;
  assign n3012 = n3011 ^ n2800 ;
  assign n3013 = n3012 ^ n696 ;
  assign n3014 = n3013 ^ n842 ;
  assign n3015 = ~n3010 & n3014 ;
  assign n3016 = n3015 ^ n3013 ;
  assign n3017 = n2804 & ~n2894 ;
  assign n3018 = n3017 ^ n2806 ;
  assign n3019 = n3018 ^ n609 ;
  assign n3020 = n3019 ^ n835 ;
  assign n3021 = ~n3016 & n3020 ;
  assign n3022 = n3021 ^ n3019 ;
  assign n3023 = ~n2911 & n3022 ;
  assign n3025 = n3024 ^ n3023 ;
  assign n3026 = n2908 & n3025 ;
  assign n3027 = n3026 ^ n750 ;
  assign n3028 = ~n2904 & n3027 ;
  assign n3029 = n3028 ^ n2903 ;
  assign n3032 = n3031 ^ n3029 ;
  assign n3033 = n3031 ^ n401 ;
  assign n3034 = ~n3032 & n3033 ;
  assign n3035 = n3034 ^ n462 ;
  assign n3036 = n2901 & n3035 ;
  assign n3037 = n3036 ^ n349 ;
  assign n3038 = n2824 & ~n2894 ;
  assign n3039 = n3038 ^ n2826 ;
  assign n3040 = n3039 ^ n291 ;
  assign n3041 = ~n3037 & n3040 ;
  assign n3042 = n3041 ^ n307 ;
  assign n3043 = n2897 & n3042 ;
  assign n3044 = n3043 ^ n2896 ;
  assign n3047 = n3046 ^ n3044 ;
  assign n3048 = n3046 ^ n188 ;
  assign n3049 = ~n3047 & n3048 ;
  assign n3050 = n3049 ^ n203 ;
  assign n3073 = n2846 ^ n188 ;
  assign n3074 = ~n2894 & n3073 ;
  assign n3075 = n3074 ^ n2848 ;
  assign n3076 = n3075 ^ n157 ;
  assign n3077 = ~n3050 & ~n3076 ;
  assign n3078 = n3077 ^ n3075 ;
  assign n3081 = n3080 ^ n3078 ;
  assign n3082 = n3078 ^ n138 ;
  assign n3083 = n3081 & ~n3082 ;
  assign n3084 = n3083 ^ n138 ;
  assign n3085 = n183 & n3084 ;
  assign n3086 = n3085 ^ n3084 ;
  assign n3087 = n3072 & ~n3086 ;
  assign n3088 = n2894 ^ n2855 ;
  assign n3089 = n3088 ^ n3051 ;
  assign n3090 = n3089 ^ n2857 ;
  assign n3091 = n3084 & n3090 ;
  assign n3092 = n3087 & n3091 ;
  assign n3093 = n3092 ^ n3087 ;
  assign n3153 = ~x72 & ~x73 ;
  assign n3195 = ~n3093 & ~n3153 ;
  assign n3196 = n2951 & n3195 ;
  assign n3154 = ~x74 & n3153 ;
  assign n3155 = n3154 ^ x75 ;
  assign n3178 = n3155 ^ n2707 ;
  assign n3179 = n3178 ^ n3093 ;
  assign n3184 = n3179 ^ n2707 ;
  assign n3185 = ~n3093 & ~n3184 ;
  assign n3187 = n3185 ^ n3184 ;
  assign n3188 = ~n3154 & ~n3187 ;
  assign n3186 = n3185 ^ x76 ;
  assign n3189 = n3188 ^ n3186 ;
  assign n3190 = n3188 ^ n3179 ;
  assign n3191 = n3189 & ~n3190 ;
  assign n3158 = n3154 ^ n2707 ;
  assign n3159 = n3158 ^ n3093 ;
  assign n3165 = n2707 ^ x75 ;
  assign n3166 = n3165 ^ n3093 ;
  assign n3167 = ~n3159 & n3166 ;
  assign n3170 = n3165 ^ n3154 ;
  assign n3171 = n3170 ^ n3093 ;
  assign n3174 = ~n3093 & n3171 ;
  assign n3175 = n3174 ^ n2931 ;
  assign n3176 = n3167 & n3175 ;
  assign n3177 = n3176 ^ n3171 ;
  assign n3192 = n3191 ^ n3177 ;
  assign n3156 = n3155 ^ n3093 ;
  assign n3157 = n3156 ^ n3093 ;
  assign n3162 = n3157 & ~n3159 ;
  assign n3163 = n3162 ^ n3156 ;
  assign n3164 = n2932 & n3163 ;
  assign n3193 = n3192 ^ n3164 ;
  assign n3197 = n3196 ^ n3193 ;
  assign n3198 = n3197 ^ n2511 ;
  assign n3200 = n2951 ^ n2932 ;
  assign n3201 = n3200 ^ n2707 ;
  assign n3202 = ~n3093 & ~n3201 ;
  assign n3199 = n2931 ^ x77 ;
  assign n3203 = n3202 ^ n3199 ;
  assign n3204 = n3203 ^ n3197 ;
  assign n3205 = ~n3198 & n3204 ;
  assign n3206 = n3205 ^ n2511 ;
  assign n3151 = n2926 ^ x78 ;
  assign n3143 = n2933 ^ n2737 ;
  assign n3144 = n3143 ^ n2958 ;
  assign n3145 = n3144 ^ n3143 ;
  assign n3146 = n3143 ^ n2936 ;
  assign n3147 = n3146 ^ n3143 ;
  assign n3148 = ~n3145 & n3147 ;
  assign n3149 = n3148 ^ n3143 ;
  assign n3150 = ~n3093 & ~n3149 ;
  assign n3152 = n3151 ^ n3150 ;
  assign n3207 = n3206 ^ n3152 ;
  assign n3208 = n3206 ^ n2366 ;
  assign n3209 = ~n3207 & n3208 ;
  assign n3210 = n3209 ^ n2399 ;
  assign n3109 = ~n3082 & ~n3093 ;
  assign n3110 = n3109 ^ n3080 ;
  assign n3098 = ~n183 & n3080 ;
  assign n3100 = n4971 ^ n3083 ;
  assign n3101 = ~n3072 & ~n3100 ;
  assign n3099 = n4971 ^ n3078 ;
  assign n3102 = n3101 ^ n3099 ;
  assign n3103 = n3098 & n3102 ;
  assign n3104 = n3103 ^ n3101 ;
  assign n3105 = n3104 ^ n3085 ;
  assign n3096 = ~n1355 & ~n3080 ;
  assign n3097 = n3078 & n3096 ;
  assign n3106 = n3105 ^ n3097 ;
  assign n3107 = n3090 & ~n3106 ;
  assign n3108 = n3107 ^ n3104 ;
  assign n3094 = n3050 & ~n3093 ;
  assign n3095 = n3094 ^ n3075 ;
  assign n3114 = ~n3042 & ~n3093 ;
  assign n3115 = n3114 ^ n2896 ;
  assign n3116 = n3115 ^ n188 ;
  assign n3283 = ~n3037 & ~n3093 ;
  assign n3284 = n3283 ^ n3039 ;
  assign n3117 = n3035 & ~n3093 ;
  assign n3118 = n3117 ^ n2900 ;
  assign n3119 = n3118 ^ n291 ;
  assign n3123 = ~n3027 & ~n3093 ;
  assign n3124 = n3123 ^ n2903 ;
  assign n3125 = n3124 ^ n401 ;
  assign n3126 = n3025 & ~n3093 ;
  assign n3127 = n3126 ^ n2907 ;
  assign n3128 = n3127 ^ n457 ;
  assign n3129 = n3016 & ~n3093 ;
  assign n3130 = n3129 ^ n3018 ;
  assign n3131 = n3130 ^ n609 ;
  assign n3132 = ~n2988 & ~n3093 ;
  assign n3133 = n3132 ^ n2990 ;
  assign n3134 = n3133 ^ n1136 ;
  assign n3219 = ~n2977 & ~n3093 ;
  assign n3220 = n3219 ^ n2979 ;
  assign n3223 = n3220 ^ n1427 ;
  assign n3135 = n2972 & ~n3093 ;
  assign n3136 = n3135 ^ n2974 ;
  assign n3137 = n3136 ^ n1739 ;
  assign n3140 = n2968 & ~n3093 ;
  assign n3141 = n3140 ^ n2929 ;
  assign n3142 = n3141 ^ n2175 ;
  assign n3211 = n3142 & n3210 ;
  assign n3212 = n3211 ^ n2175 ;
  assign n3138 = n2970 & ~n3093 ;
  assign n3139 = n3138 ^ n2921 ;
  assign n3213 = n3212 ^ n3139 ;
  assign n3214 = n3212 ^ n2008 ;
  assign n3215 = n3213 & n3214 ;
  assign n3216 = n3215 ^ n2064 ;
  assign n3217 = ~n3137 & ~n3216 ;
  assign n3218 = n3217 ^ n1763 ;
  assign n3221 = n3220 ^ n1572 ;
  assign n3222 = n3218 & ~n3221 ;
  assign n3224 = n3223 ^ n3222 ;
  assign n3225 = n2982 ^ n1572 ;
  assign n3226 = ~n3093 & ~n3225 ;
  assign n3227 = n3226 ^ n2919 ;
  assign n3228 = n3227 ^ n1427 ;
  assign n3229 = n3224 & n3228 ;
  assign n3230 = n3229 ^ n1450 ;
  assign n3231 = ~n2986 & ~n3093 ;
  assign n3232 = n3231 ^ n2916 ;
  assign n3233 = n3232 ^ n1290 ;
  assign n3234 = ~n3230 & ~n3233 ;
  assign n3235 = n3234 ^ n1461 ;
  assign n3236 = n3134 & n3235 ;
  assign n3237 = n3236 ^ n1143 ;
  assign n3238 = n2994 & ~n3093 ;
  assign n3239 = n3238 ^ n2913 ;
  assign n3242 = n3239 ^ n1034 ;
  assign n3243 = ~n3237 & ~n3242 ;
  assign n3240 = n3239 ^ n892 ;
  assign n3244 = n3243 ^ n3240 ;
  assign n3245 = n2996 & ~n3093 ;
  assign n3246 = n3245 ^ n2999 ;
  assign n3247 = n3246 ^ n786 ;
  assign n3248 = n3247 ^ n927 ;
  assign n3249 = n3244 & ~n3248 ;
  assign n3250 = n3249 ^ n3247 ;
  assign n3251 = ~n3004 & ~n3093 ;
  assign n3252 = n3251 ^ n3006 ;
  assign n3253 = n3252 ^ n696 ;
  assign n3254 = n3253 ^ n842 ;
  assign n3255 = n3250 & n3254 ;
  assign n3256 = n3255 ^ n3253 ;
  assign n3257 = n3010 & ~n3093 ;
  assign n3258 = n3257 ^ n3012 ;
  assign n3259 = n3258 ^ n609 ;
  assign n3260 = n3259 ^ n835 ;
  assign n3261 = ~n3256 & n3260 ;
  assign n3262 = n3261 ^ n3259 ;
  assign n3263 = ~n3131 & ~n3262 ;
  assign n3264 = n3263 ^ n834 ;
  assign n3265 = ~n3022 & ~n3093 ;
  assign n3266 = n3265 ^ n2910 ;
  assign n3267 = n3266 ^ n534 ;
  assign n3268 = ~n3264 & n3267 ;
  assign n3269 = n3268 ^ n750 ;
  assign n3270 = ~n3128 & n3269 ;
  assign n3271 = n3270 ^ n3127 ;
  assign n3272 = n3271 ^ n3124 ;
  assign n3273 = n3125 & ~n3272 ;
  assign n3274 = n3273 ^ n401 ;
  assign n3120 = n3029 ^ n401 ;
  assign n3121 = ~n3093 & n3120 ;
  assign n3122 = n3121 ^ n3031 ;
  assign n3275 = n3274 ^ n3122 ;
  assign n3276 = n3274 ^ n341 ;
  assign n3277 = ~n3275 & n3276 ;
  assign n3278 = n3277 ^ n349 ;
  assign n3279 = ~n3119 & ~n3278 ;
  assign n3280 = n3279 ^ n291 ;
  assign n3281 = n3280 ^ n3115 ;
  assign n3282 = n3281 ^ n245 ;
  assign n3285 = n3284 ^ n3282 ;
  assign n3286 = n3285 ^ n3281 ;
  assign n3287 = n3281 ^ n3280 ;
  assign n3288 = n3287 ^ n245 ;
  assign n3289 = n3288 ^ n3281 ;
  assign n3290 = n3286 & ~n3289 ;
  assign n3291 = n3290 ^ n3281 ;
  assign n3292 = n3116 & n3291 ;
  assign n3293 = n3292 ^ n203 ;
  assign n3294 = n3044 ^ n188 ;
  assign n3295 = ~n3093 & n3294 ;
  assign n3296 = n3295 ^ n3046 ;
  assign n3297 = n3296 ^ n157 ;
  assign n3298 = ~n3293 & n3297 ;
  assign n3299 = n3298 ^ n3296 ;
  assign n3304 = n3095 & ~n3299 ;
  assign n3300 = n3299 ^ n3095 ;
  assign n3309 = n3304 ^ n3300 ;
  assign n3301 = n138 & n3300 ;
  assign n3310 = n3309 ^ n3301 ;
  assign n3311 = n3310 ^ n138 ;
  assign n3316 = ~n3108 & n3311 ;
  assign n3317 = n183 & n3316 ;
  assign n3318 = ~n3110 & n3317 ;
  assign n3319 = n3318 ^ n3316 ;
  assign n3320 = n3319 ^ n3108 ;
  assign n3344 = n3210 & n3320 ;
  assign n3345 = n3344 ^ n3141 ;
  assign n3346 = n3345 ^ n2008 ;
  assign n3347 = n3208 & n3320 ;
  assign n3348 = n3347 ^ n3152 ;
  assign n3349 = n3348 ^ n2175 ;
  assign n3359 = n2950 ^ x76 ;
  assign n3355 = n2950 ^ x75 ;
  assign n3356 = ~n3093 & n3355 ;
  assign n3352 = n3154 ^ n2894 ;
  assign n3353 = n3156 & n3352 ;
  assign n3354 = n3353 ^ n3165 ;
  assign n3357 = n3356 ^ n3354 ;
  assign n3358 = n3320 & ~n3357 ;
  assign n3360 = n3359 ^ n3358 ;
  assign n3350 = n2950 ^ n2894 ;
  assign n3351 = n3093 & ~n3350 ;
  assign n3361 = n3360 ^ n3351 ;
  assign n3362 = n3361 ^ n2511 ;
  assign n3373 = ~x74 & ~n3093 ;
  assign n3363 = n3093 ^ n2894 ;
  assign n3364 = n3363 ^ x74 ;
  assign n3365 = n3364 ^ n3363 ;
  assign n3366 = n3153 ^ n3093 ;
  assign n3369 = ~n3365 & ~n3366 ;
  assign n3370 = n3369 ^ n3363 ;
  assign n3371 = n3320 & n3370 ;
  assign n3372 = n3371 ^ x75 ;
  assign n3374 = n3373 ^ n3372 ;
  assign n3375 = n3374 ^ n2707 ;
  assign n3396 = n2894 ^ n2707 ;
  assign n3377 = ~n3320 & ~n3366 ;
  assign n3376 = n3153 ^ x74 ;
  assign n3378 = n3377 ^ n3376 ;
  assign n3379 = n3378 ^ n2894 ;
  assign n3381 = n3320 ^ x73 ;
  assign n3380 = ~x70 & ~x71 ;
  assign n3382 = n3381 ^ n3380 ;
  assign n3383 = n3380 ^ n3093 ;
  assign n3384 = n3382 & ~n3383 ;
  assign n3393 = n3384 ^ n3363 ;
  assign n3387 = n3320 ^ n3093 ;
  assign n3390 = n3381 & ~n3387 ;
  assign n3391 = n3390 ^ n3384 ;
  assign n3392 = x72 & n3391 ;
  assign n3394 = n3393 ^ n3392 ;
  assign n3395 = n3379 & n3394 ;
  assign n3397 = n3396 ^ n3395 ;
  assign n3398 = ~n3375 & ~n3397 ;
  assign n3399 = n3398 ^ n2707 ;
  assign n3400 = n3399 ^ n3361 ;
  assign n3401 = n3362 & n3400 ;
  assign n3402 = n3401 ^ n2530 ;
  assign n3403 = ~n3198 & n3320 ;
  assign n3404 = n3403 ^ n3203 ;
  assign n3405 = n3404 ^ n2366 ;
  assign n3406 = n3402 & n3405 ;
  assign n3407 = n3406 ^ n2399 ;
  assign n3408 = n3349 & n3407 ;
  assign n3409 = n3408 ^ n2204 ;
  assign n3410 = n3346 & n3409 ;
  assign n3411 = n3410 ^ n2008 ;
  assign n3412 = n3411 ^ n1739 ;
  assign n3507 = n3299 ^ n138 ;
  assign n3508 = n3320 & n3507 ;
  assign n3509 = n3508 ^ n3095 ;
  assign n3535 = n3509 ^ n183 ;
  assign n3111 = ~n3108 & ~n3110 ;
  assign n3112 = ~n3095 & n3111 ;
  assign n3113 = n3112 ^ n3111 ;
  assign n3305 = n3108 & n3304 ;
  assign n3302 = n3301 ^ n3110 ;
  assign n3303 = n3302 ^ n3112 ;
  assign n3306 = n3305 ^ n3303 ;
  assign n3307 = ~n183 & n3306 ;
  assign n3308 = n3307 ^ n3112 ;
  assign n3312 = n3311 ^ n3110 ;
  assign n3313 = ~n3308 & n3312 ;
  assign n3314 = n3313 ^ n183 ;
  assign n3315 = ~n3113 & ~n3314 ;
  assign n3325 = ~n3278 & n3320 ;
  assign n3326 = n3325 ^ n3118 ;
  assign n3327 = n3326 ^ n245 ;
  assign n3328 = n3276 & n3320 ;
  assign n3329 = n3328 ^ n3122 ;
  assign n3330 = n3329 ^ n291 ;
  assign n3331 = n3271 ^ n401 ;
  assign n3332 = n3320 & n3331 ;
  assign n3333 = n3332 ^ n3124 ;
  assign n3334 = n3333 ^ n341 ;
  assign n3472 = ~n3269 & n3320 ;
  assign n3473 = n3472 ^ n3127 ;
  assign n3335 = ~n3264 & n3320 ;
  assign n3336 = n3335 ^ n3266 ;
  assign n3337 = n3336 ^ n457 ;
  assign n3338 = ~n3262 & n3320 ;
  assign n3339 = n3338 ^ n3130 ;
  assign n3340 = n3339 ^ n534 ;
  assign n3341 = n3256 & n3320 ;
  assign n3342 = n3341 ^ n3258 ;
  assign n3466 = n3342 ^ n534 ;
  assign n3343 = n3342 ^ n609 ;
  assign n3429 = n3224 & n3320 ;
  assign n3430 = n3429 ^ n3227 ;
  assign n3433 = n3430 ^ n1136 ;
  assign n3418 = ~n3216 & n3320 ;
  assign n3419 = n3418 ^ n3136 ;
  assign n3422 = n3419 ^ n1427 ;
  assign n3413 = n3214 & n3320 ;
  assign n3414 = n3413 ^ n3139 ;
  assign n3415 = n3414 ^ n3411 ;
  assign n3416 = ~n3412 & n3415 ;
  assign n3417 = n3416 ^ n1763 ;
  assign n3420 = n3419 ^ n1572 ;
  assign n3421 = n3417 & n3420 ;
  assign n3423 = n3422 ^ n3421 ;
  assign n3424 = ~n3218 & n3320 ;
  assign n3425 = n3424 ^ n3220 ;
  assign n3426 = n3425 ^ n1427 ;
  assign n3427 = ~n3423 & n3426 ;
  assign n3428 = n3427 ^ n1450 ;
  assign n3431 = n3430 ^ n1290 ;
  assign n3432 = n3428 & ~n3431 ;
  assign n3434 = n3433 ^ n3432 ;
  assign n3435 = ~n3230 & n3320 ;
  assign n3436 = n3435 ^ n3232 ;
  assign n3437 = n3436 ^ n1136 ;
  assign n3438 = ~n3434 & ~n3437 ;
  assign n3439 = n3438 ^ n1143 ;
  assign n3440 = n3235 & n3320 ;
  assign n3441 = n3440 ^ n3133 ;
  assign n3444 = n3441 ^ n1034 ;
  assign n3445 = ~n3439 & n3444 ;
  assign n3442 = n3441 ^ n892 ;
  assign n3446 = n3445 ^ n3442 ;
  assign n3447 = n3237 & n3320 ;
  assign n3448 = n3447 ^ n3239 ;
  assign n3449 = n3448 ^ n786 ;
  assign n3450 = n3449 ^ n927 ;
  assign n3451 = ~n3446 & ~n3450 ;
  assign n3452 = n3451 ^ n3449 ;
  assign n3453 = ~n3244 & n3320 ;
  assign n3454 = n3453 ^ n3246 ;
  assign n3455 = n3454 ^ n696 ;
  assign n3456 = n3455 ^ n842 ;
  assign n3457 = n3452 & ~n3456 ;
  assign n3458 = n3457 ^ n3455 ;
  assign n3459 = ~n3250 & n3320 ;
  assign n3460 = n3459 ^ n3252 ;
  assign n3461 = n3460 ^ n609 ;
  assign n3462 = n3461 ^ n835 ;
  assign n3463 = n3458 & n3462 ;
  assign n3464 = n3463 ^ n3461 ;
  assign n3465 = ~n3343 & n3464 ;
  assign n3467 = n3466 ^ n3465 ;
  assign n3468 = n3340 & n3467 ;
  assign n3469 = n3468 ^ n750 ;
  assign n3470 = ~n3337 & n3469 ;
  assign n3471 = n3470 ^ n3336 ;
  assign n3474 = n3473 ^ n3471 ;
  assign n3475 = n3473 ^ n401 ;
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = n3476 ^ n462 ;
  assign n3478 = n3334 & n3477 ;
  assign n3479 = n3478 ^ n349 ;
  assign n3480 = ~n3330 & ~n3479 ;
  assign n3481 = n3480 ^ n307 ;
  assign n3482 = n3327 & n3481 ;
  assign n3483 = n3482 ^ n3326 ;
  assign n3484 = n3483 ^ n188 ;
  assign n3485 = n3280 ^ n245 ;
  assign n3486 = n3320 & ~n3485 ;
  assign n3487 = n3486 ^ n3284 ;
  assign n3488 = n3487 ^ n3483 ;
  assign n3489 = n3484 & n3488 ;
  assign n3490 = n3489 ^ n203 ;
  assign n3491 = n3280 ^ n188 ;
  assign n3492 = n3491 ^ n245 ;
  assign n3493 = n3492 ^ n3284 ;
  assign n3494 = n3493 ^ n3491 ;
  assign n3495 = n3491 ^ n246 ;
  assign n3496 = n3494 & ~n3495 ;
  assign n3497 = n3496 ^ n3491 ;
  assign n3498 = n3320 & ~n3497 ;
  assign n3499 = n3498 ^ n3115 ;
  assign n3500 = n3499 ^ n157 ;
  assign n3501 = ~n3490 & n3500 ;
  assign n3502 = n3501 ^ n3499 ;
  assign n3321 = n3293 & n3320 ;
  assign n3322 = n3321 ^ n3296 ;
  assign n3503 = n3502 ^ n3322 ;
  assign n3521 = n3322 ^ n138 ;
  assign n3522 = ~n3503 & n3521 ;
  assign n3523 = n3522 ^ n138 ;
  assign n3536 = ~n3315 & n3523 ;
  assign n3537 = n3535 & n3536 ;
  assign n3538 = n3537 ^ n3315 ;
  assign n3564 = ~n3412 & n3538 ;
  assign n3565 = n3564 ^ n3414 ;
  assign n3566 = n3565 ^ n1572 ;
  assign n3567 = n3409 & n3538 ;
  assign n3568 = n3567 ^ n3345 ;
  assign n3569 = n3568 ^ n1739 ;
  assign n3572 = n3402 & n3538 ;
  assign n3573 = n3572 ^ n3404 ;
  assign n3574 = n3573 ^ n2175 ;
  assign n3575 = ~n3397 & n3538 ;
  assign n3576 = n3575 ^ n3374 ;
  assign n3577 = n3576 ^ n2511 ;
  assign n3615 = n3394 & n3538 ;
  assign n3616 = n3615 ^ n3378 ;
  assign n3579 = n3380 ^ n3320 ;
  assign n3580 = n3579 ^ n3387 ;
  assign n3581 = n3580 ^ n3387 ;
  assign n3582 = n3387 ^ x72 ;
  assign n3583 = n3582 ^ n3387 ;
  assign n3584 = n3581 & ~n3583 ;
  assign n3585 = n3584 ^ n3387 ;
  assign n3586 = n3538 & ~n3585 ;
  assign n3587 = n3586 ^ x73 ;
  assign n3578 = ~x72 & n3320 ;
  assign n3588 = n3587 ^ n3578 ;
  assign n3589 = n3588 ^ n2894 ;
  assign n3607 = n3538 & n3579 ;
  assign n3606 = n3320 ^ x72 ;
  assign n3608 = n3607 ^ n3606 ;
  assign n3611 = n3608 ^ n2894 ;
  assign n3590 = n3320 ^ x71 ;
  assign n3591 = n3590 ^ n3538 ;
  assign n3593 = ~x68 & ~x69 ;
  assign n3592 = n3320 ^ x70 ;
  assign n3594 = n3593 ^ n3592 ;
  assign n3595 = ~n3591 & n3594 ;
  assign n3604 = n3595 ^ n3387 ;
  assign n3596 = n3538 ^ n3320 ;
  assign n3597 = n3596 ^ n3595 ;
  assign n3598 = n3597 ^ n3595 ;
  assign n3601 = ~n3590 & n3598 ;
  assign n3602 = n3601 ^ n3595 ;
  assign n3603 = x70 & n3602 ;
  assign n3605 = n3604 ^ n3603 ;
  assign n3609 = n3608 ^ n3093 ;
  assign n3610 = n3605 & n3609 ;
  assign n3612 = n3611 ^ n3610 ;
  assign n3613 = n3589 & n3612 ;
  assign n3614 = n3613 ^ n2894 ;
  assign n3617 = n3616 ^ n3614 ;
  assign n3618 = n3616 ^ n2707 ;
  assign n3619 = ~n3617 & ~n3618 ;
  assign n3620 = n3619 ^ n2707 ;
  assign n3621 = n3620 ^ n3576 ;
  assign n3622 = n3577 & n3621 ;
  assign n3623 = n3622 ^ n2530 ;
  assign n3624 = n3399 ^ n2511 ;
  assign n3625 = n3538 & ~n3624 ;
  assign n3626 = n3625 ^ n3361 ;
  assign n3627 = n3626 ^ n2366 ;
  assign n3628 = n3623 & n3627 ;
  assign n3629 = n3628 ^ n2399 ;
  assign n3630 = n3574 & n3629 ;
  assign n3631 = n3630 ^ n2175 ;
  assign n3570 = n3407 & n3538 ;
  assign n3571 = n3570 ^ n3348 ;
  assign n3632 = n3631 ^ n3571 ;
  assign n3633 = n3631 ^ n2008 ;
  assign n3634 = ~n3632 & n3633 ;
  assign n3635 = n3634 ^ n2064 ;
  assign n3636 = ~n3569 & ~n3635 ;
  assign n3637 = n3636 ^ n1763 ;
  assign n3638 = ~n3566 & ~n3637 ;
  assign n3639 = n3638 ^ n1605 ;
  assign n3640 = ~n3417 & n3538 ;
  assign n3641 = n3640 ^ n3419 ;
  assign n3642 = n3641 ^ n1427 ;
  assign n3643 = ~n3639 & ~n3642 ;
  assign n3644 = n3643 ^ n1450 ;
  assign n3710 = n3502 ^ n138 ;
  assign n3711 = n3538 & n3710 ;
  assign n3712 = n3711 ^ n3322 ;
  assign n3719 = n3712 ^ n183 ;
  assign n3323 = ~n3315 & ~n3322 ;
  assign n3324 = ~n183 & ~n3323 ;
  assign n3504 = n3503 ^ n130 ;
  assign n3505 = n3324 & n3504 ;
  assign n3506 = n3505 ^ n3323 ;
  assign n3510 = n3509 ^ n3315 ;
  assign n3511 = n3510 ^ n3509 ;
  assign n3514 = n3509 ^ n3322 ;
  assign n3515 = n3514 ^ n3509 ;
  assign n3516 = ~n138 & ~n3515 ;
  assign n3517 = n3511 & n3516 ;
  assign n3518 = n3517 ^ n3511 ;
  assign n3519 = n3518 ^ n3510 ;
  assign n3520 = n3506 & n3519 ;
  assign n3524 = n3523 ^ n3509 ;
  assign n3525 = n183 & ~n3524 ;
  assign n3527 = n3323 ^ n3315 ;
  assign n3528 = n3525 & ~n3527 ;
  assign n3530 = ~n138 & ~n3502 ;
  assign n3531 = n3528 & n3530 ;
  assign n3526 = n3525 ^ n183 ;
  assign n3529 = n3528 ^ n3526 ;
  assign n3532 = n3531 ^ n3529 ;
  assign n3533 = ~n3520 & ~n3532 ;
  assign n3539 = n3490 & n3538 ;
  assign n3540 = n3539 ^ n3499 ;
  assign n3541 = n3540 ^ n138 ;
  assign n3544 = ~n3479 & n3538 ;
  assign n3545 = n3544 ^ n3329 ;
  assign n3546 = n3545 ^ n245 ;
  assign n3547 = n3477 & n3538 ;
  assign n3548 = n3547 ^ n3333 ;
  assign n3549 = n3548 ^ n291 ;
  assign n3553 = ~n3469 & n3538 ;
  assign n3554 = n3553 ^ n3336 ;
  assign n3555 = n3554 ^ n401 ;
  assign n3556 = n3467 & n3538 ;
  assign n3557 = n3556 ^ n3339 ;
  assign n3558 = n3557 ^ n457 ;
  assign n3559 = ~n3458 & n3538 ;
  assign n3560 = n3559 ^ n3460 ;
  assign n3561 = n3560 ^ n609 ;
  assign n3645 = ~n3423 & n3538 ;
  assign n3646 = n3645 ^ n3425 ;
  assign n3647 = n3646 ^ n1290 ;
  assign n3648 = n3644 & ~n3647 ;
  assign n3649 = n3648 ^ n3646 ;
  assign n3562 = ~n3428 & n3538 ;
  assign n3563 = n3562 ^ n3430 ;
  assign n3650 = n3649 ^ n3563 ;
  assign n3651 = n3649 ^ n1136 ;
  assign n3652 = ~n3650 & ~n3651 ;
  assign n3653 = n3652 ^ n1143 ;
  assign n3654 = ~n3434 & n3538 ;
  assign n3655 = n3654 ^ n3436 ;
  assign n3656 = n3655 ^ n1034 ;
  assign n3657 = n3653 & ~n3656 ;
  assign n3658 = n3657 ^ n1072 ;
  assign n3659 = n3439 & n3538 ;
  assign n3660 = n3659 ^ n3441 ;
  assign n3663 = n3660 ^ n892 ;
  assign n3664 = ~n3658 & n3663 ;
  assign n3661 = n3660 ^ n786 ;
  assign n3665 = n3664 ^ n3661 ;
  assign n3666 = n3446 & n3538 ;
  assign n3667 = n3666 ^ n3448 ;
  assign n3668 = n3667 ^ n696 ;
  assign n3669 = n3668 ^ n842 ;
  assign n3670 = ~n3665 & ~n3669 ;
  assign n3671 = n3670 ^ n3668 ;
  assign n3672 = ~n3452 & n3538 ;
  assign n3673 = n3672 ^ n3454 ;
  assign n3674 = n3673 ^ n609 ;
  assign n3675 = n3674 ^ n835 ;
  assign n3676 = n3671 & ~n3675 ;
  assign n3677 = n3676 ^ n3674 ;
  assign n3678 = ~n3561 & n3677 ;
  assign n3679 = n3678 ^ n834 ;
  assign n3680 = ~n3464 & n3538 ;
  assign n3681 = n3680 ^ n3342 ;
  assign n3682 = n3681 ^ n534 ;
  assign n3683 = ~n3679 & n3682 ;
  assign n3684 = n3683 ^ n750 ;
  assign n3685 = ~n3558 & n3684 ;
  assign n3686 = n3685 ^ n3557 ;
  assign n3687 = n3686 ^ n3554 ;
  assign n3688 = n3555 & ~n3687 ;
  assign n3689 = n3688 ^ n401 ;
  assign n3550 = n3471 ^ n401 ;
  assign n3551 = n3538 & n3550 ;
  assign n3552 = n3551 ^ n3473 ;
  assign n3690 = n3689 ^ n3552 ;
  assign n3691 = n3689 ^ n341 ;
  assign n3692 = ~n3690 & n3691 ;
  assign n3693 = n3692 ^ n349 ;
  assign n3694 = ~n3549 & ~n3693 ;
  assign n3695 = n3694 ^ n307 ;
  assign n3696 = n3546 & n3695 ;
  assign n3697 = n3696 ^ n3545 ;
  assign n3542 = ~n3481 & n3538 ;
  assign n3543 = n3542 ^ n3326 ;
  assign n3698 = n3697 ^ n3543 ;
  assign n3699 = n3697 ^ n188 ;
  assign n3700 = ~n3698 & n3699 ;
  assign n3701 = n3700 ^ n203 ;
  assign n3702 = n3484 & n3538 ;
  assign n3703 = n3702 ^ n3487 ;
  assign n3704 = n3703 ^ n157 ;
  assign n3705 = n3701 & ~n3704 ;
  assign n3706 = n3705 ^ n157 ;
  assign n3707 = n3706 ^ n3540 ;
  assign n3708 = n3541 & ~n3707 ;
  assign n3709 = n3708 ^ n138 ;
  assign n3720 = ~n3533 & n3709 ;
  assign n3721 = ~n3719 & n3720 ;
  assign n3722 = n3721 ^ n3533 ;
  assign n3753 = ~n3644 & n3722 ;
  assign n3754 = n3753 ^ n3646 ;
  assign n3755 = n3754 ^ n1136 ;
  assign n3844 = ~n3639 & n3722 ;
  assign n3845 = n3844 ^ n3641 ;
  assign n3848 = n3845 ^ n1136 ;
  assign n3756 = ~n3637 & n3722 ;
  assign n3757 = n3756 ^ n3565 ;
  assign n3758 = n3757 ^ n1427 ;
  assign n3759 = ~n3635 & n3722 ;
  assign n3760 = n3759 ^ n3568 ;
  assign n3840 = n3760 ^ n1427 ;
  assign n3761 = n3760 ^ n1572 ;
  assign n3764 = n3629 & n3722 ;
  assign n3765 = n3764 ^ n3573 ;
  assign n3766 = n3765 ^ n2008 ;
  assign n3767 = n3623 & n3722 ;
  assign n3768 = n3767 ^ n3626 ;
  assign n3769 = n3768 ^ n2175 ;
  assign n3770 = n3614 ^ n2707 ;
  assign n3771 = n3722 & ~n3770 ;
  assign n3772 = n3771 ^ n3616 ;
  assign n3773 = n3772 ^ n2511 ;
  assign n3774 = n3612 & n3722 ;
  assign n3775 = n3774 ^ n3588 ;
  assign n3776 = n3775 ^ n2707 ;
  assign n3777 = ~n3605 & n3722 ;
  assign n3778 = n3777 ^ n3608 ;
  assign n3779 = n3778 ^ n2894 ;
  assign n3792 = n3538 ^ x70 ;
  assign n3781 = n3593 ^ n3538 ;
  assign n3791 = n3722 & n3781 ;
  assign n3793 = n3792 ^ n3791 ;
  assign n3794 = n3793 ^ n3320 ;
  assign n3796 = n3538 ^ x69 ;
  assign n3797 = n3796 ^ x68 ;
  assign n3800 = n3797 ^ n3796 ;
  assign n3802 = n3796 ^ n3722 ;
  assign n3803 = ~x66 & ~x67 ;
  assign n3795 = n3722 ^ n3538 ;
  assign n3798 = n3797 ^ n3795 ;
  assign n3804 = n3803 ^ n3798 ;
  assign n3805 = ~n3802 & n3804 ;
  assign n3801 = ~n3796 & ~n3798 ;
  assign n3806 = n3805 ^ n3801 ;
  assign n3807 = ~n3800 & n3806 ;
  assign n3808 = n3807 ^ n3801 ;
  assign n3809 = n3808 ^ n3538 ;
  assign n3810 = n3809 ^ n3793 ;
  assign n3811 = ~n3794 & n3810 ;
  assign n3812 = n3811 ^ n3320 ;
  assign n3816 = n3812 ^ n2894 ;
  assign n3784 = n3596 ^ x70 ;
  assign n3785 = n3784 ^ n3596 ;
  assign n3786 = n3781 & ~n3785 ;
  assign n3787 = n3786 ^ n3596 ;
  assign n3788 = n3722 & n3787 ;
  assign n3789 = n3788 ^ x71 ;
  assign n3780 = ~x70 & n3538 ;
  assign n3790 = n3789 ^ n3780 ;
  assign n3813 = n3812 ^ n3790 ;
  assign n3814 = n3790 ^ n3093 ;
  assign n3815 = ~n3813 & ~n3814 ;
  assign n3817 = n3816 ^ n3815 ;
  assign n3818 = n3779 & ~n3817 ;
  assign n3819 = n3818 ^ n3396 ;
  assign n3820 = ~n3776 & ~n3819 ;
  assign n3821 = n3820 ^ n2707 ;
  assign n3822 = n3821 ^ n3772 ;
  assign n3823 = n3773 & n3822 ;
  assign n3824 = n3823 ^ n2530 ;
  assign n3825 = n3620 ^ n2511 ;
  assign n3826 = n3722 & ~n3825 ;
  assign n3827 = n3826 ^ n3576 ;
  assign n3828 = n3827 ^ n2366 ;
  assign n3829 = n3824 & n3828 ;
  assign n3830 = n3829 ^ n2399 ;
  assign n3831 = n3769 & n3830 ;
  assign n3832 = n3831 ^ n2204 ;
  assign n3833 = n3766 & n3832 ;
  assign n3834 = n3833 ^ n2008 ;
  assign n3762 = n3633 & n3722 ;
  assign n3763 = n3762 ^ n3571 ;
  assign n3835 = n3834 ^ n3763 ;
  assign n3836 = n3834 ^ n1739 ;
  assign n3837 = ~n3835 & ~n3836 ;
  assign n3838 = n3837 ^ n1763 ;
  assign n3839 = n3761 & n3838 ;
  assign n3841 = n3840 ^ n3839 ;
  assign n3842 = n3758 & ~n3841 ;
  assign n3843 = n3842 ^ n1450 ;
  assign n3846 = n3845 ^ n1290 ;
  assign n3847 = n3843 & n3846 ;
  assign n3849 = n3848 ^ n3847 ;
  assign n3850 = ~n3755 & n3849 ;
  assign n3851 = n3850 ^ n1143 ;
  assign n3852 = ~n3651 & n3722 ;
  assign n3853 = n3852 ^ n3563 ;
  assign n3854 = n3853 ^ n1034 ;
  assign n3855 = n3851 & ~n3854 ;
  assign n3856 = n3855 ^ n1072 ;
  assign n3857 = n3653 & n3722 ;
  assign n3858 = n3857 ^ n3655 ;
  assign n3859 = n3858 ^ n892 ;
  assign n3860 = n3856 & ~n3859 ;
  assign n3861 = n3860 ^ n927 ;
  assign n3862 = n3658 & n3722 ;
  assign n3863 = n3862 ^ n3660 ;
  assign n3866 = n3863 ^ n786 ;
  assign n3867 = ~n3861 & n3866 ;
  assign n3864 = n3863 ^ n696 ;
  assign n3868 = n3867 ^ n3864 ;
  assign n3715 = n3709 ^ n183 ;
  assign n3716 = ~n3520 & ~n3715 ;
  assign n3534 = n3533 ^ n3520 ;
  assign n3713 = n3709 & ~n3712 ;
  assign n3714 = ~n3534 & n3713 ;
  assign n3717 = n3716 ^ n3714 ;
  assign n3718 = n3717 ^ n3712 ;
  assign n3723 = n3706 ^ n138 ;
  assign n3724 = n3722 & n3723 ;
  assign n3725 = n3724 ^ n3540 ;
  assign n3726 = n3725 ^ n183 ;
  assign n3730 = n3725 ^ n138 ;
  assign n3727 = n3701 & n3722 ;
  assign n3728 = n3727 ^ n3703 ;
  assign n3729 = n3728 ^ n3725 ;
  assign n3731 = n3730 ^ n3729 ;
  assign n3732 = n3699 & n3722 ;
  assign n3733 = n3732 ^ n3543 ;
  assign n3734 = n3733 ^ n157 ;
  assign n3894 = ~n3695 & n3722 ;
  assign n3895 = n3894 ^ n3545 ;
  assign n3735 = n3691 & n3722 ;
  assign n3736 = n3735 ^ n3552 ;
  assign n3737 = n3736 ^ n291 ;
  assign n3738 = n3686 ^ n401 ;
  assign n3739 = n3722 & n3738 ;
  assign n3740 = n3739 ^ n3554 ;
  assign n3741 = n3740 ^ n341 ;
  assign n3879 = ~n3684 & n3722 ;
  assign n3880 = n3879 ^ n3557 ;
  assign n3742 = ~n3679 & n3722 ;
  assign n3743 = n3742 ^ n3681 ;
  assign n3744 = n3743 ^ n457 ;
  assign n3745 = n3677 & n3722 ;
  assign n3746 = n3745 ^ n3560 ;
  assign n3747 = n3746 ^ n534 ;
  assign n3750 = n3665 & n3722 ;
  assign n3751 = n3750 ^ n3667 ;
  assign n3752 = n3751 ^ n696 ;
  assign n3869 = ~n3752 & ~n3868 ;
  assign n3870 = n3869 ^ n3751 ;
  assign n3748 = ~n3671 & n3722 ;
  assign n3749 = n3748 ^ n3673 ;
  assign n3871 = n3870 ^ n3749 ;
  assign n3872 = n3749 ^ n609 ;
  assign n3873 = ~n3871 & n3872 ;
  assign n3874 = n3873 ^ n834 ;
  assign n3875 = n3747 & ~n3874 ;
  assign n3876 = n3875 ^ n750 ;
  assign n3877 = ~n3744 & n3876 ;
  assign n3878 = n3877 ^ n3743 ;
  assign n3881 = n3880 ^ n3878 ;
  assign n3882 = n3880 ^ n401 ;
  assign n3883 = ~n3881 & n3882 ;
  assign n3884 = n3883 ^ n462 ;
  assign n3885 = n3741 & n3884 ;
  assign n3886 = n3885 ^ n349 ;
  assign n3887 = ~n3737 & ~n3886 ;
  assign n3888 = n3887 ^ n307 ;
  assign n3889 = ~n3693 & n3722 ;
  assign n3890 = n3889 ^ n3548 ;
  assign n3891 = n3890 ^ n245 ;
  assign n3892 = n3888 & n3891 ;
  assign n3893 = n3892 ^ n3890 ;
  assign n3896 = n3895 ^ n3893 ;
  assign n3897 = n3895 ^ n188 ;
  assign n3898 = ~n3896 & n3897 ;
  assign n3899 = n3898 ^ n203 ;
  assign n3900 = n3734 & ~n3899 ;
  assign n3901 = n3900 ^ n3733 ;
  assign n3902 = n3901 ^ n3725 ;
  assign n3903 = n3902 ^ n3730 ;
  assign n3904 = ~n3731 & n3903 ;
  assign n3905 = n3904 ^ n3730 ;
  assign n3906 = ~n3726 & ~n3905 ;
  assign n3907 = n3906 ^ n183 ;
  assign n3908 = ~n3718 & n3907 ;
  assign n3934 = n3868 & ~n3908 ;
  assign n3935 = n3934 ^ n3751 ;
  assign n3937 = n3935 ^ n609 ;
  assign n3938 = n3856 & ~n3908 ;
  assign n3939 = n3938 ^ n3858 ;
  assign n3940 = n3939 ^ n786 ;
  assign n3941 = ~n3838 & ~n3908 ;
  assign n3942 = n3941 ^ n3760 ;
  assign n3943 = n3942 ^ n1427 ;
  assign n4026 = ~n3836 & ~n3908 ;
  assign n4027 = n4026 ^ n3763 ;
  assign n4031 = n4027 ^ n1427 ;
  assign n3944 = n3830 & ~n3908 ;
  assign n3945 = n3944 ^ n3768 ;
  assign n3946 = n3945 ^ n2008 ;
  assign n3947 = n3824 & ~n3908 ;
  assign n3948 = n3947 ^ n3827 ;
  assign n3949 = n3948 ^ n2175 ;
  assign n3950 = ~n3819 & ~n3908 ;
  assign n3951 = n3950 ^ n3775 ;
  assign n3952 = n3951 ^ n2511 ;
  assign n3953 = n3812 ^ n3093 ;
  assign n3954 = ~n3908 & ~n3953 ;
  assign n3955 = n3954 ^ n3790 ;
  assign n3956 = n3955 ^ n2894 ;
  assign n3957 = n3809 ^ n3320 ;
  assign n3958 = ~n3908 & n3957 ;
  assign n3959 = n3958 ^ n3793 ;
  assign n3999 = n3959 ^ n2894 ;
  assign n3960 = n3959 ^ n3093 ;
  assign n3977 = n3803 ^ n3722 ;
  assign n3987 = n3795 ^ x68 ;
  assign n3988 = n3987 ^ n3795 ;
  assign n3989 = n3977 & ~n3988 ;
  assign n3990 = n3989 ^ n3795 ;
  assign n3991 = ~n3908 & n3990 ;
  assign n3992 = n3991 ^ x69 ;
  assign n3984 = ~x68 & n3722 ;
  assign n3993 = n3992 ^ n3984 ;
  assign n3978 = ~n3908 & n3977 ;
  assign n3976 = n3722 ^ x68 ;
  assign n3979 = n3978 ^ n3976 ;
  assign n3962 = n3722 ^ x67 ;
  assign n3963 = n3962 ^ x66 ;
  assign n3966 = n3963 ^ n3962 ;
  assign n3968 = n3962 ^ n3908 ;
  assign n3969 = ~x64 & ~x65 ;
  assign n3961 = n3908 ^ n3722 ;
  assign n3964 = n3963 ^ n3961 ;
  assign n3970 = n3969 ^ n3964 ;
  assign n3971 = n3968 & ~n3970 ;
  assign n3967 = ~n3962 & n3964 ;
  assign n3972 = n3971 ^ n3967 ;
  assign n3973 = ~n3966 & n3972 ;
  assign n3974 = n3973 ^ n3967 ;
  assign n3975 = n3974 ^ n3722 ;
  assign n3980 = n3979 ^ n3975 ;
  assign n3981 = n3979 ^ n3538 ;
  assign n3982 = n3980 & ~n3981 ;
  assign n3983 = n3982 ^ n3538 ;
  assign n3994 = n3993 ^ n3983 ;
  assign n3995 = n3993 ^ n3320 ;
  assign n3996 = n3994 & ~n3995 ;
  assign n3997 = n3996 ^ n3387 ;
  assign n3998 = n3960 & n3997 ;
  assign n4000 = n3999 ^ n3998 ;
  assign n4001 = n3956 & n4000 ;
  assign n4002 = n4001 ^ n3396 ;
  assign n4003 = ~n3817 & ~n3908 ;
  assign n4004 = n4003 ^ n3778 ;
  assign n4005 = n4004 ^ n2707 ;
  assign n4006 = ~n4002 & ~n4005 ;
  assign n4007 = n4006 ^ n2707 ;
  assign n4008 = n4007 ^ n3951 ;
  assign n4009 = n3952 & n4008 ;
  assign n4010 = n4009 ^ n2530 ;
  assign n4011 = n3821 ^ n2511 ;
  assign n4012 = ~n3908 & ~n4011 ;
  assign n4013 = n4012 ^ n3772 ;
  assign n4014 = n4013 ^ n2366 ;
  assign n4015 = n4010 & n4014 ;
  assign n4016 = n4015 ^ n2399 ;
  assign n4017 = n3949 & n4016 ;
  assign n4018 = n4017 ^ n2204 ;
  assign n4019 = n3946 & n4018 ;
  assign n4020 = n4019 ^ n2064 ;
  assign n4021 = n3832 & ~n3908 ;
  assign n4022 = n4021 ^ n3765 ;
  assign n4023 = n4022 ^ n1739 ;
  assign n4024 = ~n4020 & ~n4023 ;
  assign n4025 = n4024 ^ n1739 ;
  assign n4028 = n4027 ^ n4025 ;
  assign n4029 = n4025 ^ n1572 ;
  assign n4030 = ~n4028 & n4029 ;
  assign n4032 = n4031 ^ n4030 ;
  assign n4033 = ~n3943 & ~n4032 ;
  assign n4034 = n4033 ^ n1450 ;
  assign n4035 = ~n3841 & ~n3908 ;
  assign n4036 = n4035 ^ n3757 ;
  assign n4037 = n4036 ^ n1290 ;
  assign n4038 = ~n4034 & ~n4037 ;
  assign n4039 = n4038 ^ n1461 ;
  assign n4040 = ~n3843 & ~n3908 ;
  assign n4041 = n4040 ^ n3845 ;
  assign n4042 = n4041 ^ n1136 ;
  assign n4043 = n4039 & n4042 ;
  assign n4044 = n4043 ^ n1143 ;
  assign n4045 = n3849 & ~n3908 ;
  assign n4046 = n4045 ^ n3754 ;
  assign n4049 = n4046 ^ n1034 ;
  assign n4050 = ~n4044 & ~n4049 ;
  assign n4047 = n4046 ^ n892 ;
  assign n4051 = n4050 ^ n4047 ;
  assign n4052 = n3851 & ~n3908 ;
  assign n4053 = n4052 ^ n3853 ;
  assign n4054 = n4053 ^ n786 ;
  assign n4055 = n4054 ^ n927 ;
  assign n4056 = n4051 & ~n4055 ;
  assign n4057 = n4056 ^ n4054 ;
  assign n4058 = ~n3940 & ~n4057 ;
  assign n4059 = n4058 ^ n842 ;
  assign n4060 = n3861 & ~n3908 ;
  assign n4061 = n4060 ^ n3863 ;
  assign n4064 = n4061 ^ n696 ;
  assign n4065 = ~n4059 & n4064 ;
  assign n4062 = n4061 ^ n609 ;
  assign n4066 = n4065 ^ n4062 ;
  assign n4067 = n3937 & n4066 ;
  assign n3936 = n3935 ^ n534 ;
  assign n4068 = n4067 ^ n3936 ;
  assign n4108 = ~n183 & ~n3728 ;
  assign n4109 = ~n3725 & ~n4108 ;
  assign n4121 = n3901 ^ n3730 ;
  assign n4122 = n4121 ^ n3728 ;
  assign n4123 = n4122 ^ n183 ;
  assign n4117 = n4108 ^ n183 ;
  assign n4118 = ~n3901 & ~n4117 ;
  assign n4126 = n4123 ^ n4118 ;
  assign n4127 = n4108 ^ n3901 ;
  assign n4128 = n4971 ^ n4127 ;
  assign n4129 = n4126 & ~n4128 ;
  assign n4094 = n3901 ^ n138 ;
  assign n4114 = n183 & ~n3725 ;
  assign n4115 = n4970 ^ n4114 ;
  assign n4116 = ~n4094 & n4115 ;
  assign n4130 = n4129 ^ n4116 ;
  assign n4131 = ~n3718 & ~n4130 ;
  assign n4132 = n4109 & n4131 ;
  assign n4133 = n4132 ^ n4130 ;
  assign n3911 = n3893 ^ n188 ;
  assign n3912 = ~n3908 & n3911 ;
  assign n3913 = n3912 ^ n3895 ;
  assign n3915 = n3913 ^ n157 ;
  assign n3918 = ~n3886 & ~n3908 ;
  assign n3919 = n3918 ^ n3736 ;
  assign n3920 = n3919 ^ n245 ;
  assign n3921 = n3884 & ~n3908 ;
  assign n3922 = n3921 ^ n3740 ;
  assign n3923 = n3922 ^ n291 ;
  assign n4076 = n3878 ^ n401 ;
  assign n4077 = ~n3908 & n4076 ;
  assign n4078 = n4077 ^ n3880 ;
  assign n3924 = ~n3876 & ~n3908 ;
  assign n3925 = n3924 ^ n3743 ;
  assign n3926 = n3925 ^ n401 ;
  assign n3927 = ~n3874 & ~n3908 ;
  assign n3928 = n3927 ^ n3746 ;
  assign n3929 = n3928 ^ n457 ;
  assign n3930 = n3870 ^ n609 ;
  assign n3931 = ~n3908 & n3930 ;
  assign n3932 = n3931 ^ n3749 ;
  assign n3933 = n3932 ^ n534 ;
  assign n4069 = ~n3933 & ~n4068 ;
  assign n4070 = n4069 ^ n750 ;
  assign n4071 = ~n3929 & n4070 ;
  assign n4072 = n4071 ^ n3928 ;
  assign n4073 = n4072 ^ n3925 ;
  assign n4074 = n3926 & ~n4073 ;
  assign n4075 = n4074 ^ n401 ;
  assign n4079 = n4078 ^ n4075 ;
  assign n4080 = n4078 ^ n341 ;
  assign n4081 = ~n4079 & n4080 ;
  assign n4082 = n4081 ^ n349 ;
  assign n4083 = ~n3923 & ~n4082 ;
  assign n4084 = n4083 ^ n307 ;
  assign n4085 = n3920 & n4084 ;
  assign n4086 = n4085 ^ n3919 ;
  assign n3916 = ~n3888 & ~n3908 ;
  assign n3917 = n3916 ^ n3890 ;
  assign n4087 = n4086 ^ n3917 ;
  assign n4088 = n4086 ^ n188 ;
  assign n4089 = ~n4087 & n4088 ;
  assign n4090 = n4089 ^ n203 ;
  assign n4091 = n3915 & ~n4090 ;
  assign n3914 = n3913 ^ n138 ;
  assign n4092 = n4091 ^ n3914 ;
  assign n3909 = n3899 & ~n3908 ;
  assign n3910 = n3909 ^ n3733 ;
  assign n4098 = n3910 ^ n138 ;
  assign n4099 = n4092 & n4098 ;
  assign n4100 = n4099 ^ n138 ;
  assign n4095 = ~n3908 & n4094 ;
  assign n4096 = n4095 ^ n3728 ;
  assign n4145 = n183 & n4096 ;
  assign n4151 = n4100 & ~n4145 ;
  assign n4152 = n4133 & n4151 ;
  assign n4153 = n4152 ^ n4133 ;
  assign n4165 = ~n4068 & ~n4153 ;
  assign n4166 = n4165 ^ n3932 ;
  assign n4167 = n4166 ^ n457 ;
  assign n4168 = ~n4057 & ~n4153 ;
  assign n4169 = n4168 ^ n3939 ;
  assign n4170 = n4169 ^ n696 ;
  assign n4275 = ~n4034 & ~n4153 ;
  assign n4276 = n4275 ^ n4036 ;
  assign n4259 = ~n4020 & ~n4153 ;
  assign n4260 = n4259 ^ n4022 ;
  assign n4263 = n4260 ^ n1427 ;
  assign n4171 = n4016 & ~n4153 ;
  assign n4172 = n4171 ^ n3948 ;
  assign n4173 = n4172 ^ n2008 ;
  assign n4174 = n4010 & ~n4153 ;
  assign n4175 = n4174 ^ n4013 ;
  assign n4176 = n4175 ^ n2175 ;
  assign n4177 = ~n4002 & ~n4153 ;
  assign n4178 = n4177 ^ n4004 ;
  assign n4179 = n4178 ^ n2511 ;
  assign n4180 = n4000 & ~n4153 ;
  assign n4181 = n4180 ^ n3955 ;
  assign n4182 = n4181 ^ n2707 ;
  assign n4233 = ~n3997 & ~n4153 ;
  assign n4234 = n4233 ^ n3959 ;
  assign n4183 = n3983 ^ n3320 ;
  assign n4184 = ~n4153 & n4183 ;
  assign n4185 = n4184 ^ n3993 ;
  assign n4186 = n4185 ^ n3093 ;
  assign n4224 = n3975 ^ n3538 ;
  assign n4225 = ~n4153 & n4224 ;
  assign n4226 = n4225 ^ n3979 ;
  assign n4188 = n3969 ^ n3908 ;
  assign n4189 = ~n4153 & ~n4188 ;
  assign n4187 = n3908 ^ x66 ;
  assign n4190 = n4189 ^ n4187 ;
  assign n4191 = n4190 ^ n3722 ;
  assign n4194 = n4153 ^ n3908 ;
  assign n4192 = n3908 ^ x65 ;
  assign n4193 = n4192 ^ x64 ;
  assign n4195 = n4194 ^ n4193 ;
  assign n4196 = n4195 ^ n4194 ;
  assign n4197 = n4196 ^ n4192 ;
  assign n4199 = n4192 ^ n4153 ;
  assign n4200 = ~x62 & ~x63 ;
  assign n4201 = n4200 ^ n4195 ;
  assign n4202 = ~n4199 & ~n4201 ;
  assign n4198 = n4192 & n4194 ;
  assign n4203 = n4202 ^ n4198 ;
  assign n4204 = ~n4197 & n4203 ;
  assign n4205 = n4204 ^ n4198 ;
  assign n4206 = n4205 ^ n3908 ;
  assign n4207 = n4206 ^ n4190 ;
  assign n4208 = n4191 & n4207 ;
  assign n4209 = n4208 ^ n3722 ;
  assign n4210 = n4209 ^ n3538 ;
  assign n4212 = n4188 ^ n3961 ;
  assign n4213 = n4212 ^ n3961 ;
  assign n4214 = n3961 ^ x66 ;
  assign n4215 = n4214 ^ n3961 ;
  assign n4216 = ~n4213 & ~n4215 ;
  assign n4217 = n4216 ^ n3961 ;
  assign n4218 = ~n4153 & ~n4217 ;
  assign n4219 = n4218 ^ x67 ;
  assign n4211 = ~x66 & ~n3908 ;
  assign n4220 = n4219 ^ n4211 ;
  assign n4221 = n4220 ^ n4209 ;
  assign n4222 = n4210 & n4221 ;
  assign n4223 = n4222 ^ n3538 ;
  assign n4227 = n4226 ^ n4223 ;
  assign n4228 = n4226 ^ n3320 ;
  assign n4229 = n4227 & ~n4228 ;
  assign n4230 = n4229 ^ n3387 ;
  assign n4231 = n4186 & n4230 ;
  assign n4232 = n4231 ^ n4185 ;
  assign n4235 = n4234 ^ n4232 ;
  assign n4236 = n4234 ^ n2894 ;
  assign n4237 = ~n4235 & n4236 ;
  assign n4238 = n4237 ^ n3396 ;
  assign n4239 = ~n4182 & ~n4238 ;
  assign n4240 = n4239 ^ n2707 ;
  assign n4241 = n4240 ^ n4178 ;
  assign n4242 = n4179 & n4241 ;
  assign n4243 = n4242 ^ n2530 ;
  assign n4244 = n4007 ^ n2511 ;
  assign n4245 = ~n4153 & ~n4244 ;
  assign n4246 = n4245 ^ n3951 ;
  assign n4247 = n4246 ^ n2366 ;
  assign n4248 = n4243 & n4247 ;
  assign n4249 = n4248 ^ n2399 ;
  assign n4250 = n4176 & n4249 ;
  assign n4251 = n4250 ^ n2204 ;
  assign n4252 = n4173 & n4251 ;
  assign n4253 = n4252 ^ n2064 ;
  assign n4254 = n4018 & ~n4153 ;
  assign n4255 = n4254 ^ n3945 ;
  assign n4256 = n4255 ^ n1739 ;
  assign n4257 = ~n4253 & ~n4256 ;
  assign n4258 = n4257 ^ n1763 ;
  assign n4261 = n4260 ^ n1572 ;
  assign n4262 = n4258 & n4261 ;
  assign n4264 = n4263 ^ n4262 ;
  assign n4265 = ~n4029 & ~n4153 ;
  assign n4266 = n4265 ^ n4027 ;
  assign n4267 = n4266 ^ n1427 ;
  assign n4268 = ~n4264 & ~n4267 ;
  assign n4269 = n4268 ^ n1450 ;
  assign n4270 = ~n4032 & ~n4153 ;
  assign n4271 = n4270 ^ n3942 ;
  assign n4272 = n4271 ^ n1290 ;
  assign n4273 = n4269 & n4272 ;
  assign n4274 = n4273 ^ n4271 ;
  assign n4277 = n4276 ^ n4274 ;
  assign n4278 = n4276 ^ n1136 ;
  assign n4279 = n4277 & ~n4278 ;
  assign n4280 = n4279 ^ n1143 ;
  assign n4281 = n4039 & ~n4153 ;
  assign n4282 = n4281 ^ n4041 ;
  assign n4285 = n4282 ^ n1034 ;
  assign n4286 = ~n4280 & n4285 ;
  assign n4283 = n4282 ^ n892 ;
  assign n4287 = n4286 ^ n4283 ;
  assign n4288 = n4044 & ~n4153 ;
  assign n4289 = n4288 ^ n4046 ;
  assign n4290 = n4289 ^ n786 ;
  assign n4291 = n4290 ^ n927 ;
  assign n4292 = ~n4287 & ~n4291 ;
  assign n4293 = n4292 ^ n4290 ;
  assign n4294 = ~n4051 & ~n4153 ;
  assign n4295 = n4294 ^ n4053 ;
  assign n4296 = n4295 ^ n696 ;
  assign n4297 = n4296 ^ n842 ;
  assign n4298 = n4293 & ~n4297 ;
  assign n4299 = n4298 ^ n4296 ;
  assign n4300 = ~n4170 & ~n4299 ;
  assign n4301 = n4300 ^ n835 ;
  assign n4302 = n4059 & ~n4153 ;
  assign n4303 = n4302 ^ n4061 ;
  assign n4304 = n4303 ^ n609 ;
  assign n4305 = ~n4301 & ~n4304 ;
  assign n4306 = n4305 ^ n834 ;
  assign n4307 = ~n4066 & ~n4153 ;
  assign n4308 = n4307 ^ n3935 ;
  assign n4309 = n4308 ^ n534 ;
  assign n4310 = ~n4306 & ~n4309 ;
  assign n4311 = n4310 ^ n750 ;
  assign n4312 = n4167 & n4311 ;
  assign n4313 = n4312 ^ n4166 ;
  assign n4314 = n4313 ^ n401 ;
  assign n4093 = n4092 ^ n3910 ;
  assign n4097 = n4096 ^ n183 ;
  assign n4101 = n4100 ^ n4097 ;
  assign n4102 = ~n138 & ~n3910 ;
  assign n4103 = n4102 ^ n4098 ;
  assign n4104 = n4103 ^ n4096 ;
  assign n4105 = ~n4101 & n4104 ;
  assign n4106 = n4093 & n4105 ;
  assign n4107 = n4106 ^ n4101 ;
  assign n4134 = n4107 ^ n4096 ;
  assign n4135 = n4134 ^ n4107 ;
  assign n4136 = n4107 ^ n4102 ;
  assign n4137 = n4136 ^ n4107 ;
  assign n4138 = ~n4135 & n4137 ;
  assign n4139 = n4138 ^ n4107 ;
  assign n4140 = n4133 & n4139 ;
  assign n4141 = n4140 ^ n4107 ;
  assign n4142 = n4107 & ~n4141 ;
  assign n4143 = n3910 ^ n183 ;
  assign n4144 = n4097 ^ n3910 ;
  assign n4146 = n4145 ^ n4144 ;
  assign n4147 = n4143 & ~n4146 ;
  assign n4148 = n4147 ^ n4096 ;
  assign n4149 = n4142 & ~n4148 ;
  assign n4150 = n4149 ^ n4141 ;
  assign n4347 = n4092 & ~n4153 ;
  assign n4348 = n4347 ^ n3910 ;
  assign n4341 = n4090 & ~n4153 ;
  assign n4342 = n4341 ^ n3913 ;
  assign n4154 = n4088 & ~n4153 ;
  assign n4155 = n4154 ^ n3917 ;
  assign n4156 = n4155 ^ n157 ;
  assign n4333 = ~n4084 & ~n4153 ;
  assign n4334 = n4333 ^ n3919 ;
  assign n4157 = ~n4082 & ~n4153 ;
  assign n4158 = n4157 ^ n3922 ;
  assign n4159 = n4158 ^ n245 ;
  assign n4160 = n4075 ^ n341 ;
  assign n4161 = ~n4153 & n4160 ;
  assign n4162 = n4161 ^ n4078 ;
  assign n4163 = n4162 ^ n245 ;
  assign n4164 = n4163 ^ n307 ;
  assign n4315 = ~n4070 & ~n4153 ;
  assign n4316 = n4315 ^ n3928 ;
  assign n4317 = n4316 ^ n4313 ;
  assign n4318 = ~n4314 & n4317 ;
  assign n4319 = n4318 ^ n462 ;
  assign n4320 = n4072 ^ n401 ;
  assign n4321 = ~n4153 & n4320 ;
  assign n4322 = n4321 ^ n3925 ;
  assign n4323 = n4322 ^ n341 ;
  assign n4324 = n4319 & n4323 ;
  assign n4325 = n4324 ^ n341 ;
  assign n4326 = n4325 ^ n291 ;
  assign n4329 = ~n4164 & ~n4326 ;
  assign n4330 = n4329 ^ n307 ;
  assign n4331 = n4159 & n4330 ;
  assign n4332 = n4331 ^ n4158 ;
  assign n4335 = n4334 ^ n4332 ;
  assign n4336 = n4334 ^ n188 ;
  assign n4337 = ~n4335 & n4336 ;
  assign n4338 = n4337 ^ n203 ;
  assign n4339 = n4156 & ~n4338 ;
  assign n4340 = n4339 ^ n4155 ;
  assign n4343 = n4342 ^ n4340 ;
  assign n4344 = n4342 ^ n138 ;
  assign n4345 = ~n4343 & n4344 ;
  assign n4346 = n4345 ^ n138 ;
  assign n4351 = n183 & n4346 ;
  assign n4354 = ~n4348 & n4351 ;
  assign n4355 = n4354 ^ n4346 ;
  assign n4356 = ~n4150 & ~n4355 ;
  assign n4373 = ~n4314 & ~n4356 ;
  assign n4374 = n4373 ^ n4316 ;
  assign n4375 = n4374 ^ n341 ;
  assign n4529 = ~n4311 & ~n4356 ;
  assign n4530 = n4529 ^ n4166 ;
  assign n4376 = ~n4306 & ~n4356 ;
  assign n4377 = n4376 ^ n4308 ;
  assign n4378 = n4377 ^ n457 ;
  assign n4379 = ~n4301 & ~n4356 ;
  assign n4380 = n4379 ^ n4303 ;
  assign n4381 = n4380 ^ n534 ;
  assign n4382 = ~n4299 & ~n4356 ;
  assign n4383 = n4382 ^ n4169 ;
  assign n4384 = n4383 ^ n609 ;
  assign n4385 = n4274 ^ n1136 ;
  assign n4386 = ~n4356 & n4385 ;
  assign n4387 = n4386 ^ n4276 ;
  assign n4388 = n4387 ^ n1034 ;
  assign n4491 = ~n4264 & ~n4356 ;
  assign n4492 = n4491 ^ n4266 ;
  assign n4495 = n4492 ^ n1136 ;
  assign n4480 = ~n4253 & ~n4356 ;
  assign n4481 = n4480 ^ n4255 ;
  assign n4484 = n4481 ^ n1427 ;
  assign n4389 = n4251 & ~n4356 ;
  assign n4390 = n4389 ^ n4172 ;
  assign n4391 = n4390 ^ n1739 ;
  assign n4394 = n4243 & ~n4356 ;
  assign n4395 = n4394 ^ n4246 ;
  assign n4396 = n4395 ^ n2175 ;
  assign n4397 = ~n4238 & ~n4356 ;
  assign n4398 = n4397 ^ n4181 ;
  assign n4399 = n4398 ^ n2511 ;
  assign n4456 = n4232 ^ n2894 ;
  assign n4457 = ~n4356 & n4456 ;
  assign n4458 = n4457 ^ n4234 ;
  assign n4400 = ~n4230 & ~n4356 ;
  assign n4401 = n4400 ^ n4185 ;
  assign n4402 = n4401 ^ n2894 ;
  assign n4447 = n4223 ^ n3320 ;
  assign n4448 = ~n4356 & n4447 ;
  assign n4449 = n4448 ^ n4226 ;
  assign n4452 = n4449 ^ n2894 ;
  assign n4403 = n4206 ^ n3722 ;
  assign n4404 = ~n4356 & ~n4403 ;
  assign n4405 = n4404 ^ n4190 ;
  assign n4406 = n4405 ^ n3538 ;
  assign n4407 = n4200 ^ n4153 ;
  assign n4408 = ~n4356 & ~n4407 ;
  assign n4409 = n4408 ^ n4153 ;
  assign n4410 = n4409 ^ x64 ;
  assign n4411 = n4410 ^ n3908 ;
  assign n4414 = n4356 ^ n4153 ;
  assign n4412 = n4153 ^ x63 ;
  assign n4413 = n4412 ^ x62 ;
  assign n4415 = n4414 ^ n4413 ;
  assign n4416 = n4415 ^ n4414 ;
  assign n4417 = n4416 ^ n4412 ;
  assign n4419 = n4412 ^ n4356 ;
  assign n4420 = ~x60 & ~x61 ;
  assign n4421 = n4420 ^ n4415 ;
  assign n4422 = ~n4419 & ~n4421 ;
  assign n4418 = n4412 & n4414 ;
  assign n4423 = n4422 ^ n4418 ;
  assign n4424 = ~n4417 & n4423 ;
  assign n4425 = n4424 ^ n4418 ;
  assign n4426 = n4425 ^ n4153 ;
  assign n4427 = n4426 ^ n4410 ;
  assign n4428 = ~n4411 & n4427 ;
  assign n4429 = n4428 ^ n3908 ;
  assign n4430 = n4429 ^ n3722 ;
  assign n4434 = n4153 ^ x65 ;
  assign n4432 = n4200 ^ n3908 ;
  assign n4433 = ~n4356 & ~n4432 ;
  assign n4435 = n4434 ^ n4433 ;
  assign n4431 = x64 & ~n4409 ;
  assign n4436 = n4435 ^ n4431 ;
  assign n4437 = n4436 ^ n4429 ;
  assign n4438 = ~n4430 & n4437 ;
  assign n4439 = n4438 ^ n3795 ;
  assign n4440 = n4406 & n4439 ;
  assign n4441 = n4440 ^ n3596 ;
  assign n4442 = n4210 & ~n4356 ;
  assign n4443 = n4442 ^ n4220 ;
  assign n4444 = n4443 ^ n3320 ;
  assign n4445 = n4441 & ~n4444 ;
  assign n4446 = n4445 ^ n3387 ;
  assign n4450 = n4449 ^ n3093 ;
  assign n4451 = n4446 & n4450 ;
  assign n4453 = n4452 ^ n4451 ;
  assign n4454 = n4402 & n4453 ;
  assign n4455 = n4454 ^ n2894 ;
  assign n4459 = n4458 ^ n4455 ;
  assign n4460 = n4458 ^ n2707 ;
  assign n4461 = ~n4459 & ~n4460 ;
  assign n4462 = n4461 ^ n2707 ;
  assign n4463 = n4462 ^ n4398 ;
  assign n4464 = n4399 & n4463 ;
  assign n4465 = n4464 ^ n2530 ;
  assign n4466 = n4240 ^ n2511 ;
  assign n4467 = ~n4356 & ~n4466 ;
  assign n4468 = n4467 ^ n4178 ;
  assign n4469 = n4468 ^ n2366 ;
  assign n4470 = n4465 & n4469 ;
  assign n4471 = n4470 ^ n2399 ;
  assign n4472 = n4396 & n4471 ;
  assign n4473 = n4472 ^ n2175 ;
  assign n4392 = n4249 & ~n4356 ;
  assign n4393 = n4392 ^ n4175 ;
  assign n4474 = n4473 ^ n4393 ;
  assign n4475 = n4473 ^ n2008 ;
  assign n4476 = ~n4474 & n4475 ;
  assign n4477 = n4476 ^ n2064 ;
  assign n4478 = ~n4391 & ~n4477 ;
  assign n4479 = n4478 ^ n1763 ;
  assign n4482 = n4481 ^ n1572 ;
  assign n4483 = n4479 & n4482 ;
  assign n4485 = n4484 ^ n4483 ;
  assign n4486 = ~n4258 & ~n4356 ;
  assign n4487 = n4486 ^ n4260 ;
  assign n4488 = n4487 ^ n1427 ;
  assign n4489 = ~n4485 & ~n4488 ;
  assign n4490 = n4489 ^ n1450 ;
  assign n4493 = n4492 ^ n1290 ;
  assign n4494 = n4490 & n4493 ;
  assign n4496 = n4495 ^ n4494 ;
  assign n4497 = ~n4269 & ~n4356 ;
  assign n4498 = n4497 ^ n4271 ;
  assign n4499 = n4498 ^ n1136 ;
  assign n4500 = n4496 & n4499 ;
  assign n4501 = n4500 ^ n1143 ;
  assign n4502 = ~n4388 & n4501 ;
  assign n4503 = n4502 ^ n1072 ;
  assign n4504 = n4280 & ~n4356 ;
  assign n4505 = n4504 ^ n4282 ;
  assign n4508 = n4505 ^ n892 ;
  assign n4509 = ~n4503 & n4508 ;
  assign n4506 = n4505 ^ n786 ;
  assign n4510 = n4509 ^ n4506 ;
  assign n4511 = n4287 & ~n4356 ;
  assign n4512 = n4511 ^ n4289 ;
  assign n4513 = n4512 ^ n696 ;
  assign n4514 = n4513 ^ n842 ;
  assign n4515 = ~n4510 & ~n4514 ;
  assign n4516 = n4515 ^ n4513 ;
  assign n4517 = ~n4293 & ~n4356 ;
  assign n4518 = n4517 ^ n4295 ;
  assign n4519 = n4518 ^ n609 ;
  assign n4520 = n4519 ^ n835 ;
  assign n4521 = n4516 & ~n4520 ;
  assign n4522 = n4521 ^ n4519 ;
  assign n4523 = n4384 & n4522 ;
  assign n4524 = n4523 ^ n834 ;
  assign n4525 = n4381 & ~n4524 ;
  assign n4526 = n4525 ^ n750 ;
  assign n4527 = n4378 & n4526 ;
  assign n4528 = n4527 ^ n4377 ;
  assign n4531 = n4530 ^ n4528 ;
  assign n4532 = n4530 ^ n401 ;
  assign n4533 = ~n4531 & ~n4532 ;
  assign n4534 = n4533 ^ n462 ;
  assign n4535 = n4375 & n4534 ;
  assign n4536 = n4535 ^ n341 ;
  assign n4537 = n4536 ^ n291 ;
  assign n4548 = ~n4150 & ~n4342 ;
  assign n4560 = n4548 ^ n4342 ;
  assign n4561 = ~n1355 & ~n4340 ;
  assign n4562 = ~n4560 & n4561 ;
  assign n4563 = n4562 ^ n4351 ;
  assign n4549 = n4340 ^ n138 ;
  assign n4550 = n4549 ^ n4342 ;
  assign n4551 = ~n4548 & n4550 ;
  assign n4552 = ~n183 & n4551 ;
  assign n4553 = n4552 ^ n4351 ;
  assign n4554 = n4553 ^ n4552 ;
  assign n4557 = ~n4150 & n4554 ;
  assign n4558 = n4557 ^ n4552 ;
  assign n4559 = ~n4348 & ~n4558 ;
  assign n4564 = n4563 ^ n4559 ;
  assign n4565 = n4338 & ~n4356 ;
  assign n4566 = n4565 ^ n4155 ;
  assign n4567 = n4566 ^ n138 ;
  assign n4366 = ~n4326 & ~n4356 ;
  assign n4367 = n4366 ^ n4162 ;
  assign n4368 = n4367 ^ n245 ;
  assign n4369 = n4319 & ~n4356 ;
  assign n4370 = n4369 ^ n4322 ;
  assign n4371 = n4370 ^ n245 ;
  assign n4372 = n4371 ^ n307 ;
  assign n4540 = ~n4372 & ~n4537 ;
  assign n4541 = n4540 ^ n307 ;
  assign n4542 = n4368 & n4541 ;
  assign n4543 = n4542 ^ n4367 ;
  assign n4357 = n4162 ^ n307 ;
  assign n4358 = n4357 ^ n4325 ;
  assign n4359 = n4358 ^ n307 ;
  assign n4362 = ~n4164 & ~n4359 ;
  assign n4363 = n4362 ^ n307 ;
  assign n4364 = ~n4356 & ~n4363 ;
  assign n4365 = n4364 ^ n4158 ;
  assign n4544 = n4543 ^ n4365 ;
  assign n4545 = n4543 ^ n188 ;
  assign n4546 = ~n4544 & n4545 ;
  assign n4547 = n4546 ^ n203 ;
  assign n4568 = n4332 ^ n188 ;
  assign n4569 = ~n4356 & n4568 ;
  assign n4570 = n4569 ^ n4334 ;
  assign n4571 = n4570 ^ n157 ;
  assign n4572 = ~n4547 & n4571 ;
  assign n4573 = n4572 ^ n4570 ;
  assign n4574 = n4573 ^ n4566 ;
  assign n4575 = n4567 & ~n4574 ;
  assign n4576 = n4575 ^ n138 ;
  assign n4577 = n4564 & n4576 ;
  assign n4580 = n4552 ^ n183 ;
  assign n4578 = ~n4356 & n4549 ;
  assign n4579 = n4578 ^ n4342 ;
  assign n4581 = n4580 ^ n4579 ;
  assign n4582 = n4577 & ~n4581 ;
  assign n4583 = n4582 ^ n4564 ;
  assign n4590 = ~n4537 & ~n4583 ;
  assign n4591 = n4590 ^ n4370 ;
  assign n4592 = n4591 ^ n245 ;
  assign n4593 = n4534 & ~n4583 ;
  assign n4594 = n4593 ^ n4374 ;
  assign n4595 = n4594 ^ n291 ;
  assign n4596 = n4528 ^ n401 ;
  assign n4597 = ~n4583 & ~n4596 ;
  assign n4598 = n4597 ^ n4530 ;
  assign n4599 = n4598 ^ n341 ;
  assign n4757 = ~n4526 & ~n4583 ;
  assign n4758 = n4757 ^ n4377 ;
  assign n4600 = ~n4524 & ~n4583 ;
  assign n4601 = n4600 ^ n4380 ;
  assign n4602 = n4601 ^ n457 ;
  assign n4603 = ~n4516 & ~n4583 ;
  assign n4604 = n4603 ^ n4518 ;
  assign n4605 = n4604 ^ n609 ;
  assign n4606 = n4501 & ~n4583 ;
  assign n4607 = n4606 ^ n4387 ;
  assign n4608 = n4607 ^ n892 ;
  assign n4720 = ~n4490 & ~n4583 ;
  assign n4721 = n4720 ^ n4492 ;
  assign n4609 = ~n4477 & ~n4583 ;
  assign n4610 = n4609 ^ n4390 ;
  assign n4708 = n4610 ^ n1427 ;
  assign n4611 = n4610 ^ n1572 ;
  assign n4614 = n4471 & ~n4583 ;
  assign n4615 = n4614 ^ n4395 ;
  assign n4616 = n4615 ^ n2008 ;
  assign n4617 = n4465 & ~n4583 ;
  assign n4618 = n4617 ^ n4468 ;
  assign n4619 = n4618 ^ n2175 ;
  assign n4620 = n4455 ^ n2707 ;
  assign n4621 = ~n4583 & ~n4620 ;
  assign n4622 = n4621 ^ n4458 ;
  assign n4623 = n4622 ^ n2511 ;
  assign n4624 = n4453 & ~n4583 ;
  assign n4625 = n4624 ^ n4401 ;
  assign n4626 = n4625 ^ n2707 ;
  assign n4627 = ~n4446 & ~n4583 ;
  assign n4628 = n4627 ^ n4449 ;
  assign n4629 = n4628 ^ n2894 ;
  assign n4630 = n4441 & ~n4583 ;
  assign n4631 = n4630 ^ n4443 ;
  assign n4684 = n4631 ^ n2894 ;
  assign n4632 = n4631 ^ n3093 ;
  assign n4677 = n4439 & ~n4583 ;
  assign n4678 = n4677 ^ n4405 ;
  assign n4633 = n4426 ^ n3908 ;
  assign n4634 = ~n4583 & n4633 ;
  assign n4635 = n4634 ^ n4410 ;
  assign n4636 = n4635 ^ n3722 ;
  assign n4653 = n4420 ^ n4356 ;
  assign n4654 = n4583 & ~n4653 ;
  assign n4655 = n4654 ^ n4420 ;
  assign n4664 = x62 & n4655 ;
  assign n4661 = n4420 ^ n4153 ;
  assign n4662 = ~n4583 & ~n4661 ;
  assign n4660 = n4356 ^ x63 ;
  assign n4663 = n4662 ^ n4660 ;
  assign n4665 = n4664 ^ n4663 ;
  assign n4638 = ~x58 & ~x59 ;
  assign n4639 = n4638 ^ x60 ;
  assign n4637 = n4583 ^ x61 ;
  assign n4640 = n4639 ^ n4637 ;
  assign n4641 = n4637 ^ n4356 ;
  assign n4642 = ~n4640 & ~n4641 ;
  assign n4651 = n4642 ^ n4414 ;
  assign n4643 = n4642 ^ n4637 ;
  assign n4644 = n4643 ^ n4642 ;
  assign n4645 = n4583 ^ n4356 ;
  assign n4646 = n4645 ^ n4642 ;
  assign n4647 = n4646 ^ n4642 ;
  assign n4648 = ~n4644 & n4647 ;
  assign n4649 = n4648 ^ n4642 ;
  assign n4650 = x60 & n4649 ;
  assign n4652 = n4651 ^ n4650 ;
  assign n4656 = n4655 ^ x62 ;
  assign n4657 = n4656 ^ n4153 ;
  assign n4658 = n4652 & n4657 ;
  assign n4659 = n4658 ^ n4153 ;
  assign n4666 = n4665 ^ n4659 ;
  assign n4667 = n4665 ^ n3908 ;
  assign n4668 = n4666 & ~n4667 ;
  assign n4669 = n4668 ^ n3961 ;
  assign n4670 = n4636 & ~n4669 ;
  assign n4671 = n4670 ^ n3795 ;
  assign n4672 = ~n4430 & ~n4583 ;
  assign n4673 = n4672 ^ n4436 ;
  assign n4674 = n4673 ^ n3538 ;
  assign n4675 = n4671 & n4674 ;
  assign n4676 = n4675 ^ n3538 ;
  assign n4679 = n4678 ^ n4676 ;
  assign n4680 = n4678 ^ n3320 ;
  assign n4681 = ~n4679 & n4680 ;
  assign n4682 = n4681 ^ n3387 ;
  assign n4683 = n4632 & n4682 ;
  assign n4685 = n4684 ^ n4683 ;
  assign n4686 = n4629 & n4685 ;
  assign n4687 = n4686 ^ n3396 ;
  assign n4688 = ~n4626 & ~n4687 ;
  assign n4689 = n4688 ^ n2707 ;
  assign n4690 = n4689 ^ n4622 ;
  assign n4691 = n4623 & n4690 ;
  assign n4692 = n4691 ^ n2530 ;
  assign n4693 = n4462 ^ n2511 ;
  assign n4694 = ~n4583 & ~n4693 ;
  assign n4695 = n4694 ^ n4398 ;
  assign n4696 = n4695 ^ n2366 ;
  assign n4697 = n4692 & n4696 ;
  assign n4698 = n4697 ^ n2399 ;
  assign n4699 = n4619 & n4698 ;
  assign n4700 = n4699 ^ n2204 ;
  assign n4701 = n4616 & n4700 ;
  assign n4702 = n4701 ^ n2008 ;
  assign n4612 = n4475 & ~n4583 ;
  assign n4613 = n4612 ^ n4393 ;
  assign n4703 = n4702 ^ n4613 ;
  assign n4704 = n4702 ^ n1739 ;
  assign n4705 = ~n4703 & ~n4704 ;
  assign n4706 = n4705 ^ n1763 ;
  assign n4707 = n4611 & n4706 ;
  assign n4709 = n4708 ^ n4707 ;
  assign n4710 = ~n4479 & ~n4583 ;
  assign n4711 = n4710 ^ n4481 ;
  assign n4712 = n4711 ^ n1427 ;
  assign n4713 = ~n4709 & ~n4712 ;
  assign n4714 = n4713 ^ n1450 ;
  assign n4715 = ~n4485 & ~n4583 ;
  assign n4716 = n4715 ^ n4487 ;
  assign n4717 = n4716 ^ n1290 ;
  assign n4718 = n4714 & n4717 ;
  assign n4719 = n4718 ^ n4716 ;
  assign n4722 = n4721 ^ n4719 ;
  assign n4723 = n4721 ^ n1136 ;
  assign n4724 = ~n4722 & n4723 ;
  assign n4725 = n4724 ^ n1143 ;
  assign n4726 = n4496 & ~n4583 ;
  assign n4727 = n4726 ^ n4498 ;
  assign n4730 = n4727 ^ n1034 ;
  assign n4731 = ~n4725 & n4730 ;
  assign n4728 = n4727 ^ n892 ;
  assign n4732 = n4731 ^ n4728 ;
  assign n4733 = ~n4608 & n4732 ;
  assign n4734 = n4733 ^ n927 ;
  assign n4735 = n4503 & ~n4583 ;
  assign n4736 = n4735 ^ n4505 ;
  assign n4737 = n4736 ^ n696 ;
  assign n4738 = n4737 ^ n696 ;
  assign n4739 = n4738 ^ n786 ;
  assign n4740 = ~n4734 & n4739 ;
  assign n4741 = n4740 ^ n4737 ;
  assign n4742 = n4510 & ~n4583 ;
  assign n4743 = n4742 ^ n4512 ;
  assign n4744 = n4743 ^ n609 ;
  assign n4745 = n4744 ^ n835 ;
  assign n4746 = ~n4741 & ~n4745 ;
  assign n4747 = n4746 ^ n4744 ;
  assign n4748 = n4605 & n4747 ;
  assign n4749 = n4748 ^ n834 ;
  assign n4750 = n4522 & ~n4583 ;
  assign n4751 = n4750 ^ n4383 ;
  assign n4752 = n4751 ^ n534 ;
  assign n4753 = ~n4749 & ~n4752 ;
  assign n4754 = n4753 ^ n750 ;
  assign n4755 = ~n4602 & n4754 ;
  assign n4756 = n4755 ^ n4601 ;
  assign n4759 = n4758 ^ n4756 ;
  assign n4760 = n4758 ^ n401 ;
  assign n4761 = n4759 & ~n4760 ;
  assign n4762 = n4761 ^ n462 ;
  assign n4763 = ~n4599 & n4762 ;
  assign n4764 = n4763 ^ n349 ;
  assign n4765 = ~n4595 & ~n4764 ;
  assign n4766 = n4765 ^ n307 ;
  assign n4767 = n4592 & n4766 ;
  assign n4768 = n4767 ^ n4591 ;
  assign n4769 = n4768 ^ n188 ;
  assign n4801 = n4579 ^ n4576 ;
  assign n4802 = n4579 ^ n183 ;
  assign n4805 = n4564 & n4802 ;
  assign n4806 = n4805 ^ n183 ;
  assign n4807 = n4801 & n4806 ;
  assign n4584 = n4547 & ~n4583 ;
  assign n4585 = n4584 ^ n4570 ;
  assign n4586 = n4585 ^ n138 ;
  assign n4587 = n4545 & ~n4583 ;
  assign n4588 = n4587 ^ n4365 ;
  assign n4589 = n4588 ^ n157 ;
  assign n4770 = n4370 ^ n307 ;
  assign n4771 = n4770 ^ n4536 ;
  assign n4772 = n4771 ^ n307 ;
  assign n4775 = ~n4372 & ~n4772 ;
  assign n4776 = n4775 ^ n307 ;
  assign n4777 = ~n4583 & ~n4776 ;
  assign n4778 = n4777 ^ n4367 ;
  assign n4779 = n4778 ^ n4768 ;
  assign n4780 = n4769 & ~n4779 ;
  assign n4781 = n4780 ^ n203 ;
  assign n4782 = n4589 & ~n4781 ;
  assign n4783 = n4782 ^ n4588 ;
  assign n4784 = n4783 ^ n4585 ;
  assign n4785 = n4586 & ~n4784 ;
  assign n4786 = n4785 ^ n138 ;
  assign n4788 = n4573 ^ n138 ;
  assign n4789 = n4788 ^ n4566 ;
  assign n4790 = ~n4786 & ~n4789 ;
  assign n4791 = n4579 ^ n4573 ;
  assign n4792 = n4791 ^ n4579 ;
  assign n4795 = ~n4788 & ~n4792 ;
  assign n4796 = n4795 ^ n4579 ;
  assign n4797 = n4790 & n4796 ;
  assign n4798 = n4797 ^ n4788 ;
  assign n4799 = ~n4583 & n4798 ;
  assign n4787 = n4786 ^ n4566 ;
  assign n4800 = n4799 ^ n4787 ;
  assign n4808 = n4786 ^ n183 ;
  assign n4809 = n4808 ^ n4807 ;
  assign n4810 = n4800 & ~n4809 ;
  assign n4811 = n4810 ^ n4786 ;
  assign n4812 = ~n4807 & ~n4811 ;
  assign n4998 = n4769 & ~n4812 ;
  assign n4999 = n4998 ^ n4778 ;
  assign n5000 = n4999 ^ n157 ;
  assign n5001 = ~n4766 & ~n4812 ;
  assign n5002 = n5001 ^ n4591 ;
  assign n5003 = n5002 ^ n188 ;
  assign n5046 = ~n4764 & ~n4812 ;
  assign n5047 = n5046 ^ n4594 ;
  assign n5004 = n4762 & ~n4812 ;
  assign n5005 = n5004 ^ n4598 ;
  assign n5006 = n5005 ^ n291 ;
  assign n5036 = n4756 ^ n401 ;
  assign n5037 = ~n4812 & n5036 ;
  assign n5038 = n5037 ^ n4758 ;
  assign n5007 = ~n4754 & ~n4812 ;
  assign n5008 = n5007 ^ n4601 ;
  assign n5009 = n5008 ^ n401 ;
  assign n5010 = n4747 & ~n4812 ;
  assign n5011 = n5010 ^ n4604 ;
  assign n5012 = n5011 ^ n534 ;
  assign n5013 = n4741 & ~n4812 ;
  assign n5014 = n5013 ^ n4743 ;
  assign n5024 = n5014 ^ n534 ;
  assign n5015 = n5014 ^ n609 ;
  assign n4813 = n4732 & ~n4812 ;
  assign n4814 = n4813 ^ n4607 ;
  assign n4815 = n4814 ^ n786 ;
  assign n4816 = ~n4714 & ~n4812 ;
  assign n4817 = n4816 ^ n4716 ;
  assign n4818 = n4817 ^ n1136 ;
  assign n4933 = ~n4709 & ~n4812 ;
  assign n4934 = n4933 ^ n4711 ;
  assign n4937 = n4934 ^ n1136 ;
  assign n4819 = ~n4706 & ~n4812 ;
  assign n4820 = n4819 ^ n4610 ;
  assign n4821 = n4820 ^ n1427 ;
  assign n4924 = ~n4704 & ~n4812 ;
  assign n4925 = n4924 ^ n4613 ;
  assign n4929 = n4925 ^ n1427 ;
  assign n4822 = n4698 & ~n4812 ;
  assign n4823 = n4822 ^ n4618 ;
  assign n4824 = n4823 ^ n2008 ;
  assign n4825 = n4692 & ~n4812 ;
  assign n4826 = n4825 ^ n4695 ;
  assign n4827 = n4826 ^ n2175 ;
  assign n4828 = ~n4687 & ~n4812 ;
  assign n4829 = n4828 ^ n4625 ;
  assign n4830 = n4829 ^ n2511 ;
  assign n4900 = n4685 & ~n4812 ;
  assign n4901 = n4900 ^ n4628 ;
  assign n4831 = ~n4682 & ~n4812 ;
  assign n4832 = n4831 ^ n4631 ;
  assign n4833 = n4832 ^ n2894 ;
  assign n4837 = ~n4669 & ~n4812 ;
  assign n4838 = n4837 ^ n4635 ;
  assign n4839 = n4838 ^ n3538 ;
  assign n4875 = n4652 & ~n4812 ;
  assign n4876 = n4875 ^ n4656 ;
  assign n4841 = n4638 ^ n4583 ;
  assign n4851 = n4812 & ~n4841 ;
  assign n4852 = n4851 ^ n4639 ;
  assign n4853 = n4852 ^ n4356 ;
  assign n4856 = n4812 ^ x59 ;
  assign n4855 = ~x56 & ~x57 ;
  assign n4857 = n4856 ^ n4855 ;
  assign n4858 = n4855 ^ n4583 ;
  assign n4859 = ~n4857 & ~n4858 ;
  assign n4867 = n4859 ^ n4645 ;
  assign n4854 = n4812 ^ n4583 ;
  assign n4860 = n4859 ^ n4854 ;
  assign n4861 = n4860 ^ n4859 ;
  assign n4862 = n4859 ^ n4856 ;
  assign n4863 = n4862 ^ n4859 ;
  assign n4864 = n4861 & ~n4863 ;
  assign n4865 = n4864 ^ n4859 ;
  assign n4866 = x58 & n4865 ;
  assign n4868 = n4867 ^ n4866 ;
  assign n4869 = n4853 & ~n4868 ;
  assign n4870 = n4869 ^ n4852 ;
  assign n4844 = n4645 ^ x60 ;
  assign n4845 = n4844 ^ n4645 ;
  assign n4846 = ~n4841 & ~n4845 ;
  assign n4847 = n4846 ^ n4645 ;
  assign n4848 = ~n4812 & n4847 ;
  assign n4849 = n4848 ^ x61 ;
  assign n4840 = ~x60 & ~n4583 ;
  assign n4850 = n4849 ^ n4840 ;
  assign n4871 = n4870 ^ n4850 ;
  assign n4872 = n4870 ^ n4153 ;
  assign n4873 = ~n4871 & n4872 ;
  assign n4874 = n4873 ^ n4153 ;
  assign n4877 = n4876 ^ n4874 ;
  assign n4878 = n4876 ^ n3908 ;
  assign n4879 = ~n4877 & n4878 ;
  assign n4880 = n4879 ^ n3961 ;
  assign n4881 = n4659 ^ n3908 ;
  assign n4882 = ~n4812 & n4881 ;
  assign n4883 = n4882 ^ n4665 ;
  assign n4884 = n4883 ^ n3722 ;
  assign n4885 = ~n4880 & n4884 ;
  assign n4886 = n4885 ^ n3795 ;
  assign n4887 = n4839 & n4886 ;
  assign n4888 = n4887 ^ n3596 ;
  assign n4889 = n4671 & ~n4812 ;
  assign n4890 = n4889 ^ n4673 ;
  assign n4891 = n4890 ^ n3320 ;
  assign n4892 = n4888 & n4891 ;
  assign n4893 = n4892 ^ n3320 ;
  assign n4834 = n4676 ^ n3320 ;
  assign n4835 = ~n4812 & n4834 ;
  assign n4836 = n4835 ^ n4678 ;
  assign n4894 = n4893 ^ n4836 ;
  assign n4895 = n4836 ^ n3093 ;
  assign n4896 = ~n4894 & ~n4895 ;
  assign n4897 = n4896 ^ n3363 ;
  assign n4898 = n4833 & n4897 ;
  assign n4899 = n4898 ^ n2894 ;
  assign n4902 = n4901 ^ n4899 ;
  assign n4903 = n4901 ^ n2707 ;
  assign n4904 = ~n4902 & ~n4903 ;
  assign n4905 = n4904 ^ n2707 ;
  assign n4906 = n4905 ^ n4829 ;
  assign n4907 = n4830 & n4906 ;
  assign n4908 = n4907 ^ n2530 ;
  assign n4909 = n4689 ^ n2511 ;
  assign n4910 = ~n4812 & ~n4909 ;
  assign n4911 = n4910 ^ n4622 ;
  assign n4912 = n4911 ^ n2366 ;
  assign n4913 = n4908 & n4912 ;
  assign n4914 = n4913 ^ n2399 ;
  assign n4915 = n4827 & n4914 ;
  assign n4916 = n4915 ^ n2204 ;
  assign n4917 = n4824 & n4916 ;
  assign n4918 = n4917 ^ n2064 ;
  assign n4919 = n4700 & ~n4812 ;
  assign n4920 = n4919 ^ n4615 ;
  assign n4921 = n4920 ^ n1739 ;
  assign n4922 = ~n4918 & ~n4921 ;
  assign n4923 = n4922 ^ n1739 ;
  assign n4926 = n4925 ^ n4923 ;
  assign n4927 = n4923 ^ n1572 ;
  assign n4928 = ~n4926 & n4927 ;
  assign n4930 = n4929 ^ n4928 ;
  assign n4931 = ~n4821 & ~n4930 ;
  assign n4932 = n4931 ^ n1450 ;
  assign n4935 = n4934 ^ n1290 ;
  assign n4936 = n4932 & n4935 ;
  assign n4938 = n4937 ^ n4936 ;
  assign n4939 = n4818 & n4938 ;
  assign n4940 = n4939 ^ n1143 ;
  assign n4941 = n4719 ^ n1136 ;
  assign n4942 = ~n4812 & n4941 ;
  assign n4943 = n4942 ^ n4721 ;
  assign n4946 = n4943 ^ n1034 ;
  assign n4947 = ~n4940 & n4946 ;
  assign n4944 = n4943 ^ n892 ;
  assign n4948 = n4947 ^ n4944 ;
  assign n4949 = n4725 & ~n4812 ;
  assign n4950 = n4949 ^ n4727 ;
  assign n4951 = n4950 ^ n786 ;
  assign n4952 = n4951 ^ n927 ;
  assign n4953 = ~n4948 & n4952 ;
  assign n4954 = n4953 ^ n4951 ;
  assign n4955 = ~n4815 & n4954 ;
  assign n4956 = n4955 ^ n842 ;
  assign n5016 = n4734 & ~n4812 ;
  assign n5017 = n5016 ^ n4736 ;
  assign n5020 = n5017 ^ n696 ;
  assign n5021 = ~n4956 & n5020 ;
  assign n5018 = n5017 ^ n609 ;
  assign n5022 = n5021 ^ n5018 ;
  assign n5023 = n5015 & n5022 ;
  assign n5025 = n5024 ^ n5023 ;
  assign n5026 = ~n5012 & ~n5025 ;
  assign n5027 = n5026 ^ n750 ;
  assign n5028 = ~n4749 & ~n4812 ;
  assign n5029 = n5028 ^ n4751 ;
  assign n5030 = n5029 ^ n457 ;
  assign n5031 = n5027 & n5030 ;
  assign n5032 = n5031 ^ n5029 ;
  assign n5033 = n5032 ^ n5008 ;
  assign n5034 = n5009 & n5033 ;
  assign n5035 = n5034 ^ n401 ;
  assign n5039 = n5038 ^ n5035 ;
  assign n5040 = n5038 ^ n341 ;
  assign n5041 = n5039 & ~n5040 ;
  assign n5042 = n5041 ^ n349 ;
  assign n5043 = n5006 & ~n5042 ;
  assign n5044 = n5043 ^ n291 ;
  assign n5045 = n5044 ^ n5002 ;
  assign n5048 = n5047 ^ n5045 ;
  assign n5049 = n5048 ^ n245 ;
  assign n5050 = n5049 ^ n5045 ;
  assign n5051 = n5045 ^ n5044 ;
  assign n5052 = n5051 ^ n5047 ;
  assign n5053 = n5052 ^ n5045 ;
  assign n5054 = ~n5050 & ~n5053 ;
  assign n5055 = n5054 ^ n5045 ;
  assign n5056 = n5003 & n5055 ;
  assign n5057 = n5056 ^ n203 ;
  assign n5058 = n5000 & ~n5057 ;
  assign n5059 = n5058 ^ n4999 ;
  assign n5060 = n5059 ^ n138 ;
  assign n5061 = n4781 & ~n4812 ;
  assign n5062 = n5061 ^ n4588 ;
  assign n5063 = n5062 ^ n5059 ;
  assign n5064 = n5060 & ~n5063 ;
  assign n5065 = n5064 ^ n138 ;
  assign n5239 = n183 & n5065 ;
  assign n4957 = ~n4585 & n4812 ;
  assign n4985 = n4812 ^ n183 ;
  assign n4964 = n138 & ~n4812 ;
  assign n4962 = n4812 ^ n1003 ;
  assign n4963 = n4783 & ~n4962 ;
  assign n4965 = n4964 ^ n4963 ;
  assign n4966 = ~n4784 & n4965 ;
  assign n4967 = n4966 ^ n4964 ;
  assign n4968 = n4967 ^ n4812 ;
  assign n4986 = n4985 ^ n4968 ;
  assign n4972 = n4971 ^ n4783 ;
  assign n4973 = ~n4784 & ~n4972 ;
  assign n4974 = n4973 ^ n4970 ;
  assign n4975 = n4974 ^ n1355 ;
  assign n4980 = ~x127 & n4973 ;
  assign n4981 = ~n4975 & n4980 ;
  assign n4982 = n4981 ^ n4975 ;
  assign n4983 = n4982 ^ n1355 ;
  assign n4984 = ~n4812 & n4983 ;
  assign n4987 = n4986 ^ n4984 ;
  assign n4988 = n4987 ^ n4968 ;
  assign n4989 = n4957 & n4988 ;
  assign n4990 = n4989 ^ n4987 ;
  assign n4992 = n4789 ^ n4583 ;
  assign n4993 = n4992 ^ n4789 ;
  assign n4994 = n4788 & n4993 ;
  assign n4995 = n4994 ^ n4789 ;
  assign n4996 = n4990 & ~n4995 ;
  assign n4997 = n4996 ^ n4984 ;
  assign n5240 = ~n4997 & ~n5062 ;
  assign n5241 = ~n1355 & ~n5059 ;
  assign n5242 = n5240 & n5241 ;
  assign n5066 = n4783 ^ n138 ;
  assign n5067 = ~n4812 & n5066 ;
  assign n5068 = n5067 ^ n4585 ;
  assign n5243 = n5242 ^ n5068 ;
  assign n5069 = ~n183 & ~n5068 ;
  assign n5070 = n5069 ^ n5068 ;
  assign n5246 = n5243 ^ n5070 ;
  assign n5247 = n5246 ^ n5243 ;
  assign n5248 = ~n4997 & ~n5247 ;
  assign n5249 = n5248 ^ n5243 ;
  assign n5250 = n5239 & n5249 ;
  assign n5251 = n5250 ^ n5243 ;
  assign n5253 = n5059 & ~n5240 ;
  assign n5252 = n4997 ^ n138 ;
  assign n5254 = n5253 ^ n5252 ;
  assign n5255 = n5062 ^ n5060 ;
  assign n5256 = n5255 ^ n4997 ;
  assign n5257 = n5254 & ~n5256 ;
  assign n5258 = n5257 ^ n4997 ;
  assign n5259 = n5069 & ~n5258 ;
  assign n5260 = ~n5251 & n5259 ;
  assign n5261 = n5260 ^ n5251 ;
  assign n5071 = n5065 & n5070 ;
  assign n5072 = n4997 & n5071 ;
  assign n5073 = n5072 ^ n4997 ;
  assign n5308 = n5060 & ~n5073 ;
  assign n5309 = n5308 ^ n5062 ;
  assign n5302 = n5057 & ~n5073 ;
  assign n5303 = n5302 ^ n4999 ;
  assign n5262 = n5044 ^ n188 ;
  assign n5263 = n5262 ^ n246 ;
  assign n5264 = n5047 ^ n188 ;
  assign n5265 = n5264 ^ n5262 ;
  assign n5266 = ~n5263 & ~n5265 ;
  assign n5267 = n5266 ^ n5262 ;
  assign n5268 = ~n5073 & ~n5267 ;
  assign n5269 = n5268 ^ n5002 ;
  assign n5270 = n5269 ^ n157 ;
  assign n5274 = ~n5042 & ~n5073 ;
  assign n5275 = n5274 ^ n5005 ;
  assign n5276 = n5275 ^ n245 ;
  assign n5277 = n5032 ^ n401 ;
  assign n5278 = ~n5073 & ~n5277 ;
  assign n5279 = n5278 ^ n5008 ;
  assign n5280 = n5279 ^ n341 ;
  assign n5076 = n4954 & ~n5073 ;
  assign n5077 = n5076 ^ n4814 ;
  assign n5078 = n5077 ^ n696 ;
  assign n5079 = ~n4932 & ~n5073 ;
  assign n5080 = n5079 ^ n4934 ;
  assign n5081 = n5080 ^ n1136 ;
  assign n5195 = ~n4930 & ~n5073 ;
  assign n5196 = n5195 ^ n4820 ;
  assign n5199 = n5196 ^ n1136 ;
  assign n5184 = ~n4918 & ~n5073 ;
  assign n5185 = n5184 ^ n4920 ;
  assign n5188 = n5185 ^ n1427 ;
  assign n5082 = n4914 & ~n5073 ;
  assign n5083 = n5082 ^ n4826 ;
  assign n5084 = n5083 ^ n2008 ;
  assign n5085 = n4908 & ~n5073 ;
  assign n5086 = n5085 ^ n4911 ;
  assign n5087 = n5086 ^ n2175 ;
  assign n5088 = n4899 ^ n2707 ;
  assign n5089 = ~n5073 & ~n5088 ;
  assign n5090 = n5089 ^ n4901 ;
  assign n5091 = n5090 ^ n2511 ;
  assign n5092 = n4897 & ~n5073 ;
  assign n5093 = n5092 ^ n4832 ;
  assign n5094 = n5093 ^ n2707 ;
  assign n5095 = n4893 ^ n3093 ;
  assign n5096 = ~n5073 & ~n5095 ;
  assign n5097 = n5096 ^ n4836 ;
  assign n5098 = n5097 ^ n2894 ;
  assign n5099 = ~n4880 & ~n5073 ;
  assign n5100 = n5099 ^ n4883 ;
  assign n5101 = n5100 ^ n3538 ;
  assign n5102 = n4874 ^ n3908 ;
  assign n5103 = ~n5073 & n5102 ;
  assign n5104 = n5103 ^ n4876 ;
  assign n5105 = n5104 ^ n3722 ;
  assign n5142 = n4872 & ~n5073 ;
  assign n5143 = n5142 ^ n4850 ;
  assign n5106 = n4868 & ~n5073 ;
  assign n5107 = n5106 ^ n4852 ;
  assign n5108 = n5107 ^ n4153 ;
  assign n5125 = n4855 ^ n4812 ;
  assign n5126 = ~n5073 & ~n5125 ;
  assign n5127 = n5126 ^ n4812 ;
  assign n5133 = x58 & ~n5127 ;
  assign n5132 = ~n4858 & ~n5073 ;
  assign n5134 = n5133 ^ n5132 ;
  assign n5135 = n5134 ^ n4856 ;
  assign n5138 = n5135 ^ n4153 ;
  assign n5109 = n4812 ^ x57 ;
  assign n5110 = n5109 ^ n5073 ;
  assign n5112 = ~x54 & ~x55 ;
  assign n5111 = n4812 ^ x56 ;
  assign n5113 = n5112 ^ n5111 ;
  assign n5114 = ~n5110 & ~n5113 ;
  assign n5123 = n5114 ^ n4854 ;
  assign n5115 = n5073 ^ n4812 ;
  assign n5116 = n5115 ^ n5114 ;
  assign n5117 = n5116 ^ n5114 ;
  assign n5120 = n5109 & n5117 ;
  assign n5121 = n5120 ^ n5114 ;
  assign n5122 = x56 & n5121 ;
  assign n5124 = n5123 ^ n5122 ;
  assign n5128 = n5127 ^ x58 ;
  assign n5129 = n5128 ^ n4583 ;
  assign n5130 = n5124 & ~n5129 ;
  assign n5131 = n5130 ^ n4645 ;
  assign n5136 = n5135 ^ n4356 ;
  assign n5137 = ~n5131 & ~n5136 ;
  assign n5139 = n5138 ^ n5137 ;
  assign n5140 = n5108 & ~n5139 ;
  assign n5141 = n5140 ^ n4153 ;
  assign n5144 = n5143 ^ n5141 ;
  assign n5145 = n5143 ^ n3908 ;
  assign n5146 = ~n5144 & n5145 ;
  assign n5147 = n5146 ^ n3961 ;
  assign n5148 = ~n5105 & ~n5147 ;
  assign n5149 = n5148 ^ n3795 ;
  assign n5150 = n5101 & n5149 ;
  assign n5151 = n5150 ^ n3596 ;
  assign n5152 = n4886 & ~n5073 ;
  assign n5153 = n5152 ^ n4838 ;
  assign n5154 = n5153 ^ n3320 ;
  assign n5155 = n5151 & n5154 ;
  assign n5156 = n5155 ^ n3387 ;
  assign n5157 = n4888 & ~n5073 ;
  assign n5158 = n5157 ^ n4890 ;
  assign n5159 = n5158 ^ n3093 ;
  assign n5160 = ~n5156 & ~n5159 ;
  assign n5161 = n5160 ^ n3363 ;
  assign n5162 = ~n5098 & n5161 ;
  assign n5163 = n5162 ^ n3396 ;
  assign n5164 = ~n5094 & ~n5163 ;
  assign n5165 = n5164 ^ n2707 ;
  assign n5166 = n5165 ^ n5090 ;
  assign n5167 = n5091 & n5166 ;
  assign n5168 = n5167 ^ n2530 ;
  assign n5169 = n4905 ^ n2511 ;
  assign n5170 = ~n5073 & ~n5169 ;
  assign n5171 = n5170 ^ n4829 ;
  assign n5172 = n5171 ^ n2366 ;
  assign n5173 = n5168 & n5172 ;
  assign n5174 = n5173 ^ n2399 ;
  assign n5175 = n5087 & n5174 ;
  assign n5176 = n5175 ^ n2204 ;
  assign n5177 = n5084 & n5176 ;
  assign n5178 = n5177 ^ n2064 ;
  assign n5179 = n4916 & ~n5073 ;
  assign n5180 = n5179 ^ n4823 ;
  assign n5181 = n5180 ^ n1739 ;
  assign n5182 = ~n5178 & ~n5181 ;
  assign n5183 = n5182 ^ n1763 ;
  assign n5186 = n5185 ^ n1572 ;
  assign n5187 = n5183 & n5186 ;
  assign n5189 = n5188 ^ n5187 ;
  assign n5190 = ~n4927 & ~n5073 ;
  assign n5191 = n5190 ^ n4925 ;
  assign n5192 = n5191 ^ n1427 ;
  assign n5193 = ~n5189 & ~n5192 ;
  assign n5194 = n5193 ^ n1450 ;
  assign n5197 = n5196 ^ n1290 ;
  assign n5198 = n5194 & n5197 ;
  assign n5200 = n5199 ^ n5198 ;
  assign n5201 = n5081 & n5200 ;
  assign n5202 = n5201 ^ n1143 ;
  assign n5203 = n4938 & ~n5073 ;
  assign n5204 = n5203 ^ n4817 ;
  assign n5207 = n5204 ^ n1034 ;
  assign n5208 = ~n5202 & n5207 ;
  assign n5205 = n5204 ^ n892 ;
  assign n5209 = n5208 ^ n5205 ;
  assign n5210 = n4940 & ~n5073 ;
  assign n5211 = n5210 ^ n4943 ;
  assign n5212 = n5211 ^ n786 ;
  assign n5213 = n5212 ^ n927 ;
  assign n5214 = ~n5209 & n5213 ;
  assign n5215 = n5214 ^ n5212 ;
  assign n5216 = n4948 & ~n5073 ;
  assign n5217 = n5216 ^ n4950 ;
  assign n5218 = n5217 ^ n696 ;
  assign n5219 = n5218 ^ n842 ;
  assign n5220 = ~n5215 & n5219 ;
  assign n5221 = n5220 ^ n5218 ;
  assign n5222 = ~n5078 & ~n5221 ;
  assign n5223 = n5222 ^ n5077 ;
  assign n5074 = n4956 & ~n5073 ;
  assign n5075 = n5074 ^ n5017 ;
  assign n5224 = n5223 ^ n5075 ;
  assign n5225 = n5075 ^ n609 ;
  assign n5226 = n5224 & ~n5225 ;
  assign n5227 = n5226 ^ n834 ;
  assign n5228 = ~n5022 & ~n5073 ;
  assign n5229 = n5228 ^ n5014 ;
  assign n5230 = n5229 ^ n534 ;
  assign n5231 = ~n5227 & ~n5230 ;
  assign n5232 = n5231 ^ n750 ;
  assign n5233 = ~n5025 & ~n5073 ;
  assign n5234 = n5233 ^ n5011 ;
  assign n5235 = n5234 ^ n457 ;
  assign n5236 = n5232 & n5235 ;
  assign n5237 = n5236 ^ n5234 ;
  assign n5238 = n5237 ^ n401 ;
  assign n5281 = ~n5027 & ~n5073 ;
  assign n5282 = n5281 ^ n5029 ;
  assign n5283 = n5282 ^ n5237 ;
  assign n5284 = ~n5238 & ~n5283 ;
  assign n5285 = n5284 ^ n462 ;
  assign n5286 = n5280 & n5285 ;
  assign n5287 = n5286 ^ n349 ;
  assign n5288 = n5035 ^ n341 ;
  assign n5289 = ~n5073 & n5288 ;
  assign n5290 = n5289 ^ n5038 ;
  assign n5291 = n5290 ^ n291 ;
  assign n5292 = ~n5287 & n5291 ;
  assign n5293 = n5292 ^ n307 ;
  assign n5294 = ~n5276 & n5293 ;
  assign n5295 = n5294 ^ n5275 ;
  assign n5271 = n5044 ^ n245 ;
  assign n5272 = ~n5073 & ~n5271 ;
  assign n5273 = n5272 ^ n5047 ;
  assign n5296 = n5295 ^ n5273 ;
  assign n5297 = n5295 ^ n188 ;
  assign n5298 = n5296 & ~n5297 ;
  assign n5299 = n5298 ^ n203 ;
  assign n5300 = n5270 & ~n5299 ;
  assign n5301 = n5300 ^ n5269 ;
  assign n5304 = n5303 ^ n5301 ;
  assign n5305 = n5303 ^ n138 ;
  assign n5306 = ~n5304 & n5305 ;
  assign n5307 = n5306 ^ n138 ;
  assign n5312 = n183 & n5307 ;
  assign n5315 = ~n5309 & n5312 ;
  assign n5316 = n5315 ^ n5307 ;
  assign n5317 = ~n5261 & ~n5316 ;
  assign n5506 = n5301 ^ n138 ;
  assign n5507 = ~n5317 & n5506 ;
  assign n5508 = n5507 ^ n5303 ;
  assign n5532 = n5299 & ~n5317 ;
  assign n5533 = n5532 ^ n5269 ;
  assign n5770 = ~n5508 & ~n5533 ;
  assign n5793 = n5770 ^ n183 ;
  assign n5771 = ~n183 & n5770 ;
  assign n5794 = n5793 ^ n5771 ;
  assign n5534 = ~n5297 & ~n5317 ;
  assign n5535 = n5534 ^ n5273 ;
  assign n5536 = n5535 ^ n157 ;
  assign n5547 = ~n5293 & ~n5317 ;
  assign n5548 = n5547 ^ n5275 ;
  assign n5318 = ~n5238 & ~n5317 ;
  assign n5319 = n5318 ^ n5282 ;
  assign n5320 = n5319 ^ n341 ;
  assign n5498 = ~n5232 & ~n5317 ;
  assign n5499 = n5498 ^ n5234 ;
  assign n5321 = ~n5227 & ~n5317 ;
  assign n5322 = n5321 ^ n5229 ;
  assign n5323 = n5322 ^ n457 ;
  assign n5324 = n5223 ^ n609 ;
  assign n5325 = ~n5317 & n5324 ;
  assign n5326 = n5325 ^ n5075 ;
  assign n5327 = n5326 ^ n534 ;
  assign n5330 = n5215 & ~n5317 ;
  assign n5331 = n5330 ^ n5217 ;
  assign n5332 = n5331 ^ n696 ;
  assign n5333 = ~n5194 & ~n5317 ;
  assign n5334 = n5333 ^ n5196 ;
  assign n5335 = n5334 ^ n1136 ;
  assign n5461 = ~n5189 & ~n5317 ;
  assign n5462 = n5461 ^ n5191 ;
  assign n5465 = n5462 ^ n1136 ;
  assign n5450 = ~n5178 & ~n5317 ;
  assign n5451 = n5450 ^ n5180 ;
  assign n5454 = n5451 ^ n1427 ;
  assign n5336 = n5176 & ~n5317 ;
  assign n5337 = n5336 ^ n5083 ;
  assign n5338 = n5337 ^ n1739 ;
  assign n5341 = n5168 & ~n5317 ;
  assign n5342 = n5341 ^ n5171 ;
  assign n5343 = n5342 ^ n2175 ;
  assign n5344 = n5165 ^ n2511 ;
  assign n5345 = ~n5317 & ~n5344 ;
  assign n5346 = n5345 ^ n5090 ;
  assign n5347 = n5346 ^ n2366 ;
  assign n5434 = ~n5163 & ~n5317 ;
  assign n5435 = n5434 ^ n5093 ;
  assign n5348 = n5161 & ~n5317 ;
  assign n5349 = n5348 ^ n5097 ;
  assign n5350 = n5349 ^ n2707 ;
  assign n5421 = n5151 & ~n5317 ;
  assign n5422 = n5421 ^ n5153 ;
  assign n5425 = n5422 ^ n2894 ;
  assign n5351 = ~n5147 & ~n5317 ;
  assign n5352 = n5351 ^ n5104 ;
  assign n5353 = n5352 ^ n3538 ;
  assign n5354 = ~n5139 & ~n5317 ;
  assign n5355 = n5354 ^ n5107 ;
  assign n5356 = n5355 ^ n3908 ;
  assign n5357 = n5131 & ~n5317 ;
  assign n5358 = n5357 ^ n5135 ;
  assign n5359 = n5358 ^ n4153 ;
  assign n5397 = n5124 & ~n5317 ;
  assign n5398 = n5397 ^ n5128 ;
  assign n5401 = n5398 ^ n4153 ;
  assign n5376 = n5112 ^ n5073 ;
  assign n5384 = n5115 ^ x56 ;
  assign n5385 = n5384 ^ n5115 ;
  assign n5388 = ~n5376 & ~n5385 ;
  assign n5389 = n5388 ^ n5115 ;
  assign n5390 = ~n5317 & n5389 ;
  assign n5391 = n5390 ^ x57 ;
  assign n5383 = ~x56 & ~n5073 ;
  assign n5392 = n5391 ^ n5383 ;
  assign n5377 = ~n5317 & ~n5376 ;
  assign n5375 = n5073 ^ x56 ;
  assign n5378 = n5377 ^ n5375 ;
  assign n5361 = n5073 ^ x55 ;
  assign n5362 = n5361 ^ x54 ;
  assign n5365 = n5362 ^ n5361 ;
  assign n5367 = ~x52 & ~x53 ;
  assign n5360 = n5317 ^ n5073 ;
  assign n5363 = n5362 ^ n5360 ;
  assign n5368 = n5367 ^ n5363 ;
  assign n5369 = n5361 ^ n5317 ;
  assign n5370 = ~n5368 & ~n5369 ;
  assign n5366 = n5361 & n5363 ;
  assign n5371 = n5370 ^ n5366 ;
  assign n5372 = ~n5365 & n5371 ;
  assign n5373 = n5372 ^ n5366 ;
  assign n5374 = n5373 ^ n5073 ;
  assign n5379 = n5378 ^ n5374 ;
  assign n5380 = n5378 ^ n4812 ;
  assign n5381 = n5379 & ~n5380 ;
  assign n5382 = n5381 ^ n4812 ;
  assign n5393 = n5392 ^ n5382 ;
  assign n5394 = n5392 ^ n4583 ;
  assign n5395 = ~n5393 & n5394 ;
  assign n5396 = n5395 ^ n4645 ;
  assign n5399 = n5398 ^ n4356 ;
  assign n5400 = ~n5396 & ~n5399 ;
  assign n5402 = n5401 ^ n5400 ;
  assign n5403 = ~n5359 & ~n5402 ;
  assign n5404 = n5403 ^ n4153 ;
  assign n5405 = n5404 ^ n5355 ;
  assign n5406 = n5356 & ~n5405 ;
  assign n5407 = n5406 ^ n3961 ;
  assign n5408 = n5141 ^ n3908 ;
  assign n5409 = ~n5317 & n5408 ;
  assign n5410 = n5409 ^ n5143 ;
  assign n5411 = n5410 ^ n3722 ;
  assign n5412 = ~n5407 & ~n5411 ;
  assign n5413 = n5412 ^ n3795 ;
  assign n5414 = ~n5353 & n5413 ;
  assign n5415 = n5414 ^ n3596 ;
  assign n5416 = n5149 & ~n5317 ;
  assign n5417 = n5416 ^ n5100 ;
  assign n5418 = n5417 ^ n3320 ;
  assign n5419 = n5415 & n5418 ;
  assign n5420 = n5419 ^ n3387 ;
  assign n5423 = n5422 ^ n3093 ;
  assign n5424 = n5420 & ~n5423 ;
  assign n5426 = n5425 ^ n5424 ;
  assign n5427 = ~n5156 & ~n5317 ;
  assign n5428 = n5427 ^ n5158 ;
  assign n5429 = n5428 ^ n2894 ;
  assign n5430 = ~n5426 & ~n5429 ;
  assign n5431 = n5430 ^ n3396 ;
  assign n5432 = n5350 & ~n5431 ;
  assign n5433 = n5432 ^ n2707 ;
  assign n5436 = n5435 ^ n5433 ;
  assign n5437 = n5435 ^ n2511 ;
  assign n5438 = n5436 & n5437 ;
  assign n5439 = n5438 ^ n2530 ;
  assign n5440 = n5347 & n5439 ;
  assign n5441 = n5440 ^ n2399 ;
  assign n5442 = n5343 & n5441 ;
  assign n5443 = n5442 ^ n2175 ;
  assign n5339 = n5174 & ~n5317 ;
  assign n5340 = n5339 ^ n5086 ;
  assign n5444 = n5443 ^ n5340 ;
  assign n5445 = n5443 ^ n2008 ;
  assign n5446 = ~n5444 & n5445 ;
  assign n5447 = n5446 ^ n2064 ;
  assign n5448 = ~n5338 & ~n5447 ;
  assign n5449 = n5448 ^ n1763 ;
  assign n5452 = n5451 ^ n1572 ;
  assign n5453 = n5449 & n5452 ;
  assign n5455 = n5454 ^ n5453 ;
  assign n5456 = ~n5183 & ~n5317 ;
  assign n5457 = n5456 ^ n5185 ;
  assign n5458 = n5457 ^ n1427 ;
  assign n5459 = ~n5455 & ~n5458 ;
  assign n5460 = n5459 ^ n1450 ;
  assign n5463 = n5462 ^ n1290 ;
  assign n5464 = n5460 & n5463 ;
  assign n5466 = n5465 ^ n5464 ;
  assign n5467 = n5335 & n5466 ;
  assign n5468 = n5467 ^ n1143 ;
  assign n5469 = n5200 & ~n5317 ;
  assign n5470 = n5469 ^ n5080 ;
  assign n5473 = n5470 ^ n1034 ;
  assign n5474 = ~n5468 & n5473 ;
  assign n5471 = n5470 ^ n892 ;
  assign n5475 = n5474 ^ n5471 ;
  assign n5476 = n5202 & ~n5317 ;
  assign n5477 = n5476 ^ n5204 ;
  assign n5478 = n5477 ^ n786 ;
  assign n5479 = n5478 ^ n927 ;
  assign n5480 = ~n5475 & n5479 ;
  assign n5481 = n5480 ^ n5478 ;
  assign n5482 = n5209 & ~n5317 ;
  assign n5483 = n5482 ^ n5211 ;
  assign n5484 = n5483 ^ n696 ;
  assign n5485 = n5484 ^ n842 ;
  assign n5486 = ~n5481 & n5485 ;
  assign n5487 = n5486 ^ n5484 ;
  assign n5488 = n5332 & ~n5487 ;
  assign n5489 = n5488 ^ n5331 ;
  assign n5328 = n5221 & ~n5317 ;
  assign n5329 = n5328 ^ n5077 ;
  assign n5490 = n5489 ^ n5329 ;
  assign n5491 = n5329 ^ n609 ;
  assign n5492 = n5490 & n5491 ;
  assign n5493 = n5492 ^ n834 ;
  assign n5494 = n5327 & ~n5493 ;
  assign n5495 = n5494 ^ n750 ;
  assign n5496 = n5323 & n5495 ;
  assign n5497 = n5496 ^ n5322 ;
  assign n5500 = n5499 ^ n5497 ;
  assign n5501 = n5499 ^ n401 ;
  assign n5502 = ~n5500 & ~n5501 ;
  assign n5503 = n5502 ^ n462 ;
  assign n5504 = ~n5320 & n5503 ;
  assign n5505 = n5504 ^ n349 ;
  assign n5537 = n5285 & ~n5317 ;
  assign n5538 = n5537 ^ n5279 ;
  assign n5539 = n5538 ^ n291 ;
  assign n5540 = ~n5505 & ~n5539 ;
  assign n5541 = n5540 ^ n307 ;
  assign n5542 = ~n5287 & ~n5317 ;
  assign n5543 = n5542 ^ n5290 ;
  assign n5544 = n5543 ^ n245 ;
  assign n5545 = n5541 & ~n5544 ;
  assign n5546 = n5545 ^ n5543 ;
  assign n5549 = n5548 ^ n5546 ;
  assign n5550 = n5548 ^ n188 ;
  assign n5551 = ~n5549 & ~n5550 ;
  assign n5552 = n5551 ^ n203 ;
  assign n5553 = n5536 & ~n5552 ;
  assign n5554 = n5553 ^ n5535 ;
  assign n5555 = n5533 & n5554 ;
  assign n5556 = n5554 ^ n5533 ;
  assign n5557 = n5556 ^ n5555 ;
  assign n5558 = n138 & n5557 ;
  assign n5559 = ~n5555 & ~n5558 ;
  assign n5795 = n5770 ^ n5559 ;
  assign n5796 = ~n5794 & n5795 ;
  assign n5774 = n5558 ^ n138 ;
  assign n5797 = n5796 ^ n5774 ;
  assign n5787 = n1355 ^ n138 ;
  assign n5788 = n5770 ^ n138 ;
  assign n5789 = ~n5787 & ~n5788 ;
  assign n5524 = ~n1355 & n5261 ;
  assign n5525 = ~n5301 & ~n5303 ;
  assign n5526 = n5524 & n5525 ;
  assign n5527 = n5526 ^ n5312 ;
  assign n5510 = n5303 ^ n4971 ;
  assign n5511 = n5510 ^ n5261 ;
  assign n5512 = n5511 ^ n5301 ;
  assign n5513 = n5512 ^ n5304 ;
  assign n5514 = n5513 ^ n5512 ;
  assign n5515 = n5512 ^ n5506 ;
  assign n5516 = n5515 ^ n5512 ;
  assign n5517 = ~n5514 & ~n5516 ;
  assign n5518 = n5517 ^ n5512 ;
  assign n5519 = n5261 & ~n5518 ;
  assign n5528 = n5527 ^ n5519 ;
  assign n5520 = n5512 ^ n5261 ;
  assign n5521 = n5520 ^ n5519 ;
  assign n5522 = ~n183 & n5303 ;
  assign n5523 = n5521 & n5522 ;
  assign n5529 = n5528 ^ n5523 ;
  assign n5530 = ~n5309 & ~n5529 ;
  assign n5531 = n5530 ^ n5527 ;
  assign n5790 = ~n5531 & ~n5557 ;
  assign n5791 = n5790 ^ n138 ;
  assign n5792 = n5789 & n5791 ;
  assign n5798 = n5797 ^ n5792 ;
  assign n5777 = n138 & ~n5508 ;
  assign n5778 = n5555 & n5777 ;
  assign n5779 = n5778 ^ n5508 ;
  assign n5799 = n5798 ^ n5779 ;
  assign n5775 = n5774 ^ n5559 ;
  assign n5776 = n5775 ^ n183 ;
  assign n5769 = ~n5508 & ~n5531 ;
  assign n5780 = n5779 ^ n5769 ;
  assign n5781 = n5780 ^ n5779 ;
  assign n5782 = n5779 ^ n5775 ;
  assign n5783 = n5782 ^ n5779 ;
  assign n5784 = n5781 & ~n5783 ;
  assign n5785 = n5784 ^ n5779 ;
  assign n5786 = n5776 & n5785 ;
  assign n5800 = n5799 ^ n5786 ;
  assign n5772 = ~n138 & n5771 ;
  assign n5773 = n5769 & n5772 ;
  assign n5801 = n5800 ^ n5773 ;
  assign n5509 = n5508 ^ n183 ;
  assign n5560 = n5531 & ~n5559 ;
  assign n5561 = ~n5509 & n5560 ;
  assign n5562 = n5561 ^ n5531 ;
  assign n5802 = ~n5541 & ~n5562 ;
  assign n5803 = n5802 ^ n5543 ;
  assign n5804 = n5803 ^ n188 ;
  assign n5563 = ~n5505 & ~n5562 ;
  assign n5564 = n5563 ^ n5538 ;
  assign n5565 = n5564 ^ n245 ;
  assign n5566 = n5497 ^ n401 ;
  assign n5567 = ~n5562 & ~n5566 ;
  assign n5568 = n5567 ^ n5499 ;
  assign n5569 = n5568 ^ n341 ;
  assign n5574 = ~n5493 & ~n5562 ;
  assign n5575 = n5574 ^ n5326 ;
  assign n5576 = n5575 ^ n457 ;
  assign n5577 = n5489 ^ n609 ;
  assign n5578 = ~n5562 & ~n5577 ;
  assign n5579 = n5578 ^ n5329 ;
  assign n5580 = n5579 ^ n534 ;
  assign n5581 = n5487 & ~n5562 ;
  assign n5582 = n5581 ^ n5331 ;
  assign n5583 = n5582 ^ n609 ;
  assign n5716 = ~n5460 & ~n5562 ;
  assign n5717 = n5716 ^ n5462 ;
  assign n5584 = ~n5447 & ~n5562 ;
  assign n5585 = n5584 ^ n5337 ;
  assign n5704 = n5585 ^ n1427 ;
  assign n5586 = n5585 ^ n1572 ;
  assign n5589 = n5441 & ~n5562 ;
  assign n5590 = n5589 ^ n5342 ;
  assign n5591 = n5590 ^ n2008 ;
  assign n5592 = n5439 & ~n5562 ;
  assign n5593 = n5592 ^ n5346 ;
  assign n5594 = n5593 ^ n2175 ;
  assign n5595 = n5433 ^ n2511 ;
  assign n5596 = ~n5562 & ~n5595 ;
  assign n5597 = n5596 ^ n5435 ;
  assign n5598 = n5597 ^ n2366 ;
  assign n5687 = ~n5431 & ~n5562 ;
  assign n5688 = n5687 ^ n5349 ;
  assign n5599 = ~n5420 & ~n5562 ;
  assign n5600 = n5599 ^ n5422 ;
  assign n5601 = n5600 ^ n2894 ;
  assign n5674 = n5415 & ~n5562 ;
  assign n5675 = n5674 ^ n5417 ;
  assign n5678 = n5675 ^ n2894 ;
  assign n5602 = ~n5407 & ~n5562 ;
  assign n5603 = n5602 ^ n5410 ;
  assign n5604 = n5603 ^ n3538 ;
  assign n5660 = n5404 ^ n3908 ;
  assign n5661 = ~n5562 & n5660 ;
  assign n5662 = n5661 ^ n5355 ;
  assign n5605 = ~n5402 & ~n5562 ;
  assign n5606 = n5605 ^ n5358 ;
  assign n5607 = n5606 ^ n3908 ;
  assign n5608 = n5396 & ~n5562 ;
  assign n5609 = n5608 ^ n5398 ;
  assign n5610 = n5609 ^ n4153 ;
  assign n5648 = n5382 ^ n4583 ;
  assign n5649 = ~n5562 & n5648 ;
  assign n5650 = n5649 ^ n5392 ;
  assign n5653 = n5650 ^ n4153 ;
  assign n5611 = n5374 ^ n4812 ;
  assign n5612 = ~n5562 & n5611 ;
  assign n5613 = n5612 ^ n5378 ;
  assign n5614 = n5613 ^ n4583 ;
  assign n5615 = n5367 ^ n5317 ;
  assign n5627 = n5562 & ~n5615 ;
  assign n5626 = n5367 ^ x54 ;
  assign n5628 = n5627 ^ n5626 ;
  assign n5629 = n5628 ^ n5073 ;
  assign n5634 = ~x50 & ~x51 ;
  assign n5635 = ~x52 & n5634 ;
  assign n5633 = n5562 ^ x53 ;
  assign n5636 = n5635 ^ n5633 ;
  assign n5630 = ~x52 & ~n5562 ;
  assign n5631 = n5630 ^ x53 ;
  assign n5637 = n5631 ^ n5317 ;
  assign n5638 = n5636 & n5637 ;
  assign n5632 = n5631 ^ n5073 ;
  assign n5639 = n5638 ^ n5632 ;
  assign n5640 = n5629 & n5639 ;
  assign n5641 = n5640 ^ n5073 ;
  assign n5624 = ~x54 & ~n5317 ;
  assign n5618 = n5360 ^ x54 ;
  assign n5619 = n5618 ^ n5360 ;
  assign n5620 = ~n5615 & ~n5619 ;
  assign n5621 = n5620 ^ n5360 ;
  assign n5622 = ~n5562 & n5621 ;
  assign n5623 = n5622 ^ x55 ;
  assign n5625 = n5624 ^ n5623 ;
  assign n5642 = n5641 ^ n5625 ;
  assign n5643 = n5641 ^ n4812 ;
  assign n5644 = ~n5642 & n5643 ;
  assign n5645 = n5644 ^ n4854 ;
  assign n5646 = ~n5614 & n5645 ;
  assign n5647 = n5646 ^ n4645 ;
  assign n5651 = n5650 ^ n4356 ;
  assign n5652 = ~n5647 & n5651 ;
  assign n5654 = n5653 ^ n5652 ;
  assign n5655 = ~n5610 & n5654 ;
  assign n5656 = n5655 ^ n4153 ;
  assign n5657 = n5656 ^ n5606 ;
  assign n5658 = ~n5607 & n5657 ;
  assign n5659 = n5658 ^ n3908 ;
  assign n5663 = n5662 ^ n5659 ;
  assign n5664 = n5662 ^ n3722 ;
  assign n5665 = ~n5663 & ~n5664 ;
  assign n5666 = n5665 ^ n3795 ;
  assign n5667 = ~n5604 & n5666 ;
  assign n5668 = n5667 ^ n3596 ;
  assign n5669 = n5413 & ~n5562 ;
  assign n5670 = n5669 ^ n5352 ;
  assign n5671 = n5670 ^ n3320 ;
  assign n5672 = n5668 & ~n5671 ;
  assign n5673 = n5672 ^ n3387 ;
  assign n5676 = n5675 ^ n3093 ;
  assign n5677 = n5673 & ~n5676 ;
  assign n5679 = n5678 ^ n5677 ;
  assign n5680 = ~n5601 & ~n5679 ;
  assign n5681 = n5680 ^ n3396 ;
  assign n5682 = ~n5426 & ~n5562 ;
  assign n5683 = n5682 ^ n5428 ;
  assign n5684 = n5683 ^ n2707 ;
  assign n5685 = ~n5681 & n5684 ;
  assign n5686 = n5685 ^ n2707 ;
  assign n5689 = n5688 ^ n5686 ;
  assign n5690 = n5688 ^ n2511 ;
  assign n5691 = ~n5689 & ~n5690 ;
  assign n5692 = n5691 ^ n2530 ;
  assign n5693 = n5598 & n5692 ;
  assign n5694 = n5693 ^ n2399 ;
  assign n5695 = n5594 & n5694 ;
  assign n5696 = n5695 ^ n2204 ;
  assign n5697 = n5591 & n5696 ;
  assign n5698 = n5697 ^ n2008 ;
  assign n5587 = n5445 & ~n5562 ;
  assign n5588 = n5587 ^ n5340 ;
  assign n5699 = n5698 ^ n5588 ;
  assign n5700 = n5698 ^ n1739 ;
  assign n5701 = ~n5699 & ~n5700 ;
  assign n5702 = n5701 ^ n1763 ;
  assign n5703 = n5586 & n5702 ;
  assign n5705 = n5704 ^ n5703 ;
  assign n5706 = ~n5449 & ~n5562 ;
  assign n5707 = n5706 ^ n5451 ;
  assign n5708 = n5707 ^ n1427 ;
  assign n5709 = ~n5705 & ~n5708 ;
  assign n5710 = n5709 ^ n1450 ;
  assign n5711 = ~n5455 & ~n5562 ;
  assign n5712 = n5711 ^ n5457 ;
  assign n5713 = n5712 ^ n1290 ;
  assign n5714 = n5710 & n5713 ;
  assign n5715 = n5714 ^ n5712 ;
  assign n5718 = n5717 ^ n5715 ;
  assign n5719 = n5717 ^ n1136 ;
  assign n5720 = ~n5718 & n5719 ;
  assign n5721 = n5720 ^ n1143 ;
  assign n5722 = n5466 & ~n5562 ;
  assign n5723 = n5722 ^ n5334 ;
  assign n5726 = n5723 ^ n1034 ;
  assign n5727 = ~n5721 & n5726 ;
  assign n5724 = n5723 ^ n892 ;
  assign n5728 = n5727 ^ n5724 ;
  assign n5729 = n5468 & ~n5562 ;
  assign n5730 = n5729 ^ n5470 ;
  assign n5731 = n5730 ^ n786 ;
  assign n5732 = n5731 ^ n927 ;
  assign n5733 = ~n5728 & n5732 ;
  assign n5734 = n5733 ^ n5731 ;
  assign n5735 = n5475 & ~n5562 ;
  assign n5736 = n5735 ^ n5477 ;
  assign n5737 = n5736 ^ n696 ;
  assign n5738 = n5737 ^ n842 ;
  assign n5739 = ~n5734 & n5738 ;
  assign n5740 = n5739 ^ n5737 ;
  assign n5741 = n5481 & ~n5562 ;
  assign n5742 = n5741 ^ n5483 ;
  assign n5743 = n5742 ^ n609 ;
  assign n5744 = n5743 ^ n835 ;
  assign n5745 = ~n5740 & n5744 ;
  assign n5746 = n5745 ^ n5743 ;
  assign n5747 = ~n5583 & ~n5746 ;
  assign n5748 = n5747 ^ n834 ;
  assign n5749 = ~n5580 & ~n5748 ;
  assign n5750 = n5749 ^ n750 ;
  assign n5751 = ~n5576 & n5750 ;
  assign n5752 = n5751 ^ n5575 ;
  assign n5572 = n5568 ^ n401 ;
  assign n5570 = ~n5495 & ~n5562 ;
  assign n5571 = n5570 ^ n5322 ;
  assign n5573 = n5572 ^ n5571 ;
  assign n5753 = n5752 ^ n5573 ;
  assign n5754 = n5753 ^ n5572 ;
  assign n5755 = n5571 ^ n5568 ;
  assign n5756 = n5755 ^ n5572 ;
  assign n5757 = n5754 & ~n5756 ;
  assign n5758 = n5757 ^ n5572 ;
  assign n5759 = ~n5569 & n5758 ;
  assign n5760 = n5759 ^ n349 ;
  assign n5761 = n5503 & ~n5562 ;
  assign n5762 = n5761 ^ n5319 ;
  assign n5763 = n5762 ^ n291 ;
  assign n5764 = ~n5760 & n5763 ;
  assign n5765 = n5764 ^ n307 ;
  assign n5766 = n5565 & n5765 ;
  assign n5767 = n5766 ^ n5564 ;
  assign n5805 = n5803 ^ n5767 ;
  assign n5806 = ~n5804 & n5805 ;
  assign n5807 = n5806 ^ n203 ;
  assign n5808 = n5546 ^ n188 ;
  assign n5809 = ~n5562 & ~n5808 ;
  assign n5810 = n5809 ^ n5548 ;
  assign n5811 = n5810 ^ n157 ;
  assign n5812 = ~n5807 & ~n5811 ;
  assign n5813 = n5812 ^ n5810 ;
  assign n5814 = n5813 ^ n138 ;
  assign n5815 = n5552 & ~n5562 ;
  assign n5816 = n5815 ^ n5535 ;
  assign n5817 = n5816 ^ n5813 ;
  assign n5818 = ~n5814 & n5817 ;
  assign n5819 = n5818 ^ n138 ;
  assign n5820 = n183 & n5819 ;
  assign n5823 = n5554 ^ n138 ;
  assign n5824 = ~n5562 & n5823 ;
  assign n5825 = n5824 ^ n5533 ;
  assign n5828 = n5820 & ~n5825 ;
  assign n5829 = n5828 ^ n5819 ;
  assign n5830 = ~n5801 & ~n5829 ;
  assign n5876 = n5656 ^ n3908 ;
  assign n5877 = ~n5830 & n5876 ;
  assign n5878 = n5877 ^ n5606 ;
  assign n5879 = n5878 ^ n3722 ;
  assign n5940 = n5654 & ~n5830 ;
  assign n5941 = n5940 ^ n5609 ;
  assign n5880 = n5647 & ~n5830 ;
  assign n5881 = n5880 ^ n5650 ;
  assign n5882 = n5881 ^ n4153 ;
  assign n5932 = n5645 & ~n5830 ;
  assign n5933 = n5932 ^ n5613 ;
  assign n5936 = n5933 ^ n4153 ;
  assign n5885 = n5562 ^ n5317 ;
  assign n5886 = n5885 ^ x52 ;
  assign n5887 = n5886 ^ n5885 ;
  assign n5888 = n5634 ^ n5562 ;
  assign n5891 = ~n5887 & ~n5888 ;
  assign n5892 = n5891 ^ n5885 ;
  assign n5893 = ~n5830 & n5892 ;
  assign n5894 = n5893 ^ n5631 ;
  assign n5895 = n5894 ^ n5073 ;
  assign n5901 = n5562 ^ x51 ;
  assign n5902 = n5901 ^ n5830 ;
  assign n5903 = x48 & ~x49 ;
  assign n5904 = n5903 ^ x49 ;
  assign n5905 = n5904 ^ n5562 ;
  assign n5906 = n5905 ^ x50 ;
  assign n5907 = ~n5902 & n5906 ;
  assign n5915 = n5907 ^ n5562 ;
  assign n5916 = n5915 ^ n5317 ;
  assign n5900 = n5830 ^ n5562 ;
  assign n5908 = n5907 ^ n5900 ;
  assign n5909 = n5908 ^ n5907 ;
  assign n5912 = n5901 & n5909 ;
  assign n5913 = n5912 ^ n5907 ;
  assign n5914 = x50 & n5913 ;
  assign n5917 = n5916 ^ n5914 ;
  assign n5897 = ~n5830 & ~n5888 ;
  assign n5896 = n5562 ^ x52 ;
  assign n5898 = n5897 ^ n5896 ;
  assign n5918 = n5898 ^ n5317 ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5899 = n5898 ^ n5073 ;
  assign n5920 = n5919 ^ n5899 ;
  assign n5921 = n5895 & ~n5920 ;
  assign n5922 = n5921 ^ n5073 ;
  assign n5883 = n5639 & ~n5830 ;
  assign n5884 = n5883 ^ n5628 ;
  assign n5923 = n5922 ^ n5884 ;
  assign n5924 = n5922 ^ n4812 ;
  assign n5925 = ~n5923 & n5924 ;
  assign n5926 = n5925 ^ n4854 ;
  assign n5927 = n5643 & ~n5830 ;
  assign n5928 = n5927 ^ n5625 ;
  assign n5929 = n5928 ^ n4583 ;
  assign n5930 = n5926 & n5929 ;
  assign n5931 = n5930 ^ n4645 ;
  assign n5934 = n5933 ^ n4356 ;
  assign n5935 = ~n5931 & ~n5934 ;
  assign n5937 = n5936 ^ n5935 ;
  assign n5938 = n5882 & ~n5937 ;
  assign n5939 = n5938 ^ n4153 ;
  assign n5942 = n5941 ^ n5939 ;
  assign n5943 = n5941 ^ n3908 ;
  assign n5944 = n5942 & ~n5943 ;
  assign n5945 = n5944 ^ n3961 ;
  assign n5946 = n5879 & ~n5945 ;
  assign n5947 = n5946 ^ n3795 ;
  assign n6069 = ~n5814 & ~n5830 ;
  assign n6070 = n6069 ^ n5816 ;
  assign n6112 = n6070 ^ n183 ;
  assign n6063 = n5807 & ~n5830 ;
  assign n6064 = n6063 ^ n5810 ;
  assign n5768 = n5767 ^ n188 ;
  assign n5831 = n5768 & ~n5830 ;
  assign n5832 = n5831 ^ n5803 ;
  assign n5833 = n5832 ^ n157 ;
  assign n5834 = ~n5765 & ~n5830 ;
  assign n5835 = n5834 ^ n5564 ;
  assign n5836 = n5835 ^ n188 ;
  assign n5837 = ~n5760 & ~n5830 ;
  assign n5838 = n5837 ^ n5762 ;
  assign n5839 = n5838 ^ n245 ;
  assign n6044 = n5752 ^ n341 ;
  assign n6045 = n6044 ^ n462 ;
  assign n6046 = n5571 ^ n341 ;
  assign n6047 = n6046 ^ n462 ;
  assign n6048 = n6045 & ~n6047 ;
  assign n6049 = n6048 ^ n462 ;
  assign n6050 = ~n5830 & n6049 ;
  assign n6051 = n6050 ^ n5568 ;
  assign n6037 = n5752 ^ n401 ;
  assign n6038 = ~n5830 & n6037 ;
  assign n6039 = n6038 ^ n5571 ;
  assign n5840 = ~n5750 & ~n5830 ;
  assign n5841 = n5840 ^ n5575 ;
  assign n5842 = n5841 ^ n401 ;
  assign n5843 = ~n5748 & ~n5830 ;
  assign n5844 = n5843 ^ n5579 ;
  assign n5845 = n5844 ^ n457 ;
  assign n5846 = ~n5746 & ~n5830 ;
  assign n5847 = n5846 ^ n5582 ;
  assign n5848 = n5847 ^ n534 ;
  assign n5849 = n5740 & ~n5830 ;
  assign n5850 = n5849 ^ n5742 ;
  assign n5851 = n5850 ^ n609 ;
  assign n5852 = ~n5710 & ~n5830 ;
  assign n5853 = n5852 ^ n5712 ;
  assign n5854 = n5853 ^ n1136 ;
  assign n5994 = ~n5705 & ~n5830 ;
  assign n5995 = n5994 ^ n5707 ;
  assign n5998 = n5995 ^ n1136 ;
  assign n5855 = ~n5702 & ~n5830 ;
  assign n5856 = n5855 ^ n5585 ;
  assign n5857 = n5856 ^ n1427 ;
  assign n5985 = ~n5700 & ~n5830 ;
  assign n5986 = n5985 ^ n5588 ;
  assign n5990 = n5986 ^ n1427 ;
  assign n5858 = n5696 & ~n5830 ;
  assign n5859 = n5858 ^ n5590 ;
  assign n5860 = n5859 ^ n1739 ;
  assign n5863 = n5692 & ~n5830 ;
  assign n5864 = n5863 ^ n5597 ;
  assign n5865 = n5864 ^ n2175 ;
  assign n5866 = ~n5679 & ~n5830 ;
  assign n5867 = n5866 ^ n5600 ;
  assign n5868 = n5867 ^ n2707 ;
  assign n5869 = ~n5673 & ~n5830 ;
  assign n5870 = n5869 ^ n5675 ;
  assign n5871 = n5870 ^ n2894 ;
  assign n5955 = n5668 & ~n5830 ;
  assign n5956 = n5955 ^ n5670 ;
  assign n5959 = n5956 ^ n2894 ;
  assign n5872 = n5659 ^ n3722 ;
  assign n5873 = ~n5830 & ~n5872 ;
  assign n5874 = n5873 ^ n5662 ;
  assign n5875 = n5874 ^ n3538 ;
  assign n5948 = ~n5875 & n5947 ;
  assign n5949 = n5948 ^ n3596 ;
  assign n5950 = n5666 & ~n5830 ;
  assign n5951 = n5950 ^ n5603 ;
  assign n5952 = n5951 ^ n3320 ;
  assign n5953 = n5949 & ~n5952 ;
  assign n5954 = n5953 ^ n3387 ;
  assign n5957 = n5956 ^ n3093 ;
  assign n5958 = n5954 & n5957 ;
  assign n5960 = n5959 ^ n5958 ;
  assign n5961 = ~n5871 & n5960 ;
  assign n5962 = n5961 ^ n3396 ;
  assign n5963 = n5868 & ~n5962 ;
  assign n5964 = n5963 ^ n2707 ;
  assign n5965 = n5964 ^ n2511 ;
  assign n5966 = ~n5681 & ~n5830 ;
  assign n5967 = n5966 ^ n5683 ;
  assign n5968 = n5967 ^ n5964 ;
  assign n5969 = ~n5965 & ~n5968 ;
  assign n5970 = n5969 ^ n2530 ;
  assign n5971 = n5686 ^ n2511 ;
  assign n5972 = ~n5830 & ~n5971 ;
  assign n5973 = n5972 ^ n5688 ;
  assign n5974 = n5973 ^ n2366 ;
  assign n5975 = n5970 & ~n5974 ;
  assign n5976 = n5975 ^ n2399 ;
  assign n5977 = n5865 & n5976 ;
  assign n5978 = n5977 ^ n2175 ;
  assign n5861 = n5694 & ~n5830 ;
  assign n5862 = n5861 ^ n5593 ;
  assign n5979 = n5978 ^ n5862 ;
  assign n5980 = n5978 ^ n2008 ;
  assign n5981 = ~n5979 & n5980 ;
  assign n5982 = n5981 ^ n2064 ;
  assign n5983 = ~n5860 & ~n5982 ;
  assign n5984 = n5983 ^ n1739 ;
  assign n5987 = n5986 ^ n5984 ;
  assign n5988 = n5984 ^ n1572 ;
  assign n5989 = ~n5987 & n5988 ;
  assign n5991 = n5990 ^ n5989 ;
  assign n5992 = ~n5857 & ~n5991 ;
  assign n5993 = n5992 ^ n1450 ;
  assign n5996 = n5995 ^ n1290 ;
  assign n5997 = n5993 & n5996 ;
  assign n5999 = n5998 ^ n5997 ;
  assign n6000 = n5854 & n5999 ;
  assign n6001 = n6000 ^ n1143 ;
  assign n6002 = n5715 ^ n1136 ;
  assign n6003 = ~n5830 & n6002 ;
  assign n6004 = n6003 ^ n5717 ;
  assign n6007 = n6004 ^ n1034 ;
  assign n6008 = ~n6001 & n6007 ;
  assign n6005 = n6004 ^ n892 ;
  assign n6009 = n6008 ^ n6005 ;
  assign n6010 = n5721 & ~n5830 ;
  assign n6011 = n6010 ^ n5723 ;
  assign n6012 = n6011 ^ n786 ;
  assign n6013 = n6012 ^ n927 ;
  assign n6014 = ~n6009 & n6013 ;
  assign n6015 = n6014 ^ n6012 ;
  assign n6016 = n5728 & ~n5830 ;
  assign n6017 = n6016 ^ n5730 ;
  assign n6018 = n6017 ^ n696 ;
  assign n6019 = n6018 ^ n842 ;
  assign n6020 = ~n6015 & n6019 ;
  assign n6021 = n6020 ^ n6018 ;
  assign n6022 = n5734 & ~n5830 ;
  assign n6023 = n6022 ^ n5736 ;
  assign n6024 = n6023 ^ n609 ;
  assign n6025 = n6024 ^ n835 ;
  assign n6026 = ~n6021 & n6025 ;
  assign n6027 = n6026 ^ n6024 ;
  assign n6028 = ~n5851 & ~n6027 ;
  assign n6029 = n6028 ^ n834 ;
  assign n6030 = n5848 & ~n6029 ;
  assign n6031 = n6030 ^ n750 ;
  assign n6032 = n5845 & n6031 ;
  assign n6033 = n6032 ^ n5844 ;
  assign n6034 = n6033 ^ n5841 ;
  assign n6035 = n5842 & n6034 ;
  assign n6036 = n6035 ^ n401 ;
  assign n6040 = n6039 ^ n6036 ;
  assign n6041 = n6039 ^ n341 ;
  assign n6042 = n6040 & ~n6041 ;
  assign n6043 = n6042 ^ n341 ;
  assign n6052 = n6051 ^ n6043 ;
  assign n6053 = n6051 ^ n291 ;
  assign n6054 = n6052 & n6053 ;
  assign n6055 = n6054 ^ n307 ;
  assign n6056 = ~n5839 & n6055 ;
  assign n6057 = n6056 ^ n5838 ;
  assign n6058 = n6057 ^ n5835 ;
  assign n6059 = n5836 & n6058 ;
  assign n6060 = n6059 ^ n203 ;
  assign n6061 = ~n5833 & ~n6060 ;
  assign n6062 = n6061 ^ n5832 ;
  assign n6065 = n6064 ^ n6062 ;
  assign n6066 = n6064 ^ n138 ;
  assign n6067 = ~n6065 & ~n6066 ;
  assign n6068 = n6067 ^ n138 ;
  assign n6087 = n5555 ^ n138 ;
  assign n6090 = n6087 ^ n5791 ;
  assign n6091 = n6087 ^ n5508 ;
  assign n6092 = n6091 ^ n6087 ;
  assign n6093 = n6090 & n6092 ;
  assign n6094 = n6093 ^ n6087 ;
  assign n6095 = ~n1355 & ~n6094 ;
  assign n6096 = ~n5816 & n6095 ;
  assign n6097 = n5813 & n6096 ;
  assign n6099 = n5531 & n5770 ;
  assign n6100 = n6097 & n6099 ;
  assign n6098 = n6097 ^ n5820 ;
  assign n6101 = n6100 ^ n6098 ;
  assign n6073 = n5816 ^ n4971 ;
  assign n6074 = n6073 ^ n5801 ;
  assign n6075 = n6074 ^ n5813 ;
  assign n6076 = n6075 ^ n5814 ;
  assign n6077 = n6076 ^ n6075 ;
  assign n6078 = n6075 ^ n5817 ;
  assign n6079 = n6078 ^ n6075 ;
  assign n6080 = n6077 & n6079 ;
  assign n6081 = n6080 ^ n6075 ;
  assign n6082 = n5801 & n6081 ;
  assign n6102 = n6101 ^ n6082 ;
  assign n6083 = n6075 ^ n5801 ;
  assign n6084 = n6083 ^ n6082 ;
  assign n6085 = ~n183 & n5816 ;
  assign n6086 = ~n6084 & n6085 ;
  assign n6103 = n6102 ^ n6086 ;
  assign n6104 = ~n5825 & ~n6103 ;
  assign n6105 = n6104 ^ n6101 ;
  assign n6113 = n6068 & n6105 ;
  assign n6114 = ~n6112 & n6113 ;
  assign n6115 = n6114 ^ n6105 ;
  assign n6230 = n5947 & ~n6115 ;
  assign n6231 = n6230 ^ n5874 ;
  assign n6154 = ~n5945 & ~n6115 ;
  assign n6155 = n6154 ^ n5878 ;
  assign n6156 = n6155 ^ n3538 ;
  assign n6221 = n5939 ^ n3908 ;
  assign n6222 = ~n6115 & n6221 ;
  assign n6223 = n6222 ^ n5941 ;
  assign n6157 = ~n5937 & ~n6115 ;
  assign n6158 = n6157 ^ n5881 ;
  assign n6159 = n6158 ^ n3908 ;
  assign n6212 = n5931 & ~n6115 ;
  assign n6213 = n6212 ^ n5933 ;
  assign n6160 = n5926 & ~n6115 ;
  assign n6161 = n6160 ^ n5928 ;
  assign n6162 = n6161 ^ n4356 ;
  assign n6163 = n5917 & ~n6115 ;
  assign n6164 = n6163 ^ n5898 ;
  assign n6165 = n6164 ^ n5073 ;
  assign n6166 = n5904 ^ n5830 ;
  assign n6177 = n6115 & n6166 ;
  assign n6176 = n5904 ^ x50 ;
  assign n6178 = n6177 ^ n6176 ;
  assign n6179 = n6178 ^ n5562 ;
  assign n6181 = ~x46 & ~x47 ;
  assign n6182 = ~x48 & n6181 ;
  assign n6180 = n6115 ^ x49 ;
  assign n6183 = n6182 ^ n6180 ;
  assign n6185 = n6182 ^ n5830 ;
  assign n6188 = n6183 & n6185 ;
  assign n6184 = n6183 ^ n5830 ;
  assign n6186 = n6185 ^ n6184 ;
  assign n6187 = ~n5903 & ~n6186 ;
  assign n6189 = n6188 ^ n6187 ;
  assign n6190 = n6189 ^ n6178 ;
  assign n6191 = ~n6179 & n6190 ;
  assign n6192 = n6191 ^ n5562 ;
  assign n6196 = n6192 ^ n5073 ;
  assign n6174 = ~x50 & ~n5830 ;
  assign n6167 = n6166 ^ n5905 ;
  assign n6168 = n6167 ^ n5905 ;
  assign n6169 = n5906 ^ n5905 ;
  assign n6170 = n6168 & n6169 ;
  assign n6171 = n6170 ^ n5905 ;
  assign n6172 = ~n6115 & n6171 ;
  assign n6173 = n6172 ^ x51 ;
  assign n6175 = n6174 ^ n6173 ;
  assign n6193 = n6192 ^ n6175 ;
  assign n6194 = n6175 ^ n5317 ;
  assign n6195 = n6193 & ~n6194 ;
  assign n6197 = n6196 ^ n6195 ;
  assign n6198 = ~n6165 & n6197 ;
  assign n6199 = n6198 ^ n5115 ;
  assign n6200 = ~n5920 & ~n6115 ;
  assign n6201 = n6200 ^ n5894 ;
  assign n6202 = n6201 ^ n4812 ;
  assign n6203 = n6199 & n6202 ;
  assign n6204 = n6203 ^ n4854 ;
  assign n6205 = n5924 & ~n6115 ;
  assign n6206 = n6205 ^ n5884 ;
  assign n6207 = n6206 ^ n4583 ;
  assign n6208 = n6204 & n6207 ;
  assign n6209 = n6208 ^ n4645 ;
  assign n6210 = n6162 & ~n6209 ;
  assign n6211 = n6210 ^ n6161 ;
  assign n6214 = n6213 ^ n6211 ;
  assign n6215 = n6213 ^ n4153 ;
  assign n6216 = n6214 & ~n6215 ;
  assign n6217 = n6216 ^ n4153 ;
  assign n6218 = n6217 ^ n6158 ;
  assign n6219 = n6159 & ~n6218 ;
  assign n6220 = n6219 ^ n3908 ;
  assign n6224 = n6223 ^ n6220 ;
  assign n6225 = n6223 ^ n3722 ;
  assign n6226 = n6224 & n6225 ;
  assign n6227 = n6226 ^ n3795 ;
  assign n6228 = n6156 & n6227 ;
  assign n6229 = n6228 ^ n3538 ;
  assign n6232 = n6231 ^ n6229 ;
  assign n6233 = n6231 ^ n3320 ;
  assign n6234 = n6232 & ~n6233 ;
  assign n6235 = n6234 ^ n3387 ;
  assign n6071 = n6070 ^ n6068 ;
  assign n6072 = n6068 ^ n183 ;
  assign n6108 = ~n6072 & n6105 ;
  assign n6109 = n6108 ^ n183 ;
  assign n6110 = n6071 & n6109 ;
  assign n6111 = n6062 ^ n138 ;
  assign n6116 = ~n6111 & ~n6115 ;
  assign n6117 = n6116 ^ n6064 ;
  assign n6118 = n6033 ^ n401 ;
  assign n6119 = ~n6115 & ~n6118 ;
  assign n6120 = n6119 ^ n5841 ;
  assign n6121 = n6120 ^ n341 ;
  assign n6310 = ~n6031 & ~n6115 ;
  assign n6311 = n6310 ^ n5844 ;
  assign n6122 = ~n6027 & ~n6115 ;
  assign n6123 = n6122 ^ n5850 ;
  assign n6124 = n6123 ^ n534 ;
  assign n6125 = n6021 & ~n6115 ;
  assign n6126 = n6125 ^ n6023 ;
  assign n6301 = n6126 ^ n534 ;
  assign n6127 = n6126 ^ n609 ;
  assign n6128 = ~n5993 & ~n6115 ;
  assign n6129 = n6128 ^ n5995 ;
  assign n6130 = n6129 ^ n1136 ;
  assign n6267 = ~n5991 & ~n6115 ;
  assign n6268 = n6267 ^ n5856 ;
  assign n6271 = n6268 ^ n1136 ;
  assign n6131 = ~n5982 & ~n6115 ;
  assign n6132 = n6131 ^ n5859 ;
  assign n6260 = n6132 ^ n1427 ;
  assign n6133 = n6132 ^ n1572 ;
  assign n6136 = n5976 & ~n6115 ;
  assign n6137 = n6136 ^ n5864 ;
  assign n6138 = n6137 ^ n2008 ;
  assign n6139 = n5970 & ~n6115 ;
  assign n6140 = n6139 ^ n5973 ;
  assign n6141 = n6140 ^ n2175 ;
  assign n6142 = ~n5965 & ~n6115 ;
  assign n6143 = n6142 ^ n5967 ;
  assign n6144 = n6143 ^ n2366 ;
  assign n6243 = ~n5962 & ~n6115 ;
  assign n6244 = n6243 ^ n5867 ;
  assign n6145 = n5960 & ~n6115 ;
  assign n6146 = n6145 ^ n5870 ;
  assign n6147 = n6146 ^ n2707 ;
  assign n6148 = ~n5954 & ~n6115 ;
  assign n6149 = n6148 ^ n5956 ;
  assign n6150 = n6149 ^ n2894 ;
  assign n6151 = n5949 & ~n6115 ;
  assign n6152 = n6151 ^ n5951 ;
  assign n6237 = n6152 ^ n2894 ;
  assign n6153 = n6152 ^ n3093 ;
  assign n6236 = n6153 & n6235 ;
  assign n6238 = n6237 ^ n6236 ;
  assign n6239 = n6150 & n6238 ;
  assign n6240 = n6239 ^ n3396 ;
  assign n6241 = n6147 & ~n6240 ;
  assign n6242 = n6241 ^ n2707 ;
  assign n6245 = n6244 ^ n6242 ;
  assign n6246 = n6244 ^ n2511 ;
  assign n6247 = ~n6245 & ~n6246 ;
  assign n6248 = n6247 ^ n2530 ;
  assign n6249 = ~n6144 & n6248 ;
  assign n6250 = n6249 ^ n2399 ;
  assign n6251 = ~n6141 & n6250 ;
  assign n6252 = n6251 ^ n2204 ;
  assign n6253 = n6138 & n6252 ;
  assign n6254 = n6253 ^ n2008 ;
  assign n6134 = n5980 & ~n6115 ;
  assign n6135 = n6134 ^ n5862 ;
  assign n6255 = n6254 ^ n6135 ;
  assign n6256 = n6254 ^ n1739 ;
  assign n6257 = ~n6255 & ~n6256 ;
  assign n6258 = n6257 ^ n1763 ;
  assign n6259 = n6133 & n6258 ;
  assign n6261 = n6260 ^ n6259 ;
  assign n6262 = ~n5988 & ~n6115 ;
  assign n6263 = n6262 ^ n5986 ;
  assign n6264 = n6263 ^ n1427 ;
  assign n6265 = ~n6261 & ~n6264 ;
  assign n6266 = n6265 ^ n1450 ;
  assign n6269 = n6268 ^ n1290 ;
  assign n6270 = n6266 & n6269 ;
  assign n6272 = n6271 ^ n6270 ;
  assign n6273 = n6130 & n6272 ;
  assign n6274 = n6273 ^ n1143 ;
  assign n6275 = n5999 & ~n6115 ;
  assign n6276 = n6275 ^ n5853 ;
  assign n6279 = n6276 ^ n1034 ;
  assign n6280 = ~n6274 & n6279 ;
  assign n6277 = n6276 ^ n892 ;
  assign n6281 = n6280 ^ n6277 ;
  assign n6282 = n6001 & ~n6115 ;
  assign n6283 = n6282 ^ n6004 ;
  assign n6284 = n6283 ^ n786 ;
  assign n6285 = n6284 ^ n927 ;
  assign n6286 = ~n6281 & n6285 ;
  assign n6287 = n6286 ^ n6284 ;
  assign n6288 = n6009 & ~n6115 ;
  assign n6289 = n6288 ^ n6011 ;
  assign n6290 = n6289 ^ n696 ;
  assign n6291 = n6290 ^ n842 ;
  assign n6292 = ~n6287 & n6291 ;
  assign n6293 = n6292 ^ n6290 ;
  assign n6294 = n6015 & ~n6115 ;
  assign n6295 = n6294 ^ n6017 ;
  assign n6296 = n6295 ^ n609 ;
  assign n6297 = n6296 ^ n835 ;
  assign n6298 = ~n6293 & n6297 ;
  assign n6299 = n6298 ^ n6296 ;
  assign n6300 = ~n6127 & n6299 ;
  assign n6302 = n6301 ^ n6300 ;
  assign n6303 = n6124 & n6302 ;
  assign n6304 = n6303 ^ n750 ;
  assign n6305 = ~n6029 & ~n6115 ;
  assign n6306 = n6305 ^ n5847 ;
  assign n6307 = n6306 ^ n457 ;
  assign n6308 = n6304 & ~n6307 ;
  assign n6309 = n6308 ^ n6306 ;
  assign n6312 = n6311 ^ n6309 ;
  assign n6313 = n6311 ^ n401 ;
  assign n6314 = n6312 & ~n6313 ;
  assign n6315 = n6314 ^ n462 ;
  assign n6316 = n6121 & n6315 ;
  assign n6317 = n6316 ^ n349 ;
  assign n6318 = n6036 ^ n341 ;
  assign n6319 = ~n6115 & n6318 ;
  assign n6320 = n6319 ^ n6039 ;
  assign n6321 = n6320 ^ n291 ;
  assign n6322 = ~n6317 & n6321 ;
  assign n6323 = n6322 ^ n307 ;
  assign n6324 = n6043 ^ n291 ;
  assign n6325 = ~n6115 & ~n6324 ;
  assign n6326 = n6325 ^ n6051 ;
  assign n6327 = n6326 ^ n245 ;
  assign n6328 = n6323 & ~n6327 ;
  assign n6329 = n6328 ^ n6326 ;
  assign n6330 = n6329 ^ n188 ;
  assign n6331 = ~n6055 & ~n6115 ;
  assign n6332 = n6331 ^ n5838 ;
  assign n6333 = n6332 ^ n6329 ;
  assign n6334 = ~n6330 & ~n6333 ;
  assign n6335 = n6334 ^ n203 ;
  assign n6336 = n6057 ^ n188 ;
  assign n6337 = ~n6115 & ~n6336 ;
  assign n6338 = n6337 ^ n5835 ;
  assign n6339 = n6338 ^ n157 ;
  assign n6340 = ~n6335 & n6339 ;
  assign n6341 = n6340 ^ n6338 ;
  assign n6342 = n138 & n6341 ;
  assign n6343 = n6060 & ~n6115 ;
  assign n6344 = n6343 ^ n5832 ;
  assign n6345 = n6341 ^ n138 ;
  assign n6346 = n6345 ^ n6342 ;
  assign n6347 = ~n6344 & n6346 ;
  assign n6348 = ~n6342 & ~n6347 ;
  assign n6349 = ~n6117 & ~n6348 ;
  assign n6350 = ~n6110 & n6349 ;
  assign n6351 = n6350 ^ n6110 ;
  assign n6352 = ~n183 & ~n6351 ;
  assign n6353 = n6066 ^ n6062 ;
  assign n6354 = n6341 ^ n6064 ;
  assign n6356 = n138 & n6354 ;
  assign n6357 = n6356 ^ n6064 ;
  assign n6358 = ~n6353 & ~n6357 ;
  assign n6359 = n6358 ^ n6115 ;
  assign n6368 = n6062 & n6115 ;
  assign n6369 = n6368 ^ n6070 ;
  assign n6370 = n6369 ^ n6359 ;
  assign n6367 = n6070 ^ n138 ;
  assign n6371 = n6370 ^ n6367 ;
  assign n6360 = n6115 ^ n6062 ;
  assign n6364 = n6115 & n6341 ;
  assign n6365 = n6364 ^ n138 ;
  assign n6366 = ~n6360 & ~n6365 ;
  assign n6372 = n6371 ^ n6366 ;
  assign n6373 = n6372 ^ n6370 ;
  assign n6374 = n6373 ^ n6366 ;
  assign n6375 = n6070 ^ n6062 ;
  assign n6376 = n6366 ^ n6062 ;
  assign n6377 = n6375 & n6376 ;
  assign n6378 = ~n6374 & n6377 ;
  assign n6379 = n6378 ^ n6372 ;
  assign n6380 = n6379 ^ n6359 ;
  assign n6381 = n6064 & ~n6347 ;
  assign n6382 = ~n6380 & n6381 ;
  assign n6383 = n6382 ^ n6347 ;
  assign n6385 = ~n6369 & ~n6383 ;
  assign n6386 = n6359 & n6385 ;
  assign n6387 = n6386 ^ n6382 ;
  assign n6388 = n6352 & ~n6387 ;
  assign n6389 = n6388 ^ n6351 ;
  assign n6390 = ~n6235 & n6389 ;
  assign n6391 = n6390 ^ n6152 ;
  assign n6392 = n6391 ^ n2894 ;
  assign n6490 = n6229 ^ n3320 ;
  assign n6491 = n6389 & n6490 ;
  assign n6492 = n6491 ^ n6231 ;
  assign n6495 = n6492 ^ n2894 ;
  assign n6393 = n6220 ^ n3722 ;
  assign n6394 = n6389 & ~n6393 ;
  assign n6395 = n6394 ^ n6223 ;
  assign n6396 = n6395 ^ n3538 ;
  assign n6476 = n6217 ^ n3908 ;
  assign n6477 = n6389 & n6476 ;
  assign n6478 = n6477 ^ n6158 ;
  assign n6469 = n6211 ^ n4153 ;
  assign n6470 = n6389 & n6469 ;
  assign n6471 = n6470 ^ n6213 ;
  assign n6397 = n6209 & n6389 ;
  assign n6398 = n6397 ^ n6161 ;
  assign n6399 = n6398 ^ n4153 ;
  assign n6461 = n6204 & n6389 ;
  assign n6462 = n6461 ^ n6206 ;
  assign n6465 = n6462 ^ n4153 ;
  assign n6400 = n6199 & n6389 ;
  assign n6401 = n6400 ^ n6201 ;
  assign n6402 = n6401 ^ n4583 ;
  assign n6405 = n6192 ^ n5317 ;
  assign n6406 = n6389 & n6405 ;
  assign n6407 = n6406 ^ n6175 ;
  assign n6408 = n6407 ^ n5073 ;
  assign n6415 = n6185 ^ n6115 ;
  assign n6420 = n6415 ^ x49 ;
  assign n6413 = n6185 ^ x48 ;
  assign n6414 = n6413 ^ n6185 ;
  assign n6416 = n6415 ^ n6185 ;
  assign n6417 = n6414 & ~n6416 ;
  assign n6418 = n6417 ^ n6185 ;
  assign n6419 = ~n6389 & ~n6418 ;
  assign n6421 = n6420 ^ n6419 ;
  assign n6422 = n6421 ^ n5562 ;
  assign n6429 = n6115 ^ n5830 ;
  assign n6425 = n6389 ^ x47 ;
  assign n6424 = ~x44 & ~x45 ;
  assign n6426 = n6425 ^ n6424 ;
  assign n6427 = n6425 ^ n6115 ;
  assign n6428 = n6426 & n6427 ;
  assign n6430 = n6429 ^ n6428 ;
  assign n6431 = n6430 ^ n6429 ;
  assign n6423 = n6389 ^ n6115 ;
  assign n6432 = n6431 ^ n6423 ;
  assign n6433 = n6432 ^ n6431 ;
  assign n6434 = n6431 ^ n6425 ;
  assign n6435 = n6434 ^ n6431 ;
  assign n6436 = ~n6433 & n6435 ;
  assign n6437 = n6436 ^ n6431 ;
  assign n6438 = x46 & n6437 ;
  assign n6439 = n6438 ^ n6430 ;
  assign n6441 = n6181 ^ n6115 ;
  assign n6442 = n6389 & ~n6441 ;
  assign n6440 = n6115 ^ x48 ;
  assign n6443 = n6442 ^ n6440 ;
  assign n6444 = n6443 ^ n5830 ;
  assign n6445 = ~n6439 & ~n6444 ;
  assign n6446 = n6445 ^ n6443 ;
  assign n6447 = n6446 ^ n6421 ;
  assign n6448 = n6422 & n6447 ;
  assign n6449 = n6448 ^ n5885 ;
  assign n6409 = n6189 ^ n5562 ;
  assign n6410 = n6389 & n6409 ;
  assign n6411 = n6410 ^ n6178 ;
  assign n6450 = n6411 ^ n5317 ;
  assign n6451 = ~n6449 & ~n6450 ;
  assign n6412 = n6411 ^ n5073 ;
  assign n6452 = n6451 ^ n6412 ;
  assign n6453 = n6408 & ~n6452 ;
  assign n6454 = n6453 ^ n5073 ;
  assign n6403 = n6197 & n6389 ;
  assign n6404 = n6403 ^ n6164 ;
  assign n6455 = n6454 ^ n6404 ;
  assign n6456 = n6454 ^ n4812 ;
  assign n6457 = n6455 & n6456 ;
  assign n6458 = n6457 ^ n4854 ;
  assign n6459 = n6402 & n6458 ;
  assign n6460 = n6459 ^ n4645 ;
  assign n6463 = n6462 ^ n4356 ;
  assign n6464 = ~n6460 & n6463 ;
  assign n6466 = n6465 ^ n6464 ;
  assign n6467 = n6399 & n6466 ;
  assign n6468 = n6467 ^ n4153 ;
  assign n6472 = n6471 ^ n6468 ;
  assign n6473 = n6471 ^ n3908 ;
  assign n6474 = n6472 & ~n6473 ;
  assign n6475 = n6474 ^ n3908 ;
  assign n6479 = n6478 ^ n6475 ;
  assign n6480 = n6478 ^ n3722 ;
  assign n6481 = ~n6479 & ~n6480 ;
  assign n6482 = n6481 ^ n3795 ;
  assign n6483 = n6396 & n6482 ;
  assign n6484 = n6483 ^ n3596 ;
  assign n6485 = n6227 & n6389 ;
  assign n6486 = n6485 ^ n6155 ;
  assign n6487 = n6486 ^ n3320 ;
  assign n6488 = n6484 & n6487 ;
  assign n6489 = n6488 ^ n3387 ;
  assign n6493 = n6492 ^ n3093 ;
  assign n6494 = n6489 & n6493 ;
  assign n6496 = n6495 ^ n6494 ;
  assign n6497 = n6392 & n6496 ;
  assign n6498 = n6497 ^ n3396 ;
  assign n6499 = n6345 & n6389 ;
  assign n6500 = n6499 ^ n6344 ;
  assign n6501 = n6500 ^ n183 ;
  assign n6515 = n6347 ^ n6342 ;
  assign n6516 = n6389 & n6515 ;
  assign n6519 = n6516 ^ n6348 ;
  assign n6520 = n6519 ^ n6516 ;
  assign n6523 = n6351 & ~n6520 ;
  assign n6524 = n6523 ^ n6516 ;
  assign n6525 = n183 & ~n6524 ;
  assign n6502 = n6344 ^ n6341 ;
  assign n6503 = n6341 ^ n4971 ;
  assign n6504 = ~n6502 & n6503 ;
  assign n6511 = n6504 ^ n1355 ;
  assign n6508 = n138 & n6504 ;
  assign n6509 = n6508 ^ n1003 ;
  assign n6510 = ~n6344 & ~n6509 ;
  assign n6512 = n6511 ^ n6510 ;
  assign n6513 = n6389 & ~n6512 ;
  assign n6517 = n6516 ^ n6513 ;
  assign n6526 = n6525 ^ n6517 ;
  assign n6527 = n6117 & ~n6526 ;
  assign n6529 = n6344 & ~n6389 ;
  assign n6530 = n6527 & n6529 ;
  assign n6514 = n6513 ^ n6117 ;
  assign n6528 = n6527 ^ n6514 ;
  assign n6531 = n6530 ^ n6528 ;
  assign n6532 = n6335 & n6389 ;
  assign n6533 = n6532 ^ n6338 ;
  assign n6534 = n6533 ^ n138 ;
  assign n6537 = ~n6317 & n6389 ;
  assign n6538 = n6537 ^ n6320 ;
  assign n6539 = n6538 ^ n245 ;
  assign n6540 = n6315 & n6389 ;
  assign n6541 = n6540 ^ n6120 ;
  assign n6542 = n6541 ^ n291 ;
  assign n6543 = ~n6304 & n6389 ;
  assign n6544 = n6543 ^ n6306 ;
  assign n6545 = n6544 ^ n401 ;
  assign n6546 = n6302 & n6389 ;
  assign n6547 = n6546 ^ n6123 ;
  assign n6548 = n6547 ^ n457 ;
  assign n6549 = n6293 & n6389 ;
  assign n6550 = n6549 ^ n6295 ;
  assign n6551 = n6550 ^ n609 ;
  assign n6552 = ~n6266 & n6389 ;
  assign n6553 = n6552 ^ n6268 ;
  assign n6554 = n6553 ^ n1136 ;
  assign n6603 = ~n6261 & n6389 ;
  assign n6604 = n6603 ^ n6263 ;
  assign n6607 = n6604 ^ n1136 ;
  assign n6592 = ~n6256 & n6389 ;
  assign n6593 = n6592 ^ n6135 ;
  assign n6596 = n6593 ^ n1427 ;
  assign n6555 = n6252 & n6389 ;
  assign n6556 = n6555 ^ n6137 ;
  assign n6557 = n6556 ^ n1739 ;
  assign n6562 = ~n6240 & n6389 ;
  assign n6563 = n6562 ^ n6146 ;
  assign n6564 = n6563 ^ n2511 ;
  assign n6565 = n6238 & n6389 ;
  assign n6566 = n6565 ^ n6149 ;
  assign n6567 = n6566 ^ n2707 ;
  assign n6568 = ~n6498 & ~n6567 ;
  assign n6569 = n6568 ^ n2707 ;
  assign n6570 = n6569 ^ n6563 ;
  assign n6571 = ~n6564 & ~n6570 ;
  assign n6572 = n6571 ^ n2530 ;
  assign n6573 = n6242 ^ n2511 ;
  assign n6574 = n6389 & ~n6573 ;
  assign n6575 = n6574 ^ n6244 ;
  assign n6576 = n6575 ^ n2366 ;
  assign n6577 = n6572 & ~n6576 ;
  assign n6578 = n6577 ^ n2399 ;
  assign n6579 = n6248 & n6389 ;
  assign n6580 = n6579 ^ n6143 ;
  assign n6581 = n6580 ^ n2175 ;
  assign n6582 = n6578 & ~n6581 ;
  assign n6583 = n6582 ^ n2175 ;
  assign n6560 = n6556 ^ n2008 ;
  assign n6558 = n6250 & n6389 ;
  assign n6559 = n6558 ^ n6140 ;
  assign n6561 = n6560 ^ n6559 ;
  assign n6584 = n6583 ^ n6561 ;
  assign n6585 = n6584 ^ n6560 ;
  assign n6586 = n6559 ^ n6556 ;
  assign n6587 = n6586 ^ n6560 ;
  assign n6588 = n6585 & ~n6587 ;
  assign n6589 = n6588 ^ n6560 ;
  assign n6590 = ~n6557 & ~n6589 ;
  assign n6591 = n6590 ^ n1763 ;
  assign n6594 = n6593 ^ n1572 ;
  assign n6595 = n6591 & n6594 ;
  assign n6597 = n6596 ^ n6595 ;
  assign n6598 = ~n6258 & n6389 ;
  assign n6599 = n6598 ^ n6132 ;
  assign n6600 = n6599 ^ n1427 ;
  assign n6601 = ~n6597 & ~n6600 ;
  assign n6602 = n6601 ^ n1450 ;
  assign n6605 = n6604 ^ n1290 ;
  assign n6606 = n6602 & n6605 ;
  assign n6608 = n6607 ^ n6606 ;
  assign n6609 = n6554 & n6608 ;
  assign n6610 = n6609 ^ n1143 ;
  assign n6611 = n6272 & n6389 ;
  assign n6612 = n6611 ^ n6129 ;
  assign n6615 = n6612 ^ n1034 ;
  assign n6616 = ~n6610 & n6615 ;
  assign n6613 = n6612 ^ n892 ;
  assign n6617 = n6616 ^ n6613 ;
  assign n6618 = n6274 & n6389 ;
  assign n6619 = n6618 ^ n6276 ;
  assign n6620 = n6619 ^ n786 ;
  assign n6621 = n6620 ^ n927 ;
  assign n6622 = ~n6617 & n6621 ;
  assign n6623 = n6622 ^ n6620 ;
  assign n6624 = n6281 & n6389 ;
  assign n6625 = n6624 ^ n6283 ;
  assign n6626 = n6625 ^ n696 ;
  assign n6627 = n6626 ^ n842 ;
  assign n6628 = ~n6623 & n6627 ;
  assign n6629 = n6628 ^ n6626 ;
  assign n6630 = n6287 & n6389 ;
  assign n6631 = n6630 ^ n6289 ;
  assign n6632 = n6631 ^ n609 ;
  assign n6633 = n6632 ^ n835 ;
  assign n6634 = ~n6629 & n6633 ;
  assign n6635 = n6634 ^ n6632 ;
  assign n6636 = ~n6551 & ~n6635 ;
  assign n6637 = n6636 ^ n834 ;
  assign n6638 = ~n6299 & n6389 ;
  assign n6639 = n6638 ^ n6126 ;
  assign n6640 = n6639 ^ n534 ;
  assign n6641 = ~n6637 & n6640 ;
  assign n6642 = n6641 ^ n750 ;
  assign n6643 = ~n6548 & n6642 ;
  assign n6644 = n6643 ^ n6547 ;
  assign n6645 = n6644 ^ n6544 ;
  assign n6646 = n6545 & ~n6645 ;
  assign n6647 = n6646 ^ n401 ;
  assign n6648 = n6647 ^ n341 ;
  assign n6649 = n6309 ^ n401 ;
  assign n6650 = n6389 & n6649 ;
  assign n6651 = n6650 ^ n6311 ;
  assign n6652 = n6651 ^ n6647 ;
  assign n6653 = n6648 & n6652 ;
  assign n6654 = n6653 ^ n349 ;
  assign n6655 = ~n6542 & ~n6654 ;
  assign n6656 = n6655 ^ n307 ;
  assign n6657 = ~n6539 & n6656 ;
  assign n6658 = n6657 ^ n6538 ;
  assign n6535 = ~n6323 & n6389 ;
  assign n6536 = n6535 ^ n6326 ;
  assign n6659 = n6658 ^ n6536 ;
  assign n6660 = n6658 ^ n188 ;
  assign n6661 = ~n6659 & ~n6660 ;
  assign n6662 = n6661 ^ n203 ;
  assign n6663 = ~n6330 & n6389 ;
  assign n6664 = n6663 ^ n6332 ;
  assign n6665 = n6664 ^ n157 ;
  assign n6666 = ~n6662 & ~n6665 ;
  assign n6667 = n6666 ^ n6664 ;
  assign n6668 = n6667 ^ n138 ;
  assign n6669 = n6534 & ~n6668 ;
  assign n6670 = n6669 ^ n138 ;
  assign n6671 = n6531 & n6670 ;
  assign n6672 = n6501 & n6671 ;
  assign n6673 = n6672 ^ n6531 ;
  assign n6674 = ~n6498 & ~n6673 ;
  assign n6675 = n6674 ^ n6566 ;
  assign n6676 = n6675 ^ n2511 ;
  assign n6677 = n6496 & ~n6673 ;
  assign n6678 = n6677 ^ n6391 ;
  assign n6679 = n6678 ^ n2707 ;
  assign n6782 = ~n6489 & ~n6673 ;
  assign n6783 = n6782 ^ n6492 ;
  assign n6680 = n6484 & ~n6673 ;
  assign n6681 = n6680 ^ n6486 ;
  assign n6682 = n6681 ^ n3093 ;
  assign n6683 = n6475 ^ n3722 ;
  assign n6684 = ~n6673 & ~n6683 ;
  assign n6685 = n6684 ^ n6478 ;
  assign n6686 = n6685 ^ n3538 ;
  assign n6760 = n6466 & ~n6673 ;
  assign n6761 = n6760 ^ n6398 ;
  assign n6754 = n6460 & ~n6673 ;
  assign n6755 = n6754 ^ n6462 ;
  assign n6687 = n6458 & ~n6673 ;
  assign n6688 = n6687 ^ n6401 ;
  assign n6689 = n6688 ^ n4356 ;
  assign n6690 = ~n6452 & ~n6673 ;
  assign n6691 = n6690 ^ n6407 ;
  assign n6692 = n6691 ^ n4812 ;
  assign n6693 = n6449 & ~n6673 ;
  assign n6694 = n6693 ^ n6411 ;
  assign n6695 = n6694 ^ n5073 ;
  assign n6696 = n6446 ^ n5562 ;
  assign n6697 = ~n6673 & ~n6696 ;
  assign n6698 = n6697 ^ n6421 ;
  assign n6700 = n6698 ^ n5317 ;
  assign n6734 = n6439 & ~n6673 ;
  assign n6735 = n6734 ^ n6443 ;
  assign n6704 = n6424 ^ n6389 ;
  assign n6705 = ~n6673 & n6704 ;
  assign n6706 = n6705 ^ n6389 ;
  assign n6707 = x46 & n6706 ;
  assign n6701 = n6424 ^ n6115 ;
  assign n6702 = ~n6673 & ~n6701 ;
  assign n6703 = n6702 ^ n6425 ;
  assign n6708 = n6707 ^ n6703 ;
  assign n6709 = n6708 ^ n5830 ;
  assign n6717 = n6115 ^ x45 ;
  assign n6711 = ~x42 & ~x43 ;
  assign n6710 = n6389 ^ x44 ;
  assign n6712 = n6711 ^ n6710 ;
  assign n6713 = n6673 ^ n6389 ;
  assign n6714 = n6713 ^ x45 ;
  assign n6715 = n6712 & n6714 ;
  assign n6716 = n6715 ^ n6423 ;
  assign n6718 = n6717 ^ n6716 ;
  assign n6719 = n6718 ^ x45 ;
  assign n6720 = n6719 ^ n6673 ;
  assign n6721 = n6720 ^ n6718 ;
  assign n6722 = n6718 ^ n6713 ;
  assign n6723 = n6722 ^ n6718 ;
  assign n6724 = n6721 & n6723 ;
  assign n6725 = n6724 ^ n6718 ;
  assign n6726 = x44 & ~n6725 ;
  assign n6727 = n6726 ^ n6716 ;
  assign n6728 = n6706 ^ x46 ;
  assign n6729 = n6728 ^ n6115 ;
  assign n6730 = ~n6727 & n6729 ;
  assign n6731 = n6730 ^ n6429 ;
  assign n6732 = n6709 & n6731 ;
  assign n6733 = n6732 ^ n5830 ;
  assign n6736 = n6735 ^ n6733 ;
  assign n6737 = n6735 ^ n5562 ;
  assign n6738 = n6736 & ~n6737 ;
  assign n6739 = n6738 ^ n5885 ;
  assign n6740 = n6700 & ~n6739 ;
  assign n6699 = n6698 ^ n5073 ;
  assign n6741 = n6740 ^ n6699 ;
  assign n6742 = ~n6695 & n6741 ;
  assign n6743 = n6742 ^ n5115 ;
  assign n6744 = n6692 & n6743 ;
  assign n6745 = n6744 ^ n4812 ;
  assign n6746 = n6745 ^ n4583 ;
  assign n6747 = n6456 & ~n6673 ;
  assign n6748 = n6747 ^ n6404 ;
  assign n6749 = n6748 ^ n6745 ;
  assign n6750 = n6746 & n6749 ;
  assign n6751 = n6750 ^ n4645 ;
  assign n6752 = n6689 & ~n6751 ;
  assign n6753 = n6752 ^ n6688 ;
  assign n6756 = n6755 ^ n6753 ;
  assign n6757 = n6755 ^ n4153 ;
  assign n6758 = ~n6756 & n6757 ;
  assign n6759 = n6758 ^ n4153 ;
  assign n6762 = n6761 ^ n6759 ;
  assign n6763 = n6761 ^ n3908 ;
  assign n6764 = ~n6762 & n6763 ;
  assign n6765 = n6764 ^ n3908 ;
  assign n6766 = n6765 ^ n3722 ;
  assign n6767 = n6468 ^ n3908 ;
  assign n6768 = ~n6673 & n6767 ;
  assign n6769 = n6768 ^ n6471 ;
  assign n6770 = n6769 ^ n6765 ;
  assign n6771 = ~n6766 & n6770 ;
  assign n6772 = n6771 ^ n3795 ;
  assign n6773 = ~n6686 & n6772 ;
  assign n6774 = n6773 ^ n3596 ;
  assign n6775 = n6482 & ~n6673 ;
  assign n6776 = n6775 ^ n6395 ;
  assign n6777 = n6776 ^ n3320 ;
  assign n6778 = n6774 & n6777 ;
  assign n6779 = n6778 ^ n3387 ;
  assign n6780 = ~n6682 & n6779 ;
  assign n6781 = n6780 ^ n6681 ;
  assign n6784 = n6783 ^ n6781 ;
  assign n6785 = n6783 ^ n2894 ;
  assign n6786 = n6784 & n6785 ;
  assign n6787 = n6786 ^ n3396 ;
  assign n6788 = ~n6679 & ~n6787 ;
  assign n6789 = n6788 ^ n2707 ;
  assign n6790 = n6789 ^ n6675 ;
  assign n6791 = n6676 & n6790 ;
  assign n6792 = n6791 ^ n2530 ;
  assign n6793 = n6569 ^ n2511 ;
  assign n6794 = ~n6673 & ~n6793 ;
  assign n6795 = n6794 ^ n6563 ;
  assign n6796 = n6795 ^ n2366 ;
  assign n6797 = n6792 & ~n6796 ;
  assign n6798 = n6797 ^ n2399 ;
  assign n6812 = n6500 ^ n138 ;
  assign n6814 = n6500 ^ n130 ;
  assign n6813 = n6533 ^ n6500 ;
  assign n6815 = n6814 ^ n6813 ;
  assign n6818 = n183 & n6815 ;
  assign n6819 = n6818 ^ n6814 ;
  assign n6820 = n6812 & n6819 ;
  assign n6803 = n6534 ^ n6500 ;
  assign n6799 = n6667 ^ n183 ;
  assign n6800 = ~n138 & n6799 ;
  assign n6801 = n6667 & n6800 ;
  assign n6802 = n6801 ^ n6799 ;
  assign n6804 = n6803 ^ n6802 ;
  assign n6809 = ~n183 & n6667 ;
  assign n6810 = n6809 ^ n6534 ;
  assign n6811 = ~n6804 & n6810 ;
  assign n6821 = n6820 ^ n6811 ;
  assign n6822 = n6531 & ~n6821 ;
  assign n6823 = n6802 ^ n4971 ;
  assign n6824 = n6802 ^ n6534 ;
  assign n6825 = n6824 ^ n6802 ;
  assign n6826 = ~n6823 & ~n6825 ;
  assign n6827 = n6826 ^ n6802 ;
  assign n6828 = n6822 & n6827 ;
  assign n6829 = n6828 ^ n6821 ;
  assign n6830 = ~n6660 & ~n6673 ;
  assign n6831 = n6830 ^ n6536 ;
  assign n6832 = n6831 ^ n157 ;
  assign n6940 = ~n6656 & ~n6673 ;
  assign n6941 = n6940 ^ n6538 ;
  assign n6833 = n6648 & ~n6673 ;
  assign n6834 = n6833 ^ n6651 ;
  assign n6835 = n6834 ^ n291 ;
  assign n6836 = n6644 ^ n401 ;
  assign n6837 = ~n6673 & n6836 ;
  assign n6838 = n6837 ^ n6544 ;
  assign n6839 = n6838 ^ n341 ;
  assign n6925 = ~n6642 & ~n6673 ;
  assign n6926 = n6925 ^ n6547 ;
  assign n6840 = ~n6637 & ~n6673 ;
  assign n6841 = n6840 ^ n6639 ;
  assign n6842 = n6841 ^ n457 ;
  assign n6843 = ~n6635 & ~n6673 ;
  assign n6844 = n6843 ^ n6550 ;
  assign n6845 = n6844 ^ n534 ;
  assign n6846 = n6629 & ~n6673 ;
  assign n6847 = n6846 ^ n6631 ;
  assign n6848 = n6847 ^ n609 ;
  assign n6888 = ~n6602 & ~n6673 ;
  assign n6889 = n6888 ^ n6604 ;
  assign n6866 = n6583 ^ n1739 ;
  assign n6867 = n6866 ^ n2064 ;
  assign n6868 = n6559 ^ n1739 ;
  assign n6869 = n6868 ^ n2064 ;
  assign n6870 = n6867 & ~n6869 ;
  assign n6871 = n6870 ^ n2064 ;
  assign n6872 = ~n6673 & ~n6871 ;
  assign n6873 = n6872 ^ n6556 ;
  assign n6876 = n6873 ^ n1427 ;
  assign n6849 = n6572 & ~n6673 ;
  assign n6850 = n6849 ^ n6575 ;
  assign n6851 = n6850 ^ n2175 ;
  assign n6852 = n6798 & ~n6851 ;
  assign n6853 = n6852 ^ n2204 ;
  assign n6854 = n6578 & ~n6673 ;
  assign n6855 = n6854 ^ n6580 ;
  assign n6856 = n6855 ^ n2008 ;
  assign n6857 = n6853 & ~n6856 ;
  assign n6858 = n6857 ^ n2008 ;
  assign n6859 = n6858 ^ n1739 ;
  assign n6860 = n6583 ^ n2008 ;
  assign n6861 = ~n6673 & n6860 ;
  assign n6862 = n6861 ^ n6559 ;
  assign n6863 = n6862 ^ n6858 ;
  assign n6864 = ~n6859 & n6863 ;
  assign n6865 = n6864 ^ n1763 ;
  assign n6874 = n6873 ^ n1572 ;
  assign n6875 = n6865 & n6874 ;
  assign n6877 = n6876 ^ n6875 ;
  assign n6878 = ~n6591 & ~n6673 ;
  assign n6879 = n6878 ^ n6593 ;
  assign n6880 = n6879 ^ n1427 ;
  assign n6881 = ~n6877 & ~n6880 ;
  assign n6882 = n6881 ^ n1450 ;
  assign n6883 = ~n6597 & ~n6673 ;
  assign n6884 = n6883 ^ n6599 ;
  assign n6885 = n6884 ^ n1290 ;
  assign n6886 = n6882 & n6885 ;
  assign n6887 = n6886 ^ n6884 ;
  assign n6890 = n6889 ^ n6887 ;
  assign n6891 = n6889 ^ n1136 ;
  assign n6892 = ~n6890 & n6891 ;
  assign n6893 = n6892 ^ n1143 ;
  assign n6894 = n6608 & ~n6673 ;
  assign n6895 = n6894 ^ n6553 ;
  assign n6898 = n6895 ^ n1034 ;
  assign n6899 = ~n6893 & n6898 ;
  assign n6896 = n6895 ^ n892 ;
  assign n6900 = n6899 ^ n6896 ;
  assign n6901 = n6610 & ~n6673 ;
  assign n6902 = n6901 ^ n6612 ;
  assign n6903 = n6902 ^ n786 ;
  assign n6904 = n6903 ^ n927 ;
  assign n6905 = ~n6900 & n6904 ;
  assign n6906 = n6905 ^ n6903 ;
  assign n6907 = n6617 & ~n6673 ;
  assign n6908 = n6907 ^ n6619 ;
  assign n6909 = n6908 ^ n696 ;
  assign n6910 = n6909 ^ n842 ;
  assign n6911 = ~n6906 & n6910 ;
  assign n6912 = n6911 ^ n6909 ;
  assign n6913 = n6623 & ~n6673 ;
  assign n6914 = n6913 ^ n6625 ;
  assign n6915 = n6914 ^ n609 ;
  assign n6916 = n6915 ^ n835 ;
  assign n6917 = ~n6912 & n6916 ;
  assign n6918 = n6917 ^ n6915 ;
  assign n6919 = ~n6848 & ~n6918 ;
  assign n6920 = n6919 ^ n834 ;
  assign n6921 = n6845 & ~n6920 ;
  assign n6922 = n6921 ^ n750 ;
  assign n6923 = ~n6842 & n6922 ;
  assign n6924 = n6923 ^ n6841 ;
  assign n6927 = n6926 ^ n6924 ;
  assign n6928 = n6926 ^ n401 ;
  assign n6929 = ~n6927 & n6928 ;
  assign n6930 = n6929 ^ n462 ;
  assign n6931 = n6839 & n6930 ;
  assign n6932 = n6931 ^ n349 ;
  assign n6933 = n6835 & ~n6932 ;
  assign n6934 = n6933 ^ n307 ;
  assign n6935 = ~n6654 & ~n6673 ;
  assign n6936 = n6935 ^ n6541 ;
  assign n6937 = n6936 ^ n245 ;
  assign n6938 = n6934 & n6937 ;
  assign n6939 = n6938 ^ n6936 ;
  assign n6942 = n6941 ^ n6939 ;
  assign n6943 = n6941 ^ n188 ;
  assign n6944 = n6942 & ~n6943 ;
  assign n6945 = n6944 ^ n203 ;
  assign n6946 = ~n6832 & ~n6945 ;
  assign n6947 = n6946 ^ n6831 ;
  assign n6948 = n6947 ^ n138 ;
  assign n6949 = n6662 & ~n6673 ;
  assign n6950 = n6949 ^ n6664 ;
  assign n6951 = n6950 ^ n6947 ;
  assign n6952 = ~n6948 & ~n6951 ;
  assign n6953 = n6952 ^ n138 ;
  assign n6954 = ~n6668 & ~n6673 ;
  assign n6955 = n6954 ^ n6533 ;
  assign n6956 = n183 & ~n6955 ;
  assign n6957 = n6953 & ~n6956 ;
  assign n6958 = n6829 & n6957 ;
  assign n6959 = n6958 ^ n6829 ;
  assign n6960 = n6798 & ~n6959 ;
  assign n6961 = n6960 ^ n6850 ;
  assign n6962 = n6961 ^ n2008 ;
  assign n6963 = n6792 & ~n6959 ;
  assign n6964 = n6963 ^ n6795 ;
  assign n6965 = n6964 ^ n2175 ;
  assign n6966 = n6789 ^ n2511 ;
  assign n6967 = ~n6959 & ~n6966 ;
  assign n6968 = n6967 ^ n6675 ;
  assign n6969 = n6968 ^ n2366 ;
  assign n7092 = ~n6787 & ~n6959 ;
  assign n7093 = n7092 ^ n6678 ;
  assign n7085 = n6781 ^ n2894 ;
  assign n7086 = ~n6959 & ~n7085 ;
  assign n7087 = n7086 ^ n6783 ;
  assign n6970 = ~n6779 & ~n6959 ;
  assign n6971 = n6970 ^ n6681 ;
  assign n6972 = n6971 ^ n2894 ;
  assign n7077 = n6774 & ~n6959 ;
  assign n7078 = n7077 ^ n6776 ;
  assign n7081 = n7078 ^ n2894 ;
  assign n6973 = n6759 ^ n3908 ;
  assign n6974 = ~n6959 & n6973 ;
  assign n6975 = n6974 ^ n6761 ;
  assign n6976 = n6975 ^ n3722 ;
  assign n7058 = n6753 ^ n4153 ;
  assign n7059 = ~n6959 & n7058 ;
  assign n7060 = n7059 ^ n6755 ;
  assign n6977 = n6746 & ~n6959 ;
  assign n6978 = n6977 ^ n6748 ;
  assign n6979 = n6978 ^ n4356 ;
  assign n6980 = n6741 & ~n6959 ;
  assign n6981 = n6980 ^ n6694 ;
  assign n6982 = n6981 ^ n4812 ;
  assign n6983 = n6739 & ~n6959 ;
  assign n6984 = n6983 ^ n6698 ;
  assign n6985 = n6984 ^ n5073 ;
  assign n6986 = n6733 ^ n5562 ;
  assign n6987 = ~n6959 & n6986 ;
  assign n6988 = n6987 ^ n6735 ;
  assign n7040 = n6988 ^ n5073 ;
  assign n6989 = n6988 ^ n5317 ;
  assign n7033 = n6731 & ~n6959 ;
  assign n7034 = n7033 ^ n6708 ;
  assign n6990 = ~n6727 & ~n6959 ;
  assign n6991 = n6990 ^ n6728 ;
  assign n6992 = n6991 ^ n5830 ;
  assign n6993 = n6711 ^ n6673 ;
  assign n7005 = ~n6959 & ~n6993 ;
  assign n7004 = n6673 ^ x44 ;
  assign n7006 = n7005 ^ n7004 ;
  assign n7007 = n7006 ^ n6389 ;
  assign n7011 = n6959 ^ n6673 ;
  assign n7009 = n6673 ^ x43 ;
  assign n7010 = n7009 ^ x42 ;
  assign n7012 = n7011 ^ n7010 ;
  assign n7008 = ~x40 & ~x41 ;
  assign n7013 = n7012 ^ n7008 ;
  assign n7014 = n7011 ^ x43 ;
  assign n7015 = ~n7013 & ~n7014 ;
  assign n7023 = n7015 ^ n6713 ;
  assign n7016 = n7015 ^ n7011 ;
  assign n7017 = n7016 ^ n7015 ;
  assign n7018 = n7015 ^ n7012 ;
  assign n7019 = n7018 ^ n7015 ;
  assign n7020 = n7017 & n7019 ;
  assign n7021 = n7020 ^ n7015 ;
  assign n7022 = x42 & n7021 ;
  assign n7024 = n7023 ^ n7022 ;
  assign n7025 = n7007 & ~n7024 ;
  assign n7026 = n7025 ^ n6389 ;
  assign n7002 = ~x44 & ~n6673 ;
  assign n6996 = n6713 ^ x44 ;
  assign n6997 = n6996 ^ n6713 ;
  assign n6998 = ~n6993 & ~n6997 ;
  assign n6999 = n6998 ^ n6713 ;
  assign n7000 = ~n6959 & ~n6999 ;
  assign n7001 = n7000 ^ x45 ;
  assign n7003 = n7002 ^ n7001 ;
  assign n7027 = n7026 ^ n7003 ;
  assign n7028 = n7026 ^ n6115 ;
  assign n7029 = n7027 & ~n7028 ;
  assign n7030 = n7029 ^ n6429 ;
  assign n7031 = n6992 & ~n7030 ;
  assign n7032 = n7031 ^ n6991 ;
  assign n7035 = n7034 ^ n7032 ;
  assign n7036 = n7034 ^ n5562 ;
  assign n7037 = ~n7035 & n7036 ;
  assign n7038 = n7037 ^ n5885 ;
  assign n7039 = ~n6989 & ~n7038 ;
  assign n7041 = n7040 ^ n7039 ;
  assign n7042 = n6985 & ~n7041 ;
  assign n7043 = n7042 ^ n5115 ;
  assign n7044 = ~n6982 & n7043 ;
  assign n7045 = n7044 ^ n4854 ;
  assign n7046 = n6743 & ~n6959 ;
  assign n7047 = n7046 ^ n6691 ;
  assign n7048 = n7047 ^ n4583 ;
  assign n7049 = n7045 & n7048 ;
  assign n7050 = n7049 ^ n4645 ;
  assign n7051 = ~n6979 & n7050 ;
  assign n7052 = n7051 ^ n4414 ;
  assign n7053 = n6751 & ~n6959 ;
  assign n7054 = n7053 ^ n6688 ;
  assign n7055 = n7054 ^ n4153 ;
  assign n7056 = n7052 & n7055 ;
  assign n7057 = n7056 ^ n4153 ;
  assign n7061 = n7060 ^ n7057 ;
  assign n7062 = n7060 ^ n3908 ;
  assign n7063 = ~n7061 & n7062 ;
  assign n7064 = n7063 ^ n3961 ;
  assign n7065 = ~n6976 & ~n7064 ;
  assign n7066 = n7065 ^ n3795 ;
  assign n7067 = ~n6766 & ~n6959 ;
  assign n7068 = n7067 ^ n6769 ;
  assign n7069 = n7068 ^ n3538 ;
  assign n7070 = n7066 & n7069 ;
  assign n7071 = n7070 ^ n3596 ;
  assign n7072 = n6772 & ~n6959 ;
  assign n7073 = n7072 ^ n6685 ;
  assign n7074 = n7073 ^ n3320 ;
  assign n7075 = n7071 & ~n7074 ;
  assign n7076 = n7075 ^ n3387 ;
  assign n7079 = n7078 ^ n3093 ;
  assign n7080 = n7076 & ~n7079 ;
  assign n7082 = n7081 ^ n7080 ;
  assign n7083 = ~n6972 & ~n7082 ;
  assign n7084 = n7083 ^ n2894 ;
  assign n7088 = n7087 ^ n7084 ;
  assign n7089 = n7087 ^ n2707 ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = n7090 ^ n2707 ;
  assign n7094 = n7093 ^ n7091 ;
  assign n7095 = n7093 ^ n2511 ;
  assign n7096 = n7094 & n7095 ;
  assign n7097 = n7096 ^ n2530 ;
  assign n7098 = n6969 & n7097 ;
  assign n7099 = n7098 ^ n2399 ;
  assign n7100 = ~n6965 & n7099 ;
  assign n7101 = n7100 ^ n2204 ;
  assign n7102 = ~n6962 & n7101 ;
  assign n7103 = n7102 ^ n2064 ;
  assign n7104 = n6853 & ~n6959 ;
  assign n7105 = n7104 ^ n6855 ;
  assign n7106 = n7105 ^ n1739 ;
  assign n7107 = ~n7103 & n7106 ;
  assign n7108 = n7107 ^ n1763 ;
  assign n7196 = ~n6859 & ~n6959 ;
  assign n7197 = n7196 ^ n6862 ;
  assign n7198 = n7197 ^ n1572 ;
  assign n7199 = ~n7108 & ~n7198 ;
  assign n7200 = n7199 ^ n1605 ;
  assign n7201 = ~n6865 & ~n6959 ;
  assign n7202 = n7201 ^ n6873 ;
  assign n7203 = n7202 ^ n1427 ;
  assign n7204 = ~n7200 & ~n7203 ;
  assign n7205 = n7204 ^ n1450 ;
  assign n7109 = ~n6948 & n6950 ;
  assign n7152 = ~n4970 & ~n6956 ;
  assign n7156 = n7152 ^ n6829 ;
  assign n7157 = n7156 ^ n7152 ;
  assign n7160 = ~n6955 & ~n7157 ;
  assign n7161 = n7160 ^ n7152 ;
  assign n7162 = n6953 & n7161 ;
  assign n7110 = n6948 ^ n6829 ;
  assign n7111 = n6955 ^ n6950 ;
  assign n7112 = n7111 ^ n138 ;
  assign n7113 = n7112 ^ n6947 ;
  assign n7114 = n7113 ^ n6829 ;
  assign n7143 = n7114 ^ n6955 ;
  assign n7144 = ~n7110 & ~n7143 ;
  assign n7145 = n7144 ^ n6829 ;
  assign n7146 = n6955 ^ n138 ;
  assign n7147 = n7144 ^ n7143 ;
  assign n7148 = n7146 & ~n7147 ;
  assign n7149 = n7148 ^ n6955 ;
  assign n7150 = ~n7145 & ~n7149 ;
  assign n7151 = n7150 ^ n6955 ;
  assign n7153 = n7152 ^ n7151 ;
  assign n7154 = n7153 ^ n7152 ;
  assign n7163 = n7162 ^ n7154 ;
  assign n7164 = n183 & ~n7163 ;
  assign n7165 = n7164 ^ n7153 ;
  assign n7166 = n6955 & n7165 ;
  assign n7167 = n7109 & n7166 ;
  assign n7168 = n7167 ^ n7165 ;
  assign n7169 = ~n6934 & ~n6959 ;
  assign n7170 = n7169 ^ n6936 ;
  assign n7171 = n7170 ^ n188 ;
  assign n7172 = ~n6932 & ~n6959 ;
  assign n7173 = n7172 ^ n6834 ;
  assign n7174 = n7173 ^ n245 ;
  assign n7175 = n6930 & ~n6959 ;
  assign n7176 = n7175 ^ n6838 ;
  assign n7177 = n7176 ^ n291 ;
  assign n7181 = ~n6922 & ~n6959 ;
  assign n7182 = n7181 ^ n6841 ;
  assign n7183 = n7182 ^ n401 ;
  assign n7184 = ~n6920 & ~n6959 ;
  assign n7185 = n7184 ^ n6844 ;
  assign n7186 = n7185 ^ n457 ;
  assign n7187 = ~n6918 & ~n6959 ;
  assign n7188 = n7187 ^ n6847 ;
  assign n7189 = n7188 ^ n534 ;
  assign n7190 = n6912 & ~n6959 ;
  assign n7191 = n7190 ^ n6914 ;
  assign n7192 = n7191 ^ n609 ;
  assign n7193 = ~n6882 & ~n6959 ;
  assign n7194 = n7193 ^ n6884 ;
  assign n7195 = n7194 ^ n1136 ;
  assign n7206 = ~n6877 & ~n6959 ;
  assign n7207 = n7206 ^ n6879 ;
  assign n7210 = n7207 ^ n1136 ;
  assign n7208 = n7207 ^ n1290 ;
  assign n7209 = n7205 & n7208 ;
  assign n7211 = n7210 ^ n7209 ;
  assign n7212 = n7195 & n7211 ;
  assign n7213 = n7212 ^ n1143 ;
  assign n7214 = n6887 ^ n1136 ;
  assign n7215 = ~n6959 & n7214 ;
  assign n7216 = n7215 ^ n6889 ;
  assign n7219 = n7216 ^ n1034 ;
  assign n7220 = ~n7213 & n7219 ;
  assign n7217 = n7216 ^ n892 ;
  assign n7221 = n7220 ^ n7217 ;
  assign n7222 = n6893 & ~n6959 ;
  assign n7223 = n7222 ^ n6895 ;
  assign n7224 = n7223 ^ n786 ;
  assign n7225 = n7224 ^ n927 ;
  assign n7226 = ~n7221 & n7225 ;
  assign n7227 = n7226 ^ n7224 ;
  assign n7228 = n6900 & ~n6959 ;
  assign n7229 = n7228 ^ n6902 ;
  assign n7230 = n7229 ^ n696 ;
  assign n7231 = n7230 ^ n842 ;
  assign n7232 = ~n7227 & n7231 ;
  assign n7233 = n7232 ^ n7230 ;
  assign n7234 = n6906 & ~n6959 ;
  assign n7235 = n7234 ^ n6908 ;
  assign n7236 = n7235 ^ n609 ;
  assign n7237 = n7236 ^ n835 ;
  assign n7238 = ~n7233 & n7237 ;
  assign n7239 = n7238 ^ n7236 ;
  assign n7240 = ~n7192 & ~n7239 ;
  assign n7241 = n7240 ^ n834 ;
  assign n7242 = n7189 & ~n7241 ;
  assign n7243 = n7242 ^ n750 ;
  assign n7244 = ~n7186 & n7243 ;
  assign n7245 = n7244 ^ n7185 ;
  assign n7246 = n7245 ^ n7182 ;
  assign n7247 = n7183 & ~n7246 ;
  assign n7248 = n7247 ^ n401 ;
  assign n7178 = n6924 ^ n401 ;
  assign n7179 = ~n6959 & n7178 ;
  assign n7180 = n7179 ^ n6926 ;
  assign n7249 = n7248 ^ n7180 ;
  assign n7250 = n7248 ^ n341 ;
  assign n7251 = ~n7249 & n7250 ;
  assign n7252 = n7251 ^ n349 ;
  assign n7253 = ~n7177 & ~n7252 ;
  assign n7254 = n7253 ^ n307 ;
  assign n7255 = ~n7174 & n7254 ;
  assign n7256 = n7255 ^ n7173 ;
  assign n7257 = n7256 ^ n7170 ;
  assign n7258 = n7171 & n7257 ;
  assign n7259 = n7258 ^ n203 ;
  assign n7260 = n6939 ^ n188 ;
  assign n7261 = ~n6959 & n7260 ;
  assign n7262 = n7261 ^ n6941 ;
  assign n7263 = n7262 ^ n157 ;
  assign n7264 = ~n7259 & ~n7263 ;
  assign n7265 = n7264 ^ n7262 ;
  assign n7266 = n7265 ^ n138 ;
  assign n7267 = n6945 & ~n6959 ;
  assign n7268 = n7267 ^ n6831 ;
  assign n7269 = n7268 ^ n7265 ;
  assign n7270 = ~n7266 & ~n7269 ;
  assign n7271 = n7270 ^ n138 ;
  assign n7272 = n7168 & n7271 ;
  assign n7273 = ~n6948 & ~n6959 ;
  assign n7274 = n7273 ^ n6950 ;
  assign n7275 = n7274 ^ n183 ;
  assign n7276 = n7272 & n7275 ;
  assign n7277 = n7276 ^ n7168 ;
  assign n7460 = ~n7205 & ~n7277 ;
  assign n7461 = n7460 ^ n7207 ;
  assign n7278 = ~n7108 & ~n7277 ;
  assign n7279 = n7278 ^ n7197 ;
  assign n7280 = n7279 ^ n1427 ;
  assign n7281 = n7099 & ~n7277 ;
  assign n7282 = n7281 ^ n6964 ;
  assign n7283 = n7282 ^ n2008 ;
  assign n7284 = n7097 & ~n7277 ;
  assign n7285 = n7284 ^ n6968 ;
  assign n7286 = n7285 ^ n2175 ;
  assign n7287 = n7091 ^ n2511 ;
  assign n7288 = ~n7277 & ~n7287 ;
  assign n7289 = n7288 ^ n7093 ;
  assign n7290 = n7289 ^ n2366 ;
  assign n7430 = n7084 ^ n2707 ;
  assign n7431 = ~n7277 & ~n7430 ;
  assign n7432 = n7431 ^ n7087 ;
  assign n7291 = ~n7082 & ~n7277 ;
  assign n7292 = n7291 ^ n6971 ;
  assign n7293 = n7292 ^ n2707 ;
  assign n7294 = ~n7076 & ~n7277 ;
  assign n7295 = n7294 ^ n7078 ;
  assign n7296 = n7295 ^ n2894 ;
  assign n7420 = n7071 & ~n7277 ;
  assign n7421 = n7420 ^ n7073 ;
  assign n7424 = n7421 ^ n2894 ;
  assign n7297 = ~n7064 & ~n7277 ;
  assign n7298 = n7297 ^ n6975 ;
  assign n7299 = n7298 ^ n3538 ;
  assign n7300 = n7057 ^ n3908 ;
  assign n7301 = ~n7277 & n7300 ;
  assign n7302 = n7301 ^ n7060 ;
  assign n7303 = n7302 ^ n3722 ;
  assign n7310 = n7045 & ~n7277 ;
  assign n7311 = n7310 ^ n7047 ;
  assign n7312 = n7311 ^ n4356 ;
  assign n7313 = ~n7041 & ~n7277 ;
  assign n7314 = n7313 ^ n6984 ;
  assign n7315 = n7314 ^ n4812 ;
  assign n7316 = n7038 & ~n7277 ;
  assign n7317 = n7316 ^ n6988 ;
  assign n7318 = n7317 ^ n5073 ;
  assign n7323 = ~n7028 & ~n7277 ;
  assign n7324 = n7323 ^ n7003 ;
  assign n7379 = n7324 ^ n5562 ;
  assign n7325 = n7324 ^ n5830 ;
  assign n7326 = ~n7024 & ~n7277 ;
  assign n7327 = n7326 ^ n7006 ;
  assign n7328 = n7327 ^ n6115 ;
  assign n7356 = n6959 ^ x42 ;
  assign n7339 = n7277 ^ n6959 ;
  assign n7347 = ~x38 & ~x39 ;
  assign n7358 = ~x40 & n7347 ;
  assign n7361 = n7358 ^ n7277 ;
  assign n7362 = ~n7339 & n7361 ;
  assign n7359 = n7358 ^ n7339 ;
  assign n7360 = x41 & n7359 ;
  assign n7363 = n7362 ^ n7360 ;
  assign n7364 = ~n7356 & n7363 ;
  assign n7335 = ~x42 & ~n7277 ;
  assign n7336 = n7008 & n7335 ;
  assign n7365 = n7364 ^ n7336 ;
  assign n7354 = n7008 ^ n6959 ;
  assign n7355 = ~n7277 & ~n7354 ;
  assign n7357 = n7356 ^ n7355 ;
  assign n7366 = n7365 ^ n7357 ;
  assign n7341 = n6959 ^ x41 ;
  assign n7340 = n7339 ^ x40 ;
  assign n7342 = n7341 ^ n7340 ;
  assign n7343 = n7342 ^ n7339 ;
  assign n7344 = n7343 ^ n7341 ;
  assign n7346 = n7341 ^ n7277 ;
  assign n7348 = n7347 ^ n7342 ;
  assign n7349 = ~n7346 & ~n7348 ;
  assign n7345 = n7341 & n7342 ;
  assign n7350 = n7349 ^ n7345 ;
  assign n7351 = ~n7344 & n7350 ;
  assign n7352 = n7351 ^ n7345 ;
  assign n7353 = n7352 ^ n6959 ;
  assign n7367 = n7366 ^ n7353 ;
  assign n7368 = ~n6673 & ~n7367 ;
  assign n7369 = n7357 ^ n7353 ;
  assign n7370 = n7368 & ~n7369 ;
  assign n7371 = n7370 ^ n7367 ;
  assign n7337 = n7336 ^ n7014 ;
  assign n7329 = n6673 ^ x42 ;
  assign n7330 = n7329 ^ n6673 ;
  assign n7332 = ~n6959 & n7330 ;
  assign n7333 = n7332 ^ n6673 ;
  assign n7334 = n7277 & ~n7333 ;
  assign n7338 = n7337 ^ n7334 ;
  assign n7372 = n7371 ^ n7338 ;
  assign n7373 = n7371 ^ n6389 ;
  assign n7374 = n7372 & n7373 ;
  assign n7375 = n7374 ^ n6423 ;
  assign n7376 = ~n7328 & ~n7375 ;
  assign n7377 = n7376 ^ n6429 ;
  assign n7378 = n7325 & ~n7377 ;
  assign n7380 = n7379 ^ n7378 ;
  assign n7381 = n7030 & ~n7277 ;
  assign n7382 = n7381 ^ n6991 ;
  assign n7383 = n7382 ^ n5562 ;
  assign n7384 = n7380 & n7383 ;
  assign n7385 = n7384 ^ n5885 ;
  assign n7319 = n7032 ^ n5562 ;
  assign n7320 = ~n7277 & n7319 ;
  assign n7321 = n7320 ^ n7034 ;
  assign n7386 = n7321 ^ n5317 ;
  assign n7387 = ~n7385 & n7386 ;
  assign n7322 = n7321 ^ n5073 ;
  assign n7388 = n7387 ^ n7322 ;
  assign n7389 = ~n7318 & n7388 ;
  assign n7390 = n7389 ^ n5115 ;
  assign n7391 = n7315 & n7390 ;
  assign n7392 = n7391 ^ n4854 ;
  assign n7393 = n7043 & ~n7277 ;
  assign n7394 = n7393 ^ n6981 ;
  assign n7395 = n7394 ^ n4583 ;
  assign n7396 = n7392 & ~n7395 ;
  assign n7397 = n7396 ^ n4645 ;
  assign n7398 = n7312 & ~n7397 ;
  assign n7399 = n7398 ^ n7311 ;
  assign n7308 = n7050 & ~n7277 ;
  assign n7309 = n7308 ^ n6978 ;
  assign n7400 = n7399 ^ n7309 ;
  assign n7401 = n7399 ^ n4153 ;
  assign n7402 = n7400 & n7401 ;
  assign n7403 = n7402 ^ n4153 ;
  assign n7306 = n7302 ^ n3908 ;
  assign n7304 = n7052 & ~n7277 ;
  assign n7305 = n7304 ^ n7054 ;
  assign n7307 = n7306 ^ n7305 ;
  assign n7404 = n7403 ^ n7307 ;
  assign n7405 = n7404 ^ n7306 ;
  assign n7406 = n7305 ^ n7302 ;
  assign n7407 = n7406 ^ n7306 ;
  assign n7408 = ~n7405 & n7407 ;
  assign n7409 = n7408 ^ n7306 ;
  assign n7410 = ~n7303 & ~n7409 ;
  assign n7411 = n7410 ^ n3795 ;
  assign n7412 = ~n7299 & n7411 ;
  assign n7413 = n7412 ^ n3538 ;
  assign n7414 = n7413 ^ n3320 ;
  assign n7415 = n7066 & ~n7277 ;
  assign n7416 = n7415 ^ n7068 ;
  assign n7417 = n7416 ^ n7413 ;
  assign n7418 = n7414 & ~n7417 ;
  assign n7419 = n7418 ^ n3387 ;
  assign n7422 = n7421 ^ n3093 ;
  assign n7423 = n7419 & n7422 ;
  assign n7425 = n7424 ^ n7423 ;
  assign n7426 = ~n7296 & n7425 ;
  assign n7427 = n7426 ^ n3396 ;
  assign n7428 = n7293 & ~n7427 ;
  assign n7429 = n7428 ^ n2707 ;
  assign n7433 = n7432 ^ n7429 ;
  assign n7434 = n7432 ^ n2511 ;
  assign n7435 = n7433 & n7434 ;
  assign n7436 = n7435 ^ n2530 ;
  assign n7437 = n7290 & n7436 ;
  assign n7438 = n7437 ^ n2399 ;
  assign n7439 = n7286 & n7438 ;
  assign n7440 = n7439 ^ n2204 ;
  assign n7441 = ~n7283 & n7440 ;
  assign n7442 = n7441 ^ n2064 ;
  assign n7443 = n7101 & ~n7277 ;
  assign n7444 = n7443 ^ n6961 ;
  assign n7445 = n7444 ^ n1739 ;
  assign n7446 = ~n7442 & n7445 ;
  assign n7447 = n7446 ^ n1763 ;
  assign n7448 = ~n7103 & ~n7277 ;
  assign n7449 = n7448 ^ n7105 ;
  assign n7450 = n7449 ^ n1572 ;
  assign n7451 = ~n7447 & ~n7450 ;
  assign n7452 = n7451 ^ n1605 ;
  assign n7453 = n7280 & ~n7452 ;
  assign n7454 = n7453 ^ n1450 ;
  assign n7455 = ~n7200 & ~n7277 ;
  assign n7456 = n7455 ^ n7202 ;
  assign n7457 = n7456 ^ n1290 ;
  assign n7458 = n7454 & n7457 ;
  assign n7459 = n7458 ^ n7456 ;
  assign n7462 = n7461 ^ n7459 ;
  assign n7463 = n7461 ^ n1136 ;
  assign n7464 = ~n7462 & n7463 ;
  assign n7465 = n7464 ^ n1143 ;
  assign n7466 = n7211 & ~n7277 ;
  assign n7467 = n7466 ^ n7194 ;
  assign n7470 = n7467 ^ n1034 ;
  assign n7471 = ~n7465 & n7470 ;
  assign n7468 = n7467 ^ n892 ;
  assign n7472 = n7471 ^ n7468 ;
  assign n7473 = n7213 & ~n7277 ;
  assign n7474 = n7473 ^ n7216 ;
  assign n7475 = n7474 ^ n786 ;
  assign n7476 = n7475 ^ n927 ;
  assign n7477 = ~n7472 & n7476 ;
  assign n7478 = n7477 ^ n7475 ;
  assign n7479 = n7221 & ~n7277 ;
  assign n7480 = n7479 ^ n7223 ;
  assign n7481 = n7480 ^ n696 ;
  assign n7482 = n7481 ^ n842 ;
  assign n7483 = ~n7478 & n7482 ;
  assign n7484 = n7483 ^ n7481 ;
  assign n7486 = ~n7272 & n7274 ;
  assign n7487 = n7486 ^ n7271 ;
  assign n7485 = n7274 ^ n7271 ;
  assign n7488 = n7487 ^ n7485 ;
  assign n7489 = n7487 ^ n7268 ;
  assign n7490 = n7489 ^ n7487 ;
  assign n7491 = n7488 & n7490 ;
  assign n7492 = n7491 ^ n7487 ;
  assign n7493 = ~n138 & n7268 ;
  assign n7494 = ~n7168 & n7493 ;
  assign n7495 = n7494 ^ n7274 ;
  assign n7496 = n7265 ^ n130 ;
  assign n7497 = n7496 ^ n7268 ;
  assign n7498 = n7497 ^ n7168 ;
  assign n7499 = ~n183 & n7498 ;
  assign n7500 = n7499 ^ n7168 ;
  assign n7501 = n7500 ^ n183 ;
  assign n7502 = n7500 ^ n7168 ;
  assign n7503 = n7502 ^ n7500 ;
  assign n7504 = n7500 ^ n7268 ;
  assign n7505 = n7503 & n7504 ;
  assign n7506 = ~n7501 & n7505 ;
  assign n7507 = n7506 ^ n7501 ;
  assign n7508 = n7507 ^ n183 ;
  assign n7509 = n7495 & n7508 ;
  assign n7510 = n183 & ~n7509 ;
  assign n7511 = n7492 & n7510 ;
  assign n7512 = n7511 ^ n7509 ;
  assign n7515 = n7256 ^ n188 ;
  assign n7516 = ~n7277 & ~n7515 ;
  assign n7517 = n7516 ^ n7170 ;
  assign n7518 = n7517 ^ n157 ;
  assign n7563 = ~n7254 & ~n7277 ;
  assign n7564 = n7563 ^ n7173 ;
  assign n7519 = ~n7252 & ~n7277 ;
  assign n7520 = n7519 ^ n7176 ;
  assign n7521 = n7520 ^ n245 ;
  assign n7522 = n7245 ^ n401 ;
  assign n7523 = ~n7277 & n7522 ;
  assign n7524 = n7523 ^ n7182 ;
  assign n7525 = n7524 ^ n341 ;
  assign n7548 = ~n7243 & ~n7277 ;
  assign n7549 = n7548 ^ n7185 ;
  assign n7526 = ~n7241 & ~n7277 ;
  assign n7527 = n7526 ^ n7188 ;
  assign n7528 = n7527 ^ n457 ;
  assign n7529 = ~n7239 & ~n7277 ;
  assign n7530 = n7529 ^ n7191 ;
  assign n7531 = n7530 ^ n534 ;
  assign n7532 = n7233 & ~n7277 ;
  assign n7533 = n7532 ^ n7235 ;
  assign n7542 = n7533 ^ n534 ;
  assign n7534 = n7533 ^ n609 ;
  assign n7535 = n7227 & ~n7277 ;
  assign n7536 = n7535 ^ n7229 ;
  assign n7537 = n7536 ^ n609 ;
  assign n7538 = n7537 ^ n835 ;
  assign n7539 = ~n7484 & n7538 ;
  assign n7540 = n7539 ^ n7537 ;
  assign n7541 = ~n7534 & n7540 ;
  assign n7543 = n7542 ^ n7541 ;
  assign n7544 = n7531 & n7543 ;
  assign n7545 = n7544 ^ n750 ;
  assign n7546 = ~n7528 & n7545 ;
  assign n7547 = n7546 ^ n7527 ;
  assign n7550 = n7549 ^ n7547 ;
  assign n7551 = n7549 ^ n401 ;
  assign n7552 = ~n7550 & n7551 ;
  assign n7553 = n7552 ^ n462 ;
  assign n7554 = n7525 & n7553 ;
  assign n7555 = n7554 ^ n349 ;
  assign n7556 = n7250 & ~n7277 ;
  assign n7557 = n7556 ^ n7180 ;
  assign n7558 = n7557 ^ n291 ;
  assign n7559 = ~n7555 & ~n7558 ;
  assign n7560 = n7559 ^ n307 ;
  assign n7561 = n7521 & n7560 ;
  assign n7562 = n7561 ^ n7520 ;
  assign n7565 = n7564 ^ n7562 ;
  assign n7566 = n7564 ^ n188 ;
  assign n7567 = n7565 & ~n7566 ;
  assign n7568 = n7567 ^ n203 ;
  assign n7569 = n7518 & ~n7568 ;
  assign n7570 = n7569 ^ n7517 ;
  assign n7571 = n7570 ^ n138 ;
  assign n7572 = n7259 & ~n7277 ;
  assign n7573 = n7572 ^ n7262 ;
  assign n7574 = n7573 ^ n7570 ;
  assign n7575 = n7571 & n7574 ;
  assign n7576 = n7575 ^ n138 ;
  assign n7513 = ~n7266 & ~n7277 ;
  assign n7514 = n7513 ^ n7268 ;
  assign n7577 = n7576 ^ n7514 ;
  assign n7578 = n7577 ^ n7576 ;
  assign n7579 = n183 & n7576 ;
  assign n7582 = n7578 & n7579 ;
  assign n7583 = n7582 ^ n7576 ;
  assign n7584 = n7512 & ~n7583 ;
  assign n7585 = n7484 & ~n7584 ;
  assign n7586 = n7585 ^ n7536 ;
  assign n7587 = n7586 ^ n609 ;
  assign n7759 = ~n7442 & ~n7584 ;
  assign n7760 = n7759 ^ n7444 ;
  assign n7763 = n7760 ^ n1427 ;
  assign n7588 = n7438 & ~n7584 ;
  assign n7589 = n7588 ^ n7285 ;
  assign n7590 = n7589 ^ n2008 ;
  assign n7591 = n7436 & ~n7584 ;
  assign n7592 = n7591 ^ n7289 ;
  assign n7593 = n7592 ^ n2175 ;
  assign n7594 = ~n7427 & ~n7584 ;
  assign n7595 = n7594 ^ n7292 ;
  assign n7596 = n7595 ^ n2511 ;
  assign n7597 = n7425 & ~n7584 ;
  assign n7598 = n7597 ^ n7295 ;
  assign n7599 = n7598 ^ n2707 ;
  assign n7600 = ~n7419 & ~n7584 ;
  assign n7601 = n7600 ^ n7421 ;
  assign n7602 = n7601 ^ n2894 ;
  assign n7605 = n7411 & ~n7584 ;
  assign n7606 = n7605 ^ n7298 ;
  assign n7607 = n7606 ^ n3320 ;
  assign n7608 = n7403 ^ n3722 ;
  assign n7609 = n7608 ^ n3961 ;
  assign n7610 = n7305 ^ n3722 ;
  assign n7611 = n7610 ^ n3961 ;
  assign n7612 = n7609 & n7611 ;
  assign n7613 = n7612 ^ n3961 ;
  assign n7614 = ~n7584 & ~n7613 ;
  assign n7615 = n7614 ^ n7302 ;
  assign n7616 = n7615 ^ n3538 ;
  assign n7617 = n7403 ^ n3908 ;
  assign n7618 = ~n7584 & n7617 ;
  assign n7619 = n7618 ^ n7305 ;
  assign n7620 = n7619 ^ n3722 ;
  assign n7720 = n7401 & ~n7584 ;
  assign n7721 = n7720 ^ n7309 ;
  assign n7621 = n7397 & ~n7584 ;
  assign n7622 = n7621 ^ n7311 ;
  assign n7623 = n7622 ^ n4153 ;
  assign n7712 = n7392 & ~n7584 ;
  assign n7713 = n7712 ^ n7394 ;
  assign n7716 = n7713 ^ n4153 ;
  assign n7706 = n7390 & ~n7584 ;
  assign n7707 = n7706 ^ n7314 ;
  assign n7624 = n7388 & ~n7584 ;
  assign n7625 = n7624 ^ n7317 ;
  assign n7626 = n7625 ^ n4812 ;
  assign n7697 = n7385 & ~n7584 ;
  assign n7698 = n7697 ^ n7321 ;
  assign n7627 = n7380 & ~n7584 ;
  assign n7628 = n7627 ^ n7382 ;
  assign n7629 = n7628 ^ n5317 ;
  assign n7630 = n7377 & ~n7584 ;
  assign n7631 = n7630 ^ n7324 ;
  assign n7632 = n7631 ^ n5562 ;
  assign n7633 = ~n7375 & ~n7584 ;
  assign n7634 = n7633 ^ n7327 ;
  assign n7635 = n7634 ^ n5830 ;
  assign n7640 = n7584 ^ n7338 ;
  assign n7636 = ~n7373 & ~n7584 ;
  assign n7637 = n7365 & n7636 ;
  assign n7638 = n6389 & n7637 ;
  assign n7639 = n7638 ^ n7636 ;
  assign n7641 = n7640 ^ n7639 ;
  assign n7642 = n7641 ^ n6115 ;
  assign n7643 = n7353 ^ n6673 ;
  assign n7644 = ~n7584 & n7643 ;
  assign n7645 = n7644 ^ n7357 ;
  assign n7646 = n7645 ^ n6389 ;
  assign n7676 = n7277 ^ x40 ;
  assign n7674 = n7347 ^ n7277 ;
  assign n7675 = ~n7584 & ~n7674 ;
  assign n7677 = n7676 ^ n7675 ;
  assign n7660 = n7584 ^ n7277 ;
  assign n7658 = n7277 ^ x39 ;
  assign n7659 = n7658 ^ x38 ;
  assign n7661 = n7660 ^ n7659 ;
  assign n7662 = n7661 ^ n7660 ;
  assign n7663 = n7662 ^ n7658 ;
  assign n7665 = x36 & ~x37 ;
  assign n7666 = n7665 ^ x37 ;
  assign n7667 = n7666 ^ n7661 ;
  assign n7668 = n7658 ^ n7584 ;
  assign n7669 = n7667 & ~n7668 ;
  assign n7664 = n7658 & n7660 ;
  assign n7670 = n7669 ^ n7664 ;
  assign n7671 = ~n7663 & n7670 ;
  assign n7672 = n7671 ^ n7664 ;
  assign n7673 = n7672 ^ n7277 ;
  assign n7678 = n7677 ^ n7673 ;
  assign n7679 = n7677 ^ n6959 ;
  assign n7680 = n7678 & ~n7679 ;
  assign n7681 = n7680 ^ n6959 ;
  assign n7655 = n7277 ^ x41 ;
  assign n7647 = n7358 ^ n6959 ;
  assign n7656 = n7655 ^ n7647 ;
  assign n7648 = n7647 ^ x40 ;
  assign n7649 = n7648 ^ n7647 ;
  assign n7650 = n7647 ^ n7277 ;
  assign n7651 = n7650 ^ n7647 ;
  assign n7652 = n7649 & ~n7651 ;
  assign n7653 = n7652 ^ n7647 ;
  assign n7654 = n7584 & ~n7653 ;
  assign n7657 = n7656 ^ n7654 ;
  assign n7682 = n7681 ^ n7657 ;
  assign n7683 = n7681 ^ n6673 ;
  assign n7684 = ~n7682 & n7683 ;
  assign n7685 = n7684 ^ n6713 ;
  assign n7686 = n7646 & ~n7685 ;
  assign n7687 = n7686 ^ n6423 ;
  assign n7688 = ~n7642 & ~n7687 ;
  assign n7689 = n7688 ^ n6429 ;
  assign n7690 = ~n7635 & ~n7689 ;
  assign n7691 = n7690 ^ n7634 ;
  assign n7692 = n7691 ^ n7631 ;
  assign n7693 = n7632 & n7692 ;
  assign n7694 = n7693 ^ n5885 ;
  assign n7695 = n7629 & ~n7694 ;
  assign n7696 = n7695 ^ n7628 ;
  assign n7699 = n7698 ^ n7696 ;
  assign n7700 = n7698 ^ n5073 ;
  assign n7701 = ~n7699 & n7700 ;
  assign n7702 = n7701 ^ n5073 ;
  assign n7703 = n7702 ^ n7625 ;
  assign n7704 = ~n7626 & n7703 ;
  assign n7705 = n7704 ^ n4812 ;
  assign n7708 = n7707 ^ n7705 ;
  assign n7709 = n7707 ^ n4583 ;
  assign n7710 = ~n7708 & n7709 ;
  assign n7711 = n7710 ^ n4645 ;
  assign n7714 = n7713 ^ n4356 ;
  assign n7715 = ~n7711 & ~n7714 ;
  assign n7717 = n7716 ^ n7715 ;
  assign n7718 = n7623 & ~n7717 ;
  assign n7719 = n7718 ^ n4153 ;
  assign n7722 = n7721 ^ n7719 ;
  assign n7723 = n7721 ^ n3908 ;
  assign n7724 = n7722 & ~n7723 ;
  assign n7725 = n7724 ^ n3961 ;
  assign n7726 = ~n7620 & ~n7725 ;
  assign n7727 = n7726 ^ n3795 ;
  assign n7728 = ~n7616 & n7727 ;
  assign n7729 = n7728 ^ n3596 ;
  assign n7730 = ~n7607 & n7729 ;
  assign n7731 = n7730 ^ n3320 ;
  assign n7735 = n7731 ^ n2894 ;
  assign n7603 = n7414 & ~n7584 ;
  assign n7604 = n7603 ^ n7416 ;
  assign n7732 = n7731 ^ n7604 ;
  assign n7733 = n7604 ^ n3093 ;
  assign n7734 = n7732 & n7733 ;
  assign n7736 = n7735 ^ n7734 ;
  assign n7737 = n7602 & ~n7736 ;
  assign n7738 = n7737 ^ n3396 ;
  assign n7739 = n7599 & ~n7738 ;
  assign n7740 = n7739 ^ n2707 ;
  assign n7741 = n7740 ^ n7595 ;
  assign n7742 = ~n7596 & ~n7741 ;
  assign n7743 = n7742 ^ n2530 ;
  assign n7744 = n7429 ^ n2511 ;
  assign n7745 = ~n7584 & ~n7744 ;
  assign n7746 = n7745 ^ n7432 ;
  assign n7747 = n7746 ^ n2366 ;
  assign n7748 = n7743 & n7747 ;
  assign n7749 = n7748 ^ n2399 ;
  assign n7750 = n7593 & n7749 ;
  assign n7751 = n7750 ^ n2204 ;
  assign n7752 = n7590 & n7751 ;
  assign n7753 = n7752 ^ n2064 ;
  assign n7754 = n7440 & ~n7584 ;
  assign n7755 = n7754 ^ n7282 ;
  assign n7756 = n7755 ^ n1739 ;
  assign n7757 = ~n7753 & n7756 ;
  assign n7758 = n7757 ^ n1763 ;
  assign n7761 = n7760 ^ n1572 ;
  assign n7762 = n7758 & ~n7761 ;
  assign n7764 = n7763 ^ n7762 ;
  assign n7765 = ~n7447 & ~n7584 ;
  assign n7766 = n7765 ^ n7449 ;
  assign n7767 = n7766 ^ n1427 ;
  assign n7768 = n7764 & n7767 ;
  assign n7769 = n7768 ^ n1450 ;
  assign n7770 = ~n7452 & ~n7584 ;
  assign n7771 = n7770 ^ n7279 ;
  assign n7772 = n7771 ^ n1290 ;
  assign n7773 = ~n7769 & ~n7772 ;
  assign n7774 = n7773 ^ n1461 ;
  assign n7775 = ~n7454 & ~n7584 ;
  assign n7776 = n7775 ^ n7456 ;
  assign n7777 = n7776 ^ n1136 ;
  assign n7778 = n7774 & n7777 ;
  assign n7779 = n7778 ^ n1143 ;
  assign n7780 = n7459 ^ n1136 ;
  assign n7781 = ~n7584 & n7780 ;
  assign n7782 = n7781 ^ n7461 ;
  assign n7785 = n7782 ^ n1034 ;
  assign n7786 = ~n7779 & n7785 ;
  assign n7783 = n7782 ^ n892 ;
  assign n7787 = n7786 ^ n7783 ;
  assign n7788 = n7465 & ~n7584 ;
  assign n7789 = n7788 ^ n7467 ;
  assign n7790 = n7789 ^ n786 ;
  assign n7791 = n7790 ^ n927 ;
  assign n7792 = ~n7787 & n7791 ;
  assign n7793 = n7792 ^ n7790 ;
  assign n7794 = n7472 & ~n7584 ;
  assign n7795 = n7794 ^ n7474 ;
  assign n7796 = n7795 ^ n696 ;
  assign n7797 = n7796 ^ n842 ;
  assign n7798 = ~n7793 & n7797 ;
  assign n7799 = n7798 ^ n7796 ;
  assign n7800 = n7478 & ~n7584 ;
  assign n7801 = n7800 ^ n7480 ;
  assign n7802 = n7801 ^ n609 ;
  assign n7803 = n7802 ^ n835 ;
  assign n7804 = ~n7799 & n7803 ;
  assign n7805 = n7804 ^ n7802 ;
  assign n7806 = ~n7587 & ~n7805 ;
  assign n7807 = n7806 ^ n834 ;
  assign n7834 = n7568 & ~n7584 ;
  assign n7835 = n7834 ^ n7517 ;
  assign n7836 = ~n138 & ~n7835 ;
  assign n7837 = n7835 ^ n138 ;
  assign n7838 = n7837 ^ n7836 ;
  assign n7839 = n7562 ^ n188 ;
  assign n7840 = ~n7584 & n7839 ;
  assign n7841 = n7840 ^ n7564 ;
  assign n7842 = n7841 ^ n157 ;
  assign n7843 = ~n7555 & ~n7584 ;
  assign n7844 = n7843 ^ n7557 ;
  assign n7845 = n7844 ^ n245 ;
  assign n7846 = n7553 & ~n7584 ;
  assign n7847 = n7846 ^ n7524 ;
  assign n7848 = n7847 ^ n291 ;
  assign n7865 = n7547 ^ n401 ;
  assign n7866 = ~n7584 & n7865 ;
  assign n7867 = n7866 ^ n7549 ;
  assign n7849 = ~n7545 & ~n7584 ;
  assign n7850 = n7849 ^ n7527 ;
  assign n7851 = n7850 ^ n401 ;
  assign n7852 = n7543 & ~n7584 ;
  assign n7853 = n7852 ^ n7530 ;
  assign n7854 = n7853 ^ n457 ;
  assign n7855 = ~n7540 & ~n7584 ;
  assign n7856 = n7855 ^ n7533 ;
  assign n7857 = n7856 ^ n534 ;
  assign n7858 = ~n7807 & n7857 ;
  assign n7859 = n7858 ^ n750 ;
  assign n7860 = ~n7854 & n7859 ;
  assign n7861 = n7860 ^ n7853 ;
  assign n7862 = n7861 ^ n7850 ;
  assign n7863 = n7851 & ~n7862 ;
  assign n7864 = n7863 ^ n401 ;
  assign n7868 = n7867 ^ n7864 ;
  assign n7869 = n7867 ^ n341 ;
  assign n7870 = ~n7868 & n7869 ;
  assign n7871 = n7870 ^ n349 ;
  assign n7872 = ~n7848 & ~n7871 ;
  assign n7873 = n7872 ^ n307 ;
  assign n7874 = n7845 & n7873 ;
  assign n7875 = n7874 ^ n7844 ;
  assign n7876 = n7875 ^ n188 ;
  assign n7877 = ~n7560 & ~n7584 ;
  assign n7878 = n7877 ^ n7520 ;
  assign n7879 = n7878 ^ n7875 ;
  assign n7880 = n7876 & ~n7879 ;
  assign n7881 = n7880 ^ n203 ;
  assign n7882 = ~n7842 & ~n7881 ;
  assign n7883 = n7882 ^ n7841 ;
  assign n7884 = n7838 & n7883 ;
  assign n7885 = ~n7836 & ~n7884 ;
  assign n7808 = ~n7570 & n7573 ;
  assign n7811 = n7514 ^ n7512 ;
  assign n7812 = n7811 ^ n7514 ;
  assign n7813 = n7514 ^ n1355 ;
  assign n7814 = n7813 ^ n7514 ;
  assign n7815 = ~n7812 & ~n7814 ;
  assign n7816 = n7808 & n7815 ;
  assign n7817 = n7816 ^ n7808 ;
  assign n7809 = n7808 ^ n7514 ;
  assign n7818 = n7817 ^ n7809 ;
  assign n7819 = n7574 ^ n138 ;
  assign n7820 = n7819 ^ n7487 ;
  assign n7821 = n7820 ^ n7808 ;
  assign n7822 = ~n183 & ~n7821 ;
  assign n7823 = n7822 ^ n7487 ;
  assign n7824 = n7576 & ~n7823 ;
  assign n7825 = n7824 ^ n183 ;
  assign n7828 = n7573 & n7812 ;
  assign n7829 = n7828 ^ n7514 ;
  assign n7830 = ~n7825 & n7829 ;
  assign n7831 = ~n7579 & ~n7830 ;
  assign n7832 = ~n7818 & n7831 ;
  assign n7833 = n7832 ^ n7830 ;
  assign n7886 = n7571 & ~n7584 ;
  assign n7887 = n7886 ^ n7573 ;
  assign n7888 = n7887 ^ n183 ;
  assign n7889 = ~n7833 & n7888 ;
  assign n7890 = n7885 & n7889 ;
  assign n7891 = n7890 ^ n7833 ;
  assign n7892 = ~n7807 & n7891 ;
  assign n7893 = n7892 ^ n7856 ;
  assign n7894 = n7893 ^ n457 ;
  assign n7895 = ~n7805 & n7891 ;
  assign n7896 = n7895 ^ n7586 ;
  assign n7897 = n7896 ^ n534 ;
  assign n7898 = n7799 & n7891 ;
  assign n7899 = n7898 ^ n7801 ;
  assign n7900 = n7899 ^ n609 ;
  assign n7901 = ~n7769 & n7891 ;
  assign n7902 = n7901 ^ n7771 ;
  assign n7903 = n7902 ^ n1136 ;
  assign n8123 = n7764 & n7891 ;
  assign n8124 = n8123 ^ n7766 ;
  assign n8127 = n8124 ^ n1136 ;
  assign n8112 = ~n7753 & n7891 ;
  assign n8113 = n8112 ^ n7755 ;
  assign n8116 = n8113 ^ n1427 ;
  assign n7904 = n7749 & n7891 ;
  assign n7905 = n7904 ^ n7592 ;
  assign n7906 = n7905 ^ n2008 ;
  assign n7907 = n7743 & n7891 ;
  assign n7908 = n7907 ^ n7746 ;
  assign n7909 = n7908 ^ n2175 ;
  assign n7910 = ~n7738 & n7891 ;
  assign n7911 = n7910 ^ n7598 ;
  assign n7912 = n7911 ^ n2511 ;
  assign n7913 = ~n7736 & n7891 ;
  assign n7914 = n7913 ^ n7601 ;
  assign n7915 = n7914 ^ n2707 ;
  assign n7916 = n7729 & n7891 ;
  assign n7917 = n7916 ^ n7606 ;
  assign n7918 = n7917 ^ n3093 ;
  assign n7919 = n7727 & n7891 ;
  assign n7920 = n7919 ^ n7615 ;
  assign n7921 = n7920 ^ n3320 ;
  assign n7922 = ~n7725 & n7891 ;
  assign n7923 = n7922 ^ n7619 ;
  assign n7924 = n7923 ^ n3538 ;
  assign n8071 = n7719 ^ n3908 ;
  assign n8072 = n7891 & n8071 ;
  assign n8073 = n8072 ^ n7721 ;
  assign n7925 = ~n7717 & n7891 ;
  assign n7926 = n7925 ^ n7622 ;
  assign n7927 = n7926 ^ n3908 ;
  assign n7928 = n7711 & n7891 ;
  assign n7929 = n7928 ^ n7713 ;
  assign n7930 = n7929 ^ n4153 ;
  assign n8059 = n7705 ^ n4583 ;
  assign n8060 = n7891 & n8059 ;
  assign n8061 = n8060 ^ n7707 ;
  assign n8064 = n8061 ^ n4153 ;
  assign n7931 = n7696 ^ n5073 ;
  assign n7932 = n7891 & n7931 ;
  assign n7933 = n7932 ^ n7698 ;
  assign n7934 = n7933 ^ n4812 ;
  assign n7935 = n7694 & n7891 ;
  assign n7936 = n7935 ^ n7628 ;
  assign n7937 = n7936 ^ n5073 ;
  assign n7938 = n7691 ^ n5562 ;
  assign n7939 = n7891 & ~n7938 ;
  assign n7940 = n7939 ^ n7631 ;
  assign n7942 = n7940 ^ n5317 ;
  assign n8039 = n7689 & n7891 ;
  assign n8040 = n8039 ^ n7634 ;
  assign n7943 = ~n7687 & n7891 ;
  assign n7944 = n7943 ^ n7641 ;
  assign n7945 = n7944 ^ n5830 ;
  assign n7956 = ~x38 & ~n7584 ;
  assign n7957 = n7956 ^ x39 ;
  assign n7948 = n7666 ^ n7584 ;
  assign n7951 = n7660 ^ x38 ;
  assign n7952 = n7951 ^ n7660 ;
  assign n7953 = n7948 & ~n7952 ;
  assign n7954 = n7953 ^ n7660 ;
  assign n7955 = n7891 & n7954 ;
  assign n7958 = n7957 ^ n7955 ;
  assign n7959 = n7958 ^ n6959 ;
  assign n7963 = ~x34 & ~x35 ;
  assign n7966 = ~n7666 & n7963 ;
  assign n7964 = ~x36 & n7963 ;
  assign n7977 = n7966 ^ n7964 ;
  assign n7978 = n7977 ^ x37 ;
  assign n7979 = n7956 ^ n7584 ;
  assign n7980 = ~n7978 & ~n7979 ;
  assign n7981 = n7891 & ~n7966 ;
  assign n7982 = n7980 & ~n7981 ;
  assign n7983 = n7982 ^ n6959 ;
  assign n7960 = ~x38 & ~n7666 ;
  assign n7961 = n7891 & n7960 ;
  assign n7962 = n7961 ^ x38 ;
  assign n7965 = n7964 ^ x37 ;
  assign n7969 = n7891 & n7965 ;
  assign n7970 = n7969 ^ n7966 ;
  assign n7971 = n7891 ^ n7584 ;
  assign n7972 = n7971 ^ n7891 ;
  assign n7973 = n7972 ^ n7962 ;
  assign n7974 = n7970 & n7973 ;
  assign n7975 = n7974 ^ n7891 ;
  assign n7976 = ~n7962 & n7975 ;
  assign n7984 = n7983 ^ n7976 ;
  assign n7985 = n7984 ^ n7958 ;
  assign n7986 = n7584 ^ x38 ;
  assign n7989 = ~n7584 & ~n7977 ;
  assign n7990 = n7989 ^ n7966 ;
  assign n7991 = ~n7986 & ~n7990 ;
  assign n7992 = n7991 ^ x38 ;
  assign n7993 = n7891 & ~n7992 ;
  assign n7994 = n7964 ^ x38 ;
  assign n7996 = ~x37 & n7994 ;
  assign n7997 = n7996 ^ n7964 ;
  assign n7998 = n7993 & n7997 ;
  assign n7999 = n7998 ^ n7992 ;
  assign n8002 = n7962 ^ x37 ;
  assign n8003 = n8002 ^ n7962 ;
  assign n8004 = n7962 ^ n7584 ;
  assign n8005 = n8004 ^ n7962 ;
  assign n8006 = n8003 & ~n8005 ;
  assign n8007 = ~n7891 & n8006 ;
  assign n8008 = n8007 ^ n7891 ;
  assign n8000 = n7962 ^ n7891 ;
  assign n8009 = n8008 ^ n8000 ;
  assign n8010 = ~n7999 & n8009 ;
  assign n8013 = n7984 ^ n7277 ;
  assign n8014 = n8013 ^ n7984 ;
  assign n8015 = ~n8010 & ~n8014 ;
  assign n8016 = n7985 & n8015 ;
  assign n8017 = n8016 ^ n7985 ;
  assign n8018 = n8017 ^ n7958 ;
  assign n8019 = n7959 & ~n8018 ;
  assign n8020 = n8019 ^ n6959 ;
  assign n8021 = n8020 ^ n6673 ;
  assign n8022 = n7673 ^ n6959 ;
  assign n8023 = n7891 & n8022 ;
  assign n8024 = n8023 ^ n7677 ;
  assign n8025 = n8024 ^ n8020 ;
  assign n8026 = n8021 & n8025 ;
  assign n8027 = n8026 ^ n6713 ;
  assign n8028 = n7683 & n7891 ;
  assign n8029 = n8028 ^ n7657 ;
  assign n8030 = n8029 ^ n6389 ;
  assign n8031 = ~n8027 & ~n8030 ;
  assign n8032 = n8031 ^ n6389 ;
  assign n7946 = ~n7685 & n7891 ;
  assign n7947 = n7946 ^ n7645 ;
  assign n8033 = n8032 ^ n7947 ;
  assign n8034 = n8032 ^ n6115 ;
  assign n8035 = ~n8033 & ~n8034 ;
  assign n8036 = n8035 ^ n6429 ;
  assign n8037 = ~n7945 & ~n8036 ;
  assign n8038 = n8037 ^ n7944 ;
  assign n8041 = n8040 ^ n8038 ;
  assign n8042 = n8040 ^ n5562 ;
  assign n8043 = ~n8041 & ~n8042 ;
  assign n8044 = n8043 ^ n5885 ;
  assign n8045 = n7942 & ~n8044 ;
  assign n7941 = n7940 ^ n5073 ;
  assign n8046 = n8045 ^ n7941 ;
  assign n8047 = n7937 & n8046 ;
  assign n8048 = n8047 ^ n5073 ;
  assign n8049 = n8048 ^ n7933 ;
  assign n8050 = n7934 & ~n8049 ;
  assign n8051 = n8050 ^ n4812 ;
  assign n8052 = n8051 ^ n4583 ;
  assign n8053 = n7702 ^ n4812 ;
  assign n8054 = n7891 & n8053 ;
  assign n8055 = n8054 ^ n7625 ;
  assign n8056 = n8055 ^ n8051 ;
  assign n8057 = n8052 & n8056 ;
  assign n8058 = n8057 ^ n4645 ;
  assign n8062 = n8061 ^ n4356 ;
  assign n8063 = ~n8058 & n8062 ;
  assign n8065 = n8064 ^ n8063 ;
  assign n8066 = ~n7930 & n8065 ;
  assign n8067 = n8066 ^ n4153 ;
  assign n8068 = n8067 ^ n7926 ;
  assign n8069 = n7927 & ~n8068 ;
  assign n8070 = n8069 ^ n3908 ;
  assign n8074 = n8073 ^ n8070 ;
  assign n8075 = n8073 ^ n3722 ;
  assign n8076 = n8074 & n8075 ;
  assign n8077 = n8076 ^ n3795 ;
  assign n8078 = ~n7924 & n8077 ;
  assign n8079 = n8078 ^ n3538 ;
  assign n8080 = n8079 ^ n7920 ;
  assign n8081 = ~n7921 & n8080 ;
  assign n8082 = n8081 ^ n3387 ;
  assign n8083 = n7918 & n8082 ;
  assign n8084 = n8083 ^ n7917 ;
  assign n8085 = n8084 ^ n2894 ;
  assign n8086 = n7731 ^ n3093 ;
  assign n8087 = n7891 & ~n8086 ;
  assign n8088 = n8087 ^ n7604 ;
  assign n8089 = n8088 ^ n8084 ;
  assign n8090 = n8085 & n8089 ;
  assign n8091 = n8090 ^ n3396 ;
  assign n8092 = ~n7915 & ~n8091 ;
  assign n8093 = n8092 ^ n2707 ;
  assign n8094 = n8093 ^ n7911 ;
  assign n8095 = ~n7912 & ~n8094 ;
  assign n8096 = n8095 ^ n2530 ;
  assign n8097 = n7740 ^ n2511 ;
  assign n8098 = n7891 & ~n8097 ;
  assign n8099 = n8098 ^ n7595 ;
  assign n8100 = n8099 ^ n2366 ;
  assign n8101 = n8096 & ~n8100 ;
  assign n8102 = n8101 ^ n2399 ;
  assign n8103 = n7909 & n8102 ;
  assign n8104 = n8103 ^ n2204 ;
  assign n8105 = n7906 & n8104 ;
  assign n8106 = n8105 ^ n2064 ;
  assign n8107 = n7751 & n7891 ;
  assign n8108 = n8107 ^ n7589 ;
  assign n8109 = n8108 ^ n1739 ;
  assign n8110 = ~n8106 & ~n8109 ;
  assign n8111 = n8110 ^ n1763 ;
  assign n8114 = n8113 ^ n1572 ;
  assign n8115 = n8111 & ~n8114 ;
  assign n8117 = n8116 ^ n8115 ;
  assign n8118 = ~n7758 & n7891 ;
  assign n8119 = n8118 ^ n7760 ;
  assign n8120 = n8119 ^ n1427 ;
  assign n8121 = n8117 & n8120 ;
  assign n8122 = n8121 ^ n1450 ;
  assign n8125 = n8124 ^ n1290 ;
  assign n8126 = n8122 & ~n8125 ;
  assign n8128 = n8127 ^ n8126 ;
  assign n8129 = ~n7903 & ~n8128 ;
  assign n8130 = n8129 ^ n1143 ;
  assign n8131 = n7774 & n7891 ;
  assign n8132 = n8131 ^ n7776 ;
  assign n8135 = n8132 ^ n1034 ;
  assign n8136 = ~n8130 & n8135 ;
  assign n8133 = n8132 ^ n892 ;
  assign n8137 = n8136 ^ n8133 ;
  assign n8138 = n7779 & n7891 ;
  assign n8139 = n8138 ^ n7782 ;
  assign n8140 = n8139 ^ n786 ;
  assign n8141 = n8140 ^ n927 ;
  assign n8142 = ~n8137 & n8141 ;
  assign n8143 = n8142 ^ n8140 ;
  assign n8144 = n7787 & n7891 ;
  assign n8145 = n8144 ^ n7789 ;
  assign n8146 = n8145 ^ n696 ;
  assign n8147 = n8146 ^ n842 ;
  assign n8148 = ~n8143 & n8147 ;
  assign n8149 = n8148 ^ n8146 ;
  assign n8150 = n7793 & n7891 ;
  assign n8151 = n8150 ^ n7795 ;
  assign n8152 = n8151 ^ n609 ;
  assign n8153 = n8152 ^ n835 ;
  assign n8154 = ~n8149 & n8153 ;
  assign n8155 = n8154 ^ n8152 ;
  assign n8156 = ~n7900 & ~n8155 ;
  assign n8157 = n8156 ^ n834 ;
  assign n8158 = n7897 & ~n8157 ;
  assign n8159 = n8158 ^ n750 ;
  assign n8160 = ~n7894 & n8159 ;
  assign n8161 = n8160 ^ n7893 ;
  assign n8162 = n8161 ^ n401 ;
  assign n8163 = n7883 ^ n138 ;
  assign n8164 = n7891 & ~n8163 ;
  assign n8165 = n8164 ^ n7835 ;
  assign n8166 = n8165 ^ n183 ;
  assign n8207 = n1003 & n7835 ;
  assign n8208 = n7887 & n8207 ;
  assign n8181 = n7836 ^ n7833 ;
  assign n8182 = n8181 ^ n7887 ;
  assign n8183 = n8182 ^ n7833 ;
  assign n8187 = n8183 ^ n183 ;
  assign n8188 = n8187 ^ n8182 ;
  assign n8189 = n8188 ^ n8183 ;
  assign n8185 = n7883 ^ n183 ;
  assign n8190 = n8185 ^ n8181 ;
  assign n8191 = ~n8189 & ~n8190 ;
  assign n8200 = n8191 ^ n8187 ;
  assign n8192 = n8189 ^ n8181 ;
  assign n8193 = n8192 ^ n8191 ;
  assign n8194 = n8185 ^ n8183 ;
  assign n8195 = n8193 & n8194 ;
  assign n8201 = n8200 ^ n8195 ;
  assign n8202 = n8195 ^ n7887 ;
  assign n8203 = ~n8201 & n8202 ;
  assign n8204 = ~n8181 & n8203 ;
  assign n8197 = n8195 ^ n7836 ;
  assign n8205 = n8204 ^ n8197 ;
  assign n8167 = n7887 ^ n7884 ;
  assign n8171 = n8167 ^ n7887 ;
  assign n8168 = n8167 ^ n183 ;
  assign n8169 = n8168 ^ n7887 ;
  assign n8172 = n8169 ^ n7833 ;
  assign n8173 = n8172 ^ n8169 ;
  assign n8174 = n8171 & n8173 ;
  assign n8175 = n8174 ^ n8169 ;
  assign n8176 = n8167 ^ n138 ;
  assign n8177 = n8174 ^ n8171 ;
  assign n8178 = ~n8176 & n8177 ;
  assign n8179 = n8178 ^ n8167 ;
  assign n8180 = n8175 & ~n8179 ;
  assign n8206 = n8205 ^ n8180 ;
  assign n8209 = n8208 ^ n8206 ;
  assign n8210 = n7876 & n7891 ;
  assign n8211 = n8210 ^ n7878 ;
  assign n8212 = n8211 ^ n157 ;
  assign n8236 = ~n7873 & n7891 ;
  assign n8237 = n8236 ^ n7844 ;
  assign n8213 = ~n7871 & n7891 ;
  assign n8214 = n8213 ^ n7847 ;
  assign n8215 = n8214 ^ n245 ;
  assign n8216 = n7861 ^ n401 ;
  assign n8217 = n7891 & n8216 ;
  assign n8218 = n8217 ^ n7850 ;
  assign n8219 = n8218 ^ n341 ;
  assign n8220 = ~n7859 & n7891 ;
  assign n8221 = n8220 ^ n7853 ;
  assign n8222 = n8221 ^ n8161 ;
  assign n8223 = n8221 ^ n401 ;
  assign n8224 = ~n8222 & n8223 ;
  assign n8225 = n8224 ^ n462 ;
  assign n8226 = n8219 & n8225 ;
  assign n8227 = n8226 ^ n349 ;
  assign n8228 = n7864 ^ n341 ;
  assign n8229 = n7891 & n8228 ;
  assign n8230 = n8229 ^ n7867 ;
  assign n8231 = n8230 ^ n291 ;
  assign n8232 = ~n8227 & ~n8231 ;
  assign n8233 = n8232 ^ n307 ;
  assign n8234 = n8215 & n8233 ;
  assign n8235 = n8234 ^ n8214 ;
  assign n8238 = n8237 ^ n8235 ;
  assign n8239 = n8237 ^ n188 ;
  assign n8240 = ~n8238 & n8239 ;
  assign n8241 = n8240 ^ n203 ;
  assign n8242 = n8212 & ~n8241 ;
  assign n8243 = n8242 ^ n8211 ;
  assign n8244 = n138 & n8243 ;
  assign n8245 = n8243 ^ n138 ;
  assign n8246 = n8245 ^ n8244 ;
  assign n8247 = n7881 & n7891 ;
  assign n8248 = n8247 ^ n7841 ;
  assign n8249 = n8246 & ~n8248 ;
  assign n8250 = ~n8244 & ~n8249 ;
  assign n8251 = n8209 & ~n8250 ;
  assign n8252 = ~n8166 & n8251 ;
  assign n8253 = n8252 ^ n8209 ;
  assign n8254 = n8162 & ~n8253 ;
  assign n8255 = n8254 ^ n8221 ;
  assign n8256 = n8255 ^ n341 ;
  assign n8517 = ~n8159 & ~n8253 ;
  assign n8518 = n8517 ^ n7893 ;
  assign n8257 = ~n8157 & ~n8253 ;
  assign n8258 = n8257 ^ n7896 ;
  assign n8259 = n8258 ^ n457 ;
  assign n8260 = ~n8155 & ~n8253 ;
  assign n8261 = n8260 ^ n7899 ;
  assign n8262 = n8261 ^ n534 ;
  assign n8263 = n8149 & ~n8253 ;
  assign n8264 = n8263 ^ n8151 ;
  assign n8265 = n8264 ^ n609 ;
  assign n8266 = ~n8128 & ~n8253 ;
  assign n8267 = n8266 ^ n7902 ;
  assign n8268 = n8267 ^ n1034 ;
  assign n8478 = n8117 & ~n8253 ;
  assign n8479 = n8478 ^ n8119 ;
  assign n8482 = n8479 ^ n1136 ;
  assign n8467 = ~n8106 & ~n8253 ;
  assign n8468 = n8467 ^ n8108 ;
  assign n8471 = n8468 ^ n1427 ;
  assign n8269 = n8104 & ~n8253 ;
  assign n8270 = n8269 ^ n7905 ;
  assign n8271 = n8270 ^ n1739 ;
  assign n8272 = n8102 & ~n8253 ;
  assign n8273 = n8272 ^ n7908 ;
  assign n8274 = n8273 ^ n2008 ;
  assign n8275 = n8096 & ~n8253 ;
  assign n8276 = n8275 ^ n8099 ;
  assign n8277 = n8276 ^ n2175 ;
  assign n8278 = n8093 ^ n2511 ;
  assign n8279 = ~n8253 & ~n8278 ;
  assign n8280 = n8279 ^ n7911 ;
  assign n8281 = n8280 ^ n2366 ;
  assign n8452 = ~n8091 & ~n8253 ;
  assign n8453 = n8452 ^ n7914 ;
  assign n8282 = ~n8082 & ~n8253 ;
  assign n8283 = n8282 ^ n7917 ;
  assign n8284 = n8283 ^ n2894 ;
  assign n8285 = n8077 & ~n8253 ;
  assign n8286 = n8285 ^ n7923 ;
  assign n8287 = n8286 ^ n3320 ;
  assign n8423 = n8067 ^ n3908 ;
  assign n8424 = ~n8253 & n8423 ;
  assign n8425 = n8424 ^ n7926 ;
  assign n8293 = n8065 & ~n8253 ;
  assign n8294 = n8293 ^ n7929 ;
  assign n8295 = n8294 ^ n3908 ;
  assign n8296 = n8046 & ~n8253 ;
  assign n8297 = n8296 ^ n7936 ;
  assign n8298 = n8297 ^ n4812 ;
  assign n8299 = n8044 & ~n8253 ;
  assign n8300 = n8299 ^ n7940 ;
  assign n8301 = n8300 ^ n5073 ;
  assign n8305 = n8036 & ~n8253 ;
  assign n8306 = n8305 ^ n7944 ;
  assign n8307 = n8306 ^ n5562 ;
  assign n8388 = ~n8034 & ~n8253 ;
  assign n8389 = n8388 ^ n7947 ;
  assign n8308 = n7984 ^ n6959 ;
  assign n8309 = n8308 ^ n8010 ;
  assign n8310 = n7985 ^ n7277 ;
  assign n8311 = n8010 ^ n7277 ;
  assign n8312 = n8311 ^ n7277 ;
  assign n8313 = n8310 & n8312 ;
  assign n8314 = n8313 ^ n7277 ;
  assign n8315 = ~n8309 & ~n8314 ;
  assign n8316 = n8315 ^ n7984 ;
  assign n8317 = ~n8253 & ~n8316 ;
  assign n8318 = n8317 ^ n7958 ;
  assign n8319 = n8318 ^ n6673 ;
  assign n8332 = ~n7891 & n7948 ;
  assign n8328 = ~n7665 & n7891 ;
  assign n8321 = n7964 ^ n7584 ;
  assign n8323 = n7277 ^ x37 ;
  assign n8322 = n7891 ^ n7277 ;
  assign n8324 = n8323 ^ n8322 ;
  assign n8325 = n8324 ^ n7584 ;
  assign n8326 = n8321 & n8325 ;
  assign n8327 = n8326 ^ n8323 ;
  assign n8329 = n8328 ^ n8327 ;
  assign n8330 = ~n8253 & n8329 ;
  assign n8320 = n7666 ^ x38 ;
  assign n8331 = n8330 ^ n8320 ;
  assign n8333 = n8332 ^ n8331 ;
  assign n8334 = n8333 ^ n6959 ;
  assign n8347 = n7891 ^ x36 ;
  assign n8345 = n7963 ^ n7891 ;
  assign n8346 = ~n8253 & n8345 ;
  assign n8348 = n8347 ^ n8346 ;
  assign n8349 = n8348 ^ n7584 ;
  assign n8350 = n7891 ^ x35 ;
  assign n8351 = n8350 ^ n8253 ;
  assign n8353 = ~x32 & ~x33 ;
  assign n8352 = n7891 ^ x34 ;
  assign n8354 = n8353 ^ n8352 ;
  assign n8355 = n8351 & n8354 ;
  assign n8364 = n8355 ^ n7971 ;
  assign n8356 = n8253 ^ n7891 ;
  assign n8357 = n8356 ^ n8355 ;
  assign n8358 = n8357 ^ n8355 ;
  assign n8361 = ~n8350 & ~n8358 ;
  assign n8362 = n8361 ^ n8355 ;
  assign n8363 = x34 & n8362 ;
  assign n8365 = n8364 ^ n8363 ;
  assign n8366 = n8349 & n8365 ;
  assign n8367 = n8366 ^ n8348 ;
  assign n8342 = n7891 ^ x37 ;
  assign n8343 = n8342 ^ n8321 ;
  assign n8335 = n8321 ^ x36 ;
  assign n8336 = n8335 ^ n8321 ;
  assign n8337 = n8321 ^ n7891 ;
  assign n8338 = n8337 ^ n8321 ;
  assign n8339 = n8336 & n8338 ;
  assign n8340 = n8339 ^ n8321 ;
  assign n8341 = n8253 & ~n8340 ;
  assign n8344 = n8343 ^ n8341 ;
  assign n8368 = n8367 ^ n8344 ;
  assign n8369 = n8367 ^ n7277 ;
  assign n8370 = n8368 & n8369 ;
  assign n8371 = n8370 ^ n7277 ;
  assign n8372 = n8371 ^ n8333 ;
  assign n8373 = ~n8334 & n8372 ;
  assign n8374 = n8373 ^ n7011 ;
  assign n8375 = n8319 & n8374 ;
  assign n8376 = n8375 ^ n6673 ;
  assign n8377 = n8376 ^ n6389 ;
  assign n8378 = n8021 & ~n8253 ;
  assign n8379 = n8378 ^ n8024 ;
  assign n8380 = n8379 ^ n8376 ;
  assign n8381 = ~n8377 & n8380 ;
  assign n8382 = n8381 ^ n6423 ;
  assign n8383 = ~n8027 & ~n8253 ;
  assign n8384 = n8383 ^ n8029 ;
  assign n8385 = n8384 ^ n6115 ;
  assign n8386 = ~n8382 & n8385 ;
  assign n8387 = n8386 ^ n6115 ;
  assign n8390 = n8389 ^ n8387 ;
  assign n8391 = n8387 ^ n5830 ;
  assign n8392 = n8390 & n8391 ;
  assign n8393 = n8392 ^ n5900 ;
  assign n8394 = ~n8307 & n8393 ;
  assign n8395 = n8394 ^ n5562 ;
  assign n8302 = n8038 ^ n5562 ;
  assign n8303 = ~n8253 & ~n8302 ;
  assign n8304 = n8303 ^ n8040 ;
  assign n8396 = n8395 ^ n8304 ;
  assign n8397 = n8304 ^ n5317 ;
  assign n8398 = n8396 & ~n8397 ;
  assign n8399 = n8398 ^ n5360 ;
  assign n8400 = n8301 & n8399 ;
  assign n8401 = n8400 ^ n5115 ;
  assign n8402 = n8298 & n8401 ;
  assign n8403 = n8402 ^ n4854 ;
  assign n8404 = n8048 ^ n4812 ;
  assign n8405 = ~n8253 & n8404 ;
  assign n8406 = n8405 ^ n7933 ;
  assign n8407 = n8406 ^ n4583 ;
  assign n8408 = n8403 & n8407 ;
  assign n8409 = n8408 ^ n4645 ;
  assign n8410 = n8052 & ~n8253 ;
  assign n8411 = n8410 ^ n8055 ;
  assign n8412 = n8411 ^ n4356 ;
  assign n8413 = n8409 & ~n8412 ;
  assign n8414 = n8413 ^ n4414 ;
  assign n8415 = n8058 & ~n8253 ;
  assign n8416 = n8415 ^ n8061 ;
  assign n8417 = n8416 ^ n4153 ;
  assign n8418 = n8414 & n8417 ;
  assign n8419 = n8418 ^ n4153 ;
  assign n8420 = n8419 ^ n8294 ;
  assign n8421 = ~n8295 & n8420 ;
  assign n8422 = n8421 ^ n3908 ;
  assign n8426 = n8425 ^ n8422 ;
  assign n8427 = n8425 ^ n3722 ;
  assign n8428 = ~n8426 & ~n8427 ;
  assign n8429 = n8428 ^ n3722 ;
  assign n8291 = n8286 ^ n3538 ;
  assign n8288 = n8070 ^ n3722 ;
  assign n8289 = ~n8253 & ~n8288 ;
  assign n8290 = n8289 ^ n8073 ;
  assign n8292 = n8291 ^ n8290 ;
  assign n8430 = n8429 ^ n8292 ;
  assign n8431 = n8430 ^ n8291 ;
  assign n8432 = n8290 ^ n8286 ;
  assign n8433 = n8432 ^ n8291 ;
  assign n8434 = ~n8431 & n8433 ;
  assign n8435 = n8434 ^ n8291 ;
  assign n8436 = ~n8287 & n8435 ;
  assign n8437 = n8436 ^ n3387 ;
  assign n8438 = n8079 ^ n3320 ;
  assign n8439 = ~n8253 & n8438 ;
  assign n8440 = n8439 ^ n7920 ;
  assign n8441 = n8440 ^ n3093 ;
  assign n8442 = ~n8437 & n8441 ;
  assign n8443 = n8442 ^ n3363 ;
  assign n8444 = n8284 & n8443 ;
  assign n8445 = n8444 ^ n2894 ;
  assign n8446 = n8445 ^ n2707 ;
  assign n8447 = n8085 & ~n8253 ;
  assign n8448 = n8447 ^ n8088 ;
  assign n8449 = n8448 ^ n8445 ;
  assign n8450 = ~n8446 & n8449 ;
  assign n8451 = n8450 ^ n2707 ;
  assign n8454 = n8453 ^ n8451 ;
  assign n8455 = n8453 ^ n2511 ;
  assign n8456 = n8454 & n8455 ;
  assign n8457 = n8456 ^ n2530 ;
  assign n8458 = ~n8281 & n8457 ;
  assign n8459 = n8458 ^ n2399 ;
  assign n8460 = ~n8277 & n8459 ;
  assign n8461 = n8460 ^ n2175 ;
  assign n8462 = n8461 ^ n8273 ;
  assign n8463 = n8274 & ~n8462 ;
  assign n8464 = n8463 ^ n2064 ;
  assign n8465 = ~n8271 & ~n8464 ;
  assign n8466 = n8465 ^ n1763 ;
  assign n8469 = n8468 ^ n1572 ;
  assign n8470 = n8466 & n8469 ;
  assign n8472 = n8471 ^ n8470 ;
  assign n8473 = ~n8111 & ~n8253 ;
  assign n8474 = n8473 ^ n8113 ;
  assign n8475 = n8474 ^ n1427 ;
  assign n8476 = ~n8472 & n8475 ;
  assign n8477 = n8476 ^ n1450 ;
  assign n8480 = n8479 ^ n1290 ;
  assign n8481 = n8477 & ~n8480 ;
  assign n8483 = n8482 ^ n8481 ;
  assign n8484 = ~n8122 & ~n8253 ;
  assign n8485 = n8484 ^ n8124 ;
  assign n8486 = n8485 ^ n1143 ;
  assign n8487 = n8486 ^ n1034 ;
  assign n8488 = ~n8483 & ~n8487 ;
  assign n8489 = n8488 ^ n1143 ;
  assign n8490 = ~n8268 & n8489 ;
  assign n8491 = n8490 ^ n1072 ;
  assign n8492 = n8130 & ~n8253 ;
  assign n8493 = n8492 ^ n8132 ;
  assign n8496 = n8493 ^ n892 ;
  assign n8497 = ~n8491 & n8496 ;
  assign n8494 = n8493 ^ n786 ;
  assign n8498 = n8497 ^ n8494 ;
  assign n8499 = n8137 & ~n8253 ;
  assign n8500 = n8499 ^ n8139 ;
  assign n8501 = n8500 ^ n696 ;
  assign n8502 = n8501 ^ n842 ;
  assign n8503 = ~n8498 & n8502 ;
  assign n8504 = n8503 ^ n8501 ;
  assign n8505 = n8143 & ~n8253 ;
  assign n8506 = n8505 ^ n8145 ;
  assign n8507 = n8506 ^ n609 ;
  assign n8508 = n8507 ^ n835 ;
  assign n8509 = ~n8504 & n8508 ;
  assign n8510 = n8509 ^ n8507 ;
  assign n8511 = ~n8265 & ~n8510 ;
  assign n8512 = n8511 ^ n834 ;
  assign n8513 = n8262 & ~n8512 ;
  assign n8514 = n8513 ^ n750 ;
  assign n8515 = ~n8259 & n8514 ;
  assign n8516 = n8515 ^ n8258 ;
  assign n8519 = n8518 ^ n8516 ;
  assign n8520 = n8518 ^ n401 ;
  assign n8521 = ~n8519 & n8520 ;
  assign n8522 = n8521 ^ n462 ;
  assign n8523 = n8256 & n8522 ;
  assign n8524 = n8523 ^ n349 ;
  assign n8525 = n8225 & ~n8253 ;
  assign n8526 = n8525 ^ n8218 ;
  assign n8527 = n8526 ^ n291 ;
  assign n8528 = ~n8524 & ~n8527 ;
  assign n8529 = n8528 ^ n307 ;
  assign n8536 = n8245 & ~n8253 ;
  assign n8537 = n8536 ^ n8248 ;
  assign n8538 = n183 & ~n8537 ;
  assign n8539 = n8538 ^ n183 ;
  assign n8553 = n8243 ^ n8209 ;
  assign n8554 = n8553 ^ n8248 ;
  assign n8555 = n8554 ^ n8209 ;
  assign n8558 = ~n138 & ~n8555 ;
  assign n8559 = n8558 ^ n8209 ;
  assign n8560 = n8165 & ~n8559 ;
  assign n8561 = n8560 ^ n8250 ;
  assign n8562 = ~n183 & ~n8561 ;
  assign n8542 = ~n8165 & n8209 ;
  assign n8540 = n8244 ^ n8165 ;
  assign n8541 = n8540 ^ n8244 ;
  assign n8543 = n8542 ^ n8541 ;
  assign n8544 = n8543 ^ n8540 ;
  assign n8545 = n8540 ^ n8249 ;
  assign n8546 = n8545 ^ n8540 ;
  assign n8547 = ~n8544 & n8546 ;
  assign n8548 = n8547 ^ n8540 ;
  assign n8549 = n8248 & n8542 ;
  assign n8550 = n183 & ~n8549 ;
  assign n8551 = ~n8548 & n8550 ;
  assign n8552 = n8551 ^ n8549 ;
  assign n8563 = n8248 ^ n8245 ;
  assign n8564 = ~n8552 & n8563 ;
  assign n8565 = n8562 & n8564 ;
  assign n8566 = n8565 ^ n8552 ;
  assign n8567 = n8241 & ~n8253 ;
  assign n8568 = n8567 ^ n8211 ;
  assign n8569 = n8568 ^ n138 ;
  assign n8570 = n8235 ^ n188 ;
  assign n8571 = ~n8253 & n8570 ;
  assign n8572 = n8571 ^ n8237 ;
  assign n8574 = n8572 ^ n157 ;
  assign n8530 = ~n8227 & ~n8253 ;
  assign n8531 = n8530 ^ n8230 ;
  assign n8532 = n8531 ^ n245 ;
  assign n8533 = n8529 & n8532 ;
  assign n8534 = n8533 ^ n8531 ;
  assign n8535 = n8534 ^ n188 ;
  assign n8575 = ~n8233 & ~n8253 ;
  assign n8576 = n8575 ^ n8214 ;
  assign n8577 = n8576 ^ n8534 ;
  assign n8578 = n8535 & ~n8577 ;
  assign n8579 = n8578 ^ n203 ;
  assign n8580 = n8574 & ~n8579 ;
  assign n8573 = n8572 ^ n8568 ;
  assign n8581 = n8580 ^ n8573 ;
  assign n8582 = n8569 & ~n8581 ;
  assign n8583 = n8582 ^ n138 ;
  assign n8584 = n8566 & n8583 ;
  assign n8585 = ~n8539 & n8584 ;
  assign n8586 = n8585 ^ n8566 ;
  assign n8861 = ~n8529 & ~n8586 ;
  assign n8862 = n8861 ^ n8531 ;
  assign n8590 = ~n8524 & ~n8586 ;
  assign n8591 = n8590 ^ n8526 ;
  assign n8592 = n8591 ^ n245 ;
  assign n8593 = n8522 & ~n8586 ;
  assign n8594 = n8593 ^ n8255 ;
  assign n8595 = n8594 ^ n291 ;
  assign n8596 = n8516 ^ n401 ;
  assign n8597 = ~n8586 & n8596 ;
  assign n8598 = n8597 ^ n8518 ;
  assign n8599 = n8598 ^ n341 ;
  assign n8849 = ~n8514 & ~n8586 ;
  assign n8850 = n8849 ^ n8258 ;
  assign n8600 = ~n8512 & ~n8586 ;
  assign n8601 = n8600 ^ n8261 ;
  assign n8602 = n8601 ^ n457 ;
  assign n8603 = ~n8510 & ~n8586 ;
  assign n8604 = n8603 ^ n8264 ;
  assign n8605 = n8604 ^ n534 ;
  assign n8606 = n8504 & ~n8586 ;
  assign n8607 = n8606 ^ n8506 ;
  assign n8843 = n8607 ^ n534 ;
  assign n8608 = n8607 ^ n609 ;
  assign n8609 = n8489 & ~n8586 ;
  assign n8610 = n8609 ^ n8267 ;
  assign n8611 = n8610 ^ n892 ;
  assign n8612 = ~n8477 & ~n8586 ;
  assign n8613 = n8612 ^ n8479 ;
  assign n8614 = n8613 ^ n1136 ;
  assign n8814 = ~n8472 & ~n8586 ;
  assign n8815 = n8814 ^ n8474 ;
  assign n8818 = n8815 ^ n1136 ;
  assign n8615 = ~n8464 & ~n8586 ;
  assign n8616 = n8615 ^ n8270 ;
  assign n8807 = n8616 ^ n1427 ;
  assign n8617 = n8616 ^ n1572 ;
  assign n8621 = n8459 & ~n8586 ;
  assign n8622 = n8621 ^ n8276 ;
  assign n8623 = n8622 ^ n2008 ;
  assign n8624 = n8457 & ~n8586 ;
  assign n8625 = n8624 ^ n8280 ;
  assign n8626 = n8625 ^ n2175 ;
  assign n8627 = n8451 ^ n2511 ;
  assign n8628 = ~n8586 & ~n8627 ;
  assign n8629 = n8628 ^ n8453 ;
  assign n8630 = n8629 ^ n2366 ;
  assign n8637 = n8429 ^ n3320 ;
  assign n8638 = n8637 ^ n3596 ;
  assign n8639 = n8290 ^ n3320 ;
  assign n8640 = n8639 ^ n3596 ;
  assign n8641 = n8638 & n8640 ;
  assign n8642 = n8641 ^ n3596 ;
  assign n8643 = ~n8586 & n8642 ;
  assign n8644 = n8643 ^ n8286 ;
  assign n8645 = n8644 ^ n3093 ;
  assign n8646 = n8429 ^ n3538 ;
  assign n8647 = ~n8586 & n8646 ;
  assign n8648 = n8647 ^ n8290 ;
  assign n8649 = n8648 ^ n3320 ;
  assign n8650 = n8422 ^ n3722 ;
  assign n8651 = ~n8586 & ~n8650 ;
  assign n8652 = n8651 ^ n8425 ;
  assign n8653 = n8652 ^ n3538 ;
  assign n8654 = n8414 & ~n8586 ;
  assign n8655 = n8654 ^ n8416 ;
  assign n8656 = n8655 ^ n3908 ;
  assign n8657 = n8409 & ~n8586 ;
  assign n8658 = n8657 ^ n8411 ;
  assign n8659 = n8658 ^ n4153 ;
  assign n8760 = n8403 & ~n8586 ;
  assign n8761 = n8760 ^ n8406 ;
  assign n8764 = n8761 ^ n4153 ;
  assign n8660 = n8395 ^ n5317 ;
  assign n8661 = ~n8586 & n8660 ;
  assign n8662 = n8661 ^ n8304 ;
  assign n8663 = n8662 ^ n5073 ;
  assign n8667 = n8391 & ~n8586 ;
  assign n8668 = n8667 ^ n8389 ;
  assign n8669 = n8668 ^ n5562 ;
  assign n8670 = ~n8382 & ~n8586 ;
  assign n8671 = n8670 ^ n8384 ;
  assign n8672 = n8671 ^ n5830 ;
  assign n8673 = ~n8377 & ~n8586 ;
  assign n8674 = n8673 ^ n8379 ;
  assign n8675 = n8674 ^ n6115 ;
  assign n8731 = n8374 & ~n8586 ;
  assign n8732 = n8731 ^ n8318 ;
  assign n8676 = n8371 ^ n6959 ;
  assign n8677 = ~n8586 & n8676 ;
  assign n8678 = n8677 ^ n8333 ;
  assign n8679 = n8678 ^ n6673 ;
  assign n8680 = n8369 & ~n8586 ;
  assign n8681 = n8680 ^ n8344 ;
  assign n8682 = n8681 ^ n6959 ;
  assign n8683 = ~n8365 & ~n8586 ;
  assign n8684 = n8683 ^ n8348 ;
  assign n8685 = n8684 ^ n7277 ;
  assign n8702 = n8353 ^ n8253 ;
  assign n8712 = n8356 ^ x34 ;
  assign n8713 = n8712 ^ n8356 ;
  assign n8714 = ~n8702 & ~n8713 ;
  assign n8715 = n8714 ^ n8356 ;
  assign n8716 = ~n8586 & ~n8715 ;
  assign n8717 = n8716 ^ x35 ;
  assign n8709 = ~x34 & ~n8253 ;
  assign n8718 = n8717 ^ n8709 ;
  assign n8721 = n8718 ^ n7277 ;
  assign n8703 = ~n8586 & ~n8702 ;
  assign n8701 = n8253 ^ x34 ;
  assign n8704 = n8703 ^ n8701 ;
  assign n8688 = n8586 ^ n8253 ;
  assign n8686 = n8253 ^ x33 ;
  assign n8687 = n8686 ^ x32 ;
  assign n8689 = n8688 ^ n8687 ;
  assign n8690 = n8689 ^ n8688 ;
  assign n8691 = n8690 ^ n8686 ;
  assign n8693 = n8686 ^ n8586 ;
  assign n8694 = ~x30 & ~x31 ;
  assign n8695 = n8694 ^ n8689 ;
  assign n8696 = ~n8693 & ~n8695 ;
  assign n8692 = n8686 & n8688 ;
  assign n8697 = n8696 ^ n8692 ;
  assign n8698 = ~n8691 & n8697 ;
  assign n8699 = n8698 ^ n8692 ;
  assign n8700 = n8699 ^ n8253 ;
  assign n8705 = n8704 ^ n8700 ;
  assign n8706 = n8704 ^ n7891 ;
  assign n8707 = n8705 & n8706 ;
  assign n8708 = n8707 ^ n7971 ;
  assign n8719 = n8718 ^ n7584 ;
  assign n8720 = n8708 & n8719 ;
  assign n8722 = n8721 ^ n8720 ;
  assign n8723 = n8685 & n8722 ;
  assign n8724 = n8723 ^ n7277 ;
  assign n8725 = n8724 ^ n8681 ;
  assign n8726 = ~n8682 & n8725 ;
  assign n8727 = n8726 ^ n6959 ;
  assign n8728 = n8727 ^ n8678 ;
  assign n8729 = ~n8679 & n8728 ;
  assign n8730 = n8729 ^ n6673 ;
  assign n8733 = n8732 ^ n8730 ;
  assign n8734 = n8732 ^ n6389 ;
  assign n8735 = ~n8733 & ~n8734 ;
  assign n8736 = n8735 ^ n6389 ;
  assign n8737 = n8736 ^ n8674 ;
  assign n8738 = ~n8675 & ~n8737 ;
  assign n8739 = n8738 ^ n6429 ;
  assign n8740 = n8672 & ~n8739 ;
  assign n8741 = n8740 ^ n8671 ;
  assign n8742 = n8741 ^ n8668 ;
  assign n8743 = ~n8669 & n8742 ;
  assign n8744 = n8743 ^ n5885 ;
  assign n8664 = n8393 & ~n8586 ;
  assign n8665 = n8664 ^ n8306 ;
  assign n8745 = n8665 ^ n5317 ;
  assign n8746 = ~n8744 & ~n8745 ;
  assign n8666 = n8665 ^ n5073 ;
  assign n8747 = n8746 ^ n8666 ;
  assign n8748 = ~n8663 & ~n8747 ;
  assign n8749 = n8748 ^ n5115 ;
  assign n8750 = n8399 & ~n8586 ;
  assign n8751 = n8750 ^ n8300 ;
  assign n8752 = n8751 ^ n4812 ;
  assign n8753 = n8749 & n8752 ;
  assign n8754 = n8753 ^ n4854 ;
  assign n8755 = n8401 & ~n8586 ;
  assign n8756 = n8755 ^ n8297 ;
  assign n8757 = n8756 ^ n4583 ;
  assign n8758 = n8754 & n8757 ;
  assign n8759 = n8758 ^ n4645 ;
  assign n8762 = n8761 ^ n4356 ;
  assign n8763 = ~n8759 & n8762 ;
  assign n8765 = n8764 ^ n8763 ;
  assign n8766 = ~n8659 & n8765 ;
  assign n8767 = n8766 ^ n4153 ;
  assign n8768 = n8767 ^ n8655 ;
  assign n8769 = n8656 & ~n8768 ;
  assign n8770 = n8769 ^ n3961 ;
  assign n8771 = n8419 ^ n3908 ;
  assign n8772 = ~n8586 & n8771 ;
  assign n8773 = n8772 ^ n8294 ;
  assign n8774 = n8773 ^ n3722 ;
  assign n8775 = ~n8770 & n8774 ;
  assign n8776 = n8775 ^ n3795 ;
  assign n8777 = ~n8653 & n8776 ;
  assign n8778 = n8777 ^ n3538 ;
  assign n8779 = n8778 ^ n8648 ;
  assign n8780 = n8649 & ~n8779 ;
  assign n8781 = n8780 ^ n3387 ;
  assign n8782 = n8645 & n8781 ;
  assign n8783 = n8782 ^ n8644 ;
  assign n8635 = ~n8437 & ~n8586 ;
  assign n8636 = n8635 ^ n8440 ;
  assign n8784 = n8783 ^ n8636 ;
  assign n8785 = n8783 ^ n2894 ;
  assign n8786 = ~n8784 & n8785 ;
  assign n8787 = n8786 ^ n2894 ;
  assign n8633 = n8443 & ~n8586 ;
  assign n8634 = n8633 ^ n8283 ;
  assign n8788 = n8787 ^ n8634 ;
  assign n8789 = n8787 ^ n2707 ;
  assign n8790 = ~n8788 & ~n8789 ;
  assign n8791 = n8790 ^ n2707 ;
  assign n8631 = ~n8446 & ~n8586 ;
  assign n8632 = n8631 ^ n8448 ;
  assign n8792 = n8791 ^ n8632 ;
  assign n8793 = n8791 ^ n2511 ;
  assign n8794 = ~n8792 & ~n8793 ;
  assign n8795 = n8794 ^ n2530 ;
  assign n8796 = n8630 & n8795 ;
  assign n8797 = n8796 ^ n2399 ;
  assign n8798 = ~n8626 & n8797 ;
  assign n8799 = n8798 ^ n2204 ;
  assign n8800 = ~n8623 & n8799 ;
  assign n8801 = n8800 ^ n2008 ;
  assign n8618 = n8461 ^ n2008 ;
  assign n8619 = ~n8586 & n8618 ;
  assign n8620 = n8619 ^ n8273 ;
  assign n8802 = n8801 ^ n8620 ;
  assign n8803 = n8801 ^ n1739 ;
  assign n8804 = ~n8802 & ~n8803 ;
  assign n8805 = n8804 ^ n1763 ;
  assign n8806 = n8617 & n8805 ;
  assign n8808 = n8807 ^ n8806 ;
  assign n8809 = ~n8466 & ~n8586 ;
  assign n8810 = n8809 ^ n8468 ;
  assign n8811 = n8810 ^ n1427 ;
  assign n8812 = ~n8808 & ~n8811 ;
  assign n8813 = n8812 ^ n1450 ;
  assign n8816 = n8815 ^ n1290 ;
  assign n8817 = n8813 & ~n8816 ;
  assign n8819 = n8818 ^ n8817 ;
  assign n8820 = ~n8614 & ~n8819 ;
  assign n8821 = n8820 ^ n1143 ;
  assign n8822 = ~n8483 & ~n8586 ;
  assign n8823 = n8822 ^ n8485 ;
  assign n8824 = n8823 ^ n1034 ;
  assign n8825 = n8821 & ~n8824 ;
  assign n8826 = n8825 ^ n1072 ;
  assign n8827 = ~n8611 & n8826 ;
  assign n8828 = n8827 ^ n927 ;
  assign n8829 = n8491 & ~n8586 ;
  assign n8830 = n8829 ^ n8493 ;
  assign n8833 = n8830 ^ n786 ;
  assign n8834 = ~n8828 & n8833 ;
  assign n8831 = n8830 ^ n696 ;
  assign n8835 = n8834 ^ n8831 ;
  assign n8836 = n8498 & ~n8586 ;
  assign n8837 = n8836 ^ n8500 ;
  assign n8838 = n8837 ^ n609 ;
  assign n8839 = n8838 ^ n835 ;
  assign n8840 = ~n8835 & n8839 ;
  assign n8841 = n8840 ^ n8838 ;
  assign n8842 = ~n8608 & n8841 ;
  assign n8844 = n8843 ^ n8842 ;
  assign n8845 = n8605 & n8844 ;
  assign n8846 = n8845 ^ n750 ;
  assign n8847 = ~n8602 & n8846 ;
  assign n8848 = n8847 ^ n8601 ;
  assign n8851 = n8850 ^ n8848 ;
  assign n8852 = n8850 ^ n401 ;
  assign n8853 = ~n8851 & n8852 ;
  assign n8854 = n8853 ^ n462 ;
  assign n8855 = n8599 & n8854 ;
  assign n8856 = n8855 ^ n349 ;
  assign n8857 = ~n8595 & ~n8856 ;
  assign n8858 = n8857 ^ n307 ;
  assign n8859 = n8592 & n8858 ;
  assign n8860 = n8859 ^ n8591 ;
  assign n8863 = n8862 ^ n8860 ;
  assign n8864 = n8862 ^ n188 ;
  assign n8865 = ~n8863 & n8864 ;
  assign n8866 = n8865 ^ n203 ;
  assign n8587 = n8535 & ~n8586 ;
  assign n8588 = n8587 ^ n8576 ;
  assign n8589 = n8588 ^ n157 ;
  assign n8867 = n8589 & ~n8866 ;
  assign n8868 = n8867 ^ n8588 ;
  assign n8869 = n8868 ^ n138 ;
  assign n8870 = n8579 & ~n8586 ;
  assign n8871 = n8870 ^ n8572 ;
  assign n8872 = n8871 ^ n8868 ;
  assign n8873 = n8869 & ~n8872 ;
  assign n8874 = n8873 ^ n138 ;
  assign n8902 = n8538 & n8583 ;
  assign n8887 = n8568 ^ n137 ;
  assign n8888 = n8887 ^ x127 ;
  assign n8876 = n8580 ^ n8572 ;
  assign n8889 = n8888 ^ n8876 ;
  assign n8877 = n8876 ^ n138 ;
  assign n8878 = ~n8568 & ~n8877 ;
  assign n8890 = ~n4971 & ~n8877 ;
  assign n8891 = n8890 ^ n8537 ;
  assign n8892 = ~n8878 & n8891 ;
  assign n8893 = n8889 & n8892 ;
  assign n8894 = n8893 ^ n8537 ;
  assign n8875 = n8568 ^ n8537 ;
  assign n8879 = n8878 ^ n8875 ;
  assign n8880 = ~n183 & ~n8879 ;
  assign n8881 = n8880 ^ n8537 ;
  assign n8882 = n8566 & ~n8881 ;
  assign n8883 = ~n8568 & n8882 ;
  assign n8884 = n8880 & n8883 ;
  assign n8885 = n8884 ^ n8882 ;
  assign n8886 = n8885 ^ n8566 ;
  assign n8895 = n8893 ^ n8891 ;
  assign n8896 = ~n8886 & n8895 ;
  assign n8897 = n8893 ^ n8876 ;
  assign n8898 = n8896 & n8897 ;
  assign n8899 = ~n8894 & n8898 ;
  assign n8900 = n8899 ^ n8896 ;
  assign n8901 = n8900 ^ n8886 ;
  assign n8903 = n8902 ^ n8901 ;
  assign n8904 = ~n8586 & n8877 ;
  assign n8905 = n8904 ^ n8568 ;
  assign n8906 = ~n183 & ~n8905 ;
  assign n8907 = n8906 ^ n8905 ;
  assign n8908 = n8903 & n8907 ;
  assign n8909 = n8874 & n8908 ;
  assign n8910 = n8909 ^ n8903 ;
  assign n8915 = n8866 & ~n8910 ;
  assign n8916 = n8915 ^ n8588 ;
  assign n8917 = n8916 ^ n138 ;
  assign n8918 = n8860 ^ n188 ;
  assign n8919 = ~n8910 & n8918 ;
  assign n8920 = n8919 ^ n8862 ;
  assign n8921 = n8920 ^ n157 ;
  assign n8924 = ~n8856 & ~n8910 ;
  assign n8925 = n8924 ^ n8594 ;
  assign n8926 = n8925 ^ n245 ;
  assign n8927 = ~n8846 & ~n8910 ;
  assign n8928 = n8927 ^ n8601 ;
  assign n8929 = n8928 ^ n401 ;
  assign n8930 = n8844 & ~n8910 ;
  assign n8931 = n8930 ^ n8604 ;
  assign n8932 = n8931 ^ n457 ;
  assign n8933 = n8835 & ~n8910 ;
  assign n8934 = n8933 ^ n8837 ;
  assign n8935 = n8934 ^ n609 ;
  assign n8936 = n8826 & ~n8910 ;
  assign n8937 = n8936 ^ n8610 ;
  assign n8938 = n8937 ^ n786 ;
  assign n8939 = n8821 & ~n8910 ;
  assign n8940 = n8939 ^ n8823 ;
  assign n8941 = n8940 ^ n892 ;
  assign n8942 = ~n8813 & ~n8910 ;
  assign n8943 = n8942 ^ n8815 ;
  assign n8944 = n8943 ^ n1136 ;
  assign n9136 = ~n8808 & ~n8910 ;
  assign n9137 = n9136 ^ n8810 ;
  assign n9140 = n9137 ^ n1136 ;
  assign n8945 = ~n8805 & ~n8910 ;
  assign n8946 = n8945 ^ n8616 ;
  assign n8947 = n8946 ^ n1427 ;
  assign n9127 = ~n8803 & ~n8910 ;
  assign n9128 = n9127 ^ n8620 ;
  assign n9132 = n9128 ^ n1427 ;
  assign n8948 = n8797 & ~n8910 ;
  assign n8949 = n8948 ^ n8625 ;
  assign n8950 = n8949 ^ n2008 ;
  assign n8951 = n8795 & ~n8910 ;
  assign n8952 = n8951 ^ n8629 ;
  assign n8953 = n8952 ^ n2175 ;
  assign n8954 = ~n8789 & ~n8910 ;
  assign n8955 = n8954 ^ n8634 ;
  assign n8956 = n8955 ^ n2511 ;
  assign n9104 = n8785 & ~n8910 ;
  assign n9105 = n9104 ^ n8636 ;
  assign n8957 = ~n8781 & ~n8910 ;
  assign n8958 = n8957 ^ n8644 ;
  assign n8959 = n8958 ^ n2894 ;
  assign n8963 = n8776 & ~n8910 ;
  assign n8964 = n8963 ^ n8652 ;
  assign n8965 = n8964 ^ n3320 ;
  assign n8966 = ~n8770 & ~n8910 ;
  assign n8967 = n8966 ^ n8773 ;
  assign n8968 = n8967 ^ n3538 ;
  assign n8969 = n8767 ^ n3908 ;
  assign n8970 = ~n8910 & n8969 ;
  assign n8971 = n8970 ^ n8655 ;
  assign n8972 = n8971 ^ n3722 ;
  assign n9086 = n8765 & ~n8910 ;
  assign n9087 = n9086 ^ n8658 ;
  assign n9080 = n8759 & ~n8910 ;
  assign n9081 = n9080 ^ n8761 ;
  assign n8973 = n8754 & ~n8910 ;
  assign n8974 = n8973 ^ n8756 ;
  assign n8975 = n8974 ^ n4356 ;
  assign n8976 = ~n8747 & ~n8910 ;
  assign n8977 = n8976 ^ n8662 ;
  assign n8978 = n8977 ^ n4812 ;
  assign n8979 = n8744 & ~n8910 ;
  assign n8980 = n8979 ^ n8665 ;
  assign n8981 = n8980 ^ n5073 ;
  assign n8982 = n8739 & ~n8910 ;
  assign n8983 = n8982 ^ n8671 ;
  assign n8984 = n8983 ^ n5562 ;
  assign n8985 = n8730 ^ n6389 ;
  assign n8986 = ~n8910 & ~n8985 ;
  assign n8987 = n8986 ^ n8732 ;
  assign n8988 = n8987 ^ n6115 ;
  assign n9045 = n8727 ^ n6673 ;
  assign n9046 = ~n8910 & n9045 ;
  assign n9047 = n9046 ^ n8678 ;
  assign n8989 = n8724 ^ n6959 ;
  assign n8990 = ~n8910 & n8989 ;
  assign n8991 = n8990 ^ n8681 ;
  assign n8992 = n8991 ^ n6673 ;
  assign n8993 = n8722 & ~n8910 ;
  assign n8994 = n8993 ^ n8684 ;
  assign n8995 = n8994 ^ n6959 ;
  assign n8996 = n8700 ^ n7891 ;
  assign n8997 = ~n8910 & ~n8996 ;
  assign n8998 = n8997 ^ n8704 ;
  assign n8999 = n8998 ^ n7584 ;
  assign n9000 = n8694 ^ n8586 ;
  assign n9001 = ~n8910 & ~n9000 ;
  assign n9002 = n9001 ^ n8586 ;
  assign n9003 = n9002 ^ x32 ;
  assign n9004 = n9003 ^ n8253 ;
  assign n9006 = n8586 ^ x31 ;
  assign n9007 = n9006 ^ n8910 ;
  assign n9009 = n8586 ^ x30 ;
  assign n9008 = ~x28 & ~x29 ;
  assign n9010 = n9009 ^ n9008 ;
  assign n9011 = ~n9007 & ~n9010 ;
  assign n9019 = n9011 ^ n8688 ;
  assign n9005 = n8910 ^ n8586 ;
  assign n9012 = n9011 ^ n9005 ;
  assign n9013 = n9012 ^ n9011 ;
  assign n9016 = n9006 & n9013 ;
  assign n9017 = n9016 ^ n9011 ;
  assign n9018 = x30 & n9017 ;
  assign n9020 = n9019 ^ n9018 ;
  assign n9021 = ~n9004 & n9020 ;
  assign n9022 = n9021 ^ n8253 ;
  assign n9023 = n9022 ^ n7891 ;
  assign n9027 = n8586 ^ x33 ;
  assign n9025 = n8694 ^ n8253 ;
  assign n9026 = ~n8910 & ~n9025 ;
  assign n9028 = n9027 ^ n9026 ;
  assign n9024 = x32 & ~n9002 ;
  assign n9029 = n9028 ^ n9024 ;
  assign n9030 = n9029 ^ n9022 ;
  assign n9031 = ~n9023 & n9030 ;
  assign n9032 = n9031 ^ n7971 ;
  assign n9033 = ~n8999 & ~n9032 ;
  assign n9034 = n9033 ^ n7660 ;
  assign n9035 = ~n8708 & ~n8910 ;
  assign n9036 = n9035 ^ n8718 ;
  assign n9037 = n9036 ^ n7277 ;
  assign n9038 = n9034 & n9037 ;
  assign n9039 = n9038 ^ n7339 ;
  assign n9040 = n8995 & n9039 ;
  assign n9041 = n9040 ^ n6959 ;
  assign n9042 = n9041 ^ n8991 ;
  assign n9043 = ~n8992 & n9042 ;
  assign n9044 = n9043 ^ n6673 ;
  assign n9048 = n9047 ^ n9044 ;
  assign n9049 = n9047 ^ n6389 ;
  assign n9050 = n9048 & n9049 ;
  assign n9051 = n9050 ^ n6423 ;
  assign n9052 = n8988 & ~n9051 ;
  assign n9053 = n9052 ^ n6429 ;
  assign n9054 = n8736 ^ n6115 ;
  assign n9055 = ~n8910 & ~n9054 ;
  assign n9056 = n9055 ^ n8674 ;
  assign n9057 = n9056 ^ n5830 ;
  assign n9058 = n9053 & ~n9057 ;
  assign n9059 = n9058 ^ n5900 ;
  assign n9060 = n8984 & n9059 ;
  assign n9061 = n9060 ^ n5885 ;
  assign n9062 = n8741 ^ n5562 ;
  assign n9063 = ~n8910 & n9062 ;
  assign n9064 = n9063 ^ n8668 ;
  assign n9065 = n9064 ^ n5317 ;
  assign n9066 = n9061 & ~n9065 ;
  assign n9067 = n9066 ^ n5360 ;
  assign n9068 = ~n8981 & n9067 ;
  assign n9069 = n9068 ^ n5073 ;
  assign n9070 = n9069 ^ n8977 ;
  assign n9071 = ~n8978 & n9070 ;
  assign n9072 = n9071 ^ n4854 ;
  assign n9073 = n8749 & ~n8910 ;
  assign n9074 = n9073 ^ n8751 ;
  assign n9075 = n9074 ^ n4583 ;
  assign n9076 = n9072 & n9075 ;
  assign n9077 = n9076 ^ n4645 ;
  assign n9078 = n8975 & ~n9077 ;
  assign n9079 = n9078 ^ n8974 ;
  assign n9082 = n9081 ^ n9079 ;
  assign n9083 = n9081 ^ n4153 ;
  assign n9084 = ~n9082 & n9083 ;
  assign n9085 = n9084 ^ n4153 ;
  assign n9088 = n9087 ^ n9085 ;
  assign n9089 = n9087 ^ n3908 ;
  assign n9090 = n9088 & ~n9089 ;
  assign n9091 = n9090 ^ n3961 ;
  assign n9092 = ~n8972 & ~n9091 ;
  assign n9093 = n9092 ^ n3795 ;
  assign n9094 = n8968 & n9093 ;
  assign n9095 = n9094 ^ n3596 ;
  assign n9096 = ~n8965 & n9095 ;
  assign n9097 = n9096 ^ n3320 ;
  assign n8960 = n8778 ^ n3320 ;
  assign n8961 = ~n8910 & n8960 ;
  assign n8962 = n8961 ^ n8648 ;
  assign n9098 = n9097 ^ n8962 ;
  assign n9099 = n8962 ^ n3093 ;
  assign n9100 = ~n9098 & ~n9099 ;
  assign n9101 = n9100 ^ n3363 ;
  assign n9102 = n8959 & n9101 ;
  assign n9103 = n9102 ^ n2894 ;
  assign n9106 = n9105 ^ n9103 ;
  assign n9107 = n9105 ^ n2707 ;
  assign n9108 = ~n9106 & ~n9107 ;
  assign n9109 = n9108 ^ n2707 ;
  assign n9110 = n9109 ^ n8955 ;
  assign n9111 = n8956 & n9110 ;
  assign n9112 = n9111 ^ n2530 ;
  assign n9113 = ~n8793 & ~n8910 ;
  assign n9114 = n9113 ^ n8632 ;
  assign n9115 = n9114 ^ n2366 ;
  assign n9116 = n9112 & ~n9115 ;
  assign n9117 = n9116 ^ n2399 ;
  assign n9118 = n8953 & n9117 ;
  assign n9119 = n9118 ^ n2204 ;
  assign n9120 = ~n8950 & n9119 ;
  assign n9121 = n9120 ^ n2064 ;
  assign n9122 = n8799 & ~n8910 ;
  assign n9123 = n9122 ^ n8622 ;
  assign n9124 = n9123 ^ n1739 ;
  assign n9125 = ~n9121 & n9124 ;
  assign n9126 = n9125 ^ n1739 ;
  assign n9129 = n9128 ^ n9126 ;
  assign n9130 = n9126 ^ n1572 ;
  assign n9131 = ~n9129 & n9130 ;
  assign n9133 = n9132 ^ n9131 ;
  assign n9134 = ~n8947 & ~n9133 ;
  assign n9135 = n9134 ^ n1450 ;
  assign n9138 = n9137 ^ n1290 ;
  assign n9139 = n9135 & n9138 ;
  assign n9141 = n9140 ^ n9139 ;
  assign n9142 = ~n8944 & n9141 ;
  assign n9143 = n9142 ^ n1143 ;
  assign n9144 = ~n8819 & ~n8910 ;
  assign n9145 = n9144 ^ n8613 ;
  assign n9148 = n9145 ^ n1034 ;
  assign n9149 = ~n9143 & ~n9148 ;
  assign n9146 = n9145 ^ n892 ;
  assign n9150 = n9149 ^ n9146 ;
  assign n9151 = ~n8941 & ~n9150 ;
  assign n9152 = n9151 ^ n927 ;
  assign n9153 = ~n8938 & n9152 ;
  assign n9154 = n9153 ^ n842 ;
  assign n9155 = n8828 & ~n8910 ;
  assign n9156 = n9155 ^ n8830 ;
  assign n9159 = n9156 ^ n696 ;
  assign n9160 = ~n9154 & n9159 ;
  assign n9157 = n9156 ^ n609 ;
  assign n9161 = n9160 ^ n9157 ;
  assign n9162 = ~n8935 & ~n9161 ;
  assign n9163 = n9162 ^ n834 ;
  assign n9164 = ~n8841 & ~n8910 ;
  assign n9165 = n9164 ^ n8607 ;
  assign n9166 = n9165 ^ n534 ;
  assign n9167 = ~n9163 & n9166 ;
  assign n9168 = n9167 ^ n750 ;
  assign n9169 = ~n8932 & n9168 ;
  assign n9170 = n9169 ^ n8931 ;
  assign n9171 = n9170 ^ n8928 ;
  assign n9172 = n8929 & ~n9171 ;
  assign n9173 = n9172 ^ n462 ;
  assign n9174 = n8848 ^ n401 ;
  assign n9175 = ~n8910 & n9174 ;
  assign n9176 = n9175 ^ n8850 ;
  assign n9177 = n9176 ^ n341 ;
  assign n9178 = n9173 & n9177 ;
  assign n9179 = n9178 ^ n349 ;
  assign n9180 = n8854 & ~n8910 ;
  assign n9181 = n9180 ^ n8598 ;
  assign n9182 = n9181 ^ n291 ;
  assign n9183 = ~n9179 & ~n9182 ;
  assign n9184 = n9183 ^ n307 ;
  assign n9185 = n8926 & n9184 ;
  assign n9186 = n9185 ^ n8925 ;
  assign n8922 = ~n8858 & ~n8910 ;
  assign n8923 = n8922 ^ n8591 ;
  assign n9187 = n9186 ^ n8923 ;
  assign n9188 = n9186 ^ n188 ;
  assign n9189 = ~n9187 & n9188 ;
  assign n9190 = n9189 ^ n203 ;
  assign n9191 = n8921 & ~n9190 ;
  assign n9192 = n9191 ^ n8920 ;
  assign n9193 = n9192 ^ n8916 ;
  assign n9194 = n8917 & ~n9193 ;
  assign n9195 = n9194 ^ n138 ;
  assign n8911 = n8869 & ~n8910 ;
  assign n8912 = n8911 ^ n8871 ;
  assign n9469 = n9195 ^ n8912 ;
  assign n9474 = n9469 ^ n183 ;
  assign n9475 = ~n8912 & ~n8916 ;
  assign n9200 = ~n8903 & ~n8907 ;
  assign n9196 = ~n1355 & ~n8903 ;
  assign n9197 = ~n8868 & ~n8871 ;
  assign n9198 = n9196 & n9197 ;
  assign n9199 = n9198 ^ n8905 ;
  assign n9201 = n9200 ^ n9199 ;
  assign n9202 = n183 & n8874 ;
  assign n9203 = n9201 & n9202 ;
  assign n9204 = n9203 ^ n9199 ;
  assign n9205 = n8906 & ~n9204 ;
  assign n9207 = n8903 ^ n8869 ;
  assign n9208 = ~n8871 & ~n9207 ;
  assign n9206 = n8871 ^ n8869 ;
  assign n9209 = n9208 ^ n9206 ;
  assign n9210 = n9205 & n9209 ;
  assign n9213 = n9210 ^ n9204 ;
  assign n9211 = n8868 & n9208 ;
  assign n9212 = n9210 & n9211 ;
  assign n9214 = n9213 ^ n9212 ;
  assign n9479 = n9192 ^ n8912 ;
  assign n9471 = n8912 & ~n9214 ;
  assign n9480 = n9479 ^ n9471 ;
  assign n9476 = n9203 ^ n8907 ;
  assign n8913 = n183 & n8912 ;
  assign n9477 = n9476 ^ n8913 ;
  assign n9478 = n8916 & n9477 ;
  assign n9481 = n9480 ^ n9478 ;
  assign n9482 = ~n183 & ~n9481 ;
  assign n9483 = n9482 ^ n9477 ;
  assign n9484 = n9483 ^ n9482 ;
  assign n9485 = ~n9214 & n9484 ;
  assign n9486 = n9475 & n9485 ;
  assign n9487 = n9486 ^ n9483 ;
  assign n9488 = ~n9474 & n9487 ;
  assign n9489 = n9488 ^ n9482 ;
  assign n9470 = n8912 ^ n1355 ;
  assign n9472 = n9471 ^ n9470 ;
  assign n9473 = n9469 & ~n9472 ;
  assign n9490 = n9489 ^ n9473 ;
  assign n8914 = n8913 ^ n183 ;
  assign n9215 = n9195 & ~n9214 ;
  assign n9216 = ~n8914 & n9215 ;
  assign n9217 = n9216 ^ n9214 ;
  assign n9529 = n9190 & n9217 ;
  assign n9530 = n9529 ^ n8920 ;
  assign n9491 = n9188 & n9217 ;
  assign n9492 = n9491 ^ n8923 ;
  assign n9493 = n9492 ^ n157 ;
  assign n9521 = ~n9184 & n9217 ;
  assign n9522 = n9521 ^ n8925 ;
  assign n9494 = n9170 ^ n401 ;
  assign n9495 = n9217 & n9494 ;
  assign n9496 = n9495 ^ n8928 ;
  assign n9497 = n9496 ^ n341 ;
  assign n9503 = ~n9168 & n9217 ;
  assign n9504 = n9503 ^ n8931 ;
  assign n9218 = ~n9161 & n9217 ;
  assign n9219 = n9218 ^ n8934 ;
  assign n9220 = n9219 ^ n534 ;
  assign n9221 = n9154 & n9217 ;
  assign n9222 = n9221 ^ n9156 ;
  assign n9461 = n9222 ^ n534 ;
  assign n9223 = n9222 ^ n609 ;
  assign n9224 = n9152 & n9217 ;
  assign n9225 = n9224 ^ n8937 ;
  assign n9226 = n9225 ^ n696 ;
  assign n9227 = ~n9150 & n9217 ;
  assign n9228 = n9227 ^ n8940 ;
  assign n9229 = n9228 ^ n786 ;
  assign n9230 = ~n9135 & n9217 ;
  assign n9231 = n9230 ^ n9137 ;
  assign n9232 = n9231 ^ n1136 ;
  assign n9435 = ~n9133 & n9217 ;
  assign n9436 = n9435 ^ n8946 ;
  assign n9439 = n9436 ^ n1136 ;
  assign n9424 = ~n9121 & n9217 ;
  assign n9425 = n9424 ^ n9123 ;
  assign n9428 = n9425 ^ n1427 ;
  assign n9233 = n9117 & n9217 ;
  assign n9234 = n9233 ^ n8952 ;
  assign n9235 = n9234 ^ n2008 ;
  assign n9238 = n9103 ^ n2707 ;
  assign n9239 = n9217 & ~n9238 ;
  assign n9240 = n9239 ^ n9105 ;
  assign n9241 = n9240 ^ n2511 ;
  assign n9242 = n9097 ^ n3093 ;
  assign n9243 = n9217 & ~n9242 ;
  assign n9244 = n9243 ^ n8962 ;
  assign n9245 = n9244 ^ n2894 ;
  assign n9391 = n9095 & n9217 ;
  assign n9392 = n9391 ^ n8964 ;
  assign n9395 = n9392 ^ n2894 ;
  assign n9246 = ~n9091 & n9217 ;
  assign n9247 = n9246 ^ n8971 ;
  assign n9248 = n9247 ^ n3538 ;
  assign n9377 = n9085 ^ n3908 ;
  assign n9378 = n9217 & n9377 ;
  assign n9379 = n9378 ^ n9087 ;
  assign n9370 = n9079 ^ n4153 ;
  assign n9371 = n9217 & n9370 ;
  assign n9372 = n9371 ^ n9081 ;
  assign n9249 = n9077 & n9217 ;
  assign n9250 = n9249 ^ n8974 ;
  assign n9251 = n9250 ^ n4153 ;
  assign n9362 = n9072 & n9217 ;
  assign n9363 = n9362 ^ n9074 ;
  assign n9366 = n9363 ^ n4153 ;
  assign n9252 = n9067 & n9217 ;
  assign n9253 = n9252 ^ n8980 ;
  assign n9254 = n9253 ^ n4812 ;
  assign n9257 = ~n9051 & n9217 ;
  assign n9258 = n9257 ^ n8987 ;
  assign n9259 = n9258 ^ n5830 ;
  assign n9263 = n9041 ^ n6673 ;
  assign n9264 = n9217 & n9263 ;
  assign n9265 = n9264 ^ n8991 ;
  assign n9266 = n9265 ^ n6389 ;
  assign n9324 = n9039 & n9217 ;
  assign n9325 = n9324 ^ n8994 ;
  assign n9267 = ~n9032 & n9217 ;
  assign n9268 = n9267 ^ n8998 ;
  assign n9269 = n9268 ^ n7277 ;
  assign n9311 = ~n9023 & n9217 ;
  assign n9312 = n9311 ^ n9029 ;
  assign n9315 = n9312 ^ n7277 ;
  assign n9270 = n9020 & n9217 ;
  assign n9271 = n9270 ^ n9003 ;
  assign n9272 = n9271 ^ n7891 ;
  assign n9302 = n8910 ^ x31 ;
  assign n9300 = n9008 ^ n8586 ;
  assign n9301 = n9217 & ~n9300 ;
  assign n9303 = n9302 ^ n9301 ;
  assign n9292 = n9008 ^ n8910 ;
  assign n9293 = ~n9217 & ~n9292 ;
  assign n9294 = n9293 ^ n9008 ;
  assign n9299 = x30 & n9294 ;
  assign n9304 = n9303 ^ n9299 ;
  assign n9280 = n8586 ^ x29 ;
  assign n9273 = ~x26 & ~x27 ;
  assign n9274 = n9273 ^ x28 ;
  assign n9275 = n9274 ^ n8910 ;
  assign n9276 = n9217 ^ x29 ;
  assign n9277 = n9276 ^ n8910 ;
  assign n9278 = ~n9275 & n9277 ;
  assign n9279 = n9278 ^ n9005 ;
  assign n9281 = n9280 ^ n9279 ;
  assign n9282 = n9281 ^ x29 ;
  assign n9283 = n9282 ^ n8910 ;
  assign n9284 = n9283 ^ n9281 ;
  assign n9285 = n9217 ^ n8910 ;
  assign n9286 = n9285 ^ n9281 ;
  assign n9287 = n9286 ^ n9281 ;
  assign n9288 = n9284 & n9287 ;
  assign n9289 = n9288 ^ n9281 ;
  assign n9290 = x28 & n9289 ;
  assign n9291 = n9290 ^ n9279 ;
  assign n9295 = n9294 ^ x30 ;
  assign n9296 = n9295 ^ n8586 ;
  assign n9297 = n9291 & n9296 ;
  assign n9298 = n9297 ^ n8586 ;
  assign n9305 = n9304 ^ n9298 ;
  assign n9306 = n9304 ^ n8253 ;
  assign n9307 = n9305 & ~n9306 ;
  assign n9308 = n9307 ^ n8356 ;
  assign n9309 = n9272 & ~n9308 ;
  assign n9310 = n9309 ^ n7971 ;
  assign n9313 = n9312 ^ n7584 ;
  assign n9314 = n9310 & ~n9313 ;
  assign n9316 = n9315 ^ n9314 ;
  assign n9317 = ~n9269 & ~n9316 ;
  assign n9318 = n9317 ^ n7339 ;
  assign n9319 = n9034 & n9217 ;
  assign n9320 = n9319 ^ n9036 ;
  assign n9321 = n9320 ^ n6959 ;
  assign n9322 = n9318 & n9321 ;
  assign n9323 = n9322 ^ n6959 ;
  assign n9326 = n9325 ^ n9323 ;
  assign n9327 = n9325 ^ n6673 ;
  assign n9328 = ~n9326 & n9327 ;
  assign n9329 = n9328 ^ n6713 ;
  assign n9330 = n9266 & ~n9329 ;
  assign n9331 = n9330 ^ n6389 ;
  assign n9260 = n9044 ^ n6389 ;
  assign n9261 = n9217 & ~n9260 ;
  assign n9262 = n9261 ^ n9047 ;
  assign n9332 = n9331 ^ n9262 ;
  assign n9333 = n9331 ^ n6115 ;
  assign n9334 = ~n9332 & ~n9333 ;
  assign n9335 = n9334 ^ n6429 ;
  assign n9336 = n9259 & ~n9335 ;
  assign n9337 = n9336 ^ n9258 ;
  assign n9338 = n9337 ^ n5562 ;
  assign n9339 = n9053 & n9217 ;
  assign n9340 = n9339 ^ n9056 ;
  assign n9341 = n9340 ^ n9337 ;
  assign n9342 = n9338 & n9341 ;
  assign n9343 = n9342 ^ n5885 ;
  assign n9344 = n9059 & n9217 ;
  assign n9345 = n9344 ^ n8983 ;
  assign n9346 = n9345 ^ n5317 ;
  assign n9347 = ~n9343 & n9346 ;
  assign n9348 = n9347 ^ n9345 ;
  assign n9255 = n9061 & n9217 ;
  assign n9256 = n9255 ^ n9064 ;
  assign n9349 = n9348 ^ n9256 ;
  assign n9350 = n9348 ^ n5073 ;
  assign n9351 = n9349 & n9350 ;
  assign n9352 = n9351 ^ n5115 ;
  assign n9353 = ~n9254 & n9352 ;
  assign n9354 = n9353 ^ n4812 ;
  assign n9355 = n9354 ^ n4583 ;
  assign n9356 = n9069 ^ n4812 ;
  assign n9357 = n9217 & n9356 ;
  assign n9358 = n9357 ^ n8977 ;
  assign n9359 = n9358 ^ n9354 ;
  assign n9360 = n9355 & n9359 ;
  assign n9361 = n9360 ^ n4645 ;
  assign n9364 = n9363 ^ n4356 ;
  assign n9365 = ~n9361 & n9364 ;
  assign n9367 = n9366 ^ n9365 ;
  assign n9368 = n9251 & n9367 ;
  assign n9369 = n9368 ^ n4153 ;
  assign n9373 = n9372 ^ n9369 ;
  assign n9374 = n9372 ^ n3908 ;
  assign n9375 = ~n9373 & n9374 ;
  assign n9376 = n9375 ^ n3908 ;
  assign n9380 = n9379 ^ n9376 ;
  assign n9381 = n9379 ^ n3722 ;
  assign n9382 = n9380 & n9381 ;
  assign n9383 = n9382 ^ n3795 ;
  assign n9384 = ~n9248 & n9383 ;
  assign n9385 = n9384 ^ n3596 ;
  assign n9386 = n9093 & n9217 ;
  assign n9387 = n9386 ^ n8967 ;
  assign n9388 = n9387 ^ n3320 ;
  assign n9389 = n9385 & n9388 ;
  assign n9390 = n9389 ^ n3387 ;
  assign n9393 = n9392 ^ n3093 ;
  assign n9394 = n9390 & n9393 ;
  assign n9396 = n9395 ^ n9394 ;
  assign n9397 = ~n9245 & n9396 ;
  assign n9398 = n9397 ^ n3396 ;
  assign n9399 = n9101 & n9217 ;
  assign n9400 = n9399 ^ n8958 ;
  assign n9401 = n9400 ^ n2707 ;
  assign n9402 = ~n9398 & ~n9401 ;
  assign n9403 = n9402 ^ n2707 ;
  assign n9404 = n9403 ^ n9240 ;
  assign n9405 = n9241 & n9404 ;
  assign n9406 = n9405 ^ n2530 ;
  assign n9407 = n9109 ^ n2511 ;
  assign n9408 = n9217 & ~n9407 ;
  assign n9409 = n9408 ^ n8955 ;
  assign n9410 = n9409 ^ n2366 ;
  assign n9411 = n9406 & n9410 ;
  assign n9412 = n9411 ^ n2366 ;
  assign n9236 = n9112 & n9217 ;
  assign n9237 = n9236 ^ n9114 ;
  assign n9413 = n9412 ^ n9237 ;
  assign n9414 = n9412 ^ n2175 ;
  assign n9415 = n9413 & n9414 ;
  assign n9416 = n9415 ^ n2204 ;
  assign n9417 = n9235 & n9416 ;
  assign n9418 = n9417 ^ n2064 ;
  assign n9419 = n9119 & n9217 ;
  assign n9420 = n9419 ^ n8949 ;
  assign n9421 = n9420 ^ n1739 ;
  assign n9422 = ~n9418 & n9421 ;
  assign n9423 = n9422 ^ n1763 ;
  assign n9426 = n9425 ^ n1572 ;
  assign n9427 = n9423 & ~n9426 ;
  assign n9429 = n9428 ^ n9427 ;
  assign n9430 = ~n9130 & n9217 ;
  assign n9431 = n9430 ^ n9128 ;
  assign n9432 = n9431 ^ n1427 ;
  assign n9433 = n9429 & ~n9432 ;
  assign n9434 = n9433 ^ n1450 ;
  assign n9437 = n9436 ^ n1290 ;
  assign n9438 = n9434 & n9437 ;
  assign n9440 = n9439 ^ n9438 ;
  assign n9441 = n9232 & n9440 ;
  assign n9442 = n9441 ^ n1143 ;
  assign n9443 = n9141 & n9217 ;
  assign n9444 = n9443 ^ n8943 ;
  assign n9447 = n9444 ^ n1034 ;
  assign n9448 = ~n9442 & ~n9447 ;
  assign n9445 = n9444 ^ n892 ;
  assign n9449 = n9448 ^ n9445 ;
  assign n9450 = n9143 & n9217 ;
  assign n9451 = n9450 ^ n9145 ;
  assign n9452 = n9451 ^ n786 ;
  assign n9453 = n9452 ^ n927 ;
  assign n9454 = n9449 & ~n9453 ;
  assign n9455 = n9454 ^ n9452 ;
  assign n9456 = ~n9229 & ~n9455 ;
  assign n9457 = n9456 ^ n842 ;
  assign n9458 = ~n9226 & n9457 ;
  assign n9459 = n9458 ^ n835 ;
  assign n9460 = ~n9223 & n9459 ;
  assign n9462 = n9461 ^ n9460 ;
  assign n9463 = n9220 & n9462 ;
  assign n9464 = n9463 ^ n750 ;
  assign n9498 = ~n9163 & n9217 ;
  assign n9499 = n9498 ^ n9165 ;
  assign n9500 = n9499 ^ n457 ;
  assign n9501 = n9464 & ~n9500 ;
  assign n9502 = n9501 ^ n9499 ;
  assign n9505 = n9504 ^ n9502 ;
  assign n9506 = n9504 ^ n401 ;
  assign n9507 = ~n9505 & n9506 ;
  assign n9508 = n9507 ^ n462 ;
  assign n9509 = n9497 & n9508 ;
  assign n9510 = n9509 ^ n349 ;
  assign n9511 = n9173 & n9217 ;
  assign n9512 = n9511 ^ n9176 ;
  assign n9513 = n9512 ^ n291 ;
  assign n9514 = ~n9510 & ~n9513 ;
  assign n9515 = n9514 ^ n307 ;
  assign n9516 = ~n9179 & n9217 ;
  assign n9517 = n9516 ^ n9181 ;
  assign n9518 = n9517 ^ n245 ;
  assign n9519 = n9515 & n9518 ;
  assign n9520 = n9519 ^ n9517 ;
  assign n9523 = n9522 ^ n9520 ;
  assign n9524 = n9522 ^ n188 ;
  assign n9525 = ~n9523 & n9524 ;
  assign n9526 = n9525 ^ n203 ;
  assign n9527 = n9493 & ~n9526 ;
  assign n9528 = n9527 ^ n9492 ;
  assign n9531 = n9530 ^ n9528 ;
  assign n9534 = n9530 ^ n138 ;
  assign n9537 = ~n9531 & n9534 ;
  assign n9538 = n9537 ^ n138 ;
  assign n9539 = ~n9490 & n9538 ;
  assign n9541 = n9539 ^ n9490 ;
  assign n9465 = n9192 ^ n138 ;
  assign n9466 = n9217 & n9465 ;
  assign n9467 = n9466 ^ n8916 ;
  assign n9468 = n183 & ~n9467 ;
  assign n9540 = n9468 & n9539 ;
  assign n9542 = n9541 ^ n9540 ;
  assign n9813 = n9528 ^ n138 ;
  assign n9814 = n9542 & n9813 ;
  assign n9815 = n9814 ^ n9530 ;
  assign n9816 = ~n183 & ~n9815 ;
  assign n9817 = n9816 ^ n9815 ;
  assign n9956 = n9528 ^ n9490 ;
  assign n9954 = n9528 ^ n9467 ;
  assign n9955 = n9954 ^ n9813 ;
  assign n9959 = n9956 ^ n9955 ;
  assign n9960 = n9959 ^ n138 ;
  assign n9961 = n9960 ^ n9534 ;
  assign n9855 = n9813 ^ n9467 ;
  assign n9860 = n9855 ^ n9530 ;
  assign n9857 = n9813 ^ n9534 ;
  assign n9861 = n9860 ^ n9857 ;
  assign n9856 = n9855 ^ n9490 ;
  assign n9858 = n9857 ^ n9856 ;
  assign n9936 = n9861 ^ n9858 ;
  assign n9937 = n9936 ^ n9861 ;
  assign n9938 = n9937 ^ n9857 ;
  assign n9863 = n9857 ^ n9855 ;
  assign n9942 = n9938 ^ n9863 ;
  assign n9943 = n9942 ^ n9860 ;
  assign n9944 = n9943 ^ n9813 ;
  assign n9946 = n9944 ^ n9942 ;
  assign n9868 = n9534 ^ n9490 ;
  assign n9869 = n9868 ^ n9531 ;
  assign n9873 = n9869 ^ n9530 ;
  assign n9874 = n9873 ^ n9531 ;
  assign n9870 = n9869 ^ n9467 ;
  assign n9871 = n9870 ^ n9531 ;
  assign n9919 = n9874 ^ n9871 ;
  assign n9882 = n9534 ^ n9528 ;
  assign n9883 = n9882 ^ n9530 ;
  assign n9881 = n9534 ^ n9467 ;
  assign n9884 = n9883 ^ n9881 ;
  assign n9891 = n9884 ^ n9883 ;
  assign n9888 = n9884 ^ n9530 ;
  assign n9889 = n9888 ^ n9883 ;
  assign n9885 = n9884 ^ n9490 ;
  assign n9890 = n9889 ^ n9885 ;
  assign n9892 = n9891 ^ n9890 ;
  assign n9894 = n9892 ^ n9534 ;
  assign n9899 = n9894 ^ n9891 ;
  assign n9886 = n9885 ^ n9883 ;
  assign n9897 = n9889 ^ n9886 ;
  assign n9900 = n9899 ^ n9897 ;
  assign n9901 = n9883 & ~n9900 ;
  assign n9902 = n9901 ^ n9886 ;
  assign n9903 = n9902 ^ n9891 ;
  assign n9904 = n9903 ^ n9534 ;
  assign n9905 = n9897 ^ n9891 ;
  assign n9906 = n9905 ^ n9534 ;
  assign n9907 = ~n9904 & n9906 ;
  assign n9908 = n9892 ^ n9889 ;
  assign n9909 = n9908 ^ n9894 ;
  assign n9911 = n9894 ^ n9882 ;
  assign n9912 = n9909 & ~n9911 ;
  assign n9913 = n9907 & n9912 ;
  assign n9914 = n9913 ^ n9901 ;
  assign n9915 = n9914 ^ n9897 ;
  assign n9893 = n9892 ^ n9891 ;
  assign n9895 = n9894 ^ n9893 ;
  assign n9916 = n9915 ^ n9895 ;
  assign n9917 = n9916 ^ n9490 ;
  assign n9918 = n9917 ^ n9894 ;
  assign n9920 = n9919 ^ n9918 ;
  assign n9931 = n9920 ^ n9869 ;
  assign n9875 = n9874 ^ n9870 ;
  assign n9877 = n9875 ^ n9868 ;
  assign n9879 = n9877 ^ n9534 ;
  assign n9934 = n9931 ^ n9879 ;
  assign n9947 = n9946 ^ n9934 ;
  assign n9948 = n9947 ^ n9936 ;
  assign n9949 = n9948 ^ n9944 ;
  assign n9859 = n9858 ^ n9857 ;
  assign n9862 = n9861 ^ n9859 ;
  assign n9864 = n9863 ^ n9862 ;
  assign n9866 = n9864 ^ n9534 ;
  assign n9865 = n9864 ^ n9863 ;
  assign n9867 = n9866 ^ n9865 ;
  assign n9950 = n9949 ^ n9867 ;
  assign n9951 = n9950 ^ n9855 ;
  assign n9952 = n9951 ^ n9866 ;
  assign n9962 = n9961 ^ n9952 ;
  assign n9832 = n9490 ^ n9467 ;
  assign n9833 = n9832 ^ n9528 ;
  assign n9818 = n9467 ^ n138 ;
  assign n9834 = n9833 ^ n9818 ;
  assign n9835 = n9834 ^ n9490 ;
  assign n9838 = n9835 ^ n9818 ;
  assign n9840 = n9838 ^ n9530 ;
  assign n9841 = n9840 ^ n9534 ;
  assign n9845 = n9841 ^ n9833 ;
  assign n9839 = n9838 ^ n9534 ;
  assign n9846 = n9845 ^ n9839 ;
  assign n9847 = n9846 ^ n9835 ;
  assign n9849 = n9847 ^ n9845 ;
  assign n9963 = n9962 ^ n9849 ;
  assign n9827 = n9818 ^ n9813 ;
  assign n9824 = n9818 ^ n9490 ;
  assign n9825 = n9824 ^ n9813 ;
  assign n9826 = n9825 ^ n138 ;
  assign n9828 = n9827 ^ n9826 ;
  assign n9830 = n9828 ^ n9531 ;
  assign n9968 = n9963 ^ n9830 ;
  assign n9969 = n183 & ~n9968 ;
  assign n9977 = ~n9490 & ~n9528 ;
  assign n9978 = ~n9883 & n9977 ;
  assign n9979 = n9978 ^ n9882 ;
  assign n10064 = n9979 ^ n9490 ;
  assign n9973 = n130 & ~n9528 ;
  assign n9974 = n9973 ^ n9467 ;
  assign n9975 = ~n183 & ~n9974 ;
  assign n9994 = n9979 ^ n9975 ;
  assign n10065 = n10064 ^ n9994 ;
  assign n10069 = n10065 ^ n9530 ;
  assign n10070 = n10069 ^ n9994 ;
  assign n10066 = n10065 ^ n9467 ;
  assign n10071 = n10070 ^ n10066 ;
  assign n10073 = n10071 ^ n10064 ;
  assign n10074 = n10073 ^ n9979 ;
  assign n9984 = n9530 ^ n9490 ;
  assign n10054 = n9984 ^ n9530 ;
  assign n10049 = n9979 ^ n9467 ;
  assign n10050 = n10049 ^ n9994 ;
  assign n10055 = n10054 ^ n10050 ;
  assign n10052 = n10050 ^ n9984 ;
  assign n10053 = n10052 ^ n9994 ;
  assign n10058 = n10055 ^ n10053 ;
  assign n10059 = n10058 ^ n10049 ;
  assign n10060 = n10059 ^ n9979 ;
  assign n10036 = n9979 ^ n9530 ;
  assign n10037 = n10036 ^ n9994 ;
  assign n10041 = n10037 ^ n9490 ;
  assign n10039 = n10037 ^ n9832 ;
  assign n10040 = n10039 ^ n9994 ;
  assign n10044 = n10041 ^ n10040 ;
  assign n10045 = n10044 ^ n10036 ;
  assign n10046 = n10045 ^ n9979 ;
  assign n10018 = n9979 & ~n9994 ;
  assign n9976 = n9975 ^ n9467 ;
  assign n9995 = n9994 ^ n9976 ;
  assign n10005 = n9995 ^ n9984 ;
  assign n10006 = n10005 ^ n9994 ;
  assign n10019 = n10018 ^ n10006 ;
  assign n10002 = n9995 ^ n9994 ;
  assign n10020 = n10019 ^ n10002 ;
  assign n9999 = n9995 ^ n9490 ;
  assign n10000 = n9999 ^ n9994 ;
  assign n10008 = n10005 ^ n10000 ;
  assign n10009 = n10008 ^ n10002 ;
  assign n10011 = n10009 ^ n9975 ;
  assign n10013 = n10011 ^ n10009 ;
  assign n10021 = n10020 ^ n10013 ;
  assign n10022 = n10002 ^ n9530 ;
  assign n10023 = n10022 ^ n10013 ;
  assign n10024 = ~n10021 & ~n10023 ;
  assign n10025 = n10009 ^ n10000 ;
  assign n10026 = n10025 ^ n10011 ;
  assign n10027 = n10009 ^ n10006 ;
  assign n10028 = n10027 ^ n10011 ;
  assign n10029 = ~n10026 & ~n10028 ;
  assign n10030 = n10024 & n10029 ;
  assign n10031 = n10030 ^ n10018 ;
  assign n10032 = n10031 ^ n9530 ;
  assign n10012 = n10011 ^ n10008 ;
  assign n10033 = n10032 ^ n10012 ;
  assign n10034 = n10033 ^ n9984 ;
  assign n10035 = n10034 ^ n10011 ;
  assign n10047 = n10046 ^ n10035 ;
  assign n9992 = n9530 ^ n9467 ;
  assign n9993 = n9992 ^ n9490 ;
  assign n9996 = n9995 ^ n9993 ;
  assign n10001 = n10000 ^ n9996 ;
  assign n10003 = n10002 ^ n10001 ;
  assign n10004 = n10003 ^ n9975 ;
  assign n10048 = n10047 ^ n10004 ;
  assign n10061 = n10060 ^ n10048 ;
  assign n9985 = n9984 ^ n9467 ;
  assign n10062 = n10061 ^ n9985 ;
  assign n9980 = n9979 ^ n9976 ;
  assign n9989 = n9980 ^ n9979 ;
  assign n9986 = n9985 ^ n9980 ;
  assign n9987 = n9986 ^ n9979 ;
  assign n9981 = n9980 ^ n9530 ;
  assign n9988 = n9987 ^ n9981 ;
  assign n9990 = n9989 ^ n9988 ;
  assign n9991 = n9990 ^ n9975 ;
  assign n10063 = n10062 ^ n9991 ;
  assign n10075 = n10074 ^ n10063 ;
  assign n10076 = n9969 & ~n10075 ;
  assign n10077 = n10076 ^ n10075 ;
  assign n10078 = n9520 ^ n188 ;
  assign n10079 = n9542 & n10078 ;
  assign n10080 = n10079 ^ n9522 ;
  assign n10081 = n10080 ^ n157 ;
  assign n10092 = ~n9515 & n9542 ;
  assign n10093 = n10092 ^ n9517 ;
  assign n9806 = n9502 ^ n401 ;
  assign n9807 = n9542 & n9806 ;
  assign n9808 = n9807 ^ n9504 ;
  assign n9543 = ~n9464 & n9542 ;
  assign n9544 = n9543 ^ n9499 ;
  assign n9545 = n9544 ^ n401 ;
  assign n9546 = n9462 & n9542 ;
  assign n9547 = n9546 ^ n9219 ;
  assign n9548 = n9547 ^ n457 ;
  assign n9549 = n9457 & n9542 ;
  assign n9550 = n9549 ^ n9225 ;
  assign n9551 = n9550 ^ n609 ;
  assign n9552 = ~n9455 & n9542 ;
  assign n9553 = n9552 ^ n9228 ;
  assign n9554 = n9553 ^ n696 ;
  assign n9555 = ~n9434 & n9542 ;
  assign n9556 = n9555 ^ n9436 ;
  assign n9557 = n9556 ^ n1136 ;
  assign n9765 = n9429 & n9542 ;
  assign n9766 = n9765 ^ n9431 ;
  assign n9769 = n9766 ^ n1136 ;
  assign n9754 = ~n9418 & n9542 ;
  assign n9755 = n9754 ^ n9420 ;
  assign n9758 = n9755 ^ n1427 ;
  assign n9558 = n9416 & n9542 ;
  assign n9559 = n9558 ^ n9234 ;
  assign n9560 = n9559 ^ n1739 ;
  assign n9563 = n9406 & n9542 ;
  assign n9564 = n9563 ^ n9409 ;
  assign n9565 = n9564 ^ n2175 ;
  assign n9566 = n9403 ^ n2511 ;
  assign n9567 = n9542 & ~n9566 ;
  assign n9568 = n9567 ^ n9240 ;
  assign n9569 = n9568 ^ n2366 ;
  assign n9738 = ~n9398 & n9542 ;
  assign n9739 = n9738 ^ n9400 ;
  assign n9570 = n9396 & n9542 ;
  assign n9571 = n9570 ^ n9244 ;
  assign n9572 = n9571 ^ n2707 ;
  assign n9573 = ~n9390 & n9542 ;
  assign n9574 = n9573 ^ n9392 ;
  assign n9575 = n9574 ^ n2894 ;
  assign n9728 = n9385 & n9542 ;
  assign n9729 = n9728 ^ n9387 ;
  assign n9732 = n9729 ^ n2894 ;
  assign n9576 = n9383 & n9542 ;
  assign n9577 = n9576 ^ n9247 ;
  assign n9578 = n9577 ^ n3320 ;
  assign n9719 = n9376 ^ n3722 ;
  assign n9720 = n9542 & ~n9719 ;
  assign n9721 = n9720 ^ n9379 ;
  assign n9712 = n9369 ^ n3908 ;
  assign n9713 = n9542 & n9712 ;
  assign n9714 = n9713 ^ n9372 ;
  assign n9706 = n9367 & n9542 ;
  assign n9707 = n9706 ^ n9250 ;
  assign n9579 = n9361 & n9542 ;
  assign n9580 = n9579 ^ n9363 ;
  assign n9581 = n9580 ^ n4153 ;
  assign n9698 = n9355 & n9542 ;
  assign n9699 = n9698 ^ n9358 ;
  assign n9702 = n9699 ^ n4153 ;
  assign n9582 = n9352 & n9542 ;
  assign n9583 = n9582 ^ n9253 ;
  assign n9584 = n9583 ^ n4583 ;
  assign n9587 = n9343 & n9542 ;
  assign n9588 = n9587 ^ n9345 ;
  assign n9589 = n9588 ^ n5073 ;
  assign n9590 = ~n9333 & n9542 ;
  assign n9591 = n9590 ^ n9262 ;
  assign n9678 = n9591 ^ n5562 ;
  assign n9592 = n9591 ^ n5830 ;
  assign n9598 = n9318 & n9542 ;
  assign n9599 = n9598 ^ n9320 ;
  assign n9600 = n9599 ^ n6673 ;
  assign n9601 = ~n9316 & n9542 ;
  assign n9602 = n9601 ^ n9268 ;
  assign n9603 = n9602 ^ n6959 ;
  assign n9606 = ~n9308 & n9542 ;
  assign n9607 = n9606 ^ n9271 ;
  assign n9608 = n9607 ^ n7584 ;
  assign n9609 = n9291 & n9542 ;
  assign n9610 = n9609 ^ n9295 ;
  assign n9611 = n9610 ^ n8253 ;
  assign n9621 = ~x28 & n9217 ;
  assign n9612 = n9273 ^ n9217 ;
  assign n9615 = n9285 ^ x28 ;
  assign n9616 = n9615 ^ n9285 ;
  assign n9617 = n9612 & ~n9616 ;
  assign n9618 = n9617 ^ n9285 ;
  assign n9619 = n9542 & ~n9618 ;
  assign n9620 = n9619 ^ x29 ;
  assign n9622 = n9621 ^ n9620 ;
  assign n9623 = n9622 ^ n8586 ;
  assign n9625 = n9217 ^ x28 ;
  assign n9624 = n9542 & n9612 ;
  assign n9626 = n9625 ^ n9624 ;
  assign n9627 = n9626 ^ n8910 ;
  assign n9629 = n9217 ^ x27 ;
  assign n9630 = n9629 ^ n9542 ;
  assign n9633 = n9217 ^ x26 ;
  assign n9631 = x24 & ~x25 ;
  assign n9632 = n9631 ^ x25 ;
  assign n9634 = n9633 ^ n9632 ;
  assign n9635 = ~n9630 & ~n9634 ;
  assign n9643 = n9635 ^ n9285 ;
  assign n9628 = n9542 ^ n9217 ;
  assign n9636 = n9635 ^ n9628 ;
  assign n9637 = n9636 ^ n9635 ;
  assign n9640 = ~n9629 & n9637 ;
  assign n9641 = n9640 ^ n9635 ;
  assign n9642 = x26 & n9641 ;
  assign n9644 = n9643 ^ n9642 ;
  assign n9645 = n9627 & ~n9644 ;
  assign n9646 = n9645 ^ n9005 ;
  assign n9647 = n9623 & n9646 ;
  assign n9648 = n9647 ^ n8688 ;
  assign n9649 = n9611 & n9648 ;
  assign n9650 = n9649 ^ n8253 ;
  assign n9651 = n9650 ^ n7891 ;
  assign n9652 = n9298 ^ n8253 ;
  assign n9653 = n9542 & n9652 ;
  assign n9654 = n9653 ^ n9304 ;
  assign n9655 = n9654 ^ n9650 ;
  assign n9656 = ~n9651 & n9655 ;
  assign n9657 = n9656 ^ n7971 ;
  assign n9658 = ~n9608 & n9657 ;
  assign n9659 = n9658 ^ n9607 ;
  assign n9604 = ~n9310 & n9542 ;
  assign n9605 = n9604 ^ n9312 ;
  assign n9660 = n9659 ^ n9605 ;
  assign n9661 = n9659 ^ n7277 ;
  assign n9662 = ~n9660 & ~n9661 ;
  assign n9663 = n9662 ^ n7277 ;
  assign n9664 = n9663 ^ n9602 ;
  assign n9665 = ~n9603 & n9664 ;
  assign n9666 = n9665 ^ n7011 ;
  assign n9667 = n9600 & n9666 ;
  assign n9668 = n9667 ^ n6673 ;
  assign n9595 = n9323 ^ n6673 ;
  assign n9596 = n9542 & n9595 ;
  assign n9597 = n9596 ^ n9325 ;
  assign n9669 = n9668 ^ n9597 ;
  assign n9670 = n9668 ^ n6389 ;
  assign n9671 = ~n9669 & ~n9670 ;
  assign n9672 = n9671 ^ n6389 ;
  assign n9593 = ~n9329 & n9542 ;
  assign n9594 = n9593 ^ n9265 ;
  assign n9673 = n9672 ^ n9594 ;
  assign n9674 = n9672 ^ n6115 ;
  assign n9675 = ~n9673 & ~n9674 ;
  assign n9676 = n9675 ^ n6429 ;
  assign n9677 = ~n9592 & ~n9676 ;
  assign n9679 = n9678 ^ n9677 ;
  assign n9680 = n9335 & n9542 ;
  assign n9681 = n9680 ^ n9258 ;
  assign n9682 = n9681 ^ n5562 ;
  assign n9683 = ~n9679 & n9682 ;
  assign n9684 = n9683 ^ n5885 ;
  assign n9685 = n9338 & n9542 ;
  assign n9686 = n9685 ^ n9340 ;
  assign n9687 = n9686 ^ n5317 ;
  assign n9688 = n9684 & ~n9687 ;
  assign n9689 = n9688 ^ n5360 ;
  assign n9690 = n9589 & n9689 ;
  assign n9691 = n9690 ^ n5073 ;
  assign n9585 = n9350 & n9542 ;
  assign n9586 = n9585 ^ n9256 ;
  assign n9692 = n9691 ^ n9586 ;
  assign n9693 = n9691 ^ n4812 ;
  assign n9694 = n9692 & n9693 ;
  assign n9695 = n9694 ^ n4854 ;
  assign n9696 = ~n9584 & n9695 ;
  assign n9697 = n9696 ^ n4645 ;
  assign n9700 = n9699 ^ n4356 ;
  assign n9701 = ~n9697 & ~n9700 ;
  assign n9703 = n9702 ^ n9701 ;
  assign n9704 = n9581 & ~n9703 ;
  assign n9705 = n9704 ^ n4153 ;
  assign n9708 = n9707 ^ n9705 ;
  assign n9709 = n9707 ^ n3908 ;
  assign n9710 = ~n9708 & n9709 ;
  assign n9711 = n9710 ^ n3908 ;
  assign n9715 = n9714 ^ n9711 ;
  assign n9716 = n9714 ^ n3722 ;
  assign n9717 = ~n9715 & ~n9716 ;
  assign n9718 = n9717 ^ n3722 ;
  assign n9722 = n9721 ^ n9718 ;
  assign n9723 = n9721 ^ n3538 ;
  assign n9724 = ~n9722 & n9723 ;
  assign n9725 = n9724 ^ n3596 ;
  assign n9726 = ~n9578 & n9725 ;
  assign n9727 = n9726 ^ n3387 ;
  assign n9730 = n9729 ^ n3093 ;
  assign n9731 = n9727 & ~n9730 ;
  assign n9733 = n9732 ^ n9731 ;
  assign n9734 = n9575 & ~n9733 ;
  assign n9735 = n9734 ^ n3396 ;
  assign n9736 = n9572 & ~n9735 ;
  assign n9737 = n9736 ^ n2707 ;
  assign n9740 = n9739 ^ n9737 ;
  assign n9741 = n9739 ^ n2511 ;
  assign n9742 = n9740 & n9741 ;
  assign n9743 = n9742 ^ n2530 ;
  assign n9744 = n9569 & n9743 ;
  assign n9745 = n9744 ^ n2399 ;
  assign n9746 = n9565 & n9745 ;
  assign n9747 = n9746 ^ n2175 ;
  assign n9561 = n9414 & n9542 ;
  assign n9562 = n9561 ^ n9237 ;
  assign n9748 = n9747 ^ n9562 ;
  assign n9749 = n9747 ^ n2008 ;
  assign n9750 = n9748 & n9749 ;
  assign n9751 = n9750 ^ n2064 ;
  assign n9752 = ~n9560 & ~n9751 ;
  assign n9753 = n9752 ^ n1763 ;
  assign n9756 = n9755 ^ n1572 ;
  assign n9757 = n9753 & ~n9756 ;
  assign n9759 = n9758 ^ n9757 ;
  assign n9760 = ~n9423 & n9542 ;
  assign n9761 = n9760 ^ n9425 ;
  assign n9762 = n9761 ^ n1427 ;
  assign n9763 = n9759 & n9762 ;
  assign n9764 = n9763 ^ n1450 ;
  assign n9767 = n9766 ^ n1290 ;
  assign n9768 = n9764 & n9767 ;
  assign n9770 = n9769 ^ n9768 ;
  assign n9771 = n9557 & n9770 ;
  assign n9772 = n9771 ^ n1143 ;
  assign n9773 = n9440 & n9542 ;
  assign n9774 = n9773 ^ n9231 ;
  assign n9777 = n9774 ^ n1034 ;
  assign n9778 = ~n9772 & n9777 ;
  assign n9775 = n9774 ^ n892 ;
  assign n9779 = n9778 ^ n9775 ;
  assign n9780 = n9442 & n9542 ;
  assign n9781 = n9780 ^ n9444 ;
  assign n9782 = n9781 ^ n786 ;
  assign n9783 = n9782 ^ n927 ;
  assign n9784 = ~n9779 & ~n9783 ;
  assign n9785 = n9784 ^ n9782 ;
  assign n9786 = ~n9449 & n9542 ;
  assign n9787 = n9786 ^ n9451 ;
  assign n9788 = n9787 ^ n696 ;
  assign n9789 = n9788 ^ n842 ;
  assign n9790 = n9785 & ~n9789 ;
  assign n9791 = n9790 ^ n9788 ;
  assign n9792 = ~n9554 & ~n9791 ;
  assign n9793 = n9792 ^ n835 ;
  assign n9794 = n9551 & ~n9793 ;
  assign n9795 = n9794 ^ n834 ;
  assign n9796 = ~n9459 & n9542 ;
  assign n9797 = n9796 ^ n9222 ;
  assign n9798 = n9797 ^ n534 ;
  assign n9799 = ~n9795 & n9798 ;
  assign n9800 = n9799 ^ n750 ;
  assign n9801 = ~n9548 & n9800 ;
  assign n9802 = n9801 ^ n9547 ;
  assign n9803 = n9802 ^ n9544 ;
  assign n9804 = n9545 & ~n9803 ;
  assign n9805 = n9804 ^ n401 ;
  assign n9809 = n9808 ^ n9805 ;
  assign n9810 = n9808 ^ n341 ;
  assign n9811 = ~n9809 & n9810 ;
  assign n9812 = n9811 ^ n349 ;
  assign n10082 = n9508 & n9542 ;
  assign n10083 = n10082 ^ n9496 ;
  assign n10084 = n10083 ^ n291 ;
  assign n10085 = ~n9812 & ~n10084 ;
  assign n10086 = n10085 ^ n307 ;
  assign n10087 = ~n9510 & n9542 ;
  assign n10088 = n10087 ^ n9512 ;
  assign n10089 = n10088 ^ n245 ;
  assign n10090 = n10086 & n10089 ;
  assign n10091 = n10090 ^ n10088 ;
  assign n10094 = n10093 ^ n10091 ;
  assign n10095 = n10093 ^ n188 ;
  assign n10096 = ~n10094 & n10095 ;
  assign n10097 = n10096 ^ n203 ;
  assign n10098 = n10081 & ~n10097 ;
  assign n10099 = n10098 ^ n10080 ;
  assign n10100 = n10099 ^ n138 ;
  assign n10101 = n9526 & n9542 ;
  assign n10102 = n10101 ^ n9492 ;
  assign n10103 = n10102 ^ n10099 ;
  assign n10104 = n10100 & ~n10103 ;
  assign n10105 = n10104 ^ n138 ;
  assign n10106 = n10077 & n10105 ;
  assign n10107 = n9817 & n10106 ;
  assign n10108 = n10107 ^ n10077 ;
  assign n10142 = n9718 ^ n3538 ;
  assign n10143 = ~n10108 & n10142 ;
  assign n10144 = n10143 ^ n9721 ;
  assign n10145 = n10144 ^ n3320 ;
  assign n10146 = n9711 ^ n3722 ;
  assign n10147 = ~n10108 & ~n10146 ;
  assign n10148 = n10147 ^ n9714 ;
  assign n10149 = n10148 ^ n3538 ;
  assign n10154 = n10148 ^ n3722 ;
  assign n10150 = n9705 ^ n3908 ;
  assign n10151 = ~n10108 & n10150 ;
  assign n10152 = n10151 ^ n9707 ;
  assign n10153 = n10152 ^ n10148 ;
  assign n10155 = n10154 ^ n10153 ;
  assign n10156 = ~n9703 & ~n10108 ;
  assign n10157 = n10156 ^ n9580 ;
  assign n10158 = n10157 ^ n3908 ;
  assign n10162 = n10157 ^ n4153 ;
  assign n10159 = n9697 & ~n10108 ;
  assign n10160 = n10159 ^ n9699 ;
  assign n10161 = n10160 ^ n10157 ;
  assign n10163 = n10162 ^ n10161 ;
  assign n10164 = n9695 & ~n10108 ;
  assign n10165 = n10164 ^ n9583 ;
  assign n10166 = n10165 ^ n4356 ;
  assign n10167 = n9693 & ~n10108 ;
  assign n10168 = n10167 ^ n9586 ;
  assign n10169 = n10168 ^ n4583 ;
  assign n10172 = n9689 & ~n10108 ;
  assign n10173 = n10172 ^ n9588 ;
  assign n10175 = n10173 ^ n5073 ;
  assign n10170 = n9684 & ~n10108 ;
  assign n10171 = n10170 ^ n9686 ;
  assign n10174 = n10173 ^ n10171 ;
  assign n10176 = n10175 ^ n10174 ;
  assign n10177 = ~n9679 & ~n10108 ;
  assign n10178 = n10177 ^ n9681 ;
  assign n10179 = n10178 ^ n5317 ;
  assign n10182 = ~n9674 & ~n10108 ;
  assign n10183 = n10182 ^ n9594 ;
  assign n10184 = n10183 ^ n5830 ;
  assign n10185 = n9663 ^ n6959 ;
  assign n10186 = ~n10108 & n10185 ;
  assign n10187 = n10186 ^ n9602 ;
  assign n10188 = n10187 ^ n6673 ;
  assign n10189 = ~n9661 & ~n10108 ;
  assign n10190 = n10189 ^ n9605 ;
  assign n10191 = n10190 ^ n6959 ;
  assign n10192 = ~n9651 & ~n10108 ;
  assign n10193 = n10192 ^ n9654 ;
  assign n10194 = n10193 ^ n7584 ;
  assign n10195 = ~n9644 & ~n10108 ;
  assign n10196 = n10195 ^ n9626 ;
  assign n10197 = n10196 ^ n8586 ;
  assign n10236 = ~n9631 & ~n10108 ;
  assign n10209 = ~x22 & ~x23 ;
  assign n10210 = ~x24 & n10209 ;
  assign n10211 = n10210 ^ x25 ;
  assign n10233 = n10211 ^ n10108 ;
  assign n10234 = n10210 ^ n9542 ;
  assign n10235 = n10233 & ~n10234 ;
  assign n10237 = n10236 ^ n10235 ;
  assign n10238 = n10237 ^ x25 ;
  assign n10230 = n9632 ^ n9542 ;
  assign n10231 = ~n10108 & ~n10230 ;
  assign n10212 = n9542 ^ x26 ;
  assign n10232 = n10231 ^ n10212 ;
  assign n10239 = n10238 ^ n10232 ;
  assign n10208 = n10108 ^ x25 ;
  assign n10215 = n9542 & n10212 ;
  assign n10216 = n10211 & n10215 ;
  assign n10217 = ~n10208 & n10216 ;
  assign n10218 = n10217 ^ n10215 ;
  assign n10199 = x26 & n10108 ;
  assign n10198 = n10108 ^ x26 ;
  assign n10200 = n10199 ^ n10198 ;
  assign n10201 = ~n9632 & ~n10200 ;
  assign n10213 = n10212 ^ n10201 ;
  assign n10219 = n10218 ^ n10213 ;
  assign n10220 = n10210 ^ n10198 ;
  assign n10223 = n10208 & n10220 ;
  assign n10224 = n10223 ^ n10198 ;
  assign n10225 = n10219 & n10224 ;
  assign n10227 = ~x26 & n10108 ;
  assign n10228 = n10225 & n10227 ;
  assign n10226 = n10225 ^ n10219 ;
  assign n10229 = n10228 ^ n10226 ;
  assign n10240 = n10239 ^ n10229 ;
  assign n10241 = n9217 & ~n10229 ;
  assign n10242 = n10240 & n10241 ;
  assign n10243 = n10242 ^ n10240 ;
  assign n10206 = ~n9217 & ~n10108 ;
  assign n10203 = n10108 ^ n9542 ;
  assign n10204 = ~n10199 & ~n10203 ;
  assign n10202 = n10201 ^ x27 ;
  assign n10205 = n10204 ^ n10202 ;
  assign n10207 = n10206 ^ n10205 ;
  assign n10244 = n10243 ^ n10207 ;
  assign n10245 = n10207 ^ n8910 ;
  assign n10246 = ~n10244 & n10245 ;
  assign n10247 = n10246 ^ n9005 ;
  assign n10248 = n10197 & n10247 ;
  assign n10249 = n10248 ^ n8688 ;
  assign n10250 = n9646 & ~n10108 ;
  assign n10251 = n10250 ^ n9622 ;
  assign n10252 = n10251 ^ n8253 ;
  assign n10253 = n10249 & n10252 ;
  assign n10254 = n10253 ^ n8356 ;
  assign n10255 = n9648 & ~n10108 ;
  assign n10256 = n10255 ^ n9610 ;
  assign n10257 = n10256 ^ n7891 ;
  assign n10258 = ~n10254 & ~n10257 ;
  assign n10259 = n10258 ^ n7971 ;
  assign n10260 = ~n10194 & ~n10259 ;
  assign n10261 = n10260 ^ n7660 ;
  assign n10262 = ~n9657 & ~n10108 ;
  assign n10263 = n10262 ^ n9607 ;
  assign n10264 = n10263 ^ n7277 ;
  assign n10265 = n10261 & ~n10264 ;
  assign n10266 = n10265 ^ n7277 ;
  assign n10267 = n10266 ^ n10190 ;
  assign n10268 = ~n10191 & n10267 ;
  assign n10269 = n10268 ^ n6959 ;
  assign n10270 = n10269 ^ n10187 ;
  assign n10271 = ~n10188 & n10270 ;
  assign n10272 = n10271 ^ n6673 ;
  assign n10273 = n10272 ^ n6389 ;
  assign n10274 = n9666 & ~n10108 ;
  assign n10275 = n10274 ^ n9599 ;
  assign n10276 = n10275 ^ n10272 ;
  assign n10277 = ~n10273 & ~n10276 ;
  assign n10278 = n10277 ^ n6423 ;
  assign n10279 = ~n9670 & ~n10108 ;
  assign n10280 = n10279 ^ n9597 ;
  assign n10281 = n10280 ^ n6115 ;
  assign n10282 = ~n10278 & n10281 ;
  assign n10283 = n10282 ^ n6429 ;
  assign n10284 = ~n10184 & ~n10283 ;
  assign n10285 = n10284 ^ n10183 ;
  assign n10180 = n9676 & ~n10108 ;
  assign n10181 = n10180 ^ n9591 ;
  assign n10286 = n10285 ^ n10181 ;
  assign n10287 = n10285 ^ n5562 ;
  assign n10288 = ~n10286 & ~n10287 ;
  assign n10289 = n10288 ^ n5885 ;
  assign n10290 = n10179 & ~n10289 ;
  assign n10291 = n10290 ^ n10178 ;
  assign n10292 = n10291 ^ n10173 ;
  assign n10293 = n10292 ^ n10175 ;
  assign n10294 = ~n10176 & n10293 ;
  assign n10295 = n10294 ^ n10175 ;
  assign n10297 = n10168 ^ n4812 ;
  assign n10296 = n10173 ^ n10168 ;
  assign n10298 = n10297 ^ n10296 ;
  assign n10299 = ~n10295 & n10298 ;
  assign n10300 = n10299 ^ n10297 ;
  assign n10301 = ~n10169 & n10300 ;
  assign n10302 = n10301 ^ n4645 ;
  assign n10303 = ~n10166 & ~n10302 ;
  assign n10304 = n10303 ^ n10165 ;
  assign n10305 = n10304 ^ n10157 ;
  assign n10306 = n10305 ^ n10162 ;
  assign n10307 = ~n10163 & ~n10306 ;
  assign n10308 = n10307 ^ n10162 ;
  assign n10309 = n10158 & ~n10308 ;
  assign n10310 = n10309 ^ n3908 ;
  assign n10311 = n10310 ^ n10148 ;
  assign n10312 = n10311 ^ n10154 ;
  assign n10313 = ~n10155 & ~n10312 ;
  assign n10314 = n10313 ^ n10154 ;
  assign n10315 = ~n10149 & n10314 ;
  assign n10316 = n10315 ^ n3538 ;
  assign n10317 = n10316 ^ n10144 ;
  assign n10318 = n10145 & ~n10317 ;
  assign n10319 = n10318 ^ n3387 ;
  assign n10422 = n10100 & ~n10108 ;
  assign n10423 = n10422 ^ n10102 ;
  assign n10424 = n183 & n10423 ;
  assign n10425 = n10424 ^ n183 ;
  assign n10426 = n183 & n10105 ;
  assign n10427 = ~n1355 & ~n10099 ;
  assign n10428 = ~n10077 & ~n10102 ;
  assign n10429 = n10427 & n10428 ;
  assign n10430 = n10429 ^ n9815 ;
  assign n10431 = n10430 ^ n10077 ;
  assign n10432 = n10431 ^ n10430 ;
  assign n10433 = n10430 ^ n9817 ;
  assign n10434 = n10433 ^ n10430 ;
  assign n10435 = ~n10432 & ~n10434 ;
  assign n10436 = n10435 ^ n10430 ;
  assign n10437 = n10426 & n10436 ;
  assign n10438 = n10437 ^ n10430 ;
  assign n10439 = n10099 ^ n10077 ;
  assign n10440 = ~n10428 & n10439 ;
  assign n10441 = n10440 ^ n138 ;
  assign n10442 = n10102 ^ n10100 ;
  assign n10443 = n10442 ^ n10077 ;
  assign n10444 = n10441 & ~n10443 ;
  assign n10445 = n10444 ^ n10077 ;
  assign n10446 = n9816 & ~n10445 ;
  assign n10447 = ~n10438 & n10446 ;
  assign n10448 = n10447 ^ n10438 ;
  assign n10449 = n10091 ^ n188 ;
  assign n10450 = ~n10108 & n10449 ;
  assign n10451 = n10450 ^ n10093 ;
  assign n10452 = n10451 ^ n157 ;
  assign n10109 = ~n9812 & ~n10108 ;
  assign n10110 = n10109 ^ n10083 ;
  assign n10111 = n10110 ^ n245 ;
  assign n10112 = n9805 ^ n341 ;
  assign n10113 = ~n10108 & n10112 ;
  assign n10114 = n10113 ^ n9808 ;
  assign n10115 = n10114 ^ n291 ;
  assign n10405 = ~n9800 & ~n10108 ;
  assign n10406 = n10405 ^ n9547 ;
  assign n10121 = ~n9795 & ~n10108 ;
  assign n10122 = n10121 ^ n9797 ;
  assign n10123 = n10122 ^ n457 ;
  assign n10124 = ~n9793 & ~n10108 ;
  assign n10125 = n10124 ^ n9550 ;
  assign n10126 = n10125 ^ n534 ;
  assign n10127 = ~n9791 & ~n10108 ;
  assign n10128 = n10127 ^ n9553 ;
  assign n10129 = n10128 ^ n609 ;
  assign n10368 = ~n9764 & ~n10108 ;
  assign n10369 = n10368 ^ n9766 ;
  assign n10352 = ~n9751 & ~n10108 ;
  assign n10353 = n10352 ^ n9559 ;
  assign n10356 = n10353 ^ n1427 ;
  assign n10130 = n9743 & ~n10108 ;
  assign n10131 = n10130 ^ n9568 ;
  assign n10132 = n10131 ^ n2175 ;
  assign n10133 = ~n9735 & ~n10108 ;
  assign n10134 = n10133 ^ n9571 ;
  assign n10135 = n10134 ^ n2511 ;
  assign n10136 = ~n9733 & ~n10108 ;
  assign n10137 = n10136 ^ n9574 ;
  assign n10138 = n10137 ^ n2707 ;
  assign n10139 = ~n9727 & ~n10108 ;
  assign n10140 = n10139 ^ n9729 ;
  assign n10141 = n10140 ^ n2894 ;
  assign n10320 = n9725 & ~n10108 ;
  assign n10321 = n10320 ^ n9577 ;
  assign n10324 = n10321 ^ n2894 ;
  assign n10322 = n10321 ^ n3093 ;
  assign n10323 = n10319 & n10322 ;
  assign n10325 = n10324 ^ n10323 ;
  assign n10326 = ~n10141 & n10325 ;
  assign n10327 = n10326 ^ n3396 ;
  assign n10328 = ~n10138 & ~n10327 ;
  assign n10329 = n10328 ^ n2707 ;
  assign n10330 = n10329 ^ n10134 ;
  assign n10331 = ~n10135 & ~n10330 ;
  assign n10332 = n10331 ^ n2530 ;
  assign n10333 = n9737 ^ n2511 ;
  assign n10334 = ~n10108 & ~n10333 ;
  assign n10335 = n10334 ^ n9739 ;
  assign n10336 = n10335 ^ n2366 ;
  assign n10337 = n10332 & n10336 ;
  assign n10338 = n10337 ^ n2399 ;
  assign n10339 = n10132 & n10338 ;
  assign n10340 = n10339 ^ n2204 ;
  assign n10341 = n9745 & ~n10108 ;
  assign n10342 = n10341 ^ n9564 ;
  assign n10343 = n10342 ^ n2008 ;
  assign n10344 = n10340 & n10343 ;
  assign n10345 = n10344 ^ n2008 ;
  assign n10346 = n10345 ^ n1739 ;
  assign n10347 = n9749 & ~n10108 ;
  assign n10348 = n10347 ^ n9562 ;
  assign n10349 = n10348 ^ n10345 ;
  assign n10350 = ~n10346 & n10349 ;
  assign n10351 = n10350 ^ n1763 ;
  assign n10354 = n10353 ^ n1572 ;
  assign n10355 = n10351 & n10354 ;
  assign n10357 = n10356 ^ n10355 ;
  assign n10358 = ~n9753 & ~n10108 ;
  assign n10359 = n10358 ^ n9755 ;
  assign n10360 = n10359 ^ n1427 ;
  assign n10361 = ~n10357 & n10360 ;
  assign n10362 = n10361 ^ n1450 ;
  assign n10363 = n9759 & ~n10108 ;
  assign n10364 = n10363 ^ n9761 ;
  assign n10365 = n10364 ^ n1290 ;
  assign n10366 = n10362 & ~n10365 ;
  assign n10367 = n10366 ^ n10364 ;
  assign n10370 = n10369 ^ n10367 ;
  assign n10371 = n10369 ^ n1136 ;
  assign n10372 = n10370 & n10371 ;
  assign n10373 = n10372 ^ n1143 ;
  assign n10374 = n9770 & ~n10108 ;
  assign n10375 = n10374 ^ n9556 ;
  assign n10378 = n10375 ^ n1034 ;
  assign n10379 = ~n10373 & n10378 ;
  assign n10376 = n10375 ^ n892 ;
  assign n10380 = n10379 ^ n10376 ;
  assign n10381 = n9772 & ~n10108 ;
  assign n10382 = n10381 ^ n9774 ;
  assign n10383 = n10382 ^ n786 ;
  assign n10384 = n10383 ^ n927 ;
  assign n10385 = ~n10380 & n10384 ;
  assign n10386 = n10385 ^ n10383 ;
  assign n10387 = n9779 & ~n10108 ;
  assign n10388 = n10387 ^ n9781 ;
  assign n10389 = n10388 ^ n696 ;
  assign n10390 = n10389 ^ n842 ;
  assign n10391 = ~n10386 & ~n10390 ;
  assign n10392 = n10391 ^ n10389 ;
  assign n10393 = ~n9785 & ~n10108 ;
  assign n10394 = n10393 ^ n9787 ;
  assign n10395 = n10394 ^ n609 ;
  assign n10396 = n10395 ^ n835 ;
  assign n10397 = n10392 & ~n10396 ;
  assign n10398 = n10397 ^ n10395 ;
  assign n10399 = n10129 & n10398 ;
  assign n10400 = n10399 ^ n834 ;
  assign n10401 = ~n10126 & ~n10400 ;
  assign n10402 = n10401 ^ n750 ;
  assign n10403 = ~n10123 & n10402 ;
  assign n10404 = n10403 ^ n10122 ;
  assign n10407 = n10406 ^ n10404 ;
  assign n10408 = n10406 ^ n401 ;
  assign n10409 = ~n10407 & n10408 ;
  assign n10410 = n10409 ^ n401 ;
  assign n10119 = n10114 ^ n341 ;
  assign n10116 = n9802 ^ n401 ;
  assign n10117 = ~n10108 & n10116 ;
  assign n10118 = n10117 ^ n9544 ;
  assign n10120 = n10119 ^ n10118 ;
  assign n10411 = n10410 ^ n10120 ;
  assign n10412 = n10411 ^ n10119 ;
  assign n10413 = n10118 ^ n10114 ;
  assign n10414 = n10413 ^ n10119 ;
  assign n10415 = ~n10412 & n10414 ;
  assign n10416 = n10415 ^ n10119 ;
  assign n10417 = ~n10115 & ~n10416 ;
  assign n10418 = n10417 ^ n307 ;
  assign n10419 = n10111 & n10418 ;
  assign n10420 = n10419 ^ n10110 ;
  assign n10421 = n10420 ^ n188 ;
  assign n10453 = ~n10086 & ~n10108 ;
  assign n10454 = n10453 ^ n10088 ;
  assign n10455 = n10454 ^ n10420 ;
  assign n10456 = n10421 & ~n10455 ;
  assign n10457 = n10456 ^ n203 ;
  assign n10458 = n10452 & ~n10457 ;
  assign n10459 = n10458 ^ n10451 ;
  assign n10460 = n10459 ^ n138 ;
  assign n10461 = n10097 & ~n10108 ;
  assign n10462 = n10461 ^ n10080 ;
  assign n10463 = n10462 ^ n10459 ;
  assign n10464 = n10460 & ~n10463 ;
  assign n10465 = n10464 ^ n138 ;
  assign n10466 = ~n10448 & n10465 ;
  assign n10467 = ~n10425 & n10466 ;
  assign n10468 = n10467 ^ n10448 ;
  assign n10516 = ~n10319 & n10468 ;
  assign n10517 = n10516 ^ n10321 ;
  assign n10518 = n10517 ^ n2894 ;
  assign n10519 = n10310 ^ n3538 ;
  assign n10520 = n10519 ^ n3795 ;
  assign n10521 = n10152 ^ n3538 ;
  assign n10522 = n10521 ^ n3795 ;
  assign n10523 = ~n10520 & ~n10522 ;
  assign n10524 = n10523 ^ n3795 ;
  assign n10525 = n10468 & n10524 ;
  assign n10526 = n10525 ^ n10148 ;
  assign n10527 = n10526 ^ n3320 ;
  assign n10528 = n10310 ^ n3722 ;
  assign n10529 = n10468 & ~n10528 ;
  assign n10530 = n10529 ^ n10152 ;
  assign n10531 = n10530 ^ n3538 ;
  assign n10532 = n10304 ^ n3908 ;
  assign n10533 = n10532 ^ n4194 ;
  assign n10534 = n10160 ^ n3908 ;
  assign n10535 = n10534 ^ n4194 ;
  assign n10536 = ~n10533 & ~n10535 ;
  assign n10537 = n10536 ^ n4194 ;
  assign n10538 = n10468 & n10537 ;
  assign n10539 = n10538 ^ n10157 ;
  assign n10540 = n10539 ^ n3722 ;
  assign n10713 = n10304 ^ n4153 ;
  assign n10714 = n10468 & ~n10713 ;
  assign n10715 = n10714 ^ n10160 ;
  assign n10546 = n4812 & n10173 ;
  assign n10541 = n5073 & ~n10171 ;
  assign n10542 = ~n10291 & ~n10541 ;
  assign n10543 = n10171 ^ n5073 ;
  assign n10544 = n10543 ^ n10541 ;
  assign n10545 = n10173 ^ n4812 ;
  assign n10547 = n10546 ^ n10545 ;
  assign n10548 = ~n10544 & n10547 ;
  assign n10549 = ~n10542 & n10548 ;
  assign n10554 = ~n10546 & ~n10549 ;
  assign n10555 = n10554 ^ n10168 ;
  assign n10556 = ~n10169 & ~n10555 ;
  assign n10557 = n10556 ^ n4645 ;
  assign n10558 = n10468 & n10557 ;
  assign n10559 = n10558 ^ n10165 ;
  assign n10560 = n10559 ^ n4153 ;
  assign n10573 = ~n10542 & ~n10544 ;
  assign n10574 = n10573 ^ n4812 ;
  assign n10575 = n10468 & n10574 ;
  assign n10576 = n10575 ^ n10173 ;
  assign n10577 = n10576 ^ n4583 ;
  assign n10578 = n10289 & n10468 ;
  assign n10579 = n10578 ^ n10178 ;
  assign n10580 = n10579 ^ n5073 ;
  assign n10581 = ~n10287 & n10468 ;
  assign n10582 = n10581 ^ n10181 ;
  assign n10584 = n10582 ^ n5317 ;
  assign n10587 = ~n10278 & n10468 ;
  assign n10588 = n10587 ^ n10280 ;
  assign n10589 = n10588 ^ n5830 ;
  assign n10590 = n10269 ^ n6673 ;
  assign n10591 = n10468 & n10590 ;
  assign n10592 = n10591 ^ n10187 ;
  assign n10593 = n10592 ^ n6389 ;
  assign n10674 = n10266 ^ n6959 ;
  assign n10675 = n10468 & n10674 ;
  assign n10676 = n10675 ^ n10190 ;
  assign n10594 = n10261 & n10468 ;
  assign n10595 = n10594 ^ n10263 ;
  assign n10596 = n10595 ^ n6959 ;
  assign n10666 = ~n10259 & n10468 ;
  assign n10667 = n10666 ^ n10193 ;
  assign n10597 = ~n10254 & n10468 ;
  assign n10598 = n10597 ^ n10256 ;
  assign n10599 = n10598 ^ n7584 ;
  assign n10600 = n10249 & n10468 ;
  assign n10601 = n10600 ^ n10251 ;
  assign n10602 = n10601 ^ n7891 ;
  assign n10656 = n10247 & n10468 ;
  assign n10657 = n10656 ^ n10196 ;
  assign n10603 = n10243 ^ n8910 ;
  assign n10604 = n10468 & n10603 ;
  assign n10605 = n10604 ^ n10207 ;
  assign n10606 = n10605 ^ n8586 ;
  assign n10617 = n10234 ^ x25 ;
  assign n10618 = n10617 ^ n10108 ;
  assign n10610 = n10234 ^ n10108 ;
  assign n10611 = n10610 ^ n10234 ;
  assign n10614 = x24 & ~n10611 ;
  assign n10615 = n10614 ^ n10234 ;
  assign n10616 = ~n10468 & n10615 ;
  assign n10619 = n10618 ^ n10616 ;
  assign n10620 = n10619 ^ n9217 ;
  assign n10622 = n10209 ^ n10108 ;
  assign n10623 = ~n10468 & ~n10622 ;
  assign n10621 = n10209 ^ x24 ;
  assign n10624 = n10623 ^ n10621 ;
  assign n10625 = n10624 ^ n9542 ;
  assign n10634 = n9542 ^ x23 ;
  assign n10626 = n10468 ^ x23 ;
  assign n10627 = n10626 ^ n10108 ;
  assign n10628 = x20 & ~x21 ;
  assign n10629 = n10628 ^ x21 ;
  assign n10630 = n10629 ^ x22 ;
  assign n10631 = n10630 ^ n10108 ;
  assign n10632 = n10627 & n10631 ;
  assign n10633 = n10632 ^ n10203 ;
  assign n10635 = n10634 ^ n10633 ;
  assign n10636 = n10635 ^ x23 ;
  assign n10637 = n10636 ^ n10108 ;
  assign n10638 = n10637 ^ n10635 ;
  assign n10639 = n10468 ^ n10108 ;
  assign n10642 = n10638 & n10639 ;
  assign n10643 = n10642 ^ n10635 ;
  assign n10644 = x22 & n10643 ;
  assign n10645 = n10644 ^ n10633 ;
  assign n10646 = ~n10625 & ~n10645 ;
  assign n10647 = n10646 ^ n9628 ;
  assign n10648 = n10620 & n10647 ;
  assign n10649 = n10648 ^ n9217 ;
  assign n10607 = n10238 ^ n9217 ;
  assign n10608 = n10468 & ~n10607 ;
  assign n10609 = n10608 ^ n10232 ;
  assign n10650 = n10649 ^ n10609 ;
  assign n10651 = n10609 ^ n8910 ;
  assign n10652 = n10650 & n10651 ;
  assign n10653 = n10652 ^ n9005 ;
  assign n10654 = n10606 & n10653 ;
  assign n10655 = n10654 ^ n8586 ;
  assign n10658 = n10657 ^ n10655 ;
  assign n10659 = n10657 ^ n8253 ;
  assign n10660 = ~n10658 & n10659 ;
  assign n10661 = n10660 ^ n8356 ;
  assign n10662 = ~n10602 & ~n10661 ;
  assign n10663 = n10662 ^ n7971 ;
  assign n10664 = n10599 & n10663 ;
  assign n10665 = n10664 ^ n10598 ;
  assign n10668 = n10667 ^ n10665 ;
  assign n10669 = n10667 ^ n7277 ;
  assign n10670 = n10668 & ~n10669 ;
  assign n10671 = n10670 ^ n7339 ;
  assign n10672 = ~n10596 & n10671 ;
  assign n10673 = n10672 ^ n6959 ;
  assign n10677 = n10676 ^ n10673 ;
  assign n10678 = n10676 ^ n6673 ;
  assign n10679 = n10677 & ~n10678 ;
  assign n10680 = n10679 ^ n6713 ;
  assign n10681 = n10593 & ~n10680 ;
  assign n10682 = n10681 ^ n6423 ;
  assign n10683 = ~n10273 & n10468 ;
  assign n10684 = n10683 ^ n10275 ;
  assign n10685 = n10684 ^ n6115 ;
  assign n10686 = ~n10682 & n10685 ;
  assign n10687 = n10686 ^ n6429 ;
  assign n10688 = n10589 & ~n10687 ;
  assign n10689 = n10688 ^ n10588 ;
  assign n10585 = n10283 & n10468 ;
  assign n10586 = n10585 ^ n10183 ;
  assign n10690 = n10689 ^ n10586 ;
  assign n10691 = n10689 ^ n5562 ;
  assign n10692 = n10690 & n10691 ;
  assign n10693 = n10692 ^ n5885 ;
  assign n10694 = ~n10584 & ~n10693 ;
  assign n10583 = n10582 ^ n5073 ;
  assign n10695 = n10694 ^ n10583 ;
  assign n10696 = n10580 & ~n10695 ;
  assign n10697 = n10696 ^ n5073 ;
  assign n10698 = n10697 ^ n4812 ;
  assign n10699 = n10291 ^ n5073 ;
  assign n10700 = n10468 & n10699 ;
  assign n10701 = n10700 ^ n10171 ;
  assign n10702 = n10701 ^ n10697 ;
  assign n10703 = n10698 & n10702 ;
  assign n10704 = n10703 ^ n4854 ;
  assign n10705 = n10577 & n10704 ;
  assign n10706 = n10705 ^ n4583 ;
  assign n10566 = n10554 ^ n4583 ;
  assign n10567 = n10468 & ~n10566 ;
  assign n10568 = n10567 ^ n10168 ;
  assign n10707 = n10706 ^ n10568 ;
  assign n10708 = n10568 ^ n4356 ;
  assign n10709 = n10707 & ~n10708 ;
  assign n10710 = n10709 ^ n4414 ;
  assign n10711 = ~n10560 & n10710 ;
  assign n10712 = n10711 ^ n4153 ;
  assign n10716 = n10715 ^ n10712 ;
  assign n10717 = n10715 ^ n3908 ;
  assign n10718 = n10716 & ~n10717 ;
  assign n10719 = n10718 ^ n3961 ;
  assign n10720 = ~n10540 & ~n10719 ;
  assign n10721 = n10720 ^ n3795 ;
  assign n10722 = ~n10531 & n10721 ;
  assign n10723 = n10722 ^ n3538 ;
  assign n10724 = n10723 ^ n10526 ;
  assign n10725 = ~n10527 & n10724 ;
  assign n10726 = n10725 ^ n3387 ;
  assign n10727 = n10316 ^ n3320 ;
  assign n10728 = n10468 & n10727 ;
  assign n10729 = n10728 ^ n10144 ;
  assign n10730 = n10729 ^ n3093 ;
  assign n10731 = ~n10726 & ~n10730 ;
  assign n10732 = n10731 ^ n3363 ;
  assign n10733 = n10518 & n10732 ;
  assign n10734 = n10733 ^ n3396 ;
  assign n10826 = n10460 & n10468 ;
  assign n10827 = n10826 ^ n10462 ;
  assign n10828 = n10827 ^ n183 ;
  assign n10831 = n10459 ^ n130 ;
  assign n10832 = n10462 & ~n10831 ;
  assign n10830 = n5787 & ~n10459 ;
  assign n10833 = n10832 ^ n10830 ;
  assign n10835 = n10833 ^ n10459 ;
  assign n10834 = n10833 ^ n10438 ;
  assign n10836 = n10835 ^ n10834 ;
  assign n10837 = n10835 ^ n10830 ;
  assign n10838 = n10837 ^ n10835 ;
  assign n10839 = n10836 & ~n10838 ;
  assign n10840 = n10839 ^ n10835 ;
  assign n10841 = n183 & ~n10840 ;
  assign n10842 = n10841 ^ n10833 ;
  assign n10843 = ~n10423 & n10842 ;
  assign n10829 = n10424 & n10465 ;
  assign n10844 = n10843 ^ n10829 ;
  assign n10845 = ~n10462 & ~n10844 ;
  assign n10849 = n10459 ^ n183 ;
  assign n10846 = n10448 ^ n10423 ;
  assign n10850 = n10849 ^ n10846 ;
  assign n10851 = n10850 ^ n138 ;
  assign n10858 = ~n10846 & ~n10851 ;
  assign n10861 = n10858 ^ n10423 ;
  assign n10862 = n10849 & ~n10861 ;
  assign n10852 = n10851 ^ n10448 ;
  assign n10853 = n10852 ^ n10846 ;
  assign n10859 = n10858 ^ n10853 ;
  assign n10860 = n10859 ^ n10858 ;
  assign n10863 = n10862 ^ n10860 ;
  assign n10864 = ~n10460 & n10863 ;
  assign n10865 = n10864 ^ n10859 ;
  assign n10866 = n10845 & n10865 ;
  assign n10867 = n10866 ^ n10844 ;
  assign n10469 = n10421 & n10468 ;
  assign n10470 = n10469 ^ n10454 ;
  assign n10471 = n10470 ^ n157 ;
  assign n10474 = n10410 ^ n291 ;
  assign n10475 = n10474 ^ n349 ;
  assign n10476 = n10118 ^ n291 ;
  assign n10477 = n10476 ^ n349 ;
  assign n10478 = n10475 & n10477 ;
  assign n10479 = n10478 ^ n349 ;
  assign n10480 = n10468 & ~n10479 ;
  assign n10481 = n10480 ^ n10114 ;
  assign n10482 = n10481 ^ n245 ;
  assign n10483 = n10404 ^ n401 ;
  assign n10484 = n10468 & n10483 ;
  assign n10485 = n10484 ^ n10406 ;
  assign n10486 = n10485 ^ n341 ;
  assign n10803 = ~n10402 & n10468 ;
  assign n10804 = n10803 ^ n10122 ;
  assign n10487 = ~n10400 & n10468 ;
  assign n10488 = n10487 ^ n10125 ;
  assign n10489 = n10488 ^ n457 ;
  assign n10490 = ~n10392 & n10468 ;
  assign n10491 = n10490 ^ n10394 ;
  assign n10492 = n10491 ^ n609 ;
  assign n10493 = ~n10362 & n10468 ;
  assign n10494 = n10493 ^ n10364 ;
  assign n10495 = n10494 ^ n1136 ;
  assign n10760 = ~n10357 & n10468 ;
  assign n10761 = n10760 ^ n10359 ;
  assign n10764 = n10761 ^ n1136 ;
  assign n10496 = ~n10351 & n10468 ;
  assign n10497 = n10496 ^ n10353 ;
  assign n10498 = n10497 ^ n1427 ;
  assign n10501 = n10340 & n10468 ;
  assign n10502 = n10501 ^ n10342 ;
  assign n10503 = n10502 ^ n1739 ;
  assign n10506 = n10332 & n10468 ;
  assign n10507 = n10506 ^ n10335 ;
  assign n10508 = n10507 ^ n2175 ;
  assign n10509 = n10329 ^ n2511 ;
  assign n10510 = n10468 & ~n10509 ;
  assign n10511 = n10510 ^ n10134 ;
  assign n10512 = n10511 ^ n2366 ;
  assign n10737 = ~n10327 & n10468 ;
  assign n10738 = n10737 ^ n10137 ;
  assign n10513 = n10325 & n10468 ;
  assign n10514 = n10513 ^ n10140 ;
  assign n10515 = n10514 ^ n2707 ;
  assign n10735 = n10515 & ~n10734 ;
  assign n10736 = n10735 ^ n2707 ;
  assign n10739 = n10738 ^ n10736 ;
  assign n10740 = n10738 ^ n2511 ;
  assign n10741 = n10739 & n10740 ;
  assign n10742 = n10741 ^ n2530 ;
  assign n10743 = ~n10512 & n10742 ;
  assign n10744 = n10743 ^ n2399 ;
  assign n10745 = n10508 & n10744 ;
  assign n10746 = n10745 ^ n2175 ;
  assign n10504 = n10338 & n10468 ;
  assign n10505 = n10504 ^ n10131 ;
  assign n10747 = n10746 ^ n10505 ;
  assign n10748 = n10746 ^ n2008 ;
  assign n10749 = ~n10747 & n10748 ;
  assign n10750 = n10749 ^ n2064 ;
  assign n10751 = ~n10503 & ~n10750 ;
  assign n10752 = n10751 ^ n1739 ;
  assign n10756 = n10752 ^ n1427 ;
  assign n10499 = ~n10346 & n10468 ;
  assign n10500 = n10499 ^ n10348 ;
  assign n10753 = n10752 ^ n10500 ;
  assign n10754 = n10500 ^ n1572 ;
  assign n10755 = n10753 & n10754 ;
  assign n10757 = n10756 ^ n10755 ;
  assign n10758 = ~n10498 & n10757 ;
  assign n10759 = n10758 ^ n1450 ;
  assign n10762 = n10761 ^ n1290 ;
  assign n10763 = n10759 & ~n10762 ;
  assign n10765 = n10764 ^ n10763 ;
  assign n10766 = ~n10495 & ~n10765 ;
  assign n10767 = n10766 ^ n1143 ;
  assign n10768 = n10367 ^ n1136 ;
  assign n10769 = n10468 & ~n10768 ;
  assign n10770 = n10769 ^ n10369 ;
  assign n10773 = n10770 ^ n1034 ;
  assign n10774 = ~n10767 & n10773 ;
  assign n10771 = n10770 ^ n892 ;
  assign n10775 = n10774 ^ n10771 ;
  assign n10776 = n10373 & n10468 ;
  assign n10777 = n10776 ^ n10375 ;
  assign n10778 = n10777 ^ n786 ;
  assign n10779 = n10778 ^ n927 ;
  assign n10780 = ~n10775 & n10779 ;
  assign n10781 = n10780 ^ n10778 ;
  assign n10782 = n10380 & n10468 ;
  assign n10783 = n10782 ^ n10382 ;
  assign n10784 = n10783 ^ n696 ;
  assign n10785 = n10784 ^ n842 ;
  assign n10786 = ~n10781 & n10785 ;
  assign n10787 = n10786 ^ n10784 ;
  assign n10788 = n10386 & n10468 ;
  assign n10789 = n10788 ^ n10388 ;
  assign n10790 = n10789 ^ n609 ;
  assign n10791 = n10790 ^ n835 ;
  assign n10792 = ~n10787 & ~n10791 ;
  assign n10793 = n10792 ^ n10790 ;
  assign n10794 = n10492 & n10793 ;
  assign n10795 = n10794 ^ n834 ;
  assign n10796 = n10398 & n10468 ;
  assign n10797 = n10796 ^ n10128 ;
  assign n10798 = n10797 ^ n534 ;
  assign n10799 = ~n10795 & ~n10798 ;
  assign n10800 = n10799 ^ n750 ;
  assign n10801 = n10489 & n10800 ;
  assign n10802 = n10801 ^ n10488 ;
  assign n10805 = n10804 ^ n10802 ;
  assign n10806 = n10804 ^ n401 ;
  assign n10807 = n10805 & n10806 ;
  assign n10808 = n10807 ^ n462 ;
  assign n10809 = n10486 & n10808 ;
  assign n10810 = n10809 ^ n349 ;
  assign n10811 = n10410 ^ n341 ;
  assign n10812 = n10468 & n10811 ;
  assign n10813 = n10812 ^ n10118 ;
  assign n10814 = n10813 ^ n291 ;
  assign n10815 = ~n10810 & ~n10814 ;
  assign n10816 = n10815 ^ n307 ;
  assign n10817 = n10482 & n10816 ;
  assign n10818 = n10817 ^ n10481 ;
  assign n10472 = ~n10418 & n10468 ;
  assign n10473 = n10472 ^ n10110 ;
  assign n10819 = n10818 ^ n10473 ;
  assign n10820 = n10818 ^ n188 ;
  assign n10821 = ~n10819 & n10820 ;
  assign n10822 = n10821 ^ n203 ;
  assign n10823 = n10471 & ~n10822 ;
  assign n10824 = n10823 ^ n10470 ;
  assign n10825 = n10824 ^ n138 ;
  assign n10868 = n10457 & n10468 ;
  assign n10869 = n10868 ^ n10451 ;
  assign n10870 = n10869 ^ n10824 ;
  assign n10871 = n10825 & ~n10870 ;
  assign n10872 = n10871 ^ n138 ;
  assign n10873 = n10867 & n10872 ;
  assign n10874 = ~n10828 & n10873 ;
  assign n10875 = n10874 ^ n10867 ;
  assign n10914 = ~n10734 & ~n10875 ;
  assign n10915 = n10914 ^ n10514 ;
  assign n10916 = n10915 ^ n2511 ;
  assign n10917 = n10732 & ~n10875 ;
  assign n10918 = n10917 ^ n10517 ;
  assign n10919 = n10918 ^ n2707 ;
  assign n11111 = n10723 ^ n3320 ;
  assign n11112 = ~n10875 & n11111 ;
  assign n11113 = n11112 ^ n10526 ;
  assign n11116 = n11113 ^ n2894 ;
  assign n10920 = ~n10719 & ~n10875 ;
  assign n10921 = n10920 ^ n10539 ;
  assign n10922 = n10921 ^ n3538 ;
  assign n11097 = n10712 ^ n3908 ;
  assign n11098 = ~n10875 & n11097 ;
  assign n11099 = n11098 ^ n10715 ;
  assign n10923 = n10710 & ~n10875 ;
  assign n10924 = n10923 ^ n10559 ;
  assign n10925 = n10924 ^ n3908 ;
  assign n10926 = n10706 ^ n4356 ;
  assign n10927 = ~n10875 & n10926 ;
  assign n10928 = n10927 ^ n10568 ;
  assign n10929 = n10928 ^ n4153 ;
  assign n11086 = n10704 & ~n10875 ;
  assign n11087 = n11086 ^ n10576 ;
  assign n11090 = n11087 ^ n4153 ;
  assign n10930 = ~n10695 & ~n10875 ;
  assign n10931 = n10930 ^ n10579 ;
  assign n10932 = n10931 ^ n4812 ;
  assign n10933 = n10693 & ~n10875 ;
  assign n10934 = n10933 ^ n10582 ;
  assign n10935 = n10934 ^ n5073 ;
  assign n10936 = n10691 & ~n10875 ;
  assign n10937 = n10936 ^ n10586 ;
  assign n11075 = n10937 ^ n5073 ;
  assign n10938 = n10937 ^ n5317 ;
  assign n11068 = n10687 & ~n10875 ;
  assign n11069 = n11068 ^ n10588 ;
  assign n10939 = ~n10682 & ~n10875 ;
  assign n10940 = n10939 ^ n10684 ;
  assign n10941 = n10940 ^ n5830 ;
  assign n10942 = ~n10680 & ~n10875 ;
  assign n10943 = n10942 ^ n10592 ;
  assign n10944 = n10943 ^ n6115 ;
  assign n11057 = n10673 ^ n6673 ;
  assign n11058 = ~n10875 & n11057 ;
  assign n11059 = n11058 ^ n10676 ;
  assign n10945 = n10671 & ~n10875 ;
  assign n10946 = n10945 ^ n10595 ;
  assign n10947 = n10946 ^ n6673 ;
  assign n10948 = n10665 ^ n7277 ;
  assign n10949 = ~n10875 & n10948 ;
  assign n10950 = n10949 ^ n10667 ;
  assign n10951 = n10950 ^ n6959 ;
  assign n10952 = ~n10663 & ~n10875 ;
  assign n10953 = n10952 ^ n10598 ;
  assign n10954 = n10953 ^ n7277 ;
  assign n11044 = ~n10661 & ~n10875 ;
  assign n11045 = n11044 ^ n10601 ;
  assign n11048 = n11045 ^ n7277 ;
  assign n10955 = n10649 ^ n8910 ;
  assign n10956 = ~n10875 & ~n10955 ;
  assign n10957 = n10956 ^ n10609 ;
  assign n10958 = n10957 ^ n8586 ;
  assign n10959 = n10647 & ~n10875 ;
  assign n10960 = n10959 ^ n10619 ;
  assign n10961 = n10960 ^ n8910 ;
  assign n10962 = ~x22 & ~n10629 ;
  assign n10963 = n10962 ^ n10108 ;
  assign n10971 = n10963 ^ n10626 ;
  assign n10964 = n10963 ^ n10468 ;
  assign n10965 = n10964 ^ n10963 ;
  assign n10968 = x22 & n10965 ;
  assign n10969 = n10968 ^ n10963 ;
  assign n10970 = n10875 & ~n10969 ;
  assign n10972 = n10971 ^ n10970 ;
  assign n10973 = n10972 ^ n9542 ;
  assign n10986 = n10468 ^ x22 ;
  assign n10987 = n10875 ^ x21 ;
  assign n10988 = n10987 ^ n10468 ;
  assign n10979 = ~x18 & ~x19 ;
  assign n10980 = ~x20 & n10979 ;
  assign n10989 = n10468 ^ x21 ;
  assign n10990 = ~n10980 & n10989 ;
  assign n10991 = n10990 ^ n10468 ;
  assign n10992 = ~n10988 & ~n10991 ;
  assign n10993 = n10992 ^ n10468 ;
  assign n10994 = n10986 & ~n10993 ;
  assign n10974 = n10629 ^ n10468 ;
  assign n10975 = ~n10875 & ~n10974 ;
  assign n10976 = n10975 ^ n10468 ;
  assign n10977 = n10976 ^ x22 ;
  assign n10983 = ~n10975 & ~n10980 ;
  assign n10984 = n10983 ^ n10468 ;
  assign n10985 = n10977 & ~n10984 ;
  assign n10995 = n10994 ^ n10985 ;
  assign n10996 = ~n10108 & ~n10995 ;
  assign n10981 = n10980 ^ n10468 ;
  assign n11011 = n10981 ^ x21 ;
  assign n11012 = n11011 ^ x21 ;
  assign n11013 = ~n10989 & ~n11012 ;
  assign n11014 = n11013 ^ x21 ;
  assign n11015 = ~n10986 & ~n11014 ;
  assign n10997 = x21 ^ x20 ;
  assign n10998 = n10997 ^ x20 ;
  assign n10999 = n10998 ^ x22 ;
  assign n11000 = n10986 ^ x20 ;
  assign n11001 = n10999 & n11000 ;
  assign n11002 = n11001 ^ x20 ;
  assign n11003 = n10979 ^ x22 ;
  assign n11004 = n11003 ^ x22 ;
  assign n11005 = n11001 ^ n10999 ;
  assign n11006 = n11004 & n11005 ;
  assign n11007 = n11006 ^ x22 ;
  assign n11008 = ~n11002 & ~n11007 ;
  assign n11009 = n11008 ^ x22 ;
  assign n11016 = n11015 ^ n11009 ;
  assign n11017 = n10875 & ~n11016 ;
  assign n11010 = n11009 ^ n9542 ;
  assign n11018 = n11017 ^ n11010 ;
  assign n11019 = n11018 ^ n9542 ;
  assign n11020 = n10996 & n11019 ;
  assign n11021 = n11020 ^ n11018 ;
  assign n11022 = n10973 & ~n11021 ;
  assign n11023 = n11022 ^ n9628 ;
  assign n11024 = ~n10645 & ~n10875 ;
  assign n11025 = n11024 ^ n10624 ;
  assign n11026 = n11025 ^ n9217 ;
  assign n11027 = n11023 & ~n11026 ;
  assign n11028 = n11027 ^ n9285 ;
  assign n11029 = ~n10961 & ~n11028 ;
  assign n11030 = n11029 ^ n9005 ;
  assign n11031 = n10958 & n11030 ;
  assign n11032 = n11031 ^ n8688 ;
  assign n11033 = n10653 & ~n10875 ;
  assign n11034 = n11033 ^ n10605 ;
  assign n11035 = n11034 ^ n8253 ;
  assign n11036 = n11032 & n11035 ;
  assign n11037 = n11036 ^ n8356 ;
  assign n11038 = n10655 ^ n8253 ;
  assign n11039 = ~n10875 & n11038 ;
  assign n11040 = n11039 ^ n10657 ;
  assign n11041 = n11040 ^ n7891 ;
  assign n11042 = ~n11037 & ~n11041 ;
  assign n11043 = n11042 ^ n7971 ;
  assign n11046 = n11045 ^ n7584 ;
  assign n11047 = n11043 & n11046 ;
  assign n11049 = n11048 ^ n11047 ;
  assign n11050 = n10954 & n11049 ;
  assign n11051 = n11050 ^ n7277 ;
  assign n11052 = n11051 ^ n10950 ;
  assign n11053 = ~n10951 & n11052 ;
  assign n11054 = n11053 ^ n7011 ;
  assign n11055 = ~n10947 & n11054 ;
  assign n11056 = n11055 ^ n6673 ;
  assign n11060 = n11059 ^ n11056 ;
  assign n11061 = n11059 ^ n6389 ;
  assign n11062 = n11060 & n11061 ;
  assign n11063 = n11062 ^ n6423 ;
  assign n11064 = ~n10944 & ~n11063 ;
  assign n11065 = n11064 ^ n6429 ;
  assign n11066 = n10941 & ~n11065 ;
  assign n11067 = n11066 ^ n10940 ;
  assign n11070 = n11069 ^ n11067 ;
  assign n11071 = n11069 ^ n5562 ;
  assign n11072 = ~n11070 & n11071 ;
  assign n11073 = n11072 ^ n5885 ;
  assign n11074 = ~n10938 & ~n11073 ;
  assign n11076 = n11075 ^ n11074 ;
  assign n11077 = ~n10935 & ~n11076 ;
  assign n11078 = n11077 ^ n5115 ;
  assign n11079 = n10932 & n11078 ;
  assign n11080 = n11079 ^ n4854 ;
  assign n11081 = n10698 & ~n10875 ;
  assign n11082 = n11081 ^ n10701 ;
  assign n11083 = n11082 ^ n4583 ;
  assign n11084 = n11080 & ~n11083 ;
  assign n11085 = n11084 ^ n4645 ;
  assign n11088 = n11087 ^ n4356 ;
  assign n11089 = ~n11085 & n11088 ;
  assign n11091 = n11090 ^ n11089 ;
  assign n11092 = ~n10929 & n11091 ;
  assign n11093 = n11092 ^ n4153 ;
  assign n11094 = n11093 ^ n10924 ;
  assign n11095 = ~n10925 & n11094 ;
  assign n11096 = n11095 ^ n3908 ;
  assign n11100 = n11099 ^ n11096 ;
  assign n11101 = n11099 ^ n3722 ;
  assign n11102 = n11100 & n11101 ;
  assign n11103 = n11102 ^ n3795 ;
  assign n11104 = ~n10922 & n11103 ;
  assign n11105 = n11104 ^ n3596 ;
  assign n11106 = n10721 & ~n10875 ;
  assign n11107 = n11106 ^ n10530 ;
  assign n11108 = n11107 ^ n3320 ;
  assign n11109 = n11105 & ~n11108 ;
  assign n11110 = n11109 ^ n3387 ;
  assign n11114 = n11113 ^ n3093 ;
  assign n11115 = n11110 & n11114 ;
  assign n11117 = n11116 ^ n11115 ;
  assign n11118 = ~n10726 & ~n10875 ;
  assign n11119 = n11118 ^ n10729 ;
  assign n11120 = n11119 ^ n2894 ;
  assign n11121 = n11117 & ~n11120 ;
  assign n11122 = n11121 ^ n3396 ;
  assign n11123 = ~n10919 & ~n11122 ;
  assign n11124 = n11123 ^ n2707 ;
  assign n11125 = n11124 ^ n10915 ;
  assign n11126 = ~n10916 & ~n11125 ;
  assign n11127 = n11126 ^ n2530 ;
  assign n10876 = n10825 & ~n10875 ;
  assign n10877 = n10876 ^ n10869 ;
  assign n10878 = n10877 ^ n183 ;
  assign n10879 = n10820 & ~n10875 ;
  assign n10880 = n10879 ^ n10473 ;
  assign n10882 = n10880 ^ n157 ;
  assign n10881 = n157 & n10880 ;
  assign n10883 = n10882 ^ n10881 ;
  assign n11205 = ~n10816 & ~n10875 ;
  assign n11206 = n11205 ^ n10481 ;
  assign n10884 = ~n10810 & ~n10875 ;
  assign n10885 = n10884 ^ n10813 ;
  assign n10886 = n10885 ^ n245 ;
  assign n10887 = n10808 & ~n10875 ;
  assign n10888 = n10887 ^ n10485 ;
  assign n10889 = n10888 ^ n291 ;
  assign n10890 = n10802 ^ n401 ;
  assign n10891 = ~n10875 & ~n10890 ;
  assign n10892 = n10891 ^ n10804 ;
  assign n10893 = n10892 ^ n341 ;
  assign n11193 = ~n10800 & ~n10875 ;
  assign n11194 = n11193 ^ n10488 ;
  assign n10894 = n10793 & ~n10875 ;
  assign n10895 = n10894 ^ n10491 ;
  assign n10896 = n10895 ^ n534 ;
  assign n10897 = n10787 & ~n10875 ;
  assign n10898 = n10897 ^ n10789 ;
  assign n10899 = n10898 ^ n609 ;
  assign n10900 = ~n10759 & ~n10875 ;
  assign n10901 = n10900 ^ n10761 ;
  assign n10902 = n10901 ^ n1136 ;
  assign n11151 = n10757 & ~n10875 ;
  assign n11152 = n11151 ^ n10497 ;
  assign n11155 = n11152 ^ n1136 ;
  assign n10903 = ~n10750 & ~n10875 ;
  assign n10904 = n10903 ^ n10502 ;
  assign n11143 = n10904 ^ n1427 ;
  assign n10905 = n10904 ^ n1572 ;
  assign n10908 = n10744 & ~n10875 ;
  assign n10909 = n10908 ^ n10507 ;
  assign n10910 = n10909 ^ n2008 ;
  assign n10911 = n10742 & ~n10875 ;
  assign n10912 = n10911 ^ n10511 ;
  assign n10913 = n10912 ^ n2175 ;
  assign n11128 = n10736 ^ n2511 ;
  assign n11129 = ~n10875 & ~n11128 ;
  assign n11130 = n11129 ^ n10738 ;
  assign n11131 = n11130 ^ n2366 ;
  assign n11132 = n11127 & n11131 ;
  assign n11133 = n11132 ^ n2399 ;
  assign n11134 = ~n10913 & n11133 ;
  assign n11135 = n11134 ^ n2204 ;
  assign n11136 = n10910 & n11135 ;
  assign n11137 = n11136 ^ n2008 ;
  assign n10906 = n10748 & ~n10875 ;
  assign n10907 = n10906 ^ n10505 ;
  assign n11138 = n11137 ^ n10907 ;
  assign n11139 = n11137 ^ n1739 ;
  assign n11140 = ~n11138 & ~n11139 ;
  assign n11141 = n11140 ^ n1763 ;
  assign n11142 = n10905 & n11141 ;
  assign n11144 = n11143 ^ n11142 ;
  assign n11145 = n10752 ^ n1572 ;
  assign n11146 = ~n10875 & ~n11145 ;
  assign n11147 = n11146 ^ n10500 ;
  assign n11148 = n11147 ^ n1427 ;
  assign n11149 = ~n11144 & n11148 ;
  assign n11150 = n11149 ^ n1450 ;
  assign n11153 = n11152 ^ n1290 ;
  assign n11154 = n11150 & n11153 ;
  assign n11156 = n11155 ^ n11154 ;
  assign n11157 = ~n10902 & n11156 ;
  assign n11158 = n11157 ^ n1143 ;
  assign n11159 = ~n10765 & ~n10875 ;
  assign n11160 = n11159 ^ n10494 ;
  assign n11163 = n11160 ^ n1034 ;
  assign n11164 = ~n11158 & ~n11163 ;
  assign n11161 = n11160 ^ n892 ;
  assign n11165 = n11164 ^ n11161 ;
  assign n11166 = n10767 & ~n10875 ;
  assign n11167 = n11166 ^ n10770 ;
  assign n11168 = n11167 ^ n786 ;
  assign n11169 = n11168 ^ n927 ;
  assign n11170 = n11165 & n11169 ;
  assign n11171 = n11170 ^ n11168 ;
  assign n11172 = n10775 & ~n10875 ;
  assign n11173 = n11172 ^ n10777 ;
  assign n11174 = n11173 ^ n696 ;
  assign n11175 = n11174 ^ n842 ;
  assign n11176 = ~n11171 & n11175 ;
  assign n11177 = n11176 ^ n11174 ;
  assign n11178 = n10781 & ~n10875 ;
  assign n11179 = n11178 ^ n10783 ;
  assign n11180 = n11179 ^ n609 ;
  assign n11181 = n11180 ^ n835 ;
  assign n11182 = ~n11177 & n11181 ;
  assign n11183 = n11182 ^ n11180 ;
  assign n11184 = n10899 & ~n11183 ;
  assign n11185 = n11184 ^ n834 ;
  assign n11186 = ~n10896 & ~n11185 ;
  assign n11187 = n11186 ^ n750 ;
  assign n11188 = ~n10795 & ~n10875 ;
  assign n11189 = n11188 ^ n10797 ;
  assign n11190 = n11189 ^ n457 ;
  assign n11191 = n11187 & n11190 ;
  assign n11192 = n11191 ^ n11189 ;
  assign n11195 = n11194 ^ n11192 ;
  assign n11196 = n11194 ^ n401 ;
  assign n11197 = ~n11195 & ~n11196 ;
  assign n11198 = n11197 ^ n462 ;
  assign n11199 = n10893 & n11198 ;
  assign n11200 = n11199 ^ n349 ;
  assign n11201 = ~n10889 & ~n11200 ;
  assign n11202 = n11201 ^ n307 ;
  assign n11203 = n10886 & n11202 ;
  assign n11204 = n11203 ^ n10885 ;
  assign n11207 = n11206 ^ n11204 ;
  assign n11208 = n11206 ^ n188 ;
  assign n11209 = ~n11207 & n11208 ;
  assign n11210 = n11209 ^ n188 ;
  assign n11211 = n10883 & n11210 ;
  assign n11212 = n10822 & ~n10875 ;
  assign n11213 = n11212 ^ n10470 ;
  assign n11214 = ~n10881 & ~n11213 ;
  assign n11215 = ~n11211 & n11214 ;
  assign n11216 = n138 & ~n11215 ;
  assign n11218 = n11215 ^ n11213 ;
  assign n11217 = ~n10881 & ~n11211 ;
  assign n11219 = n11218 ^ n11217 ;
  assign n11220 = ~n11216 & ~n11219 ;
  assign n11221 = ~n10827 & n10867 ;
  assign n11222 = n10872 ^ n10827 ;
  assign n11223 = ~n11221 & n11222 ;
  assign n11224 = n11223 ^ n11221 ;
  assign n11225 = n11221 ^ n10877 ;
  assign n11226 = n11225 ^ n11221 ;
  assign n11227 = n11224 & n11226 ;
  assign n11228 = n11227 ^ n11221 ;
  assign n11229 = ~n183 & ~n11228 ;
  assign n11230 = n11229 ^ n11223 ;
  assign n11231 = ~n11220 & ~n11230 ;
  assign n11232 = ~n10878 & n11231 ;
  assign n11233 = n11232 ^ n11230 ;
  assign n11259 = n11127 & n11233 ;
  assign n11260 = n11259 ^ n11130 ;
  assign n11261 = n11260 ^ n2175 ;
  assign n11262 = ~n11122 & n11233 ;
  assign n11263 = n11262 ^ n10918 ;
  assign n11264 = n11263 ^ n2511 ;
  assign n11265 = n11117 & n11233 ;
  assign n11266 = n11265 ^ n11119 ;
  assign n11267 = n11266 ^ n2707 ;
  assign n11447 = ~n11110 & n11233 ;
  assign n11448 = n11447 ^ n11113 ;
  assign n11268 = n11105 & n11233 ;
  assign n11269 = n11268 ^ n11107 ;
  assign n11270 = n11269 ^ n3093 ;
  assign n11271 = n11096 ^ n3722 ;
  assign n11272 = n11233 & ~n11271 ;
  assign n11273 = n11272 ^ n11099 ;
  assign n11274 = n11273 ^ n3538 ;
  assign n11275 = n11093 ^ n3908 ;
  assign n11276 = n11233 & n11275 ;
  assign n11277 = n11276 ^ n10924 ;
  assign n11278 = n11277 ^ n3722 ;
  assign n11429 = n11091 & n11233 ;
  assign n11430 = n11429 ^ n10928 ;
  assign n11279 = ~n11076 & n11233 ;
  assign n11280 = n11279 ^ n10934 ;
  assign n11281 = n11280 ^ n4812 ;
  assign n11282 = n11073 & n11233 ;
  assign n11283 = n11282 ^ n10937 ;
  assign n11284 = n11283 ^ n5073 ;
  assign n11289 = ~n11063 & n11233 ;
  assign n11290 = n11289 ^ n10943 ;
  assign n11291 = n11290 ^ n5830 ;
  assign n11292 = n11056 ^ n6389 ;
  assign n11293 = n11233 & ~n11292 ;
  assign n11294 = n11293 ^ n11059 ;
  assign n11295 = n11294 ^ n6115 ;
  assign n11296 = n11054 & n11233 ;
  assign n11297 = n11296 ^ n10946 ;
  assign n11298 = n11297 ^ n6389 ;
  assign n11388 = n11051 ^ n6959 ;
  assign n11389 = n11233 & n11388 ;
  assign n11390 = n11389 ^ n10950 ;
  assign n11299 = ~n11043 & n11233 ;
  assign n11300 = n11299 ^ n11045 ;
  assign n11301 = n11300 ^ n7277 ;
  assign n11375 = ~n11037 & n11233 ;
  assign n11376 = n11375 ^ n11040 ;
  assign n11379 = n11376 ^ n7277 ;
  assign n11302 = ~n11028 & n11233 ;
  assign n11303 = n11302 ^ n10960 ;
  assign n11304 = n11303 ^ n8586 ;
  assign n11305 = n11023 & n11233 ;
  assign n11306 = n11305 ^ n11025 ;
  assign n11307 = n11306 ^ n8910 ;
  assign n11308 = ~n11021 & n11233 ;
  assign n11309 = n11308 ^ n10972 ;
  assign n11310 = n11309 ^ n9217 ;
  assign n11318 = n10987 ^ n10981 ;
  assign n11313 = n10981 ^ n10875 ;
  assign n11314 = n11313 ^ n10981 ;
  assign n11315 = x20 & ~n11314 ;
  assign n11316 = n11315 ^ n10981 ;
  assign n11317 = ~n11233 & n11316 ;
  assign n11319 = n11318 ^ n11317 ;
  assign n11320 = n11319 ^ n10108 ;
  assign n11322 = n10979 ^ n10875 ;
  assign n11323 = n11233 & ~n11322 ;
  assign n11321 = n10875 ^ x20 ;
  assign n11324 = n11323 ^ n11321 ;
  assign n11325 = n11324 ^ n10468 ;
  assign n11328 = n10875 ^ x19 ;
  assign n11329 = n11328 ^ n11233 ;
  assign n11331 = n10875 ^ x18 ;
  assign n11330 = ~x16 & ~x17 ;
  assign n11332 = n11331 ^ n11330 ;
  assign n11333 = n11329 & ~n11332 ;
  assign n11326 = n11233 ^ n10875 ;
  assign n11336 = n11333 ^ n11326 ;
  assign n11337 = n11336 ^ n11333 ;
  assign n11340 = n11328 & ~n11337 ;
  assign n11341 = n11340 ^ n11333 ;
  assign n11342 = x18 & n11341 ;
  assign n11327 = n10875 ^ n10468 ;
  assign n11334 = n11333 ^ n11327 ;
  assign n11343 = n11342 ^ n11334 ;
  assign n11344 = n11325 & ~n11343 ;
  assign n11345 = n11344 ^ n10639 ;
  assign n11346 = ~n11320 & ~n11345 ;
  assign n11347 = n11346 ^ n10203 ;
  assign n11350 = n10108 ^ x21 ;
  assign n11349 = ~n10981 & n10988 ;
  assign n11351 = n11350 ^ n11349 ;
  assign n11348 = ~n10628 & ~n10875 ;
  assign n11352 = n11351 ^ n11348 ;
  assign n11353 = n11233 & n11352 ;
  assign n11354 = n11353 ^ n10977 ;
  assign n11355 = n11354 ^ n9542 ;
  assign n11356 = ~n11347 & ~n11355 ;
  assign n11357 = n11356 ^ n9628 ;
  assign n11358 = n11310 & n11357 ;
  assign n11359 = n11358 ^ n9285 ;
  assign n11360 = n11307 & ~n11359 ;
  assign n11361 = n11360 ^ n9005 ;
  assign n11362 = ~n11304 & n11361 ;
  assign n11363 = n11362 ^ n8586 ;
  assign n11364 = n11363 ^ n8253 ;
  assign n11365 = n11030 & n11233 ;
  assign n11366 = n11365 ^ n10957 ;
  assign n11367 = n11366 ^ n11363 ;
  assign n11368 = n11364 & ~n11367 ;
  assign n11369 = n11368 ^ n8356 ;
  assign n11370 = n11032 & n11233 ;
  assign n11371 = n11370 ^ n11034 ;
  assign n11372 = n11371 ^ n7891 ;
  assign n11373 = ~n11369 & ~n11372 ;
  assign n11374 = n11373 ^ n7971 ;
  assign n11377 = n11376 ^ n7584 ;
  assign n11378 = n11374 & n11377 ;
  assign n11380 = n11379 ^ n11378 ;
  assign n11381 = n11301 & n11380 ;
  assign n11382 = n11381 ^ n7339 ;
  assign n11383 = n11049 & n11233 ;
  assign n11384 = n11383 ^ n10953 ;
  assign n11385 = n11384 ^ n6959 ;
  assign n11386 = n11382 & n11385 ;
  assign n11387 = n11386 ^ n6959 ;
  assign n11391 = n11390 ^ n11387 ;
  assign n11392 = n11390 ^ n6673 ;
  assign n11393 = n11391 & ~n11392 ;
  assign n11394 = n11393 ^ n6713 ;
  assign n11395 = n11298 & ~n11394 ;
  assign n11396 = n11395 ^ n6423 ;
  assign n11397 = ~n11295 & ~n11396 ;
  assign n11398 = n11397 ^ n6429 ;
  assign n11399 = ~n11291 & n11398 ;
  assign n11400 = n11399 ^ n5900 ;
  assign n11401 = n11065 & n11233 ;
  assign n11402 = n11401 ^ n10940 ;
  assign n11403 = n11402 ^ n5562 ;
  assign n11404 = n11400 & n11403 ;
  assign n11405 = n11404 ^ n5885 ;
  assign n11285 = n11067 ^ n5562 ;
  assign n11286 = n11233 & n11285 ;
  assign n11287 = n11286 ^ n11069 ;
  assign n11406 = n11287 ^ n5317 ;
  assign n11407 = ~n11405 & n11406 ;
  assign n11288 = n11287 ^ n5073 ;
  assign n11408 = n11407 ^ n11288 ;
  assign n11409 = ~n11284 & n11408 ;
  assign n11410 = n11409 ^ n5073 ;
  assign n11411 = n11410 ^ n11280 ;
  assign n11412 = ~n11281 & n11411 ;
  assign n11413 = n11412 ^ n4854 ;
  assign n11414 = n11078 & n11233 ;
  assign n11415 = n11414 ^ n10931 ;
  assign n11416 = n11415 ^ n4583 ;
  assign n11417 = n11413 & n11416 ;
  assign n11418 = n11417 ^ n4645 ;
  assign n11419 = n11080 & n11233 ;
  assign n11420 = n11419 ^ n11082 ;
  assign n11421 = n11420 ^ n4356 ;
  assign n11422 = n11418 & ~n11421 ;
  assign n11423 = n11422 ^ n4414 ;
  assign n11424 = n11085 & n11233 ;
  assign n11425 = n11424 ^ n11087 ;
  assign n11426 = n11425 ^ n4153 ;
  assign n11427 = n11423 & n11426 ;
  assign n11428 = n11427 ^ n4153 ;
  assign n11431 = n11430 ^ n11428 ;
  assign n11432 = n11430 ^ n3908 ;
  assign n11433 = n11431 & ~n11432 ;
  assign n11434 = n11433 ^ n3961 ;
  assign n11435 = n11278 & ~n11434 ;
  assign n11436 = n11435 ^ n3722 ;
  assign n11437 = n11436 ^ n11273 ;
  assign n11438 = n11274 & ~n11437 ;
  assign n11439 = n11438 ^ n3596 ;
  assign n11440 = n11103 & n11233 ;
  assign n11441 = n11440 ^ n10921 ;
  assign n11442 = n11441 ^ n3320 ;
  assign n11443 = n11439 & ~n11442 ;
  assign n11444 = n11443 ^ n3387 ;
  assign n11445 = n11270 & n11444 ;
  assign n11446 = n11445 ^ n11269 ;
  assign n11449 = n11448 ^ n11446 ;
  assign n11450 = n11448 ^ n2894 ;
  assign n11451 = ~n11449 & n11450 ;
  assign n11452 = n11451 ^ n3396 ;
  assign n11453 = n11267 & ~n11452 ;
  assign n11454 = n11453 ^ n2707 ;
  assign n11455 = n11454 ^ n11263 ;
  assign n11456 = n11264 & n11455 ;
  assign n11457 = n11456 ^ n2530 ;
  assign n11458 = n11124 ^ n2511 ;
  assign n11459 = n11233 & ~n11458 ;
  assign n11460 = n11459 ^ n10915 ;
  assign n11461 = n11460 ^ n2366 ;
  assign n11462 = n11457 & ~n11461 ;
  assign n11463 = n11462 ^ n2399 ;
  assign n11464 = n11261 & n11463 ;
  assign n11465 = n11464 ^ n2175 ;
  assign n11257 = n11133 & n11233 ;
  assign n11258 = n11257 ^ n10912 ;
  assign n11466 = n11465 ^ n11258 ;
  assign n11467 = n11465 ^ n2008 ;
  assign n11468 = n11466 & n11467 ;
  assign n11469 = n11468 ^ n2064 ;
  assign n11543 = n11219 ^ n11216 ;
  assign n11544 = n11543 ^ n11220 ;
  assign n11545 = n11544 ^ n11223 ;
  assign n11548 = n183 & n11545 ;
  assign n11549 = n11548 ^ n11544 ;
  assign n11550 = ~n11220 & n11549 ;
  assign n11551 = n11550 ^ n183 ;
  assign n11556 = ~n11213 & ~n11230 ;
  assign n11557 = n11556 ^ n10877 ;
  assign n11558 = ~n11551 & ~n11557 ;
  assign n11538 = n130 & n11215 ;
  assign n11539 = n11538 ^ n11220 ;
  assign n11540 = ~n183 & ~n11539 ;
  assign n11541 = n11540 ^ n11220 ;
  assign n11542 = n10877 & n11541 ;
  assign n11559 = n11558 ^ n11542 ;
  assign n11560 = n11217 ^ n138 ;
  assign n11561 = n11233 & ~n11560 ;
  assign n11562 = n11561 ^ n11213 ;
  assign n11563 = n183 & ~n11562 ;
  assign n11584 = n11210 ^ n157 ;
  assign n11585 = n11233 & n11584 ;
  assign n11586 = n11585 ^ n10880 ;
  assign n11564 = n11204 ^ n188 ;
  assign n11565 = n11233 & n11564 ;
  assign n11566 = n11565 ^ n11206 ;
  assign n11567 = n11566 ^ n157 ;
  assign n11568 = ~n11202 & n11233 ;
  assign n11569 = n11568 ^ n10885 ;
  assign n11570 = n11569 ^ n157 ;
  assign n11571 = n11570 ^ n203 ;
  assign n11234 = n11198 & n11233 ;
  assign n11235 = n11234 ^ n10892 ;
  assign n11236 = n11235 ^ n291 ;
  assign n11522 = ~n11187 & n11233 ;
  assign n11523 = n11522 ^ n11189 ;
  assign n11242 = ~n11183 & n11233 ;
  assign n11243 = n11242 ^ n10898 ;
  assign n11244 = n11243 ^ n534 ;
  assign n11245 = n11177 & n11233 ;
  assign n11246 = n11245 ^ n11179 ;
  assign n11247 = n11246 ^ n609 ;
  assign n11248 = ~n11150 & n11233 ;
  assign n11249 = n11248 ^ n11152 ;
  assign n11250 = n11249 ^ n1136 ;
  assign n11251 = ~n11141 & n11233 ;
  assign n11252 = n11251 ^ n10904 ;
  assign n11253 = n11252 ^ n1427 ;
  assign n11472 = ~n11139 & n11233 ;
  assign n11473 = n11472 ^ n10907 ;
  assign n11477 = n11473 ^ n1427 ;
  assign n11254 = n11135 & n11233 ;
  assign n11255 = n11254 ^ n10909 ;
  assign n11256 = n11255 ^ n1739 ;
  assign n11470 = ~n11256 & ~n11469 ;
  assign n11471 = n11470 ^ n1739 ;
  assign n11474 = n11473 ^ n11471 ;
  assign n11475 = n11471 ^ n1572 ;
  assign n11476 = ~n11474 & n11475 ;
  assign n11478 = n11477 ^ n11476 ;
  assign n11479 = ~n11253 & ~n11478 ;
  assign n11480 = n11479 ^ n1450 ;
  assign n11481 = ~n11144 & n11233 ;
  assign n11482 = n11481 ^ n11147 ;
  assign n11483 = n11482 ^ n1290 ;
  assign n11484 = ~n11480 & ~n11483 ;
  assign n11485 = n11484 ^ n1461 ;
  assign n11486 = n11250 & n11485 ;
  assign n11487 = n11486 ^ n1143 ;
  assign n11488 = n11156 & n11233 ;
  assign n11489 = n11488 ^ n10901 ;
  assign n11492 = n11489 ^ n1034 ;
  assign n11493 = ~n11487 & ~n11492 ;
  assign n11490 = n11489 ^ n892 ;
  assign n11494 = n11493 ^ n11490 ;
  assign n11495 = n11158 & n11233 ;
  assign n11496 = n11495 ^ n11160 ;
  assign n11497 = n11496 ^ n786 ;
  assign n11498 = n11497 ^ n927 ;
  assign n11499 = n11494 & ~n11498 ;
  assign n11500 = n11499 ^ n11497 ;
  assign n11501 = ~n11165 & n11233 ;
  assign n11502 = n11501 ^ n11167 ;
  assign n11503 = n11502 ^ n696 ;
  assign n11504 = n11503 ^ n842 ;
  assign n11505 = n11500 & n11504 ;
  assign n11506 = n11505 ^ n11503 ;
  assign n11507 = n11171 & n11233 ;
  assign n11508 = n11507 ^ n11173 ;
  assign n11509 = n11508 ^ n609 ;
  assign n11510 = n11509 ^ n835 ;
  assign n11511 = ~n11506 & n11510 ;
  assign n11512 = n11511 ^ n11509 ;
  assign n11513 = ~n11247 & ~n11512 ;
  assign n11514 = n11513 ^ n834 ;
  assign n11515 = ~n11244 & ~n11514 ;
  assign n11516 = n11515 ^ n750 ;
  assign n11517 = ~n11185 & n11233 ;
  assign n11518 = n11517 ^ n10895 ;
  assign n11519 = n11518 ^ n457 ;
  assign n11520 = n11516 & n11519 ;
  assign n11521 = n11520 ^ n11518 ;
  assign n11524 = n11523 ^ n11521 ;
  assign n11525 = n11523 ^ n401 ;
  assign n11526 = ~n11524 & ~n11525 ;
  assign n11527 = n11526 ^ n401 ;
  assign n11240 = n11235 ^ n341 ;
  assign n11237 = n11192 ^ n401 ;
  assign n11238 = n11233 & ~n11237 ;
  assign n11239 = n11238 ^ n11194 ;
  assign n11241 = n11240 ^ n11239 ;
  assign n11528 = n11527 ^ n11241 ;
  assign n11529 = n11528 ^ n11240 ;
  assign n11530 = n11239 ^ n11235 ;
  assign n11531 = n11530 ^ n11240 ;
  assign n11532 = n11529 & ~n11531 ;
  assign n11533 = n11532 ^ n11240 ;
  assign n11534 = ~n11236 & ~n11533 ;
  assign n11535 = n11534 ^ n307 ;
  assign n11572 = ~n11200 & n11233 ;
  assign n11573 = n11572 ^ n10888 ;
  assign n11574 = n11573 ^ n245 ;
  assign n11575 = n11535 & n11574 ;
  assign n11576 = n11575 ^ n11573 ;
  assign n11577 = n11576 ^ n188 ;
  assign n11580 = n11571 & n11577 ;
  assign n11581 = n11580 ^ n203 ;
  assign n11582 = n11567 & ~n11581 ;
  assign n11583 = n11582 ^ n11566 ;
  assign n11589 = n11586 ^ n11583 ;
  assign n11590 = n138 & ~n11589 ;
  assign n11587 = n11583 & n11586 ;
  assign n11588 = n11587 ^ n138 ;
  assign n11591 = n11590 ^ n11588 ;
  assign n11592 = ~n11563 & n11591 ;
  assign n11593 = ~n11559 & n11592 ;
  assign n11594 = n11593 ^ n11559 ;
  assign n11614 = ~n11469 & n11594 ;
  assign n11615 = n11614 ^ n11255 ;
  assign n11843 = n11615 ^ n1427 ;
  assign n11616 = n11615 ^ n1572 ;
  assign n11619 = n11463 & n11594 ;
  assign n11620 = n11619 ^ n11260 ;
  assign n11621 = n11620 ^ n2008 ;
  assign n11622 = n11457 & n11594 ;
  assign n11623 = n11622 ^ n11460 ;
  assign n11624 = n11623 ^ n2175 ;
  assign n11625 = n11454 ^ n2511 ;
  assign n11626 = n11594 & ~n11625 ;
  assign n11627 = n11626 ^ n11263 ;
  assign n11628 = n11627 ^ n2366 ;
  assign n11826 = ~n11452 & n11594 ;
  assign n11827 = n11826 ^ n11266 ;
  assign n11819 = n11446 ^ n2894 ;
  assign n11820 = n11594 & n11819 ;
  assign n11821 = n11820 ^ n11448 ;
  assign n11629 = ~n11444 & n11594 ;
  assign n11630 = n11629 ^ n11269 ;
  assign n11631 = n11630 ^ n2894 ;
  assign n11632 = n11439 & n11594 ;
  assign n11633 = n11632 ^ n11441 ;
  assign n11815 = n11633 ^ n2894 ;
  assign n11634 = n11633 ^ n3093 ;
  assign n11807 = n11436 ^ n3538 ;
  assign n11808 = n11594 & n11807 ;
  assign n11809 = n11808 ^ n11273 ;
  assign n11635 = ~n11434 & n11594 ;
  assign n11636 = n11635 ^ n11277 ;
  assign n11637 = n11636 ^ n3538 ;
  assign n11638 = n11428 ^ n3908 ;
  assign n11639 = n11594 & n11638 ;
  assign n11640 = n11639 ^ n11430 ;
  assign n11641 = n11640 ^ n3722 ;
  assign n11796 = n11423 & n11594 ;
  assign n11797 = n11796 ^ n11425 ;
  assign n11642 = n11418 & n11594 ;
  assign n11643 = n11642 ^ n11420 ;
  assign n11644 = n11643 ^ n4153 ;
  assign n11645 = n11413 & n11594 ;
  assign n11646 = n11645 ^ n11415 ;
  assign n11647 = n11646 ^ n4356 ;
  assign n11784 = n11410 ^ n4812 ;
  assign n11785 = n11594 & n11784 ;
  assign n11786 = n11785 ^ n11280 ;
  assign n11778 = n11408 & n11594 ;
  assign n11779 = n11778 ^ n11283 ;
  assign n11772 = n11405 & n11594 ;
  assign n11773 = n11772 ^ n11287 ;
  assign n11648 = n11400 & n11594 ;
  assign n11649 = n11648 ^ n11402 ;
  assign n11650 = n11649 ^ n5317 ;
  assign n11651 = n11398 & n11594 ;
  assign n11652 = n11651 ^ n11290 ;
  assign n11653 = n11652 ^ n5562 ;
  assign n11654 = ~n11396 & n11594 ;
  assign n11655 = n11654 ^ n11294 ;
  assign n11656 = n11655 ^ n5830 ;
  assign n11657 = ~n11394 & n11594 ;
  assign n11658 = n11657 ^ n11297 ;
  assign n11659 = n11658 ^ n6115 ;
  assign n11756 = n11387 ^ n6673 ;
  assign n11757 = n11594 & n11756 ;
  assign n11758 = n11757 ^ n11390 ;
  assign n11660 = n11382 & n11594 ;
  assign n11661 = n11660 ^ n11384 ;
  assign n11662 = n11661 ^ n6673 ;
  assign n11663 = n11380 & n11594 ;
  assign n11664 = n11663 ^ n11300 ;
  assign n11665 = n11664 ^ n6959 ;
  assign n11668 = ~n11369 & n11594 ;
  assign n11669 = n11668 ^ n11371 ;
  assign n11670 = n11669 ^ n7584 ;
  assign n11673 = n11361 & n11594 ;
  assign n11674 = n11673 ^ n11303 ;
  assign n11675 = n11674 ^ n8253 ;
  assign n11676 = ~n11359 & n11594 ;
  assign n11677 = n11676 ^ n11306 ;
  assign n11678 = n11677 ^ n8586 ;
  assign n11679 = n11357 & n11594 ;
  assign n11680 = n11679 ^ n11309 ;
  assign n11681 = n11680 ^ n8910 ;
  assign n11682 = ~n11345 & n11594 ;
  assign n11683 = n11682 ^ n11319 ;
  assign n11684 = n11683 ^ n9542 ;
  assign n11685 = ~n11343 & n11594 ;
  assign n11686 = n11685 ^ n11324 ;
  assign n11687 = n11686 ^ n10108 ;
  assign n11689 = n11233 ^ x17 ;
  assign n11690 = n11689 ^ n11594 ;
  assign n11691 = ~x14 & ~x15 ;
  assign n11692 = n11691 ^ n11233 ;
  assign n11693 = n11692 ^ x16 ;
  assign n11694 = ~n11690 & n11693 ;
  assign n11702 = n11694 ^ n11326 ;
  assign n11688 = n11594 ^ n11233 ;
  assign n11695 = n11694 ^ n11688 ;
  assign n11696 = n11695 ^ n11694 ;
  assign n11697 = n11694 ^ n11689 ;
  assign n11698 = n11697 ^ n11694 ;
  assign n11699 = n11696 & ~n11698 ;
  assign n11700 = n11699 ^ n11694 ;
  assign n11701 = x16 & n11700 ;
  assign n11703 = n11702 ^ n11701 ;
  assign n11705 = n11330 ^ n11233 ;
  assign n11706 = n11594 & n11705 ;
  assign n11704 = n11233 ^ x18 ;
  assign n11707 = n11706 ^ n11704 ;
  assign n11708 = n11707 ^ n10875 ;
  assign n11709 = ~n11703 & n11708 ;
  assign n11710 = n11709 ^ n11327 ;
  assign n11711 = ~x18 & n11330 ;
  assign n11712 = n11711 ^ n11326 ;
  assign n11720 = n11712 ^ x19 ;
  assign n11717 = ~x18 & n11233 ;
  assign n11718 = n11717 ^ n11712 ;
  assign n11719 = ~n11594 & ~n11718 ;
  assign n11721 = n11720 ^ n11719 ;
  assign n11722 = n11721 ^ n10468 ;
  assign n11723 = ~n11710 & n11722 ;
  assign n11724 = n11723 ^ n10639 ;
  assign n11725 = ~n11687 & ~n11724 ;
  assign n11726 = n11725 ^ n10203 ;
  assign n11727 = n11684 & ~n11726 ;
  assign n11728 = n11727 ^ n9628 ;
  assign n11729 = ~n11347 & n11594 ;
  assign n11730 = n11729 ^ n11354 ;
  assign n11731 = n11730 ^ n9217 ;
  assign n11732 = n11728 & ~n11731 ;
  assign n11733 = n11732 ^ n9285 ;
  assign n11734 = ~n11681 & n11733 ;
  assign n11735 = n11734 ^ n11680 ;
  assign n11736 = n11735 ^ n11677 ;
  assign n11737 = n11678 & n11736 ;
  assign n11738 = n11737 ^ n8586 ;
  assign n11739 = n11738 ^ n11674 ;
  assign n11740 = ~n11675 & n11739 ;
  assign n11741 = n11740 ^ n8253 ;
  assign n11671 = n11364 & n11594 ;
  assign n11672 = n11671 ^ n11366 ;
  assign n11742 = n11741 ^ n11672 ;
  assign n11743 = n11741 ^ n7891 ;
  assign n11744 = ~n11742 & ~n11743 ;
  assign n11745 = n11744 ^ n7971 ;
  assign n11746 = n11670 & n11745 ;
  assign n11747 = n11746 ^ n11669 ;
  assign n11666 = ~n11374 & n11594 ;
  assign n11667 = n11666 ^ n11376 ;
  assign n11748 = n11747 ^ n11667 ;
  assign n11749 = n11747 ^ n7277 ;
  assign n11750 = ~n11748 & n11749 ;
  assign n11751 = n11750 ^ n7339 ;
  assign n11752 = n11665 & n11751 ;
  assign n11753 = n11752 ^ n7011 ;
  assign n11754 = n11662 & n11753 ;
  assign n11755 = n11754 ^ n6673 ;
  assign n11759 = n11758 ^ n11755 ;
  assign n11760 = n11758 ^ n6389 ;
  assign n11761 = n11759 & n11760 ;
  assign n11762 = n11761 ^ n6423 ;
  assign n11763 = ~n11659 & ~n11762 ;
  assign n11764 = n11763 ^ n6429 ;
  assign n11765 = ~n11656 & ~n11764 ;
  assign n11766 = n11765 ^ n11655 ;
  assign n11767 = n11766 ^ n11652 ;
  assign n11768 = ~n11653 & ~n11767 ;
  assign n11769 = n11768 ^ n5885 ;
  assign n11770 = n11650 & ~n11769 ;
  assign n11771 = n11770 ^ n11649 ;
  assign n11774 = n11773 ^ n11771 ;
  assign n11775 = n11773 ^ n5073 ;
  assign n11776 = ~n11774 & n11775 ;
  assign n11777 = n11776 ^ n5073 ;
  assign n11780 = n11779 ^ n11777 ;
  assign n11781 = n11779 ^ n4812 ;
  assign n11782 = n11780 & ~n11781 ;
  assign n11783 = n11782 ^ n4812 ;
  assign n11787 = n11786 ^ n11783 ;
  assign n11788 = n11786 ^ n4583 ;
  assign n11789 = n11787 & ~n11788 ;
  assign n11790 = n11789 ^ n4645 ;
  assign n11791 = n11647 & ~n11790 ;
  assign n11792 = n11791 ^ n11646 ;
  assign n11793 = n11792 ^ n11643 ;
  assign n11794 = ~n11644 & n11793 ;
  assign n11795 = n11794 ^ n4153 ;
  assign n11798 = n11797 ^ n11795 ;
  assign n11799 = n11797 ^ n3908 ;
  assign n11800 = ~n11798 & n11799 ;
  assign n11801 = n11800 ^ n3908 ;
  assign n11802 = n11801 ^ n11640 ;
  assign n11803 = n11641 & n11802 ;
  assign n11804 = n11803 ^ n3795 ;
  assign n11805 = n11637 & n11804 ;
  assign n11806 = n11805 ^ n3538 ;
  assign n11810 = n11809 ^ n11806 ;
  assign n11811 = n11809 ^ n3320 ;
  assign n11812 = ~n11810 & n11811 ;
  assign n11813 = n11812 ^ n3387 ;
  assign n11814 = n11634 & n11813 ;
  assign n11816 = n11815 ^ n11814 ;
  assign n11817 = n11631 & n11816 ;
  assign n11818 = n11817 ^ n2894 ;
  assign n11822 = n11821 ^ n11818 ;
  assign n11823 = n11821 ^ n2707 ;
  assign n11824 = ~n11822 & ~n11823 ;
  assign n11825 = n11824 ^ n2707 ;
  assign n11828 = n11827 ^ n11825 ;
  assign n11829 = n11827 ^ n2511 ;
  assign n11830 = ~n11828 & ~n11829 ;
  assign n11831 = n11830 ^ n2530 ;
  assign n11832 = n11628 & n11831 ;
  assign n11833 = n11832 ^ n2399 ;
  assign n11834 = ~n11624 & n11833 ;
  assign n11835 = n11834 ^ n2204 ;
  assign n11836 = n11621 & n11835 ;
  assign n11837 = n11836 ^ n2008 ;
  assign n11617 = n11467 & n11594 ;
  assign n11618 = n11617 ^ n11258 ;
  assign n11838 = n11837 ^ n11618 ;
  assign n11839 = n11837 ^ n1739 ;
  assign n11840 = n11838 & ~n11839 ;
  assign n11841 = n11840 ^ n1763 ;
  assign n11842 = n11616 & n11841 ;
  assign n11844 = n11843 ^ n11842 ;
  assign n11845 = ~n11475 & n11594 ;
  assign n11846 = n11845 ^ n11473 ;
  assign n11847 = n11846 ^ n1427 ;
  assign n11848 = ~n11844 & ~n11847 ;
  assign n11849 = n11848 ^ n1450 ;
  assign n11924 = n11583 ^ n138 ;
  assign n11925 = n11594 & n11924 ;
  assign n11926 = n11925 ^ n11586 ;
  assign n11927 = ~n183 & ~n11926 ;
  assign n11928 = n11927 ^ n11926 ;
  assign n11917 = n11577 & n11594 ;
  assign n11918 = n11917 ^ n11569 ;
  assign n11595 = ~n11535 & n11594 ;
  assign n11596 = n11595 ^ n11573 ;
  assign n11597 = n11596 ^ n188 ;
  assign n11598 = n11521 ^ n401 ;
  assign n11599 = n11594 & ~n11598 ;
  assign n11600 = n11599 ^ n11523 ;
  assign n11601 = n11600 ^ n341 ;
  assign n11889 = ~n11516 & n11594 ;
  assign n11890 = n11889 ^ n11518 ;
  assign n11602 = ~n11514 & n11594 ;
  assign n11603 = n11602 ^ n11243 ;
  assign n11604 = n11603 ^ n457 ;
  assign n11605 = ~n11512 & n11594 ;
  assign n11606 = n11605 ^ n11246 ;
  assign n11607 = n11606 ^ n534 ;
  assign n11608 = n11506 & n11594 ;
  assign n11609 = n11608 ^ n11508 ;
  assign n11610 = n11609 ^ n609 ;
  assign n11611 = ~n11480 & n11594 ;
  assign n11612 = n11611 ^ n11482 ;
  assign n11613 = n11612 ^ n1136 ;
  assign n11850 = ~n11478 & n11594 ;
  assign n11851 = n11850 ^ n11252 ;
  assign n11854 = n11851 ^ n1136 ;
  assign n11852 = n11851 ^ n1290 ;
  assign n11853 = n11849 & n11852 ;
  assign n11855 = n11854 ^ n11853 ;
  assign n11856 = ~n11613 & n11855 ;
  assign n11857 = n11856 ^ n1143 ;
  assign n11858 = n11485 & n11594 ;
  assign n11859 = n11858 ^ n11249 ;
  assign n11862 = n11859 ^ n1034 ;
  assign n11863 = ~n11857 & n11862 ;
  assign n11860 = n11859 ^ n892 ;
  assign n11864 = n11863 ^ n11860 ;
  assign n11865 = n11487 & n11594 ;
  assign n11866 = n11865 ^ n11489 ;
  assign n11867 = n11866 ^ n786 ;
  assign n11868 = n11867 ^ n927 ;
  assign n11869 = ~n11864 & ~n11868 ;
  assign n11870 = n11869 ^ n11867 ;
  assign n11871 = ~n11494 & n11594 ;
  assign n11872 = n11871 ^ n11496 ;
  assign n11873 = n11872 ^ n696 ;
  assign n11874 = n11873 ^ n842 ;
  assign n11875 = n11870 & ~n11874 ;
  assign n11876 = n11875 ^ n11873 ;
  assign n11877 = ~n11500 & n11594 ;
  assign n11878 = n11877 ^ n11502 ;
  assign n11879 = n11878 ^ n609 ;
  assign n11880 = n11879 ^ n835 ;
  assign n11881 = n11876 & n11880 ;
  assign n11882 = n11881 ^ n11879 ;
  assign n11883 = ~n11610 & ~n11882 ;
  assign n11884 = n11883 ^ n834 ;
  assign n11885 = n11607 & ~n11884 ;
  assign n11886 = n11885 ^ n750 ;
  assign n11887 = n11604 & n11886 ;
  assign n11888 = n11887 ^ n11603 ;
  assign n11891 = n11890 ^ n11888 ;
  assign n11892 = n11890 ^ n401 ;
  assign n11893 = ~n11891 & ~n11892 ;
  assign n11894 = n11893 ^ n462 ;
  assign n11895 = ~n11601 & n11894 ;
  assign n11896 = n11895 ^ n349 ;
  assign n11897 = n11527 ^ n341 ;
  assign n11898 = n11594 & n11897 ;
  assign n11899 = n11898 ^ n11239 ;
  assign n11900 = n11899 ^ n291 ;
  assign n11901 = ~n11896 & n11900 ;
  assign n11902 = n11901 ^ n307 ;
  assign n11903 = n11527 ^ n291 ;
  assign n11904 = n11903 ^ n349 ;
  assign n11905 = n11239 ^ n291 ;
  assign n11906 = n11905 ^ n349 ;
  assign n11907 = n11904 & ~n11906 ;
  assign n11908 = n11907 ^ n349 ;
  assign n11909 = n11594 & ~n11908 ;
  assign n11910 = n11909 ^ n11235 ;
  assign n11911 = n11910 ^ n245 ;
  assign n11912 = n11902 & n11911 ;
  assign n11913 = n11912 ^ n11910 ;
  assign n11914 = n11913 ^ n11596 ;
  assign n11915 = n11597 & ~n11914 ;
  assign n11916 = n11915 ^ n188 ;
  assign n11919 = n11918 ^ n11916 ;
  assign n11920 = n11916 ^ n157 ;
  assign n11921 = n11919 & ~n11920 ;
  assign n11922 = n11921 ^ n11918 ;
  assign n11929 = n138 & n11922 ;
  assign n11923 = n11922 ^ n138 ;
  assign n11930 = n11929 ^ n11923 ;
  assign n11931 = n11569 ^ n203 ;
  assign n11932 = n11931 ^ n11576 ;
  assign n11933 = n11932 ^ n203 ;
  assign n11936 = n11571 & ~n11933 ;
  assign n11937 = n11936 ^ n203 ;
  assign n11938 = n11594 & n11937 ;
  assign n11939 = n11938 ^ n11566 ;
  assign n11940 = n11930 & n11939 ;
  assign n11941 = ~n11929 & ~n11940 ;
  assign n11942 = ~n11559 & n11586 ;
  assign n11943 = n11942 ^ n11559 ;
  assign n11944 = ~n11562 & ~n11943 ;
  assign n11945 = n11589 ^ n138 ;
  assign n11946 = n11945 ^ n11559 ;
  assign n11947 = n11562 & n11946 ;
  assign n11948 = n11947 ^ n11588 ;
  assign n11949 = ~n183 & n11948 ;
  assign n11950 = ~n11590 & n11949 ;
  assign n11951 = ~n11944 & ~n11950 ;
  assign n11952 = n183 & n11591 ;
  assign n11953 = n11952 ^ n11563 ;
  assign n11954 = n11942 & n11952 ;
  assign n11955 = ~n11953 & n11954 ;
  assign n11956 = n11955 ^ n11953 ;
  assign n11957 = n11951 & ~n11956 ;
  assign n11958 = ~n11941 & ~n11957 ;
  assign n11959 = n11928 & n11958 ;
  assign n11960 = n11959 ^ n11957 ;
  assign n12288 = ~n11849 & n11960 ;
  assign n12289 = n12288 ^ n11851 ;
  assign n12277 = ~n11841 & n11960 ;
  assign n12278 = n12277 ^ n11615 ;
  assign n12026 = ~n11839 & n11960 ;
  assign n12027 = n12026 ^ n11618 ;
  assign n12028 = n12027 ^ n1572 ;
  assign n12029 = n11833 & n11960 ;
  assign n12030 = n12029 ^ n11623 ;
  assign n12031 = n12030 ^ n2008 ;
  assign n12032 = n11831 & n11960 ;
  assign n12033 = n12032 ^ n11627 ;
  assign n12034 = n12033 ^ n2175 ;
  assign n12035 = n11825 ^ n2511 ;
  assign n12036 = n11960 & ~n12035 ;
  assign n12037 = n12036 ^ n11827 ;
  assign n12038 = n12037 ^ n2366 ;
  assign n12257 = n11818 ^ n2707 ;
  assign n12258 = n11960 & ~n12257 ;
  assign n12259 = n12258 ^ n11821 ;
  assign n12039 = n11816 & n11960 ;
  assign n12040 = n12039 ^ n11630 ;
  assign n12041 = n12040 ^ n2707 ;
  assign n12042 = ~n11813 & n11960 ;
  assign n12043 = n12042 ^ n11633 ;
  assign n12044 = n12043 ^ n2894 ;
  assign n12048 = n11804 & n11960 ;
  assign n12049 = n12048 ^ n11636 ;
  assign n12050 = n12049 ^ n3320 ;
  assign n12051 = n11795 ^ n3908 ;
  assign n12052 = n11960 & n12051 ;
  assign n12053 = n12052 ^ n11797 ;
  assign n12054 = n12053 ^ n3722 ;
  assign n12232 = n11792 ^ n4153 ;
  assign n12233 = n11960 & n12232 ;
  assign n12234 = n12233 ^ n11643 ;
  assign n12055 = n11790 & n11960 ;
  assign n12056 = n12055 ^ n11646 ;
  assign n12057 = n12056 ^ n4153 ;
  assign n12223 = n11783 ^ n4583 ;
  assign n12224 = n11960 & n12223 ;
  assign n12225 = n12224 ^ n11786 ;
  assign n12228 = n12225 ^ n4153 ;
  assign n12208 = n4583 & ~n4854 ;
  assign n12198 = n11771 ^ n5073 ;
  assign n12199 = n11960 & n12198 ;
  assign n12200 = n12199 ^ n11773 ;
  assign n12058 = n11777 ^ n4812 ;
  assign n12059 = n11960 & n12058 ;
  assign n12060 = n12059 ^ n11779 ;
  assign n12209 = n12200 ^ n12060 ;
  assign n12210 = n12208 & ~n12209 ;
  assign n12061 = n11769 & n11960 ;
  assign n12062 = n12061 ^ n11649 ;
  assign n12063 = n12062 ^ n5073 ;
  assign n12064 = n11766 ^ n5562 ;
  assign n12065 = n11960 & ~n12064 ;
  assign n12066 = n12065 ^ n11652 ;
  assign n12068 = n12066 ^ n5317 ;
  assign n12188 = n11764 & n11960 ;
  assign n12189 = n12188 ^ n11655 ;
  assign n12069 = ~n11762 & n11960 ;
  assign n12070 = n12069 ^ n11658 ;
  assign n12071 = n12070 ^ n5830 ;
  assign n12072 = n11755 ^ n6389 ;
  assign n12073 = n11960 & ~n12072 ;
  assign n12074 = n12073 ^ n11758 ;
  assign n12075 = n12074 ^ n6115 ;
  assign n12176 = n11753 & n11960 ;
  assign n12177 = n12176 ^ n11661 ;
  assign n12077 = n11751 & n11960 ;
  assign n12078 = n12077 ^ n11664 ;
  assign n12079 = n12078 ^ n6673 ;
  assign n12080 = n11749 & n11960 ;
  assign n12081 = n12080 ^ n11667 ;
  assign n12082 = n12081 ^ n6959 ;
  assign n12083 = ~n11745 & n11960 ;
  assign n12084 = n12083 ^ n11669 ;
  assign n12085 = n12084 ^ n7277 ;
  assign n12086 = ~n11743 & n11960 ;
  assign n12087 = n12086 ^ n11672 ;
  assign n12167 = n12087 ^ n7277 ;
  assign n12088 = n12087 ^ n7584 ;
  assign n12159 = n11738 ^ n8253 ;
  assign n12160 = n11960 & n12159 ;
  assign n12161 = n12160 ^ n11674 ;
  assign n12152 = n11735 ^ n8586 ;
  assign n12153 = n11960 & ~n12152 ;
  assign n12154 = n12153 ^ n11677 ;
  assign n12089 = ~n11733 & n11960 ;
  assign n12090 = n12089 ^ n11680 ;
  assign n12091 = n12090 ^ n8586 ;
  assign n12092 = ~n11726 & n11960 ;
  assign n12093 = n12092 ^ n11683 ;
  assign n12094 = n12093 ^ n9217 ;
  assign n12137 = ~n11724 & n11960 ;
  assign n12138 = n12137 ^ n11686 ;
  assign n12095 = ~n11710 & n11960 ;
  assign n12096 = n12095 ^ n11721 ;
  assign n12097 = n12096 ^ n10108 ;
  assign n12098 = ~n11703 & n11960 ;
  assign n12099 = n12098 ^ n11707 ;
  assign n12100 = n12099 ^ n10468 ;
  assign n12101 = n11691 ^ n11594 ;
  assign n12102 = n11960 & n12101 ;
  assign n12103 = n12102 ^ n11594 ;
  assign n12127 = x16 & n12103 ;
  assign n12125 = n11692 & n11960 ;
  assign n12124 = n11594 ^ x17 ;
  assign n12126 = n12125 ^ n12124 ;
  assign n12128 = n12127 ^ n12126 ;
  assign n12104 = n12103 ^ x16 ;
  assign n12105 = n12104 ^ n11233 ;
  assign n12106 = n11594 ^ x15 ;
  assign n12107 = n12106 ^ n11960 ;
  assign n12109 = ~x12 & ~x13 ;
  assign n12108 = n11594 ^ x14 ;
  assign n12110 = n12109 ^ n12108 ;
  assign n12111 = ~n12107 & n12110 ;
  assign n12120 = n12111 ^ n11688 ;
  assign n12112 = n11960 ^ n11594 ;
  assign n12117 = ~n12106 & n12112 ;
  assign n12118 = n12117 ^ n12111 ;
  assign n12119 = x14 & n12118 ;
  assign n12121 = n12120 ^ n12119 ;
  assign n12122 = ~n12105 & n12121 ;
  assign n12123 = n12122 ^ n11233 ;
  assign n12129 = n12128 ^ n12123 ;
  assign n12130 = n12128 ^ n10875 ;
  assign n12131 = n12129 & n12130 ;
  assign n12132 = n12131 ^ n11327 ;
  assign n12133 = ~n12100 & ~n12132 ;
  assign n12134 = n12133 ^ n10639 ;
  assign n12135 = ~n12097 & n12134 ;
  assign n12136 = n12135 ^ n12096 ;
  assign n12139 = n12138 ^ n12136 ;
  assign n12140 = n12138 ^ n9542 ;
  assign n12141 = ~n12139 & n12140 ;
  assign n12142 = n12141 ^ n9628 ;
  assign n12143 = n12094 & n12142 ;
  assign n12144 = n12143 ^ n9285 ;
  assign n12145 = n11728 & n11960 ;
  assign n12146 = n12145 ^ n11730 ;
  assign n12147 = n12146 ^ n8910 ;
  assign n12148 = ~n12144 & n12147 ;
  assign n12149 = n12148 ^ n9005 ;
  assign n12150 = ~n12091 & n12149 ;
  assign n12151 = n12150 ^ n8586 ;
  assign n12155 = n12154 ^ n12151 ;
  assign n12156 = n12154 ^ n8253 ;
  assign n12157 = ~n12155 & n12156 ;
  assign n12158 = n12157 ^ n8253 ;
  assign n12162 = n12161 ^ n12158 ;
  assign n12163 = n12161 ^ n7891 ;
  assign n12164 = n12162 & n12163 ;
  assign n12165 = n12164 ^ n7971 ;
  assign n12166 = n12088 & n12165 ;
  assign n12168 = n12167 ^ n12166 ;
  assign n12169 = n12085 & n12168 ;
  assign n12170 = n12169 ^ n7339 ;
  assign n12171 = n12082 & n12170 ;
  assign n12172 = n12171 ^ n7011 ;
  assign n12173 = n12079 & n12172 ;
  assign n12174 = n12173 ^ n6673 ;
  assign n12076 = n12074 ^ n6389 ;
  assign n12175 = n12174 ^ n12076 ;
  assign n12178 = n12177 ^ n12175 ;
  assign n12179 = n12178 ^ n12076 ;
  assign n12180 = n12174 ^ n12074 ;
  assign n12181 = n12180 ^ n12076 ;
  assign n12182 = ~n12179 & ~n12181 ;
  assign n12183 = n12182 ^ n12076 ;
  assign n12184 = ~n12075 & ~n12183 ;
  assign n12185 = n12184 ^ n6429 ;
  assign n12186 = ~n12071 & ~n12185 ;
  assign n12187 = n12186 ^ n12070 ;
  assign n12190 = n12189 ^ n12187 ;
  assign n12191 = n12189 ^ n5562 ;
  assign n12192 = ~n12190 & ~n12191 ;
  assign n12193 = n12192 ^ n5885 ;
  assign n12194 = ~n12068 & ~n12193 ;
  assign n12067 = n12066 ^ n5073 ;
  assign n12195 = n12194 ^ n12067 ;
  assign n12196 = n12063 & ~n12195 ;
  assign n12197 = n12196 ^ n5073 ;
  assign n12201 = n12200 ^ n12197 ;
  assign n12202 = n12201 ^ n4583 ;
  assign n12204 = n4812 & n12202 ;
  assign n12205 = n12204 ^ n4583 ;
  assign n12206 = ~n12060 & n12205 ;
  assign n12207 = n12206 ^ n4356 ;
  assign n12211 = n12210 ^ n12207 ;
  assign n12212 = n12211 ^ n4356 ;
  assign n12213 = n12200 ^ n4583 ;
  assign n12214 = n12213 ^ n12197 ;
  assign n12215 = n12060 ^ n4812 ;
  assign n12216 = n12200 & n12215 ;
  assign n12217 = n12216 ^ n4812 ;
  assign n12218 = ~n12214 & n12217 ;
  assign n12219 = n12218 ^ n12200 ;
  assign n12220 = n12197 & n12219 ;
  assign n12221 = ~n12212 & n12220 ;
  assign n12222 = n12221 ^ n12211 ;
  assign n12226 = n12225 ^ n4356 ;
  assign n12227 = ~n12222 & ~n12226 ;
  assign n12229 = n12228 ^ n12227 ;
  assign n12230 = n12057 & ~n12229 ;
  assign n12231 = n12230 ^ n4153 ;
  assign n12235 = n12234 ^ n12231 ;
  assign n12236 = n12234 ^ n3908 ;
  assign n12237 = n12235 & ~n12236 ;
  assign n12238 = n12237 ^ n3961 ;
  assign n12239 = ~n12054 & ~n12238 ;
  assign n12240 = n12239 ^ n3795 ;
  assign n12241 = n11801 ^ n3722 ;
  assign n12242 = n11960 & ~n12241 ;
  assign n12243 = n12242 ^ n11640 ;
  assign n12244 = n12243 ^ n3538 ;
  assign n12245 = n12240 & n12244 ;
  assign n12246 = n12245 ^ n3596 ;
  assign n12247 = n12050 & n12246 ;
  assign n12248 = n12247 ^ n3320 ;
  assign n12045 = n11806 ^ n3320 ;
  assign n12046 = n11960 & n12045 ;
  assign n12047 = n12046 ^ n11809 ;
  assign n12249 = n12248 ^ n12047 ;
  assign n12250 = n12047 ^ n3093 ;
  assign n12251 = ~n12249 & ~n12250 ;
  assign n12252 = n12251 ^ n3363 ;
  assign n12253 = n12044 & n12252 ;
  assign n12254 = n12253 ^ n3396 ;
  assign n12255 = ~n12041 & ~n12254 ;
  assign n12256 = n12255 ^ n2707 ;
  assign n12260 = n12259 ^ n12256 ;
  assign n12261 = n12259 ^ n2511 ;
  assign n12262 = n12260 & n12261 ;
  assign n12263 = n12262 ^ n2530 ;
  assign n12264 = ~n12038 & n12263 ;
  assign n12265 = n12264 ^ n2399 ;
  assign n12266 = n12034 & n12265 ;
  assign n12267 = n12266 ^ n2204 ;
  assign n12268 = ~n12031 & n12267 ;
  assign n12269 = n12268 ^ n2064 ;
  assign n12270 = n11835 & n11960 ;
  assign n12271 = n12270 ^ n11620 ;
  assign n12272 = n12271 ^ n1739 ;
  assign n12273 = ~n12269 & ~n12272 ;
  assign n12274 = n12273 ^ n1763 ;
  assign n12275 = ~n12028 & n12274 ;
  assign n12276 = n12275 ^ n12027 ;
  assign n12279 = n12278 ^ n12276 ;
  assign n12280 = n12278 ^ n1427 ;
  assign n12281 = n12279 & ~n12280 ;
  assign n12282 = n12281 ^ n1450 ;
  assign n12283 = ~n11844 & n11960 ;
  assign n12284 = n12283 ^ n11846 ;
  assign n12285 = n12284 ^ n1290 ;
  assign n12286 = n12282 & n12285 ;
  assign n12287 = n12286 ^ n12284 ;
  assign n12290 = n12289 ^ n12287 ;
  assign n12291 = n12289 ^ n1136 ;
  assign n12292 = ~n12290 & n12291 ;
  assign n12293 = n12292 ^ n1143 ;
  assign n12294 = n11855 & n11960 ;
  assign n12295 = n12294 ^ n11612 ;
  assign n12296 = n12295 ^ n1034 ;
  assign n12297 = n12293 & ~n12296 ;
  assign n12298 = n12297 ^ n1072 ;
  assign n12299 = n11857 & n11960 ;
  assign n12300 = n12299 ^ n11859 ;
  assign n12303 = n12300 ^ n892 ;
  assign n12304 = ~n12298 & n12303 ;
  assign n12301 = n12300 ^ n786 ;
  assign n12305 = n12304 ^ n12301 ;
  assign n12306 = n11864 & n11960 ;
  assign n12307 = n12306 ^ n11866 ;
  assign n12308 = n12307 ^ n696 ;
  assign n12309 = n12308 ^ n842 ;
  assign n12310 = ~n12305 & ~n12309 ;
  assign n12311 = n12310 ^ n12308 ;
  assign n11961 = n11923 & n11960 ;
  assign n11962 = n11961 ^ n11939 ;
  assign n11963 = n11962 ^ n183 ;
  assign n11964 = n183 & ~n11941 ;
  assign n11965 = n11927 & ~n11939 ;
  assign n11967 = ~n11929 & n11957 ;
  assign n11968 = n11965 & n11967 ;
  assign n11966 = n11965 ^ n11926 ;
  assign n11969 = n11968 ^ n11966 ;
  assign n11971 = n11969 ^ n11957 ;
  assign n11973 = n11971 ^ n11928 ;
  assign n11970 = n11969 ^ n11929 ;
  assign n11972 = n11971 ^ n11970 ;
  assign n11974 = n11973 ^ n11972 ;
  assign n11975 = n11974 ^ n11940 ;
  assign n11976 = n11969 ^ n11940 ;
  assign n11977 = n11975 & ~n11976 ;
  assign n11978 = n11977 ^ n11940 ;
  assign n11987 = n11976 ^ n11975 ;
  assign n11988 = n11987 ^ n11940 ;
  assign n11979 = n11969 ^ n11928 ;
  assign n11980 = n11979 ^ n11940 ;
  assign n11981 = n11980 ^ n11974 ;
  assign n11982 = n11981 ^ n11971 ;
  assign n11983 = n11974 ^ n11971 ;
  assign n11984 = n11983 ^ n11969 ;
  assign n11985 = n11984 ^ n11940 ;
  assign n11986 = ~n11982 & ~n11985 ;
  assign n11989 = n11988 ^ n11986 ;
  assign n11990 = n11978 & ~n11989 ;
  assign n11991 = n11990 ^ n11940 ;
  assign n11992 = n11991 ^ n11979 ;
  assign n11993 = n11992 ^ n11940 ;
  assign n11994 = ~n1355 & ~n11939 ;
  assign n11995 = ~n11922 & n11957 ;
  assign n11996 = n11994 & n11995 ;
  assign n11997 = n11996 ^ n11926 ;
  assign n11998 = ~n11993 & ~n11997 ;
  assign n11999 = n11998 ^ n11993 ;
  assign n12000 = n11964 & ~n11999 ;
  assign n12001 = n12000 ^ n11998 ;
  assign n12002 = n11920 & n11960 ;
  assign n12003 = n12002 ^ n11918 ;
  assign n12004 = n12003 ^ n138 ;
  assign n12005 = ~n11902 & n11960 ;
  assign n12006 = n12005 ^ n11910 ;
  assign n12007 = n12006 ^ n188 ;
  assign n12008 = ~n11896 & n11960 ;
  assign n12009 = n12008 ^ n11899 ;
  assign n12010 = n12009 ^ n12006 ;
  assign n12011 = n12010 ^ n12009 ;
  assign n12012 = n12011 ^ n245 ;
  assign n12013 = n12012 ^ n12010 ;
  assign n12014 = ~n11886 & n11960 ;
  assign n12015 = n12014 ^ n11603 ;
  assign n12016 = n12015 ^ n401 ;
  assign n12017 = ~n11884 & n11960 ;
  assign n12018 = n12017 ^ n11606 ;
  assign n12019 = n12018 ^ n12015 ;
  assign n12020 = n12019 ^ n12018 ;
  assign n12021 = n12020 ^ n457 ;
  assign n12022 = n12021 ^ n12019 ;
  assign n12023 = ~n11876 & n11960 ;
  assign n12024 = n12023 ^ n11878 ;
  assign n12025 = n12024 ^ n609 ;
  assign n12312 = ~n11870 & n11960 ;
  assign n12313 = n12312 ^ n11872 ;
  assign n12314 = n12313 ^ n609 ;
  assign n12315 = n12314 ^ n835 ;
  assign n12316 = n12311 & ~n12315 ;
  assign n12317 = n12316 ^ n12314 ;
  assign n12318 = ~n12025 & n12317 ;
  assign n12319 = n12318 ^ n834 ;
  assign n12320 = ~n11882 & n11960 ;
  assign n12321 = n12320 ^ n11609 ;
  assign n12322 = n12321 ^ n534 ;
  assign n12323 = ~n12319 & n12322 ;
  assign n12324 = n12323 ^ n750 ;
  assign n12327 = ~n12022 & n12324 ;
  assign n12328 = n12327 ^ n12019 ;
  assign n12329 = ~n12016 & n12328 ;
  assign n12330 = n12329 ^ n462 ;
  assign n12331 = n11888 ^ n401 ;
  assign n12332 = n11960 & ~n12331 ;
  assign n12333 = n12332 ^ n11890 ;
  assign n12334 = n12333 ^ n341 ;
  assign n12335 = n12330 & ~n12334 ;
  assign n12336 = n12335 ^ n349 ;
  assign n12337 = n11894 & n11960 ;
  assign n12338 = n12337 ^ n11600 ;
  assign n12339 = n12338 ^ n291 ;
  assign n12340 = ~n12336 & n12339 ;
  assign n12341 = n12340 ^ n307 ;
  assign n12344 = ~n12013 & n12341 ;
  assign n12345 = n12344 ^ n12010 ;
  assign n12346 = n12007 & n12345 ;
  assign n12347 = n12346 ^ n203 ;
  assign n12348 = n11913 ^ n188 ;
  assign n12349 = n11960 & n12348 ;
  assign n12350 = n12349 ^ n11596 ;
  assign n12351 = n12350 ^ n157 ;
  assign n12352 = ~n12347 & n12351 ;
  assign n12353 = n12352 ^ n12350 ;
  assign n12354 = n12353 ^ n12003 ;
  assign n12355 = n12004 & ~n12354 ;
  assign n12356 = n12355 ^ n138 ;
  assign n12357 = n12001 & n12356 ;
  assign n12358 = ~n11963 & n12357 ;
  assign n12359 = n12358 ^ n12001 ;
  assign n12360 = ~n12311 & ~n12359 ;
  assign n12361 = n12360 ^ n12313 ;
  assign n12363 = n12361 ^ n609 ;
  assign n12364 = n12293 & ~n12359 ;
  assign n12365 = n12364 ^ n12295 ;
  assign n12366 = n12365 ^ n892 ;
  assign n12628 = ~n12282 & ~n12359 ;
  assign n12629 = n12628 ^ n12284 ;
  assign n12367 = ~n12274 & ~n12359 ;
  assign n12368 = n12367 ^ n12027 ;
  assign n12369 = n12368 ^ n1427 ;
  assign n12614 = ~n12269 & ~n12359 ;
  assign n12615 = n12614 ^ n12271 ;
  assign n12618 = n12615 ^ n1427 ;
  assign n12370 = n12265 & ~n12359 ;
  assign n12371 = n12370 ^ n12033 ;
  assign n12372 = n12371 ^ n2008 ;
  assign n12373 = n12256 ^ n2511 ;
  assign n12374 = ~n12359 & ~n12373 ;
  assign n12375 = n12374 ^ n12259 ;
  assign n12376 = n12375 ^ n2366 ;
  assign n12594 = ~n12254 & ~n12359 ;
  assign n12595 = n12594 ^ n12040 ;
  assign n12377 = n12252 & ~n12359 ;
  assign n12378 = n12377 ^ n12043 ;
  assign n12379 = n12378 ^ n2707 ;
  assign n12380 = n12248 ^ n3093 ;
  assign n12381 = ~n12359 & ~n12380 ;
  assign n12382 = n12381 ^ n12047 ;
  assign n12383 = n12382 ^ n2894 ;
  assign n12584 = n12246 & ~n12359 ;
  assign n12585 = n12584 ^ n12049 ;
  assign n12588 = n12585 ^ n2894 ;
  assign n12384 = n12240 & ~n12359 ;
  assign n12385 = n12384 ^ n12243 ;
  assign n12386 = n12385 ^ n3320 ;
  assign n12387 = ~n12238 & ~n12359 ;
  assign n12388 = n12387 ^ n12053 ;
  assign n12389 = n12388 ^ n3538 ;
  assign n12572 = n12231 ^ n3908 ;
  assign n12573 = ~n12359 & n12572 ;
  assign n12574 = n12573 ^ n12234 ;
  assign n12566 = ~n12229 & ~n12359 ;
  assign n12567 = n12566 ^ n12056 ;
  assign n12390 = n12197 ^ n4812 ;
  assign n12393 = n12213 ^ n12201 ;
  assign n12394 = n12393 ^ n12213 ;
  assign n12395 = ~n12390 & n12394 ;
  assign n12396 = n12395 ^ n12213 ;
  assign n12397 = ~n12359 & n12396 ;
  assign n12398 = n12397 ^ n12060 ;
  assign n12399 = n12398 ^ n4356 ;
  assign n12400 = ~n12195 & ~n12359 ;
  assign n12401 = n12400 ^ n12062 ;
  assign n12402 = n12401 ^ n4812 ;
  assign n12403 = n12193 & ~n12359 ;
  assign n12404 = n12403 ^ n12066 ;
  assign n12405 = n12404 ^ n5073 ;
  assign n12409 = n12185 & ~n12359 ;
  assign n12410 = n12409 ^ n12070 ;
  assign n12411 = n12410 ^ n5562 ;
  assign n12412 = n12174 ^ n6423 ;
  assign n12413 = n12412 ^ n12177 ;
  assign n12414 = n12413 ^ n6423 ;
  assign n12415 = n12174 ^ n6389 ;
  assign n12418 = ~n12414 & ~n12415 ;
  assign n12419 = n12418 ^ n6423 ;
  assign n12420 = ~n12359 & ~n12419 ;
  assign n12421 = n12420 ^ n12074 ;
  assign n12422 = n12421 ^ n5830 ;
  assign n12423 = n12172 & ~n12359 ;
  assign n12424 = n12423 ^ n12078 ;
  assign n12425 = n12424 ^ n6389 ;
  assign n12528 = n12170 & ~n12359 ;
  assign n12529 = n12528 ^ n12081 ;
  assign n12426 = ~n12165 & ~n12359 ;
  assign n12427 = n12426 ^ n12087 ;
  assign n12428 = n12427 ^ n7277 ;
  assign n12514 = n12158 ^ n7891 ;
  assign n12515 = ~n12359 & ~n12514 ;
  assign n12516 = n12515 ^ n12161 ;
  assign n12519 = n12516 ^ n7277 ;
  assign n12429 = n12136 ^ n9542 ;
  assign n12430 = ~n12359 & n12429 ;
  assign n12431 = n12430 ^ n12138 ;
  assign n12432 = n12431 ^ n9217 ;
  assign n12433 = ~n12132 & ~n12359 ;
  assign n12434 = n12433 ^ n12099 ;
  assign n12484 = n12434 ^ n9542 ;
  assign n12435 = n12434 ^ n10108 ;
  assign n12445 = ~x14 & n11960 ;
  assign n12436 = n12109 ^ n11960 ;
  assign n12439 = n12112 ^ x14 ;
  assign n12440 = n12439 ^ n12112 ;
  assign n12441 = n12436 & ~n12440 ;
  assign n12442 = n12441 ^ n12112 ;
  assign n12443 = ~n12359 & n12442 ;
  assign n12444 = n12443 ^ x15 ;
  assign n12446 = n12445 ^ n12444 ;
  assign n12447 = n12446 ^ n11233 ;
  assign n12449 = n12359 & n12436 ;
  assign n12448 = n12109 ^ x14 ;
  assign n12450 = n12449 ^ n12448 ;
  assign n12451 = n12450 ^ n11594 ;
  assign n12454 = ~x10 & ~x11 ;
  assign n12453 = n12359 ^ x13 ;
  assign n12455 = n12454 ^ n12453 ;
  assign n12456 = n12454 ^ n11960 ;
  assign n12457 = ~n12455 & n12456 ;
  assign n12465 = n12457 ^ n12112 ;
  assign n12452 = n12359 ^ n11960 ;
  assign n12458 = n12457 ^ n12452 ;
  assign n12459 = n12458 ^ n12457 ;
  assign n12460 = n12457 ^ n12453 ;
  assign n12461 = n12460 ^ n12457 ;
  assign n12462 = ~n12459 & ~n12461 ;
  assign n12463 = n12462 ^ n12457 ;
  assign n12464 = x12 & n12463 ;
  assign n12466 = n12465 ^ n12464 ;
  assign n12467 = ~n12451 & n12466 ;
  assign n12468 = n12467 ^ n11594 ;
  assign n12469 = n12468 ^ n12446 ;
  assign n12470 = ~n12447 & n12469 ;
  assign n12471 = n12470 ^ n11326 ;
  assign n12472 = n12121 & ~n12359 ;
  assign n12473 = n12472 ^ n12104 ;
  assign n12474 = n12473 ^ n10875 ;
  assign n12475 = ~n12471 & n12474 ;
  assign n12476 = n12475 ^ n11327 ;
  assign n12477 = n12123 ^ n10875 ;
  assign n12478 = ~n12359 & ~n12477 ;
  assign n12479 = n12478 ^ n12128 ;
  assign n12480 = n12479 ^ n10468 ;
  assign n12481 = ~n12476 & ~n12480 ;
  assign n12482 = n12481 ^ n10639 ;
  assign n12483 = n12435 & n12482 ;
  assign n12485 = n12484 ^ n12483 ;
  assign n12486 = ~n12134 & ~n12359 ;
  assign n12487 = n12486 ^ n12096 ;
  assign n12488 = n12487 ^ n9542 ;
  assign n12489 = ~n12485 & n12488 ;
  assign n12490 = n12489 ^ n9628 ;
  assign n12491 = n12432 & n12490 ;
  assign n12492 = n12491 ^ n9285 ;
  assign n12493 = n12142 & ~n12359 ;
  assign n12494 = n12493 ^ n12093 ;
  assign n12495 = n12494 ^ n8910 ;
  assign n12496 = ~n12492 & ~n12495 ;
  assign n12497 = n12496 ^ n9005 ;
  assign n12498 = ~n12144 & ~n12359 ;
  assign n12499 = n12498 ^ n12146 ;
  assign n12500 = n12499 ^ n8586 ;
  assign n12501 = n12497 & n12500 ;
  assign n12502 = n12501 ^ n8688 ;
  assign n12503 = n12149 & ~n12359 ;
  assign n12504 = n12503 ^ n12090 ;
  assign n12505 = n12504 ^ n8253 ;
  assign n12506 = n12502 & ~n12505 ;
  assign n12507 = n12506 ^ n8356 ;
  assign n12508 = n12151 ^ n8253 ;
  assign n12509 = ~n12359 & n12508 ;
  assign n12510 = n12509 ^ n12154 ;
  assign n12511 = n12510 ^ n7891 ;
  assign n12512 = ~n12507 & ~n12511 ;
  assign n12513 = n12512 ^ n7971 ;
  assign n12517 = n12516 ^ n7584 ;
  assign n12518 = n12513 & ~n12517 ;
  assign n12520 = n12519 ^ n12518 ;
  assign n12521 = n12428 & ~n12520 ;
  assign n12522 = n12521 ^ n7339 ;
  assign n12523 = n12168 & ~n12359 ;
  assign n12524 = n12523 ^ n12084 ;
  assign n12525 = n12524 ^ n6959 ;
  assign n12526 = n12522 & n12525 ;
  assign n12527 = n12526 ^ n6959 ;
  assign n12530 = n12529 ^ n12527 ;
  assign n12531 = n12529 ^ n6673 ;
  assign n12532 = ~n12530 & n12531 ;
  assign n12533 = n12532 ^ n6713 ;
  assign n12534 = ~n12425 & ~n12533 ;
  assign n12535 = n12534 ^ n6423 ;
  assign n12536 = ~n12359 & ~n12415 ;
  assign n12537 = n12536 ^ n12177 ;
  assign n12538 = n12537 ^ n6115 ;
  assign n12539 = ~n12535 & n12538 ;
  assign n12540 = n12539 ^ n6429 ;
  assign n12541 = ~n12422 & n12540 ;
  assign n12542 = n12541 ^ n5900 ;
  assign n12543 = ~n12411 & n12542 ;
  assign n12544 = n12543 ^ n5562 ;
  assign n12406 = n12187 ^ n5562 ;
  assign n12407 = ~n12359 & ~n12406 ;
  assign n12408 = n12407 ^ n12189 ;
  assign n12545 = n12544 ^ n12408 ;
  assign n12546 = n12408 ^ n5317 ;
  assign n12547 = n12545 & ~n12546 ;
  assign n12548 = n12547 ^ n5360 ;
  assign n12549 = ~n12405 & n12548 ;
  assign n12550 = n12549 ^ n5073 ;
  assign n12551 = n12550 ^ n12401 ;
  assign n12552 = n12402 & ~n12551 ;
  assign n12553 = n12552 ^ n4854 ;
  assign n12554 = ~n12359 & n12390 ;
  assign n12555 = n12554 ^ n12200 ;
  assign n12556 = n12555 ^ n4583 ;
  assign n12557 = n12553 & n12556 ;
  assign n12558 = n12557 ^ n4645 ;
  assign n12559 = ~n12399 & n12558 ;
  assign n12560 = n12559 ^ n4414 ;
  assign n12561 = n12222 & ~n12359 ;
  assign n12562 = n12561 ^ n12225 ;
  assign n12563 = n12562 ^ n4153 ;
  assign n12564 = n12560 & ~n12563 ;
  assign n12565 = n12564 ^ n4153 ;
  assign n12568 = n12567 ^ n12565 ;
  assign n12569 = n12567 ^ n3908 ;
  assign n12570 = ~n12568 & n12569 ;
  assign n12571 = n12570 ^ n3908 ;
  assign n12575 = n12574 ^ n12571 ;
  assign n12576 = n12574 ^ n3722 ;
  assign n12577 = n12575 & n12576 ;
  assign n12578 = n12577 ^ n3795 ;
  assign n12579 = ~n12389 & n12578 ;
  assign n12580 = n12579 ^ n3538 ;
  assign n12581 = n12580 ^ n12385 ;
  assign n12582 = n12386 & ~n12581 ;
  assign n12583 = n12582 ^ n3387 ;
  assign n12586 = n12585 ^ n3093 ;
  assign n12587 = n12583 & ~n12586 ;
  assign n12589 = n12588 ^ n12587 ;
  assign n12590 = ~n12383 & ~n12589 ;
  assign n12591 = n12590 ^ n3396 ;
  assign n12592 = ~n12379 & ~n12591 ;
  assign n12593 = n12592 ^ n2707 ;
  assign n12596 = n12595 ^ n12593 ;
  assign n12597 = n12595 ^ n2511 ;
  assign n12598 = n12596 & n12597 ;
  assign n12599 = n12598 ^ n2530 ;
  assign n12600 = n12376 & n12599 ;
  assign n12601 = n12600 ^ n2399 ;
  assign n12602 = n12263 & ~n12359 ;
  assign n12603 = n12602 ^ n12037 ;
  assign n12604 = n12603 ^ n2175 ;
  assign n12605 = n12601 & ~n12604 ;
  assign n12606 = n12605 ^ n2204 ;
  assign n12607 = n12372 & n12606 ;
  assign n12608 = n12607 ^ n2064 ;
  assign n12609 = n12267 & ~n12359 ;
  assign n12610 = n12609 ^ n12030 ;
  assign n12611 = n12610 ^ n1739 ;
  assign n12612 = ~n12608 & n12611 ;
  assign n12613 = n12612 ^ n1763 ;
  assign n12616 = n12615 ^ n1572 ;
  assign n12617 = n12613 & n12616 ;
  assign n12619 = n12618 ^ n12617 ;
  assign n12620 = n12369 & ~n12619 ;
  assign n12621 = n12620 ^ n1450 ;
  assign n12622 = n12276 ^ n1427 ;
  assign n12623 = ~n12359 & n12622 ;
  assign n12624 = n12623 ^ n12278 ;
  assign n12625 = n12624 ^ n1290 ;
  assign n12626 = n12621 & n12625 ;
  assign n12627 = n12626 ^ n12624 ;
  assign n12630 = n12629 ^ n12627 ;
  assign n12631 = n12629 ^ n1136 ;
  assign n12632 = ~n12630 & n12631 ;
  assign n12633 = n12632 ^ n1143 ;
  assign n12634 = n12287 ^ n1136 ;
  assign n12635 = ~n12359 & n12634 ;
  assign n12636 = n12635 ^ n12289 ;
  assign n12637 = n12636 ^ n892 ;
  assign n12638 = n12637 ^ n892 ;
  assign n12639 = n12638 ^ n1034 ;
  assign n12640 = ~n12633 & n12639 ;
  assign n12641 = n12640 ^ n12637 ;
  assign n12642 = ~n12366 & n12641 ;
  assign n12643 = n12642 ^ n927 ;
  assign n12644 = n12298 & ~n12359 ;
  assign n12645 = n12644 ^ n12300 ;
  assign n12646 = n12645 ^ n696 ;
  assign n12647 = n12646 ^ n696 ;
  assign n12648 = n12647 ^ n786 ;
  assign n12649 = ~n12643 & n12648 ;
  assign n12650 = n12649 ^ n12646 ;
  assign n12651 = n12305 & ~n12359 ;
  assign n12652 = n12651 ^ n12307 ;
  assign n12653 = n12652 ^ n609 ;
  assign n12654 = n12653 ^ n835 ;
  assign n12655 = ~n12650 & ~n12654 ;
  assign n12656 = n12655 ^ n12653 ;
  assign n12657 = n12363 & ~n12656 ;
  assign n12362 = n12361 ^ n534 ;
  assign n12658 = n12657 ^ n12362 ;
  assign n12659 = n12353 ^ n138 ;
  assign n12660 = ~n12359 & n12659 ;
  assign n12661 = n12660 ^ n12003 ;
  assign n12662 = n12661 ^ n183 ;
  assign n12717 = n12347 & ~n12359 ;
  assign n12718 = n12717 ^ n12350 ;
  assign n12663 = n12009 ^ n188 ;
  assign n12664 = n12663 ^ n246 ;
  assign n12667 = ~n12341 & ~n12664 ;
  assign n12668 = n12667 ^ n246 ;
  assign n12669 = ~n12359 & n12668 ;
  assign n12670 = n12669 ^ n12006 ;
  assign n12671 = n12670 ^ n157 ;
  assign n12709 = ~n12341 & ~n12359 ;
  assign n12710 = n12709 ^ n12009 ;
  assign n12672 = n12018 ^ n401 ;
  assign n12673 = n12672 ^ n461 ;
  assign n12676 = ~n12324 & ~n12673 ;
  assign n12677 = n12676 ^ n461 ;
  assign n12678 = ~n12359 & ~n12677 ;
  assign n12679 = n12678 ^ n12015 ;
  assign n12680 = n12679 ^ n341 ;
  assign n12691 = ~n12324 & ~n12359 ;
  assign n12692 = n12691 ^ n12018 ;
  assign n12681 = ~n12319 & ~n12359 ;
  assign n12682 = n12681 ^ n12321 ;
  assign n12683 = n12682 ^ n457 ;
  assign n12684 = n12317 & ~n12359 ;
  assign n12685 = n12684 ^ n12024 ;
  assign n12686 = n12685 ^ n534 ;
  assign n12687 = ~n12658 & n12686 ;
  assign n12688 = n12687 ^ n750 ;
  assign n12689 = ~n12683 & n12688 ;
  assign n12690 = n12689 ^ n12682 ;
  assign n12693 = n12692 ^ n12690 ;
  assign n12694 = n12692 ^ n401 ;
  assign n12695 = ~n12693 & n12694 ;
  assign n12696 = n12695 ^ n462 ;
  assign n12697 = ~n12680 & n12696 ;
  assign n12698 = n12697 ^ n349 ;
  assign n12699 = n12330 & ~n12359 ;
  assign n12700 = n12699 ^ n12333 ;
  assign n12701 = n12700 ^ n291 ;
  assign n12702 = ~n12698 & n12701 ;
  assign n12703 = n12702 ^ n307 ;
  assign n12704 = ~n12336 & ~n12359 ;
  assign n12705 = n12704 ^ n12338 ;
  assign n12706 = n12705 ^ n245 ;
  assign n12707 = n12703 & ~n12706 ;
  assign n12708 = n12707 ^ n12705 ;
  assign n12711 = n12710 ^ n12708 ;
  assign n12712 = n12710 ^ n188 ;
  assign n12713 = ~n12711 & ~n12712 ;
  assign n12714 = n12713 ^ n203 ;
  assign n12715 = n12671 & n12714 ;
  assign n12716 = n12715 ^ n157 ;
  assign n12719 = n12718 ^ n12716 ;
  assign n12720 = n12718 ^ n138 ;
  assign n12721 = ~n12719 & n12720 ;
  assign n12722 = n12721 ^ n4971 ;
  assign n12723 = ~n12662 & ~n12722 ;
  assign n12724 = n12723 ^ n183 ;
  assign n12725 = n12356 ^ n11962 ;
  assign n12726 = n12725 ^ n183 ;
  assign n12727 = n12724 & ~n12726 ;
  assign n12729 = ~n11962 & n12001 ;
  assign n12730 = n12727 & n12729 ;
  assign n12728 = n12727 ^ n12724 ;
  assign n12731 = n12730 ^ n12728 ;
  assign n12732 = ~n12658 & ~n12731 ;
  assign n12733 = n12732 ^ n12685 ;
  assign n12734 = n12733 ^ n457 ;
  assign n12735 = n12650 & ~n12731 ;
  assign n12736 = n12735 ^ n12652 ;
  assign n12737 = n12736 ^ n609 ;
  assign n12738 = n12641 & ~n12731 ;
  assign n12739 = n12738 ^ n12365 ;
  assign n12740 = n12739 ^ n786 ;
  assign n12979 = ~n12608 & ~n12731 ;
  assign n12980 = n12979 ^ n12610 ;
  assign n12983 = n12980 ^ n1427 ;
  assign n12741 = n12606 & ~n12731 ;
  assign n12742 = n12741 ^ n12371 ;
  assign n12743 = n12742 ^ n1739 ;
  assign n12746 = n12599 & ~n12731 ;
  assign n12747 = n12746 ^ n12375 ;
  assign n12748 = n12747 ^ n2175 ;
  assign n12749 = ~n12591 & ~n12731 ;
  assign n12750 = n12749 ^ n12378 ;
  assign n12751 = n12750 ^ n2511 ;
  assign n12752 = ~n12589 & ~n12731 ;
  assign n12753 = n12752 ^ n12382 ;
  assign n12754 = n12753 ^ n2707 ;
  assign n12755 = ~n12583 & ~n12731 ;
  assign n12756 = n12755 ^ n12585 ;
  assign n12757 = n12756 ^ n2894 ;
  assign n12951 = n12580 ^ n3320 ;
  assign n12952 = ~n12731 & n12951 ;
  assign n12953 = n12952 ^ n12385 ;
  assign n12956 = n12953 ^ n2894 ;
  assign n12758 = n12565 ^ n3908 ;
  assign n12759 = ~n12731 & n12758 ;
  assign n12760 = n12759 ^ n12567 ;
  assign n12761 = n12760 ^ n3722 ;
  assign n12762 = n12560 & ~n12731 ;
  assign n12763 = n12762 ^ n12562 ;
  assign n12764 = n12763 ^ n3908 ;
  assign n12767 = n12553 & ~n12731 ;
  assign n12768 = n12767 ^ n12555 ;
  assign n12769 = n12768 ^ n4356 ;
  assign n12922 = n12550 ^ n4812 ;
  assign n12923 = ~n12731 & n12922 ;
  assign n12924 = n12923 ^ n12401 ;
  assign n12770 = n12548 & ~n12731 ;
  assign n12771 = n12770 ^ n12404 ;
  assign n12772 = n12771 ^ n4812 ;
  assign n12773 = n12544 ^ n5317 ;
  assign n12774 = ~n12731 & n12773 ;
  assign n12775 = n12774 ^ n12408 ;
  assign n12776 = n12775 ^ n5073 ;
  assign n12777 = n12542 & ~n12731 ;
  assign n12778 = n12777 ^ n12410 ;
  assign n12780 = n12778 ^ n5317 ;
  assign n12909 = n12540 & ~n12731 ;
  assign n12910 = n12909 ^ n12421 ;
  assign n12781 = ~n12535 & ~n12731 ;
  assign n12782 = n12781 ^ n12537 ;
  assign n12783 = n12782 ^ n5830 ;
  assign n12784 = ~n12533 & ~n12731 ;
  assign n12785 = n12784 ^ n12424 ;
  assign n12786 = n12785 ^ n6115 ;
  assign n12790 = n12522 & ~n12731 ;
  assign n12791 = n12790 ^ n12524 ;
  assign n12792 = n12791 ^ n6673 ;
  assign n12793 = ~n12520 & ~n12731 ;
  assign n12794 = n12793 ^ n12427 ;
  assign n12795 = n12794 ^ n6959 ;
  assign n12800 = ~n12507 & ~n12731 ;
  assign n12801 = n12800 ^ n12510 ;
  assign n12802 = n12801 ^ n7584 ;
  assign n12803 = ~n12492 & ~n12731 ;
  assign n12804 = n12803 ^ n12494 ;
  assign n12805 = n12804 ^ n8586 ;
  assign n12806 = n12490 & ~n12731 ;
  assign n12807 = n12806 ^ n12431 ;
  assign n12808 = n12807 ^ n8910 ;
  assign n12809 = ~n12482 & ~n12731 ;
  assign n12810 = n12809 ^ n12434 ;
  assign n12811 = n12810 ^ n9542 ;
  assign n12812 = ~n12476 & ~n12731 ;
  assign n12813 = n12812 ^ n12479 ;
  assign n12815 = n12813 ^ n10108 ;
  assign n12816 = n12468 ^ n11233 ;
  assign n12817 = ~n12731 & n12816 ;
  assign n12818 = n12817 ^ n12446 ;
  assign n12819 = n12818 ^ n10875 ;
  assign n12853 = n12466 & ~n12731 ;
  assign n12854 = n12853 ^ n12450 ;
  assign n12820 = n12454 ^ n12359 ;
  assign n12821 = ~n12731 & ~n12820 ;
  assign n12822 = n12821 ^ n12359 ;
  assign n12846 = x12 & ~n12822 ;
  assign n12845 = n12456 & ~n12731 ;
  assign n12847 = n12846 ^ n12845 ;
  assign n12848 = n12847 ^ n12453 ;
  assign n12823 = n12822 ^ x12 ;
  assign n12824 = n12823 ^ n11960 ;
  assign n12832 = n11960 ^ x11 ;
  assign n12826 = ~x8 & ~x9 ;
  assign n12825 = n12359 ^ x10 ;
  assign n12827 = n12826 ^ n12825 ;
  assign n12828 = n12731 ^ n12359 ;
  assign n12829 = n12828 ^ x11 ;
  assign n12830 = ~n12827 & ~n12829 ;
  assign n12831 = n12830 ^ n12452 ;
  assign n12833 = n12832 ^ n12831 ;
  assign n12834 = n12833 ^ x11 ;
  assign n12835 = n12834 ^ n12731 ;
  assign n12836 = n12835 ^ n12833 ;
  assign n12837 = n12833 ^ n12828 ;
  assign n12838 = n12837 ^ n12833 ;
  assign n12839 = n12836 & ~n12838 ;
  assign n12840 = n12839 ^ n12833 ;
  assign n12841 = x10 & n12840 ;
  assign n12842 = n12841 ^ n12831 ;
  assign n12843 = n12824 & n12842 ;
  assign n12844 = n12843 ^ n12823 ;
  assign n12849 = n12848 ^ n12844 ;
  assign n12850 = n12848 ^ n11594 ;
  assign n12851 = ~n12849 & n12850 ;
  assign n12852 = n12851 ^ n11594 ;
  assign n12855 = n12854 ^ n12852 ;
  assign n12856 = n12854 ^ n11233 ;
  assign n12857 = n12855 & ~n12856 ;
  assign n12858 = n12857 ^ n11326 ;
  assign n12859 = n12819 & ~n12858 ;
  assign n12860 = n12859 ^ n11327 ;
  assign n12861 = ~n12471 & ~n12731 ;
  assign n12862 = n12861 ^ n12473 ;
  assign n12863 = n12862 ^ n10468 ;
  assign n12864 = ~n12860 & ~n12863 ;
  assign n12865 = n12864 ^ n10639 ;
  assign n12866 = n12815 & n12865 ;
  assign n12814 = n12813 ^ n9542 ;
  assign n12867 = n12866 ^ n12814 ;
  assign n12868 = ~n12811 & ~n12867 ;
  assign n12869 = n12868 ^ n9628 ;
  assign n12870 = ~n12485 & ~n12731 ;
  assign n12871 = n12870 ^ n12487 ;
  assign n12872 = n12871 ^ n9217 ;
  assign n12873 = n12869 & n12872 ;
  assign n12874 = n12873 ^ n9285 ;
  assign n12875 = ~n12808 & ~n12874 ;
  assign n12876 = n12875 ^ n9005 ;
  assign n12877 = ~n12805 & n12876 ;
  assign n12878 = n12877 ^ n8688 ;
  assign n12879 = n12497 & ~n12731 ;
  assign n12880 = n12879 ^ n12499 ;
  assign n12881 = n12880 ^ n8253 ;
  assign n12882 = n12878 & n12881 ;
  assign n12883 = n12882 ^ n8356 ;
  assign n12884 = n12502 & ~n12731 ;
  assign n12885 = n12884 ^ n12504 ;
  assign n12886 = n12885 ^ n7891 ;
  assign n12887 = ~n12883 & n12886 ;
  assign n12888 = n12887 ^ n7971 ;
  assign n12889 = n12802 & n12888 ;
  assign n12890 = n12889 ^ n12801 ;
  assign n12797 = ~n12513 & ~n12731 ;
  assign n12798 = n12797 ^ n12516 ;
  assign n12796 = n12794 ^ n7277 ;
  assign n12799 = n12798 ^ n12796 ;
  assign n12891 = n12890 ^ n12799 ;
  assign n12892 = n12891 ^ n12796 ;
  assign n12893 = n12798 ^ n12794 ;
  assign n12894 = n12893 ^ n12796 ;
  assign n12895 = n12892 & ~n12894 ;
  assign n12896 = n12895 ^ n12796 ;
  assign n12897 = n12795 & ~n12896 ;
  assign n12898 = n12897 ^ n7011 ;
  assign n12899 = n12792 & n12898 ;
  assign n12900 = n12899 ^ n6673 ;
  assign n12787 = n12527 ^ n6673 ;
  assign n12788 = ~n12731 & n12787 ;
  assign n12789 = n12788 ^ n12529 ;
  assign n12901 = n12900 ^ n12789 ;
  assign n12902 = n12900 ^ n6389 ;
  assign n12903 = ~n12901 & ~n12902 ;
  assign n12904 = n12903 ^ n6423 ;
  assign n12905 = n12786 & ~n12904 ;
  assign n12906 = n12905 ^ n6429 ;
  assign n12907 = n12783 & ~n12906 ;
  assign n12908 = n12907 ^ n12782 ;
  assign n12911 = n12910 ^ n12908 ;
  assign n12912 = n12910 ^ n5562 ;
  assign n12913 = n12911 & ~n12912 ;
  assign n12914 = n12913 ^ n5885 ;
  assign n12915 = ~n12780 & ~n12914 ;
  assign n12779 = n12778 ^ n5073 ;
  assign n12916 = n12915 ^ n12779 ;
  assign n12917 = ~n12776 & ~n12916 ;
  assign n12918 = n12917 ^ n5073 ;
  assign n12919 = n12918 ^ n12771 ;
  assign n12920 = ~n12772 & n12919 ;
  assign n12921 = n12920 ^ n4812 ;
  assign n12925 = n12924 ^ n12921 ;
  assign n12926 = n12924 ^ n4583 ;
  assign n12927 = ~n12925 & n12926 ;
  assign n12928 = n12927 ^ n4645 ;
  assign n12929 = n12769 & ~n12928 ;
  assign n12930 = n12929 ^ n12768 ;
  assign n12765 = n12558 & ~n12731 ;
  assign n12766 = n12765 ^ n12398 ;
  assign n12931 = n12930 ^ n12766 ;
  assign n12932 = n12930 ^ n4153 ;
  assign n12933 = n12931 & n12932 ;
  assign n12934 = n12933 ^ n4153 ;
  assign n12935 = n12934 ^ n12763 ;
  assign n12936 = ~n12764 & n12935 ;
  assign n12937 = n12936 ^ n3961 ;
  assign n12938 = ~n12761 & ~n12937 ;
  assign n12939 = n12938 ^ n3795 ;
  assign n12940 = n12571 ^ n3722 ;
  assign n12941 = ~n12731 & ~n12940 ;
  assign n12942 = n12941 ^ n12574 ;
  assign n12943 = n12942 ^ n3538 ;
  assign n12944 = n12939 & n12943 ;
  assign n12945 = n12944 ^ n3596 ;
  assign n12946 = n12578 & ~n12731 ;
  assign n12947 = n12946 ^ n12388 ;
  assign n12948 = n12947 ^ n3320 ;
  assign n12949 = n12945 & ~n12948 ;
  assign n12950 = n12949 ^ n3387 ;
  assign n12954 = n12953 ^ n3093 ;
  assign n12955 = n12950 & ~n12954 ;
  assign n12957 = n12956 ^ n12955 ;
  assign n12958 = ~n12757 & ~n12957 ;
  assign n12959 = n12958 ^ n3396 ;
  assign n12960 = n12754 & ~n12959 ;
  assign n12961 = n12960 ^ n2707 ;
  assign n12962 = n12961 ^ n12750 ;
  assign n12963 = n12751 & n12962 ;
  assign n12964 = n12963 ^ n2530 ;
  assign n12965 = n12593 ^ n2511 ;
  assign n12966 = ~n12731 & ~n12965 ;
  assign n12967 = n12966 ^ n12595 ;
  assign n12968 = n12967 ^ n2366 ;
  assign n12969 = n12964 & n12968 ;
  assign n12970 = n12969 ^ n2399 ;
  assign n12971 = n12748 & n12970 ;
  assign n12972 = n12971 ^ n2175 ;
  assign n12744 = n12601 & ~n12731 ;
  assign n12745 = n12744 ^ n12603 ;
  assign n12973 = n12972 ^ n12745 ;
  assign n12974 = n12972 ^ n2008 ;
  assign n12975 = n12973 & n12974 ;
  assign n12976 = n12975 ^ n2064 ;
  assign n12977 = ~n12743 & ~n12976 ;
  assign n12978 = n12977 ^ n1763 ;
  assign n12981 = n12980 ^ n1572 ;
  assign n12982 = n12978 & ~n12981 ;
  assign n12984 = n12983 ^ n12982 ;
  assign n12985 = ~n12613 & ~n12731 ;
  assign n12986 = n12985 ^ n12615 ;
  assign n12987 = n12986 ^ n1427 ;
  assign n12988 = n12984 & ~n12987 ;
  assign n12989 = n12988 ^ n1450 ;
  assign n12990 = ~n12619 & ~n12731 ;
  assign n12991 = n12990 ^ n12368 ;
  assign n12992 = n12991 ^ n1290 ;
  assign n12993 = ~n12989 & ~n12992 ;
  assign n12994 = n12993 ^ n1461 ;
  assign n12995 = ~n12621 & ~n12731 ;
  assign n12996 = n12995 ^ n12624 ;
  assign n12997 = n12996 ^ n1136 ;
  assign n12998 = n12994 & n12997 ;
  assign n12999 = n12998 ^ n1143 ;
  assign n13000 = n12627 ^ n1136 ;
  assign n13001 = ~n12731 & n13000 ;
  assign n13002 = n13001 ^ n12629 ;
  assign n13005 = n13002 ^ n1034 ;
  assign n13006 = ~n12999 & n13005 ;
  assign n13003 = n13002 ^ n892 ;
  assign n13007 = n13006 ^ n13003 ;
  assign n13008 = n12633 & ~n12731 ;
  assign n13009 = n13008 ^ n12636 ;
  assign n13010 = n13009 ^ n786 ;
  assign n13011 = n13010 ^ n927 ;
  assign n13012 = ~n13007 & n13011 ;
  assign n13013 = n13012 ^ n13010 ;
  assign n13014 = ~n12740 & n13013 ;
  assign n13015 = n13014 ^ n842 ;
  assign n13016 = n12643 & ~n12731 ;
  assign n13017 = n13016 ^ n12645 ;
  assign n13020 = n13017 ^ n696 ;
  assign n13021 = ~n13015 & n13020 ;
  assign n13018 = n13017 ^ n609 ;
  assign n13022 = n13021 ^ n13018 ;
  assign n13023 = n12737 & ~n13022 ;
  assign n13024 = n13023 ^ n834 ;
  assign n13025 = n12656 & ~n12731 ;
  assign n13026 = n13025 ^ n12361 ;
  assign n13027 = n13026 ^ n534 ;
  assign n13028 = ~n13024 & ~n13027 ;
  assign n13029 = n13028 ^ n750 ;
  assign n13030 = ~n12734 & n13029 ;
  assign n13031 = n13030 ^ n12733 ;
  assign n13032 = n13031 ^ n401 ;
  assign n13033 = ~n12722 & ~n12731 ;
  assign n13034 = n13033 ^ n12661 ;
  assign n13035 = n12716 ^ n138 ;
  assign n13036 = ~n12731 & n13035 ;
  assign n13037 = n13036 ^ n12718 ;
  assign n13038 = n13037 ^ n183 ;
  assign n13039 = n12714 & ~n12731 ;
  assign n13040 = n13039 ^ n12670 ;
  assign n13041 = n13040 ^ n138 ;
  assign n13069 = n12708 ^ n188 ;
  assign n13070 = ~n12731 & ~n13069 ;
  assign n13071 = n13070 ^ n12710 ;
  assign n13042 = n12690 ^ n401 ;
  assign n13043 = ~n12731 & n13042 ;
  assign n13044 = n13043 ^ n12692 ;
  assign n13045 = n13044 ^ n341 ;
  assign n13046 = ~n12688 & ~n12731 ;
  assign n13047 = n13046 ^ n12682 ;
  assign n13048 = n13047 ^ n13031 ;
  assign n13049 = n13032 & ~n13048 ;
  assign n13050 = n13049 ^ n462 ;
  assign n13051 = n13045 & n13050 ;
  assign n13052 = n13051 ^ n349 ;
  assign n13053 = n12696 & ~n12731 ;
  assign n13054 = n13053 ^ n12679 ;
  assign n13055 = n13054 ^ n291 ;
  assign n13056 = ~n13052 & n13055 ;
  assign n13057 = n13056 ^ n307 ;
  assign n13058 = ~n12698 & ~n12731 ;
  assign n13059 = n13058 ^ n12700 ;
  assign n13060 = n13059 ^ n245 ;
  assign n13061 = n13057 & ~n13060 ;
  assign n13062 = n13061 ^ n13059 ;
  assign n13063 = n13062 ^ n188 ;
  assign n13064 = ~n12703 & ~n12731 ;
  assign n13065 = n13064 ^ n12705 ;
  assign n13066 = n13065 ^ n13062 ;
  assign n13067 = ~n13063 & ~n13066 ;
  assign n13068 = n13067 ^ n188 ;
  assign n13072 = n13071 ^ n13068 ;
  assign n13073 = n13068 ^ n157 ;
  assign n13074 = ~n13072 & ~n13073 ;
  assign n13075 = n13074 ^ n13071 ;
  assign n13076 = n13075 ^ n13040 ;
  assign n13077 = n13041 & n13076 ;
  assign n13078 = n13077 ^ n138 ;
  assign n13079 = n13078 ^ n183 ;
  assign n13080 = ~n13038 & ~n13079 ;
  assign n13081 = n13080 ^ n183 ;
  assign n13082 = ~n13034 & n13081 ;
  assign n13083 = n13032 & ~n13082 ;
  assign n13084 = n13083 ^ n13047 ;
  assign n13085 = n13084 ^ n341 ;
  assign n13394 = ~n13029 & ~n13082 ;
  assign n13395 = n13394 ^ n12733 ;
  assign n13086 = ~n13024 & ~n13082 ;
  assign n13087 = n13086 ^ n13026 ;
  assign n13088 = n13087 ^ n457 ;
  assign n13089 = ~n13022 & ~n13082 ;
  assign n13090 = n13089 ^ n12736 ;
  assign n13091 = n13090 ^ n534 ;
  assign n13092 = n13013 & ~n13082 ;
  assign n13093 = n13092 ^ n12739 ;
  assign n13094 = n13093 ^ n696 ;
  assign n13097 = ~n12976 & ~n13082 ;
  assign n13098 = n13097 ^ n12742 ;
  assign n13348 = n13098 ^ n1427 ;
  assign n13099 = n13098 ^ n1572 ;
  assign n13104 = n12964 & ~n13082 ;
  assign n13105 = n13104 ^ n12967 ;
  assign n13106 = n13105 ^ n2175 ;
  assign n13107 = n12961 ^ n2511 ;
  assign n13108 = ~n13082 & ~n13107 ;
  assign n13109 = n13108 ^ n12750 ;
  assign n13110 = n13109 ^ n2366 ;
  assign n13329 = ~n12959 & ~n13082 ;
  assign n13330 = n13329 ^ n12753 ;
  assign n13111 = ~n12957 & ~n13082 ;
  assign n13112 = n13111 ^ n12756 ;
  assign n13113 = n13112 ^ n2707 ;
  assign n13114 = ~n12950 & ~n13082 ;
  assign n13115 = n13114 ^ n12953 ;
  assign n13116 = n13115 ^ n2894 ;
  assign n13319 = n12945 & ~n13082 ;
  assign n13320 = n13319 ^ n12947 ;
  assign n13323 = n13320 ^ n2894 ;
  assign n13117 = ~n12937 & ~n13082 ;
  assign n13118 = n13117 ^ n12760 ;
  assign n13119 = n13118 ^ n3538 ;
  assign n13304 = n12934 ^ n3908 ;
  assign n13305 = ~n13082 & n13304 ;
  assign n13306 = n13305 ^ n12763 ;
  assign n13298 = n12932 & ~n13082 ;
  assign n13299 = n13298 ^ n12766 ;
  assign n13292 = n12928 & ~n13082 ;
  assign n13293 = n13292 ^ n12768 ;
  assign n13120 = n12921 ^ n4583 ;
  assign n13121 = ~n13082 & n13120 ;
  assign n13122 = n13121 ^ n12924 ;
  assign n13123 = n13122 ^ n4356 ;
  assign n13124 = n12918 ^ n4812 ;
  assign n13125 = ~n13082 & n13124 ;
  assign n13126 = n13125 ^ n12771 ;
  assign n13127 = n13126 ^ n4583 ;
  assign n13128 = ~n12916 & ~n13082 ;
  assign n13129 = n13128 ^ n12775 ;
  assign n13130 = n13129 ^ n4812 ;
  assign n13131 = n12914 & ~n13082 ;
  assign n13132 = n13131 ^ n12778 ;
  assign n13133 = n13132 ^ n5073 ;
  assign n13134 = n12908 ^ n5562 ;
  assign n13135 = ~n13082 & n13134 ;
  assign n13136 = n13135 ^ n12910 ;
  assign n13137 = n13136 ^ n5317 ;
  assign n13138 = n12906 & ~n13082 ;
  assign n13139 = n13138 ^ n12782 ;
  assign n13140 = n13139 ^ n5562 ;
  assign n13141 = ~n12904 & ~n13082 ;
  assign n13142 = n13141 ^ n12785 ;
  assign n13143 = n13142 ^ n13139 ;
  assign n13144 = n13143 ^ n13142 ;
  assign n13145 = n13144 ^ n5830 ;
  assign n13146 = n13145 ^ n13143 ;
  assign n13149 = n12898 & ~n13082 ;
  assign n13150 = n13149 ^ n12791 ;
  assign n13151 = n13150 ^ n6389 ;
  assign n13152 = n12890 ^ n7277 ;
  assign n13153 = ~n13082 & n13152 ;
  assign n13154 = n13153 ^ n12798 ;
  assign n13155 = n13154 ^ n6959 ;
  assign n13248 = ~n12888 & ~n13082 ;
  assign n13249 = n13248 ^ n12801 ;
  assign n13156 = ~n12883 & ~n13082 ;
  assign n13157 = n13156 ^ n12885 ;
  assign n13158 = n13157 ^ n7584 ;
  assign n13159 = n12876 & ~n13082 ;
  assign n13160 = n13159 ^ n12804 ;
  assign n13161 = n13160 ^ n8253 ;
  assign n13162 = ~n12874 & ~n13082 ;
  assign n13163 = n13162 ^ n12807 ;
  assign n13164 = n13163 ^ n8586 ;
  assign n13165 = n12869 & ~n13082 ;
  assign n13166 = n13165 ^ n12871 ;
  assign n13167 = n13166 ^ n8910 ;
  assign n13168 = ~n12865 & ~n13082 ;
  assign n13169 = n13168 ^ n12813 ;
  assign n13170 = n13169 ^ n9542 ;
  assign n13171 = ~n12860 & ~n13082 ;
  assign n13172 = n13171 ^ n12862 ;
  assign n13173 = n13172 ^ n10108 ;
  assign n13174 = ~n12858 & ~n13082 ;
  assign n13175 = n13174 ^ n12818 ;
  assign n13176 = n13175 ^ n10468 ;
  assign n13215 = n12852 ^ n11233 ;
  assign n13216 = ~n13082 & n13215 ;
  assign n13217 = n13216 ^ n12854 ;
  assign n13177 = n12844 ^ n11594 ;
  assign n13178 = ~n13082 & n13177 ;
  assign n13179 = n13178 ^ n12848 ;
  assign n13180 = n13179 ^ n11233 ;
  assign n13181 = ~n12842 & ~n13082 ;
  assign n13182 = n13181 ^ n12823 ;
  assign n13183 = n13182 ^ n11594 ;
  assign n13184 = n12826 ^ n12731 ;
  assign n13185 = ~n13082 & ~n13184 ;
  assign n13186 = n13185 ^ n12731 ;
  assign n13204 = x10 & ~n13186 ;
  assign n13202 = n12731 ^ x11 ;
  assign n13200 = n12826 ^ n12359 ;
  assign n13201 = ~n13082 & ~n13200 ;
  assign n13203 = n13202 ^ n13201 ;
  assign n13205 = n13204 ^ n13203 ;
  assign n13208 = n13205 ^ n11594 ;
  assign n13187 = n13186 ^ x10 ;
  assign n13188 = n13187 ^ n12359 ;
  assign n13190 = ~x6 & ~x7 ;
  assign n13191 = ~x8 & n13190 ;
  assign n13189 = n13082 ^ x9 ;
  assign n13192 = n13191 ^ n13189 ;
  assign n13193 = ~x8 & ~n13082 ;
  assign n13194 = n13193 ^ x9 ;
  assign n13195 = n13194 ^ n12731 ;
  assign n13196 = ~n13192 & n13195 ;
  assign n13197 = n13196 ^ n12828 ;
  assign n13198 = ~n13188 & n13197 ;
  assign n13199 = n13198 ^ n12452 ;
  assign n13206 = n13205 ^ n11960 ;
  assign n13207 = n13199 & n13206 ;
  assign n13209 = n13208 ^ n13207 ;
  assign n13210 = n13183 & n13209 ;
  assign n13211 = n13210 ^ n11594 ;
  assign n13212 = n13211 ^ n13179 ;
  assign n13213 = n13180 & ~n13212 ;
  assign n13214 = n13213 ^ n11233 ;
  assign n13218 = n13217 ^ n13214 ;
  assign n13219 = n13217 ^ n10875 ;
  assign n13220 = n13218 & n13219 ;
  assign n13221 = n13220 ^ n11327 ;
  assign n13222 = ~n13176 & ~n13221 ;
  assign n13223 = n13222 ^ n10639 ;
  assign n13224 = n13173 & n13223 ;
  assign n13225 = n13224 ^ n13172 ;
  assign n13226 = n13225 ^ n13169 ;
  assign n13227 = ~n13170 & ~n13226 ;
  assign n13228 = n13227 ^ n9628 ;
  assign n13229 = ~n12867 & ~n13082 ;
  assign n13230 = n13229 ^ n12810 ;
  assign n13231 = n13230 ^ n9217 ;
  assign n13232 = n13228 & ~n13231 ;
  assign n13233 = n13232 ^ n9285 ;
  assign n13234 = ~n13167 & n13233 ;
  assign n13235 = n13234 ^ n13166 ;
  assign n13236 = n13235 ^ n13163 ;
  assign n13237 = ~n13164 & ~n13236 ;
  assign n13238 = n13237 ^ n8688 ;
  assign n13239 = ~n13161 & n13238 ;
  assign n13240 = n13239 ^ n8356 ;
  assign n13241 = n12878 & ~n13082 ;
  assign n13242 = n13241 ^ n12880 ;
  assign n13243 = n13242 ^ n7891 ;
  assign n13244 = ~n13240 & ~n13243 ;
  assign n13245 = n13244 ^ n7971 ;
  assign n13246 = ~n13158 & n13245 ;
  assign n13247 = n13246 ^ n13157 ;
  assign n13250 = n13249 ^ n13247 ;
  assign n13251 = n13249 ^ n7277 ;
  assign n13252 = n13250 & n13251 ;
  assign n13253 = n13252 ^ n7277 ;
  assign n13254 = n13253 ^ n13154 ;
  assign n13255 = ~n13155 & n13254 ;
  assign n13256 = n13255 ^ n6959 ;
  assign n13257 = n13256 ^ n6673 ;
  assign n13258 = n12890 ^ n6959 ;
  assign n13259 = n13258 ^ n7339 ;
  assign n13260 = n12798 ^ n6959 ;
  assign n13261 = n13260 ^ n7339 ;
  assign n13262 = n13259 & ~n13261 ;
  assign n13263 = n13262 ^ n7339 ;
  assign n13264 = ~n13082 & n13263 ;
  assign n13265 = n13264 ^ n12794 ;
  assign n13266 = n13265 ^ n13256 ;
  assign n13267 = n13257 & ~n13266 ;
  assign n13268 = n13267 ^ n6713 ;
  assign n13269 = ~n13151 & ~n13268 ;
  assign n13270 = n13269 ^ n6389 ;
  assign n13147 = ~n12902 & ~n13082 ;
  assign n13148 = n13147 ^ n12789 ;
  assign n13271 = n13270 ^ n13148 ;
  assign n13272 = n13270 ^ n6115 ;
  assign n13273 = n13271 & ~n13272 ;
  assign n13274 = n13273 ^ n6429 ;
  assign n13277 = n13146 & ~n13274 ;
  assign n13278 = n13277 ^ n13143 ;
  assign n13279 = n13140 & ~n13278 ;
  assign n13280 = n13279 ^ n5885 ;
  assign n13281 = ~n13137 & n13280 ;
  assign n13282 = n13281 ^ n5360 ;
  assign n13283 = ~n13133 & n13282 ;
  assign n13284 = n13283 ^ n5073 ;
  assign n13285 = n13284 ^ n13129 ;
  assign n13286 = ~n13130 & n13285 ;
  assign n13287 = n13286 ^ n4854 ;
  assign n13288 = ~n13127 & n13287 ;
  assign n13289 = n13288 ^ n4645 ;
  assign n13290 = n13123 & ~n13289 ;
  assign n13291 = n13290 ^ n13122 ;
  assign n13294 = n13293 ^ n13291 ;
  assign n13295 = n13293 ^ n4153 ;
  assign n13296 = ~n13294 & n13295 ;
  assign n13297 = n13296 ^ n4153 ;
  assign n13300 = n13299 ^ n13297 ;
  assign n13301 = n13299 ^ n3908 ;
  assign n13302 = n13300 & ~n13301 ;
  assign n13303 = n13302 ^ n3908 ;
  assign n13307 = n13306 ^ n13303 ;
  assign n13308 = n13306 ^ n3722 ;
  assign n13309 = n13307 & n13308 ;
  assign n13310 = n13309 ^ n3795 ;
  assign n13311 = ~n13119 & n13310 ;
  assign n13312 = n13311 ^ n3538 ;
  assign n13313 = n13312 ^ n3320 ;
  assign n13314 = n12939 & ~n13082 ;
  assign n13315 = n13314 ^ n12942 ;
  assign n13316 = n13315 ^ n13312 ;
  assign n13317 = n13313 & ~n13316 ;
  assign n13318 = n13317 ^ n3387 ;
  assign n13321 = n13320 ^ n3093 ;
  assign n13322 = n13318 & n13321 ;
  assign n13324 = n13323 ^ n13322 ;
  assign n13325 = ~n13116 & n13324 ;
  assign n13326 = n13325 ^ n3396 ;
  assign n13327 = n13113 & ~n13326 ;
  assign n13328 = n13327 ^ n2707 ;
  assign n13331 = n13330 ^ n13328 ;
  assign n13332 = n13330 ^ n2511 ;
  assign n13333 = ~n13331 & ~n13332 ;
  assign n13334 = n13333 ^ n2530 ;
  assign n13335 = n13110 & n13334 ;
  assign n13336 = n13335 ^ n2399 ;
  assign n13337 = n13106 & n13336 ;
  assign n13338 = n13337 ^ n2175 ;
  assign n13102 = n12970 & ~n13082 ;
  assign n13103 = n13102 ^ n12747 ;
  assign n13339 = n13338 ^ n13103 ;
  assign n13340 = n13338 ^ n2008 ;
  assign n13341 = ~n13339 & n13340 ;
  assign n13342 = n13341 ^ n2008 ;
  assign n13100 = n12974 & ~n13082 ;
  assign n13101 = n13100 ^ n12745 ;
  assign n13343 = n13342 ^ n13101 ;
  assign n13344 = n13342 ^ n1739 ;
  assign n13345 = n13343 & ~n13344 ;
  assign n13346 = n13345 ^ n1763 ;
  assign n13347 = n13099 & n13346 ;
  assign n13349 = n13348 ^ n13347 ;
  assign n13350 = ~n12978 & ~n13082 ;
  assign n13351 = n13350 ^ n12980 ;
  assign n13352 = n13351 ^ n1427 ;
  assign n13353 = ~n13349 & n13352 ;
  assign n13354 = n13353 ^ n1450 ;
  assign n13355 = n12984 & ~n13082 ;
  assign n13356 = n13355 ^ n12986 ;
  assign n13357 = n13356 ^ n1290 ;
  assign n13358 = n13354 & n13357 ;
  assign n13359 = n13358 ^ n13356 ;
  assign n13095 = ~n12989 & ~n13082 ;
  assign n13096 = n13095 ^ n12991 ;
  assign n13360 = n13359 ^ n13096 ;
  assign n13361 = n13359 ^ n1136 ;
  assign n13362 = n13360 & n13361 ;
  assign n13363 = n13362 ^ n1143 ;
  assign n13364 = n12994 & ~n13082 ;
  assign n13365 = n13364 ^ n12996 ;
  assign n13368 = n13365 ^ n1034 ;
  assign n13369 = ~n13363 & n13368 ;
  assign n13366 = n13365 ^ n892 ;
  assign n13370 = n13369 ^ n13366 ;
  assign n13371 = n12999 & ~n13082 ;
  assign n13372 = n13371 ^ n13002 ;
  assign n13373 = n13372 ^ n786 ;
  assign n13374 = n13373 ^ n927 ;
  assign n13375 = ~n13370 & n13374 ;
  assign n13376 = n13375 ^ n13373 ;
  assign n13377 = n13007 & ~n13082 ;
  assign n13378 = n13377 ^ n13009 ;
  assign n13379 = n13378 ^ n696 ;
  assign n13380 = n13379 ^ n842 ;
  assign n13381 = ~n13376 & n13380 ;
  assign n13382 = n13381 ^ n13379 ;
  assign n13383 = ~n13094 & n13382 ;
  assign n13384 = n13383 ^ n835 ;
  assign n13385 = n13015 & ~n13082 ;
  assign n13386 = n13385 ^ n13017 ;
  assign n13387 = n13386 ^ n609 ;
  assign n13388 = ~n13384 & ~n13387 ;
  assign n13389 = n13388 ^ n834 ;
  assign n13390 = ~n13091 & ~n13389 ;
  assign n13391 = n13390 ^ n750 ;
  assign n13392 = n13088 & n13391 ;
  assign n13393 = n13392 ^ n13087 ;
  assign n13396 = n13395 ^ n13393 ;
  assign n13397 = n13395 ^ n401 ;
  assign n13398 = n13396 & n13397 ;
  assign n13399 = n13398 ^ n462 ;
  assign n13400 = n13085 & n13399 ;
  assign n13401 = n13400 ^ n349 ;
  assign n13402 = n13075 ^ n138 ;
  assign n13403 = ~n13082 & ~n13402 ;
  assign n13404 = n13403 ^ n13040 ;
  assign n13405 = n13404 ^ n183 ;
  assign n13406 = ~n13034 & ~n13037 ;
  assign n13408 = n13406 ^ n13037 ;
  assign n13407 = ~n13078 & ~n13406 ;
  assign n13409 = n13408 ^ n13407 ;
  assign n13410 = n13409 ^ n13406 ;
  assign n13411 = n13406 ^ n13404 ;
  assign n13412 = n13411 ^ n13406 ;
  assign n13413 = ~n13410 & n13412 ;
  assign n13414 = n13413 ^ n13406 ;
  assign n13415 = ~n183 & ~n13414 ;
  assign n13416 = n13415 ^ n13409 ;
  assign n13417 = n13073 & ~n13082 ;
  assign n13418 = n13417 ^ n13071 ;
  assign n13419 = n13418 ^ n138 ;
  assign n13422 = ~n13057 & ~n13082 ;
  assign n13423 = n13422 ^ n13059 ;
  assign n13424 = n13423 ^ n188 ;
  assign n13425 = ~n13052 & ~n13082 ;
  assign n13426 = n13425 ^ n13054 ;
  assign n13427 = n13426 ^ n245 ;
  assign n13428 = n13050 & ~n13082 ;
  assign n13429 = n13428 ^ n13044 ;
  assign n13430 = n13429 ^ n291 ;
  assign n13431 = ~n13401 & ~n13430 ;
  assign n13432 = n13431 ^ n307 ;
  assign n13433 = ~n13427 & n13432 ;
  assign n13434 = n13433 ^ n13426 ;
  assign n13435 = n13434 ^ n13423 ;
  assign n13436 = ~n13424 & ~n13435 ;
  assign n13437 = n13436 ^ n188 ;
  assign n13420 = ~n13063 & ~n13082 ;
  assign n13421 = n13420 ^ n13065 ;
  assign n13438 = n13437 ^ n13421 ;
  assign n13439 = n13421 ^ n157 ;
  assign n13440 = ~n13438 & n13439 ;
  assign n13441 = n13440 ^ n13437 ;
  assign n13442 = n13441 ^ n13418 ;
  assign n13443 = ~n13419 & n13442 ;
  assign n13444 = n13443 ^ n138 ;
  assign n13445 = n13416 & n13444 ;
  assign n13446 = ~n13405 & n13445 ;
  assign n13447 = n13446 ^ n13416 ;
  assign n13448 = ~n13401 & ~n13447 ;
  assign n13449 = n13448 ^ n13429 ;
  assign n13450 = n13449 ^ n245 ;
  assign n13451 = n13393 ^ n401 ;
  assign n13452 = ~n13447 & ~n13451 ;
  assign n13453 = n13452 ^ n13395 ;
  assign n13454 = n13453 ^ n341 ;
  assign n13775 = ~n13391 & ~n13447 ;
  assign n13776 = n13775 ^ n13087 ;
  assign n13455 = ~n13389 & ~n13447 ;
  assign n13456 = n13455 ^ n13090 ;
  assign n13457 = n13456 ^ n457 ;
  assign n13458 = ~n13384 & ~n13447 ;
  assign n13459 = n13458 ^ n13386 ;
  assign n13460 = n13459 ^ n534 ;
  assign n13461 = n13382 & ~n13447 ;
  assign n13462 = n13461 ^ n13093 ;
  assign n13463 = n13462 ^ n609 ;
  assign n13464 = n13361 & ~n13447 ;
  assign n13465 = n13464 ^ n13096 ;
  assign n13466 = n13465 ^ n1034 ;
  assign n13737 = ~n13349 & ~n13447 ;
  assign n13738 = n13737 ^ n13351 ;
  assign n13741 = n13738 ^ n1136 ;
  assign n13467 = n13336 & ~n13447 ;
  assign n13468 = n13467 ^ n13105 ;
  assign n13469 = n13468 ^ n2008 ;
  assign n13470 = n13334 & ~n13447 ;
  assign n13471 = n13470 ^ n13109 ;
  assign n13472 = n13471 ^ n2175 ;
  assign n13473 = n13328 ^ n2511 ;
  assign n13474 = ~n13447 & ~n13473 ;
  assign n13475 = n13474 ^ n13330 ;
  assign n13476 = n13475 ^ n2366 ;
  assign n13710 = ~n13326 & ~n13447 ;
  assign n13711 = n13710 ^ n13112 ;
  assign n13477 = n13324 & ~n13447 ;
  assign n13478 = n13477 ^ n13115 ;
  assign n13479 = n13478 ^ n2707 ;
  assign n13480 = ~n13318 & ~n13447 ;
  assign n13481 = n13480 ^ n13320 ;
  assign n13482 = n13481 ^ n2894 ;
  assign n13698 = n13313 & ~n13447 ;
  assign n13699 = n13698 ^ n13315 ;
  assign n13703 = n13699 ^ n2894 ;
  assign n13483 = n13310 & ~n13447 ;
  assign n13484 = n13483 ^ n13118 ;
  assign n13485 = n13484 ^ n3320 ;
  assign n13689 = n13303 ^ n3722 ;
  assign n13690 = ~n13447 & ~n13689 ;
  assign n13691 = n13690 ^ n13306 ;
  assign n13682 = n13297 ^ n3908 ;
  assign n13683 = ~n13447 & n13682 ;
  assign n13684 = n13683 ^ n13299 ;
  assign n13675 = n13291 ^ n4153 ;
  assign n13676 = ~n13447 & n13675 ;
  assign n13677 = n13676 ^ n13293 ;
  assign n13486 = n13287 & ~n13447 ;
  assign n13487 = n13486 ^ n13126 ;
  assign n13488 = n13487 ^ n4356 ;
  assign n13661 = n13284 ^ n4812 ;
  assign n13662 = ~n13447 & n13661 ;
  assign n13663 = n13662 ^ n13129 ;
  assign n13489 = n13282 & ~n13447 ;
  assign n13490 = n13489 ^ n13132 ;
  assign n13491 = n13490 ^ n4812 ;
  assign n13652 = n13280 & ~n13447 ;
  assign n13653 = n13652 ^ n13136 ;
  assign n13492 = n13142 ^ n5562 ;
  assign n13493 = n13492 ^ n5900 ;
  assign n13496 = n13274 & n13493 ;
  assign n13497 = n13496 ^ n5900 ;
  assign n13498 = ~n13447 & n13497 ;
  assign n13499 = n13498 ^ n13139 ;
  assign n13500 = n13499 ^ n5317 ;
  assign n13501 = n13274 & ~n13447 ;
  assign n13502 = n13501 ^ n13142 ;
  assign n13503 = n13502 ^ n5562 ;
  assign n13504 = ~n13272 & ~n13447 ;
  assign n13505 = n13504 ^ n13148 ;
  assign n13507 = n13505 ^ n5830 ;
  assign n13508 = n13257 & ~n13447 ;
  assign n13509 = n13508 ^ n13265 ;
  assign n13510 = n13509 ^ n6389 ;
  assign n13632 = n13253 ^ n6959 ;
  assign n13633 = ~n13447 & n13632 ;
  assign n13634 = n13633 ^ n13154 ;
  assign n13511 = n13247 ^ n7277 ;
  assign n13512 = ~n13447 & ~n13511 ;
  assign n13513 = n13512 ^ n13249 ;
  assign n13514 = n13513 ^ n6959 ;
  assign n13515 = ~n13245 & ~n13447 ;
  assign n13516 = n13515 ^ n13157 ;
  assign n13517 = n13516 ^ n7277 ;
  assign n13518 = n13235 ^ n8586 ;
  assign n13519 = ~n13447 & ~n13518 ;
  assign n13520 = n13519 ^ n13163 ;
  assign n13521 = n13520 ^ n8253 ;
  assign n13522 = ~n13233 & ~n13447 ;
  assign n13523 = n13522 ^ n13166 ;
  assign n13524 = n13523 ^ n8586 ;
  assign n13525 = n13228 & ~n13447 ;
  assign n13526 = n13525 ^ n13230 ;
  assign n13527 = n13526 ^ n8910 ;
  assign n13604 = n13225 ^ n9542 ;
  assign n13605 = ~n13447 & ~n13604 ;
  assign n13606 = n13605 ^ n13169 ;
  assign n13528 = ~n13223 & ~n13447 ;
  assign n13529 = n13528 ^ n13172 ;
  assign n13530 = n13529 ^ n9542 ;
  assign n13531 = ~n13221 & ~n13447 ;
  assign n13532 = n13531 ^ n13175 ;
  assign n13600 = n13532 ^ n9542 ;
  assign n13533 = n13532 ^ n10108 ;
  assign n13537 = n13209 & ~n13447 ;
  assign n13538 = n13537 ^ n13182 ;
  assign n13539 = n13538 ^ n11233 ;
  assign n13540 = ~n13199 & ~n13447 ;
  assign n13541 = n13540 ^ n13205 ;
  assign n13542 = n13541 ^ n11594 ;
  assign n13578 = n13197 & ~n13447 ;
  assign n13579 = n13578 ^ n13187 ;
  assign n13582 = n13579 ^ n11594 ;
  assign n13544 = n13082 ^ n12731 ;
  assign n13543 = n13190 ^ n13082 ;
  assign n13545 = n13544 ^ n13543 ;
  assign n13546 = n13545 ^ n13544 ;
  assign n13547 = n13544 ^ x8 ;
  assign n13548 = n13547 ^ n13544 ;
  assign n13549 = ~n13546 & ~n13548 ;
  assign n13550 = n13549 ^ n13544 ;
  assign n13551 = ~n13447 & n13550 ;
  assign n13552 = n13551 ^ n13194 ;
  assign n13553 = n13552 ^ n12359 ;
  assign n13555 = n13447 & ~n13543 ;
  assign n13554 = n13190 ^ x8 ;
  assign n13556 = n13555 ^ n13554 ;
  assign n13557 = n13556 ^ n12731 ;
  assign n13560 = n13447 ^ x7 ;
  assign n13559 = ~x4 & ~x5 ;
  assign n13561 = n13560 ^ n13559 ;
  assign n13562 = n13559 ^ n13082 ;
  assign n13563 = ~n13561 & ~n13562 ;
  assign n13564 = n13563 ^ n13544 ;
  assign n13565 = n13564 ^ n13544 ;
  assign n13558 = n13447 ^ n13082 ;
  assign n13566 = n13565 ^ n13558 ;
  assign n13567 = n13566 ^ n13565 ;
  assign n13570 = ~n13560 & n13567 ;
  assign n13571 = n13570 ^ n13565 ;
  assign n13572 = x6 & n13571 ;
  assign n13573 = n13572 ^ n13564 ;
  assign n13574 = n13557 & n13573 ;
  assign n13575 = n13574 ^ n12828 ;
  assign n13576 = n13553 & n13575 ;
  assign n13577 = n13576 ^ n12452 ;
  assign n13580 = n13579 ^ n11960 ;
  assign n13581 = n13577 & n13580 ;
  assign n13583 = n13582 ^ n13581 ;
  assign n13584 = n13542 & n13583 ;
  assign n13585 = n13584 ^ n11688 ;
  assign n13586 = n13539 & n13585 ;
  assign n13587 = n13586 ^ n11233 ;
  assign n13588 = n13587 ^ n10875 ;
  assign n13589 = n13211 ^ n11233 ;
  assign n13590 = ~n13447 & n13589 ;
  assign n13591 = n13590 ^ n13179 ;
  assign n13592 = n13591 ^ n13587 ;
  assign n13593 = ~n13588 & ~n13592 ;
  assign n13594 = n13593 ^ n10875 ;
  assign n13534 = n13214 ^ n10875 ;
  assign n13535 = ~n13447 & ~n13534 ;
  assign n13536 = n13535 ^ n13217 ;
  assign n13595 = n13594 ^ n13536 ;
  assign n13596 = n13594 ^ n10468 ;
  assign n13597 = ~n13595 & ~n13596 ;
  assign n13598 = n13597 ^ n10639 ;
  assign n13599 = n13533 & n13598 ;
  assign n13601 = n13600 ^ n13599 ;
  assign n13602 = ~n13530 & ~n13601 ;
  assign n13603 = n13602 ^ n9542 ;
  assign n13607 = n13606 ^ n13603 ;
  assign n13608 = n13606 ^ n9217 ;
  assign n13609 = n13607 & ~n13608 ;
  assign n13610 = n13609 ^ n9285 ;
  assign n13611 = n13527 & ~n13610 ;
  assign n13612 = n13611 ^ n9005 ;
  assign n13613 = ~n13524 & n13612 ;
  assign n13614 = n13613 ^ n8586 ;
  assign n13615 = n13614 ^ n13520 ;
  assign n13616 = ~n13521 & n13615 ;
  assign n13617 = n13616 ^ n8356 ;
  assign n13618 = n13238 & ~n13447 ;
  assign n13619 = n13618 ^ n13160 ;
  assign n13620 = n13619 ^ n7891 ;
  assign n13621 = ~n13617 & n13620 ;
  assign n13622 = n13621 ^ n7971 ;
  assign n13623 = ~n13240 & ~n13447 ;
  assign n13624 = n13623 ^ n13242 ;
  assign n13625 = n13624 ^ n7584 ;
  assign n13626 = ~n13622 & n13625 ;
  assign n13627 = n13626 ^ n7660 ;
  assign n13628 = ~n13517 & n13627 ;
  assign n13629 = n13628 ^ n7339 ;
  assign n13630 = n13514 & n13629 ;
  assign n13631 = n13630 ^ n6959 ;
  assign n13635 = n13634 ^ n13631 ;
  assign n13636 = n13634 ^ n6673 ;
  assign n13637 = n13635 & ~n13636 ;
  assign n13638 = n13637 ^ n6713 ;
  assign n13639 = ~n13510 & ~n13638 ;
  assign n13640 = n13639 ^ n6423 ;
  assign n13641 = ~n13268 & ~n13447 ;
  assign n13642 = n13641 ^ n13150 ;
  assign n13643 = n13642 ^ n6115 ;
  assign n13644 = ~n13640 & n13643 ;
  assign n13645 = n13644 ^ n6429 ;
  assign n13646 = n13507 & ~n13645 ;
  assign n13506 = n13505 ^ n5562 ;
  assign n13647 = n13646 ^ n13506 ;
  assign n13648 = n13503 & n13647 ;
  assign n13649 = n13648 ^ n5885 ;
  assign n13650 = n13500 & n13649 ;
  assign n13651 = n13650 ^ n5317 ;
  assign n13654 = n13653 ^ n13651 ;
  assign n13655 = n13653 ^ n5073 ;
  assign n13656 = n13654 & ~n13655 ;
  assign n13657 = n13656 ^ n5073 ;
  assign n13658 = n13657 ^ n13490 ;
  assign n13659 = ~n13491 & n13658 ;
  assign n13660 = n13659 ^ n4812 ;
  assign n13664 = n13663 ^ n13660 ;
  assign n13665 = n13663 ^ n4583 ;
  assign n13666 = n13664 & ~n13665 ;
  assign n13667 = n13666 ^ n4645 ;
  assign n13668 = ~n13488 & n13667 ;
  assign n13669 = n13668 ^ n4414 ;
  assign n13670 = n13289 & ~n13447 ;
  assign n13671 = n13670 ^ n13122 ;
  assign n13672 = n13671 ^ n4153 ;
  assign n13673 = n13669 & n13672 ;
  assign n13674 = n13673 ^ n4153 ;
  assign n13678 = n13677 ^ n13674 ;
  assign n13679 = n13677 ^ n3908 ;
  assign n13680 = ~n13678 & n13679 ;
  assign n13681 = n13680 ^ n3908 ;
  assign n13685 = n13684 ^ n13681 ;
  assign n13686 = n13684 ^ n3722 ;
  assign n13687 = n13685 & n13686 ;
  assign n13688 = n13687 ^ n3722 ;
  assign n13692 = n13691 ^ n13688 ;
  assign n13693 = n13691 ^ n3538 ;
  assign n13694 = ~n13692 & n13693 ;
  assign n13695 = n13694 ^ n3596 ;
  assign n13696 = ~n13485 & n13695 ;
  assign n13697 = n13696 ^ n3320 ;
  assign n13700 = n13699 ^ n13697 ;
  assign n13701 = n13697 ^ n3093 ;
  assign n13702 = n13700 & n13701 ;
  assign n13704 = n13703 ^ n13702 ;
  assign n13705 = n13482 & ~n13704 ;
  assign n13706 = n13705 ^ n2894 ;
  assign n13707 = n13706 ^ n13478 ;
  assign n13708 = n13479 & n13707 ;
  assign n13709 = n13708 ^ n2707 ;
  assign n13712 = n13711 ^ n13709 ;
  assign n13713 = n13711 ^ n2511 ;
  assign n13714 = ~n13712 & ~n13713 ;
  assign n13715 = n13714 ^ n2530 ;
  assign n13716 = ~n13476 & n13715 ;
  assign n13717 = n13716 ^ n2399 ;
  assign n13718 = n13472 & n13717 ;
  assign n13719 = n13718 ^ n2204 ;
  assign n13720 = n13469 & n13719 ;
  assign n13721 = n13720 ^ n2064 ;
  assign n13722 = n13340 & ~n13447 ;
  assign n13723 = n13722 ^ n13103 ;
  assign n13724 = n13723 ^ n1739 ;
  assign n13725 = ~n13721 & ~n13724 ;
  assign n13726 = n13725 ^ n1763 ;
  assign n13727 = ~n13344 & ~n13447 ;
  assign n13728 = n13727 ^ n13101 ;
  assign n13729 = n13728 ^ n1572 ;
  assign n13730 = ~n13726 & ~n13729 ;
  assign n13731 = n13730 ^ n1605 ;
  assign n13732 = ~n13346 & ~n13447 ;
  assign n13733 = n13732 ^ n13098 ;
  assign n13734 = n13733 ^ n1427 ;
  assign n13735 = ~n13731 & ~n13734 ;
  assign n13736 = n13735 ^ n1450 ;
  assign n13739 = n13738 ^ n1290 ;
  assign n13740 = n13736 & ~n13739 ;
  assign n13742 = n13741 ^ n13740 ;
  assign n13743 = ~n13354 & ~n13447 ;
  assign n13744 = n13743 ^ n13356 ;
  assign n13745 = n13744 ^ n1136 ;
  assign n13746 = ~n13742 & n13745 ;
  assign n13747 = n13746 ^ n1143 ;
  assign n13748 = ~n13466 & n13747 ;
  assign n13749 = n13748 ^ n1072 ;
  assign n13750 = n13363 & ~n13447 ;
  assign n13751 = n13750 ^ n13365 ;
  assign n13754 = n13751 ^ n892 ;
  assign n13755 = ~n13749 & n13754 ;
  assign n13752 = n13751 ^ n786 ;
  assign n13756 = n13755 ^ n13752 ;
  assign n13757 = n13370 & ~n13447 ;
  assign n13758 = n13757 ^ n13372 ;
  assign n13759 = n13758 ^ n696 ;
  assign n13760 = n13759 ^ n842 ;
  assign n13761 = ~n13756 & n13760 ;
  assign n13762 = n13761 ^ n13759 ;
  assign n13763 = n13376 & ~n13447 ;
  assign n13764 = n13763 ^ n13378 ;
  assign n13765 = n13764 ^ n609 ;
  assign n13766 = n13765 ^ n835 ;
  assign n13767 = ~n13762 & n13766 ;
  assign n13768 = n13767 ^ n13765 ;
  assign n13769 = n13463 & ~n13768 ;
  assign n13770 = n13769 ^ n834 ;
  assign n13771 = n13460 & ~n13770 ;
  assign n13772 = n13771 ^ n750 ;
  assign n13773 = n13457 & n13772 ;
  assign n13774 = n13773 ^ n13456 ;
  assign n13777 = n13776 ^ n13774 ;
  assign n13778 = n13776 ^ n401 ;
  assign n13779 = ~n13777 & ~n13778 ;
  assign n13780 = n13779 ^ n462 ;
  assign n13781 = n13454 & n13780 ;
  assign n13782 = n13781 ^ n349 ;
  assign n13783 = n13399 & ~n13447 ;
  assign n13784 = n13783 ^ n13084 ;
  assign n13785 = n13784 ^ n291 ;
  assign n13786 = ~n13782 & ~n13785 ;
  assign n13787 = n13786 ^ n307 ;
  assign n13788 = n13450 & n13787 ;
  assign n13789 = n13788 ^ n13449 ;
  assign n13790 = n13789 ^ n188 ;
  assign n13796 = n13444 ^ n183 ;
  assign n13797 = n13444 ^ n13037 ;
  assign n13798 = n13797 ^ n13078 ;
  assign n13799 = n13798 ^ n13037 ;
  assign n13801 = ~n13406 & ~n13799 ;
  assign n13802 = n13801 ^ n13037 ;
  assign n13803 = ~n13796 & n13802 ;
  assign n13804 = n13803 ^ n13796 ;
  assign n13805 = ~n13404 & n13804 ;
  assign n13806 = n13805 ^ n13796 ;
  assign n13791 = ~n13432 & ~n13447 ;
  assign n13792 = n13791 ^ n13426 ;
  assign n13793 = n13792 ^ n13789 ;
  assign n13794 = n13790 & n13793 ;
  assign n13795 = n13794 ^ n203 ;
  assign n13807 = n13434 ^ n188 ;
  assign n13808 = ~n13447 & ~n13807 ;
  assign n13809 = n13808 ^ n13423 ;
  assign n13810 = n13809 ^ n157 ;
  assign n13811 = ~n13795 & ~n13810 ;
  assign n13812 = n13811 ^ n13809 ;
  assign n13813 = n13812 ^ n138 ;
  assign n13814 = n13437 ^ n157 ;
  assign n13815 = ~n13447 & n13814 ;
  assign n13816 = n13815 ^ n13421 ;
  assign n13817 = n13816 ^ n13812 ;
  assign n13818 = ~n13813 & ~n13817 ;
  assign n13819 = n13818 ^ n138 ;
  assign n13820 = n13819 ^ n183 ;
  assign n13821 = n13441 ^ n138 ;
  assign n13822 = ~n13447 & n13821 ;
  assign n13823 = n13822 ^ n13418 ;
  assign n13824 = n13823 ^ n13819 ;
  assign n13827 = ~n13820 & n13824 ;
  assign n13828 = n13827 ^ n183 ;
  assign n13829 = ~n13806 & n13828 ;
  assign n14182 = n13790 & ~n13829 ;
  assign n14183 = n14182 ^ n13792 ;
  assign n13833 = ~n13782 & ~n13829 ;
  assign n13834 = n13833 ^ n13784 ;
  assign n13835 = n13834 ^ n245 ;
  assign n13836 = n13780 & ~n13829 ;
  assign n13837 = n13836 ^ n13453 ;
  assign n13838 = n13837 ^ n291 ;
  assign n13839 = n13774 ^ n401 ;
  assign n13840 = ~n13829 & ~n13839 ;
  assign n13841 = n13840 ^ n13776 ;
  assign n13842 = n13841 ^ n341 ;
  assign n14164 = ~n13772 & ~n13829 ;
  assign n14165 = n14164 ^ n13456 ;
  assign n13843 = ~n13770 & ~n13829 ;
  assign n13844 = n13843 ^ n13459 ;
  assign n13845 = n13844 ^ n457 ;
  assign n13846 = ~n13768 & ~n13829 ;
  assign n13847 = n13846 ^ n13462 ;
  assign n13848 = n13847 ^ n534 ;
  assign n13849 = n13762 & ~n13829 ;
  assign n13850 = n13849 ^ n13764 ;
  assign n14158 = n13850 ^ n534 ;
  assign n13851 = n13850 ^ n609 ;
  assign n13852 = n13747 & ~n13829 ;
  assign n13853 = n13852 ^ n13465 ;
  assign n13854 = n13853 ^ n892 ;
  assign n13855 = ~n13736 & ~n13829 ;
  assign n13856 = n13855 ^ n13738 ;
  assign n13857 = n13856 ^ n1136 ;
  assign n14127 = ~n13731 & ~n13829 ;
  assign n14128 = n14127 ^ n13733 ;
  assign n14131 = n14128 ^ n1136 ;
  assign n13858 = ~n13726 & ~n13829 ;
  assign n13859 = n13858 ^ n13728 ;
  assign n13860 = n13859 ^ n1427 ;
  assign n14118 = ~n13721 & ~n13829 ;
  assign n14119 = n14118 ^ n13723 ;
  assign n14123 = n14119 ^ n1427 ;
  assign n13861 = n13715 & ~n13829 ;
  assign n13862 = n13861 ^ n13475 ;
  assign n13863 = n13862 ^ n2175 ;
  assign n13864 = n13706 ^ n2707 ;
  assign n13865 = ~n13829 & ~n13864 ;
  assign n13866 = n13865 ^ n13478 ;
  assign n13867 = n13866 ^ n2511 ;
  assign n13868 = ~n13704 & ~n13829 ;
  assign n13869 = n13868 ^ n13481 ;
  assign n13870 = n13869 ^ n2707 ;
  assign n13871 = n13695 & ~n13829 ;
  assign n13872 = n13871 ^ n13484 ;
  assign n13873 = n13872 ^ n3093 ;
  assign n14079 = n13688 ^ n3538 ;
  assign n14080 = ~n13829 & n14079 ;
  assign n14081 = n14080 ^ n13691 ;
  assign n13874 = n13681 ^ n3722 ;
  assign n13875 = ~n13829 & ~n13874 ;
  assign n13876 = n13875 ^ n13684 ;
  assign n13877 = n13876 ^ n3538 ;
  assign n13878 = n13674 ^ n3908 ;
  assign n13879 = ~n13829 & n13878 ;
  assign n13880 = n13879 ^ n13677 ;
  assign n13881 = n13880 ^ n3722 ;
  assign n13886 = n13651 ^ n5073 ;
  assign n13887 = ~n13829 & n13886 ;
  assign n13888 = n13887 ^ n13653 ;
  assign n13889 = n13888 ^ n4812 ;
  assign n13890 = n13649 & ~n13829 ;
  assign n13891 = n13890 ^ n13499 ;
  assign n13892 = n13891 ^ n5073 ;
  assign n13893 = n13647 & ~n13829 ;
  assign n13894 = n13893 ^ n13502 ;
  assign n13896 = n13894 ^ n5317 ;
  assign n14038 = n13645 & ~n13829 ;
  assign n14039 = n14038 ^ n13505 ;
  assign n13897 = ~n13640 & ~n13829 ;
  assign n13898 = n13897 ^ n13642 ;
  assign n13899 = n13898 ^ n5830 ;
  assign n13900 = ~n13638 & ~n13829 ;
  assign n13901 = n13900 ^ n13509 ;
  assign n13902 = n13901 ^ n6115 ;
  assign n13903 = n13631 ^ n6673 ;
  assign n13904 = ~n13829 & n13903 ;
  assign n13905 = n13904 ^ n13634 ;
  assign n13906 = n13905 ^ n6389 ;
  assign n14025 = n13629 & ~n13829 ;
  assign n14026 = n14025 ^ n13513 ;
  assign n13907 = ~n13622 & ~n13829 ;
  assign n13908 = n13907 ^ n13624 ;
  assign n13909 = n13908 ^ n7277 ;
  assign n14012 = ~n13617 & ~n13829 ;
  assign n14013 = n14012 ^ n13619 ;
  assign n14016 = n14013 ^ n7277 ;
  assign n13910 = n13612 & ~n13829 ;
  assign n13911 = n13910 ^ n13523 ;
  assign n13912 = n13911 ^ n8253 ;
  assign n13913 = ~n13610 & ~n13829 ;
  assign n13914 = n13913 ^ n13526 ;
  assign n13915 = n13914 ^ n8586 ;
  assign n13916 = n13603 ^ n9217 ;
  assign n13917 = ~n13829 & n13916 ;
  assign n13918 = n13917 ^ n13606 ;
  assign n13919 = n13918 ^ n8910 ;
  assign n13920 = ~n13601 & ~n13829 ;
  assign n13921 = n13920 ^ n13529 ;
  assign n13922 = n13921 ^ n9217 ;
  assign n13923 = ~n13596 & ~n13829 ;
  assign n13924 = n13923 ^ n13536 ;
  assign n13990 = n13924 ^ n9542 ;
  assign n13925 = n13924 ^ n10108 ;
  assign n13926 = n13583 & ~n13829 ;
  assign n13927 = n13926 ^ n13541 ;
  assign n13928 = n13927 ^ n11233 ;
  assign n13929 = ~n13577 & ~n13829 ;
  assign n13930 = n13929 ^ n13579 ;
  assign n13931 = n13930 ^ n11594 ;
  assign n13969 = n13575 & ~n13829 ;
  assign n13970 = n13969 ^ n13552 ;
  assign n13973 = n13970 ^ n11594 ;
  assign n13932 = n13573 & ~n13829 ;
  assign n13933 = n13932 ^ n13556 ;
  assign n13934 = n13933 ^ n12359 ;
  assign n13935 = n13559 ^ n13447 ;
  assign n13936 = ~n13829 & ~n13935 ;
  assign n13937 = n13936 ^ n13447 ;
  assign n13942 = n13937 ^ x6 ;
  assign n13943 = n13942 ^ n13082 ;
  assign n13944 = n13447 ^ x5 ;
  assign n13945 = n13944 ^ n13829 ;
  assign n13947 = ~x2 & ~x3 ;
  assign n13946 = n13447 ^ x4 ;
  assign n13948 = n13947 ^ n13946 ;
  assign n13949 = ~n13945 & ~n13948 ;
  assign n13958 = n13949 ^ n13558 ;
  assign n13950 = n13829 ^ n13447 ;
  assign n13955 = n13944 & n13950 ;
  assign n13956 = n13955 ^ n13949 ;
  assign n13957 = x4 & n13956 ;
  assign n13959 = n13958 ^ n13957 ;
  assign n13960 = ~n13943 & ~n13959 ;
  assign n13961 = n13960 ^ n13942 ;
  assign n13939 = ~n13562 & ~n13829 ;
  assign n13938 = x6 & ~n13937 ;
  assign n13940 = n13939 ^ n13938 ;
  assign n13941 = n13940 ^ n13560 ;
  assign n13962 = n13961 ^ n13941 ;
  assign n13963 = n13961 ^ n12731 ;
  assign n13964 = ~n13962 & ~n13963 ;
  assign n13965 = n13964 ^ n12731 ;
  assign n13966 = n13965 ^ n13933 ;
  assign n13967 = n13934 & ~n13966 ;
  assign n13968 = n13967 ^ n12452 ;
  assign n13971 = n13970 ^ n11960 ;
  assign n13972 = n13968 & ~n13971 ;
  assign n13974 = n13973 ^ n13972 ;
  assign n13975 = n13931 & ~n13974 ;
  assign n13976 = n13975 ^ n11688 ;
  assign n13977 = n13928 & n13976 ;
  assign n13978 = n13977 ^ n11326 ;
  assign n13979 = n13585 & ~n13829 ;
  assign n13980 = n13979 ^ n13538 ;
  assign n13981 = n13980 ^ n10875 ;
  assign n13982 = ~n13978 & ~n13981 ;
  assign n13983 = n13982 ^ n11327 ;
  assign n13984 = ~n13588 & ~n13829 ;
  assign n13985 = n13984 ^ n13591 ;
  assign n13986 = n13985 ^ n10468 ;
  assign n13987 = ~n13983 & n13986 ;
  assign n13988 = n13987 ^ n10639 ;
  assign n13989 = n13925 & n13988 ;
  assign n13991 = n13990 ^ n13989 ;
  assign n13992 = ~n13598 & ~n13829 ;
  assign n13993 = n13992 ^ n13532 ;
  assign n13994 = n13993 ^ n9542 ;
  assign n13995 = ~n13991 & ~n13994 ;
  assign n13996 = n13995 ^ n9628 ;
  assign n13997 = ~n13922 & n13996 ;
  assign n13998 = n13997 ^ n9285 ;
  assign n13999 = n13919 & ~n13998 ;
  assign n14000 = n13999 ^ n9005 ;
  assign n14001 = n13915 & n14000 ;
  assign n14002 = n14001 ^ n8688 ;
  assign n14003 = ~n13912 & n14002 ;
  assign n14004 = n14003 ^ n8253 ;
  assign n14005 = n14004 ^ n7891 ;
  assign n14006 = n13614 ^ n8253 ;
  assign n14007 = ~n13829 & n14006 ;
  assign n14008 = n14007 ^ n13520 ;
  assign n14009 = n14008 ^ n14004 ;
  assign n14010 = ~n14005 & n14009 ;
  assign n14011 = n14010 ^ n7971 ;
  assign n14014 = n14013 ^ n7584 ;
  assign n14015 = n14011 & ~n14014 ;
  assign n14017 = n14016 ^ n14015 ;
  assign n14018 = n13909 & ~n14017 ;
  assign n14019 = n14018 ^ n7339 ;
  assign n14020 = n13627 & ~n13829 ;
  assign n14021 = n14020 ^ n13516 ;
  assign n14022 = n14021 ^ n6959 ;
  assign n14023 = n14019 & ~n14022 ;
  assign n14024 = n14023 ^ n6959 ;
  assign n14027 = n14026 ^ n14024 ;
  assign n14028 = n14026 ^ n6673 ;
  assign n14029 = ~n14027 & n14028 ;
  assign n14030 = n14029 ^ n6713 ;
  assign n14031 = n13906 & ~n14030 ;
  assign n14032 = n14031 ^ n6389 ;
  assign n14033 = n14032 ^ n13901 ;
  assign n14034 = n13902 & n14033 ;
  assign n14035 = n14034 ^ n6429 ;
  assign n14036 = n13899 & ~n14035 ;
  assign n14037 = n14036 ^ n13898 ;
  assign n14040 = n14039 ^ n14037 ;
  assign n14041 = n14039 ^ n5562 ;
  assign n14042 = ~n14040 & n14041 ;
  assign n14043 = n14042 ^ n5885 ;
  assign n14044 = n13896 & ~n14043 ;
  assign n13895 = n13894 ^ n5073 ;
  assign n14045 = n14044 ^ n13895 ;
  assign n14046 = n13892 & n14045 ;
  assign n14047 = n14046 ^ n5073 ;
  assign n14048 = n14047 ^ n13888 ;
  assign n14049 = ~n13889 & n14048 ;
  assign n14050 = n14049 ^ n4854 ;
  assign n14051 = n13657 ^ n4812 ;
  assign n14052 = ~n13829 & n14051 ;
  assign n14053 = n14052 ^ n13490 ;
  assign n14054 = n14053 ^ n4583 ;
  assign n14055 = n14050 & ~n14054 ;
  assign n14056 = n14055 ^ n4645 ;
  assign n14059 = n13663 ^ n4153 ;
  assign n14057 = n13660 ^ n4583 ;
  assign n14058 = ~n13829 & n14057 ;
  assign n14060 = n14059 ^ n14058 ;
  assign n14061 = n14060 ^ n4414 ;
  assign n14062 = n14056 & ~n14061 ;
  assign n14063 = n14062 ^ n4414 ;
  assign n14064 = n13667 & ~n13829 ;
  assign n14065 = n14064 ^ n13487 ;
  assign n14066 = n14065 ^ n4153 ;
  assign n14067 = n14063 & ~n14066 ;
  assign n14068 = n14067 ^ n4153 ;
  assign n13884 = n13880 ^ n3908 ;
  assign n13882 = n13669 & ~n13829 ;
  assign n13883 = n13882 ^ n13671 ;
  assign n13885 = n13884 ^ n13883 ;
  assign n14069 = n14068 ^ n13885 ;
  assign n14070 = n14069 ^ n13884 ;
  assign n14071 = n13883 ^ n13880 ;
  assign n14072 = n14071 ^ n13884 ;
  assign n14073 = ~n14070 & n14072 ;
  assign n14074 = n14073 ^ n13884 ;
  assign n14075 = ~n13881 & ~n14074 ;
  assign n14076 = n14075 ^ n3795 ;
  assign n14077 = n13877 & n14076 ;
  assign n14078 = n14077 ^ n3538 ;
  assign n14082 = n14081 ^ n14078 ;
  assign n14083 = n14081 ^ n3320 ;
  assign n14084 = ~n14082 & n14083 ;
  assign n14085 = n14084 ^ n3387 ;
  assign n14086 = n13873 & n14085 ;
  assign n14087 = n14086 ^ n13872 ;
  assign n14088 = n14087 ^ n2894 ;
  assign n14089 = ~n13701 & ~n13829 ;
  assign n14090 = n14089 ^ n13699 ;
  assign n14091 = n14090 ^ n14087 ;
  assign n14092 = n14088 & n14091 ;
  assign n14093 = n14092 ^ n3396 ;
  assign n14094 = ~n13870 & ~n14093 ;
  assign n14095 = n14094 ^ n2707 ;
  assign n14096 = n14095 ^ n13866 ;
  assign n14097 = ~n13867 & ~n14096 ;
  assign n14098 = n14097 ^ n2530 ;
  assign n14099 = n13709 ^ n2511 ;
  assign n14100 = ~n13829 & ~n14099 ;
  assign n14101 = n14100 ^ n13711 ;
  assign n14102 = n14101 ^ n2366 ;
  assign n14103 = n14098 & ~n14102 ;
  assign n14104 = n14103 ^ n2399 ;
  assign n14105 = ~n13863 & n14104 ;
  assign n14106 = n14105 ^ n2204 ;
  assign n14108 = n13717 & ~n13829 ;
  assign n14107 = n13471 ^ n1739 ;
  assign n14109 = n14108 ^ n14107 ;
  assign n14110 = n14109 ^ n2064 ;
  assign n14111 = n14106 & n14110 ;
  assign n14112 = n14111 ^ n2064 ;
  assign n14113 = n13719 & ~n13829 ;
  assign n14114 = n14113 ^ n13468 ;
  assign n14115 = n14114 ^ n1739 ;
  assign n14116 = ~n14112 & ~n14115 ;
  assign n14117 = n14116 ^ n1739 ;
  assign n14120 = n14119 ^ n14117 ;
  assign n14121 = n14117 ^ n1572 ;
  assign n14122 = ~n14120 & n14121 ;
  assign n14124 = n14123 ^ n14122 ;
  assign n14125 = n13860 & ~n14124 ;
  assign n14126 = n14125 ^ n1450 ;
  assign n14129 = n14128 ^ n1290 ;
  assign n14130 = n14126 & n14129 ;
  assign n14132 = n14131 ^ n14130 ;
  assign n14133 = ~n13857 & n14132 ;
  assign n14134 = n14133 ^ n1143 ;
  assign n14135 = ~n13742 & ~n13829 ;
  assign n14136 = n14135 ^ n13744 ;
  assign n14139 = n14136 ^ n1034 ;
  assign n14140 = ~n14134 & n14139 ;
  assign n14137 = n14136 ^ n892 ;
  assign n14141 = n14140 ^ n14137 ;
  assign n14142 = ~n13854 & n14141 ;
  assign n14143 = n14142 ^ n927 ;
  assign n14144 = n13749 & ~n13829 ;
  assign n14145 = n14144 ^ n13751 ;
  assign n14148 = n14145 ^ n786 ;
  assign n14149 = ~n14143 & n14148 ;
  assign n14146 = n14145 ^ n696 ;
  assign n14150 = n14149 ^ n14146 ;
  assign n14151 = n13756 & ~n13829 ;
  assign n14152 = n14151 ^ n13758 ;
  assign n14153 = n14152 ^ n609 ;
  assign n14154 = n14153 ^ n835 ;
  assign n14155 = ~n14150 & n14154 ;
  assign n14156 = n14155 ^ n14153 ;
  assign n14157 = ~n13851 & n14156 ;
  assign n14159 = n14158 ^ n14157 ;
  assign n14160 = ~n13848 & n14159 ;
  assign n14161 = n14160 ^ n750 ;
  assign n14162 = ~n13845 & n14161 ;
  assign n14163 = n14162 ^ n13844 ;
  assign n14166 = n14165 ^ n14163 ;
  assign n14167 = n14165 ^ n401 ;
  assign n14168 = n14166 & ~n14167 ;
  assign n14169 = n14168 ^ n462 ;
  assign n14170 = ~n13842 & n14169 ;
  assign n14171 = n14170 ^ n349 ;
  assign n14172 = ~n13838 & ~n14171 ;
  assign n14173 = n14172 ^ n307 ;
  assign n14174 = n13835 & n14173 ;
  assign n14175 = n14174 ^ n13834 ;
  assign n14176 = n14175 ^ n188 ;
  assign n14177 = ~n13787 & ~n13829 ;
  assign n14178 = n14177 ^ n13449 ;
  assign n14179 = n14178 ^ n14175 ;
  assign n14180 = n14176 & ~n14179 ;
  assign n14181 = n14180 ^ n188 ;
  assign n14184 = n14183 ^ n14181 ;
  assign n14185 = n14181 ^ n157 ;
  assign n14186 = ~n14184 & ~n14185 ;
  assign n14187 = n14186 ^ n14183 ;
  assign n14189 = ~n138 & n14187 ;
  assign n14188 = n14187 ^ n138 ;
  assign n14190 = n14189 ^ n14188 ;
  assign n14197 = n13823 ^ n13404 ;
  assign n14198 = n14197 ^ n13803 ;
  assign n14199 = n14198 ^ n13823 ;
  assign n14200 = n13404 & n13444 ;
  assign n14201 = n13823 & n14200 ;
  assign n14202 = n14201 ^ n13823 ;
  assign n14205 = n14199 & n14202 ;
  assign n14206 = n14205 ^ n13823 ;
  assign n14207 = n13819 & ~n14206 ;
  assign n14208 = n14207 ^ n13823 ;
  assign n14209 = n183 & n14208 ;
  assign n13830 = n13795 & ~n13829 ;
  assign n13831 = n13830 ^ n13809 ;
  assign n14193 = n13831 ^ n138 ;
  assign n14194 = n14187 ^ n13831 ;
  assign n14195 = ~n14193 & ~n14194 ;
  assign n14196 = n14195 ^ n138 ;
  assign n14210 = n14209 ^ n14196 ;
  assign n14211 = ~n13813 & ~n13829 ;
  assign n14212 = n14211 ^ n13816 ;
  assign n14213 = n13416 ^ n13404 ;
  assign n14214 = ~n183 & n14202 ;
  assign n14215 = ~n13444 & n14214 ;
  assign n14216 = ~n14213 & n14215 ;
  assign n14217 = n14216 ^ n14214 ;
  assign n14218 = n14217 ^ n183 ;
  assign n14219 = n13824 & ~n14218 ;
  assign n14220 = n14219 ^ n183 ;
  assign n14221 = n14212 & ~n14220 ;
  assign n14222 = n14221 ^ n14212 ;
  assign n14223 = ~n14209 & ~n14222 ;
  assign n14224 = n14223 ^ n14212 ;
  assign n14225 = ~n14210 & ~n14224 ;
  assign n14226 = n14225 ^ n14209 ;
  assign n14227 = ~n14189 & ~n14226 ;
  assign n14230 = ~n14190 & n14227 ;
  assign n13832 = n13831 ^ n183 ;
  assign n14231 = n14230 ^ n13832 ;
  assign n14250 = n14221 ^ n14209 ;
  assign n14251 = n14250 ^ n14224 ;
  assign n14252 = n14251 ^ n183 ;
  assign n14253 = n14212 ^ n14196 ;
  assign n14254 = ~n14252 & ~n14253 ;
  assign n14234 = n14212 ^ n13831 ;
  assign n14237 = n14227 & ~n14234 ;
  assign n14232 = n14227 ^ n13831 ;
  assign n14238 = n14237 ^ n14232 ;
  assign n14239 = n14190 & n14238 ;
  assign n14240 = n14239 ^ n14232 ;
  assign n14241 = ~n183 & n14240 ;
  assign n14242 = n14212 ^ n14189 ;
  assign n14243 = n14242 ^ n14234 ;
  assign n14244 = n14234 ^ n14226 ;
  assign n14245 = n14244 ^ n14234 ;
  assign n14246 = ~n14243 & ~n14245 ;
  assign n14247 = n14246 ^ n14234 ;
  assign n14248 = n14241 & ~n14247 ;
  assign n14249 = n14248 ^ n183 ;
  assign n14255 = n14254 ^ n14249 ;
  assign n14256 = n14176 & ~n14226 ;
  assign n14257 = n14256 ^ n14178 ;
  assign n14258 = n14257 ^ n157 ;
  assign n14261 = ~n14161 & ~n14226 ;
  assign n14262 = n14261 ^ n13844 ;
  assign n14263 = n14262 ^ n401 ;
  assign n14655 = n14159 & ~n14226 ;
  assign n14656 = n14655 ^ n13847 ;
  assign n14665 = n14656 ^ n14262 ;
  assign n14264 = ~n14156 & ~n14226 ;
  assign n14265 = n14264 ^ n14158 ;
  assign n14646 = n14150 & ~n14226 ;
  assign n14647 = n14646 ^ n14152 ;
  assign n14657 = n14656 ^ n14647 ;
  assign n14593 = ~n14112 & ~n14226 ;
  assign n14594 = n14593 ^ n14114 ;
  assign n14595 = n14594 ^ n1739 ;
  assign n14266 = n14104 & ~n14226 ;
  assign n14267 = n14266 ^ n13862 ;
  assign n14268 = n14267 ^ n2008 ;
  assign n14569 = n14095 ^ n2511 ;
  assign n14570 = ~n14226 & ~n14569 ;
  assign n14269 = ~n14093 & ~n14226 ;
  assign n14270 = n14269 ^ n13869 ;
  assign n14271 = n14270 ^ n2511 ;
  assign n14279 = n14068 ^ n3908 ;
  assign n14280 = ~n14226 & n14279 ;
  assign n14281 = n14280 ^ n13883 ;
  assign n14282 = n14281 ^ n3722 ;
  assign n14283 = n14056 & ~n14226 ;
  assign n14284 = n14283 ^ n14060 ;
  assign n14505 = n14047 ^ n4812 ;
  assign n14506 = ~n14226 & n14505 ;
  assign n14288 = n14045 & ~n14226 ;
  assign n14289 = n14288 ^ n13891 ;
  assign n14290 = n14289 ^ n4812 ;
  assign n14291 = n14043 & ~n14226 ;
  assign n14292 = n14291 ^ n13894 ;
  assign n14293 = n14292 ^ n5073 ;
  assign n14294 = n14037 ^ n5562 ;
  assign n14295 = ~n14226 & n14294 ;
  assign n14296 = n14295 ^ n14039 ;
  assign n14297 = ~n5317 & ~n14296 ;
  assign n14298 = n14293 & ~n14297 ;
  assign n14299 = n14035 & ~n14226 ;
  assign n14300 = n14299 ^ n13898 ;
  assign n14301 = n14300 ^ n5562 ;
  assign n14302 = ~n14030 & ~n14226 ;
  assign n14303 = n14302 ^ n13905 ;
  assign n14304 = ~n6115 & n14303 ;
  assign n14305 = n14032 ^ n6115 ;
  assign n14306 = ~n14226 & ~n14305 ;
  assign n14307 = n14306 ^ n13901 ;
  assign n14309 = n5830 & n14307 ;
  assign n14308 = n14307 ^ n5830 ;
  assign n14310 = n14309 ^ n14308 ;
  assign n14311 = ~n14304 & n14310 ;
  assign n14312 = n14301 & n14311 ;
  assign n14313 = n14024 ^ n6673 ;
  assign n14314 = ~n14226 & n14313 ;
  assign n14315 = n14314 ^ n14026 ;
  assign n14316 = ~n6389 & n14315 ;
  assign n14317 = n14303 ^ n6115 ;
  assign n14318 = n14317 ^ n14304 ;
  assign n14319 = ~n14316 & ~n14318 ;
  assign n14320 = n14019 & ~n14226 ;
  assign n14321 = n14320 ^ n14021 ;
  assign n14322 = ~n6673 & n14321 ;
  assign n14323 = n14315 ^ n6389 ;
  assign n14324 = n14323 ^ n14316 ;
  assign n14325 = ~n14322 & ~n14324 ;
  assign n14326 = ~n14017 & ~n14226 ;
  assign n14327 = n14326 ^ n13908 ;
  assign n14328 = n6959 & n14327 ;
  assign n14329 = n14321 ^ n6673 ;
  assign n14330 = n14329 ^ n14322 ;
  assign n14331 = ~n14328 & ~n14330 ;
  assign n14332 = ~n14011 & ~n14226 ;
  assign n14333 = n14332 ^ n14013 ;
  assign n14334 = ~n7277 & n14333 ;
  assign n14335 = n14327 ^ n6959 ;
  assign n14336 = n14335 ^ n14328 ;
  assign n14337 = ~n14334 & n14336 ;
  assign n14338 = ~n14005 & ~n14226 ;
  assign n14339 = n14338 ^ n14008 ;
  assign n14340 = n7584 & ~n14339 ;
  assign n14341 = n14333 ^ n7277 ;
  assign n14342 = n14341 ^ n14334 ;
  assign n14343 = ~n14340 & ~n14342 ;
  assign n14344 = n14002 & ~n14226 ;
  assign n14345 = n14344 ^ n13911 ;
  assign n14346 = n7891 & n14345 ;
  assign n14347 = n14339 ^ n7584 ;
  assign n14348 = n14347 ^ n14340 ;
  assign n14349 = ~n14346 & ~n14348 ;
  assign n14350 = n14000 & ~n14226 ;
  assign n14351 = n14350 ^ n13914 ;
  assign n14352 = n8253 & n14351 ;
  assign n14353 = n14345 ^ n7891 ;
  assign n14354 = n14353 ^ n14346 ;
  assign n14355 = ~n14352 & n14354 ;
  assign n14356 = ~n13991 & ~n14226 ;
  assign n14357 = n14356 ^ n13993 ;
  assign n14359 = n14357 ^ n9217 ;
  assign n14358 = ~n9217 & n14357 ;
  assign n14360 = n14359 ^ n14358 ;
  assign n14362 = n13996 & ~n14226 ;
  assign n14361 = n13921 ^ n8910 ;
  assign n14363 = n14362 ^ n14361 ;
  assign n14364 = ~n14360 & n14363 ;
  assign n14365 = ~n13988 & ~n14226 ;
  assign n14366 = n14365 ^ n13924 ;
  assign n14367 = n14366 ^ n9542 ;
  assign n14368 = ~n13983 & ~n14226 ;
  assign n14369 = n14368 ^ n13985 ;
  assign n14371 = n14369 ^ n10108 ;
  assign n14452 = ~n13978 & ~n14226 ;
  assign n14453 = n14452 ^ n13980 ;
  assign n14454 = n14453 ^ n10875 ;
  assign n14372 = ~n13974 & ~n14226 ;
  assign n14373 = n14372 ^ n13930 ;
  assign n14374 = n14373 ^ n11233 ;
  assign n14379 = n13965 ^ n12359 ;
  assign n14380 = ~n14226 & n14379 ;
  assign n14378 = n13933 ^ n11960 ;
  assign n14381 = n14380 ^ n14378 ;
  assign n14382 = ~n13963 & ~n14226 ;
  assign n14383 = n14382 ^ n13941 ;
  assign n14384 = n14383 ^ n12359 ;
  assign n14389 = n13829 ^ x3 ;
  assign n14390 = n14226 ^ n13829 ;
  assign n14391 = n14389 & ~n14390 ;
  assign n14392 = n14391 ^ x3 ;
  assign n14388 = n14226 ^ x3 ;
  assign n14393 = n14392 ^ n14388 ;
  assign n14394 = n14393 ^ n13829 ;
  assign n14395 = n14394 ^ n14392 ;
  assign n14398 = ~x0 & ~x1 ;
  assign n14396 = x3 ^ x2 ;
  assign n14397 = n14396 ^ n14226 ;
  assign n14399 = n14398 ^ n14397 ;
  assign n14400 = ~n14395 & n14399 ;
  assign n14401 = n14400 ^ n14393 ;
  assign n14402 = ~x2 & ~n14401 ;
  assign n14403 = n14402 ^ n14392 ;
  assign n14387 = n13947 ^ x4 ;
  assign n14404 = n14403 ^ n14387 ;
  assign n14385 = n13947 ^ n13829 ;
  assign n14386 = n14226 & ~n14385 ;
  assign n14405 = n14404 ^ n14386 ;
  assign n14414 = ~x4 & ~n13829 ;
  assign n14406 = n13950 ^ x4 ;
  assign n14407 = n14406 ^ n13950 ;
  assign n14410 = ~n14385 & ~n14407 ;
  assign n14411 = n14410 ^ n13950 ;
  assign n14412 = ~n14226 & n14411 ;
  assign n14413 = n14412 ^ x5 ;
  assign n14415 = n14414 ^ n14413 ;
  assign n14416 = n14415 ^ n13447 ;
  assign n14417 = n14416 ^ n14403 ;
  assign n14418 = n14417 ^ n14415 ;
  assign n14419 = ~n14405 & n14418 ;
  assign n14420 = n14419 ^ n14416 ;
  assign n14421 = n13959 & ~n14226 ;
  assign n14422 = n14421 ^ n13942 ;
  assign n14424 = n14422 ^ n14415 ;
  assign n14423 = n14422 ^ n13082 ;
  assign n14425 = n14424 ^ n14423 ;
  assign n14426 = n14420 & n14425 ;
  assign n14427 = n14426 ^ n14424 ;
  assign n14429 = n14383 ^ n12731 ;
  assign n14428 = n14422 ^ n14383 ;
  assign n14430 = n14429 ^ n14428 ;
  assign n14431 = n14427 & ~n14430 ;
  assign n14432 = n14431 ^ n14429 ;
  assign n14433 = ~n14384 & n14432 ;
  assign n14434 = n14433 ^ n12452 ;
  assign n14435 = ~n14381 & ~n14434 ;
  assign n14375 = ~n13968 & ~n14226 ;
  assign n14376 = n14375 ^ n13970 ;
  assign n14377 = n14376 ^ n11960 ;
  assign n14436 = n14435 ^ n14377 ;
  assign n14438 = n14373 ^ n11594 ;
  assign n14437 = n14376 ^ n14373 ;
  assign n14439 = n14438 ^ n14437 ;
  assign n14440 = n14436 & ~n14439 ;
  assign n14441 = n14440 ^ n14438 ;
  assign n14442 = n14374 & ~n14441 ;
  assign n14443 = n14442 ^ n11326 ;
  assign n14444 = n13927 ^ n10875 ;
  assign n14445 = n14444 ^ n14226 ;
  assign n14446 = n14445 ^ n14444 ;
  assign n14447 = n14444 ^ n13976 ;
  assign n14448 = n14447 ^ n14444 ;
  assign n14449 = ~n14446 & n14448 ;
  assign n14450 = n14449 ^ n14444 ;
  assign n14451 = ~n14443 & ~n14450 ;
  assign n14455 = n14454 ^ n14451 ;
  assign n14457 = n14369 ^ n10468 ;
  assign n14456 = n14453 ^ n14369 ;
  assign n14458 = n14457 ^ n14456 ;
  assign n14459 = n14455 & n14458 ;
  assign n14460 = n14459 ^ n14457 ;
  assign n14461 = ~n14371 & n14460 ;
  assign n14370 = n14369 ^ n14366 ;
  assign n14462 = n14461 ^ n14370 ;
  assign n14463 = ~n14367 & n14462 ;
  assign n14464 = n14463 ^ n9542 ;
  assign n14465 = n14364 & ~n14464 ;
  assign n14466 = ~n13998 & ~n14226 ;
  assign n14467 = n14466 ^ n13918 ;
  assign n14468 = n14467 ^ n8586 ;
  assign n14469 = n14358 ^ n8910 ;
  assign n14472 = ~n14363 & n14469 ;
  assign n14473 = n14472 ^ n14358 ;
  assign n14474 = n14468 & ~n14473 ;
  assign n14475 = ~n14465 & n14474 ;
  assign n14476 = n14351 ^ n8253 ;
  assign n14477 = n14476 ^ n14352 ;
  assign n14478 = ~n8586 & ~n14467 ;
  assign n14479 = n14477 & n14478 ;
  assign n14480 = n14479 ^ n14477 ;
  assign n14481 = ~n14475 & n14480 ;
  assign n14482 = n14355 & ~n14481 ;
  assign n14483 = n14349 & ~n14482 ;
  assign n14484 = n14343 & ~n14483 ;
  assign n14485 = n14337 & ~n14484 ;
  assign n14486 = n14331 & ~n14485 ;
  assign n14487 = n14325 & ~n14486 ;
  assign n14488 = n14319 & ~n14487 ;
  assign n14489 = n14312 & ~n14488 ;
  assign n14490 = n14309 ^ n14300 ;
  assign n14491 = n14301 & ~n14490 ;
  assign n14492 = n14491 ^ n5562 ;
  assign n14493 = ~n14489 & ~n14492 ;
  assign n14494 = n14298 & ~n14493 ;
  assign n14495 = n14296 ^ n5317 ;
  assign n14496 = n14495 ^ n14297 ;
  assign n14497 = n14496 ^ n14292 ;
  assign n14498 = n14293 & n14497 ;
  assign n14499 = n14498 ^ n5073 ;
  assign n14500 = ~n14494 & ~n14499 ;
  assign n14501 = n14500 ^ n14289 ;
  assign n14502 = n14290 & n14501 ;
  assign n14503 = n14502 ^ n4812 ;
  assign n14504 = n14503 ^ n13888 ;
  assign n14507 = n14506 ^ n14504 ;
  assign n14508 = n14050 & ~n14226 ;
  assign n14509 = n14508 ^ n14053 ;
  assign n14510 = n14509 ^ n4583 ;
  assign n14511 = n14510 ^ n14503 ;
  assign n14512 = n14511 ^ n14509 ;
  assign n14513 = n14507 & n14512 ;
  assign n14514 = n14513 ^ n14510 ;
  assign n14285 = n14063 & ~n14226 ;
  assign n14286 = n14285 ^ n14065 ;
  assign n14516 = n14509 ^ n14286 ;
  assign n14515 = n14286 ^ n4356 ;
  assign n14517 = n14516 ^ n14515 ;
  assign n14518 = ~n14514 & ~n14517 ;
  assign n14519 = n14518 ^ n14516 ;
  assign n14287 = n14286 ^ n4153 ;
  assign n14520 = n14519 ^ n14287 ;
  assign n14521 = n14284 & ~n14520 ;
  assign n14522 = n14521 ^ n14519 ;
  assign n14524 = n14281 ^ n3908 ;
  assign n14523 = n14286 ^ n14281 ;
  assign n14525 = n14524 ^ n14523 ;
  assign n14526 = ~n14522 & ~n14525 ;
  assign n14527 = n14526 ^ n14524 ;
  assign n14528 = ~n14282 & ~n14527 ;
  assign n14529 = n14528 ^ n3722 ;
  assign n14530 = n14529 ^ n13880 ;
  assign n14272 = n14068 ^ n3722 ;
  assign n14273 = n14272 ^ n3961 ;
  assign n14274 = n13883 ^ n3722 ;
  assign n14275 = n14274 ^ n3961 ;
  assign n14276 = n14273 & n14275 ;
  assign n14277 = n14276 ^ n3961 ;
  assign n14278 = ~n14226 & ~n14277 ;
  assign n14531 = n14530 ^ n14278 ;
  assign n14532 = n14076 & ~n14226 ;
  assign n14533 = n14532 ^ n13876 ;
  assign n14534 = n14533 ^ n3538 ;
  assign n14535 = n14534 ^ n14529 ;
  assign n14536 = n14535 ^ n14533 ;
  assign n14537 = n14531 & n14536 ;
  assign n14538 = n14537 ^ n14534 ;
  assign n14539 = n14078 ^ n3320 ;
  assign n14540 = ~n14226 & n14539 ;
  assign n14541 = n14540 ^ n14081 ;
  assign n14543 = n14541 ^ n3320 ;
  assign n14542 = n14541 ^ n14533 ;
  assign n14544 = n14543 ^ n14542 ;
  assign n14545 = ~n14538 & n14544 ;
  assign n14546 = n14545 ^ n14543 ;
  assign n14547 = ~n14085 & ~n14226 ;
  assign n14548 = n14547 ^ n13872 ;
  assign n14550 = n14548 ^ n14541 ;
  assign n14549 = n14548 ^ n3093 ;
  assign n14551 = n14550 ^ n14549 ;
  assign n14552 = n14546 & ~n14551 ;
  assign n14553 = n14552 ^ n14550 ;
  assign n14554 = n14088 & ~n14226 ;
  assign n14555 = n14554 ^ n14090 ;
  assign n14557 = n14555 ^ n2894 ;
  assign n14556 = n14555 ^ n14548 ;
  assign n14558 = n14557 ^ n14556 ;
  assign n14559 = n14553 & n14558 ;
  assign n14560 = n14559 ^ n14557 ;
  assign n14562 = n14270 ^ n2707 ;
  assign n14561 = n14555 ^ n14270 ;
  assign n14563 = n14562 ^ n14561 ;
  assign n14564 = n14560 & n14563 ;
  assign n14565 = n14564 ^ n14562 ;
  assign n14566 = n14271 & n14565 ;
  assign n14567 = n14566 ^ n2511 ;
  assign n14568 = n14567 ^ n13866 ;
  assign n14571 = n14570 ^ n14568 ;
  assign n14572 = n14098 & ~n14226 ;
  assign n14573 = n14572 ^ n14101 ;
  assign n14574 = n14573 ^ n2366 ;
  assign n14575 = n14574 ^ n14567 ;
  assign n14576 = n14575 ^ n14573 ;
  assign n14577 = n14571 & n14576 ;
  assign n14578 = n14577 ^ n14574 ;
  assign n14580 = n14267 ^ n2175 ;
  assign n14579 = n14573 ^ n14267 ;
  assign n14581 = n14580 ^ n14579 ;
  assign n14582 = n14578 & ~n14581 ;
  assign n14583 = n14582 ^ n14580 ;
  assign n14584 = ~n14268 & n14583 ;
  assign n14585 = n14584 ^ n2064 ;
  assign n14588 = n14109 ^ n14106 ;
  assign n14589 = n14588 ^ n14109 ;
  assign n14590 = ~n14226 & n14589 ;
  assign n14591 = n14590 ^ n14109 ;
  assign n14592 = ~n14585 & ~n14591 ;
  assign n14596 = n14595 ^ n14592 ;
  assign n14597 = ~n14121 & ~n14226 ;
  assign n14598 = n14597 ^ n14119 ;
  assign n14599 = n14598 ^ n14594 ;
  assign n14600 = n14599 ^ n14598 ;
  assign n14601 = n14600 ^ n1572 ;
  assign n14602 = ~n14596 & n14601 ;
  assign n14603 = n14602 ^ n14599 ;
  assign n14604 = ~n14124 & ~n14226 ;
  assign n14605 = n14604 ^ n13859 ;
  assign n14607 = n14605 ^ n1427 ;
  assign n14606 = n14605 ^ n14598 ;
  assign n14608 = n14607 ^ n14606 ;
  assign n14609 = ~n14603 & ~n14608 ;
  assign n14610 = n14609 ^ n14607 ;
  assign n14611 = ~n14126 & ~n14226 ;
  assign n14612 = n14611 ^ n14128 ;
  assign n14614 = n14612 ^ n14605 ;
  assign n14613 = n14612 ^ n1290 ;
  assign n14615 = n14614 ^ n14613 ;
  assign n14616 = n14610 & ~n14615 ;
  assign n14617 = n14616 ^ n14614 ;
  assign n14618 = n14132 & ~n14226 ;
  assign n14619 = n14618 ^ n13856 ;
  assign n14621 = n14619 ^ n14612 ;
  assign n14620 = n14619 ^ n1136 ;
  assign n14622 = n14621 ^ n14620 ;
  assign n14623 = n14617 & n14622 ;
  assign n14624 = n14623 ^ n14620 ;
  assign n14625 = n14134 & ~n14226 ;
  assign n14626 = n14625 ^ n14136 ;
  assign n14628 = n14626 ^ n14619 ;
  assign n14627 = n14626 ^ n1034 ;
  assign n14629 = n14628 ^ n14627 ;
  assign n14630 = ~n14624 & ~n14629 ;
  assign n14631 = n14630 ^ n14628 ;
  assign n14632 = n14141 & ~n14226 ;
  assign n14633 = n14632 ^ n13853 ;
  assign n14635 = n14633 ^ n14626 ;
  assign n14634 = n14633 ^ n892 ;
  assign n14636 = n14635 ^ n14634 ;
  assign n14637 = ~n14631 & n14636 ;
  assign n14638 = n14637 ^ n14635 ;
  assign n14639 = n14143 & ~n14226 ;
  assign n14640 = n14639 ^ n14145 ;
  assign n14642 = n14640 ^ n14633 ;
  assign n14641 = n14640 ^ n786 ;
  assign n14643 = n14642 ^ n14641 ;
  assign n14644 = ~n14638 & ~n14643 ;
  assign n14645 = n14644 ^ n14642 ;
  assign n14649 = n14647 ^ n14640 ;
  assign n14648 = n14647 ^ n696 ;
  assign n14650 = n14649 ^ n14648 ;
  assign n14651 = ~n14645 & n14650 ;
  assign n14652 = n14651 ^ n14649 ;
  assign n14653 = n14647 ^ n609 ;
  assign n14654 = n14652 & ~n14653 ;
  assign n14658 = n14657 ^ n14654 ;
  assign n14659 = n14658 ^ n14656 ;
  assign n14660 = n14659 ^ n534 ;
  assign n14661 = ~n14265 & n14660 ;
  assign n14662 = n14661 ^ n14658 ;
  assign n14663 = n14656 ^ n457 ;
  assign n14664 = ~n14662 & n14663 ;
  assign n14666 = n14665 ^ n14664 ;
  assign n14667 = n14263 & n14666 ;
  assign n14668 = n14667 ^ n401 ;
  assign n14669 = n14668 ^ n14165 ;
  assign n14259 = n14163 ^ n401 ;
  assign n14260 = ~n14226 & n14259 ;
  assign n14670 = n14669 ^ n14260 ;
  assign n14671 = n14169 & ~n14226 ;
  assign n14672 = n14671 ^ n13841 ;
  assign n14673 = n14672 ^ n341 ;
  assign n14674 = n14673 ^ n14668 ;
  assign n14675 = n14674 ^ n14672 ;
  assign n14676 = n14670 & n14675 ;
  assign n14677 = n14676 ^ n14673 ;
  assign n14678 = ~n14171 & ~n14226 ;
  assign n14679 = n14678 ^ n13837 ;
  assign n14681 = n14679 ^ n291 ;
  assign n14680 = n14679 ^ n14672 ;
  assign n14682 = n14681 ^ n14680 ;
  assign n14683 = n14677 & n14682 ;
  assign n14684 = n14683 ^ n14681 ;
  assign n14685 = ~n14173 & ~n14226 ;
  assign n14686 = n14685 ^ n13834 ;
  assign n14688 = n14686 ^ n14679 ;
  assign n14687 = n14686 ^ n245 ;
  assign n14689 = n14688 ^ n14687 ;
  assign n14690 = ~n14684 & n14689 ;
  assign n14691 = n14690 ^ n14688 ;
  assign n14693 = n14257 ^ n188 ;
  assign n14692 = n14686 ^ n14257 ;
  assign n14694 = n14693 ^ n14692 ;
  assign n14695 = ~n14691 & n14694 ;
  assign n14696 = n14695 ^ n14693 ;
  assign n14697 = n14258 & n14696 ;
  assign n14698 = n14697 ^ n14257 ;
  assign n14699 = n14698 ^ n138 ;
  assign n14700 = n14698 ^ n14183 ;
  assign n14701 = n14700 ^ n14226 ;
  assign n14702 = n14701 ^ n14700 ;
  assign n14703 = n14700 ^ n14185 ;
  assign n14704 = n14703 ^ n14700 ;
  assign n14705 = ~n14702 & n14704 ;
  assign n14706 = n14705 ^ n14700 ;
  assign n14707 = n14699 & n14706 ;
  assign n14708 = n14707 ^ n138 ;
  assign n14709 = n14255 & n14708 ;
  assign n14710 = n14231 & n14709 ;
  assign n14711 = n14710 ^ n14255 ;
  assign y0 = ~n14711 ;
  assign y1 = ~n14226 ;
  assign y2 = ~n13829 ;
  assign y3 = ~n13447 ;
  assign y4 = ~n13082 ;
  assign y5 = ~n12731 ;
  assign y6 = ~n12359 ;
  assign y7 = n11960 ;
  assign y8 = n11594 ;
  assign y9 = n11233 ;
  assign y10 = ~n10875 ;
  assign y11 = n10468 ;
  assign y12 = ~n10108 ;
  assign y13 = n9542 ;
  assign y14 = n9217 ;
  assign y15 = ~n8910 ;
  assign y16 = ~n8586 ;
  assign y17 = ~n8253 ;
  assign y18 = n7891 ;
  assign y19 = ~n7584 ;
  assign y20 = ~n7277 ;
  assign y21 = ~n6959 ;
  assign y22 = ~n6673 ;
  assign y23 = n6389 ;
  assign y24 = ~n6115 ;
  assign y25 = ~n5830 ;
  assign y26 = ~n5562 ;
  assign y27 = ~n5317 ;
  assign y28 = ~n5073 ;
  assign y29 = ~n4812 ;
  assign y30 = ~n4583 ;
  assign y31 = ~n4356 ;
  assign y32 = ~n4153 ;
  assign y33 = ~n3908 ;
  assign y34 = n3722 ;
  assign y35 = n3538 ;
  assign y36 = n3320 ;
  assign y37 = ~n3093 ;
  assign y38 = ~n2894 ;
  assign y39 = n2707 ;
  assign y40 = ~n2511 ;
  assign y41 = ~n2366 ;
  assign y42 = ~n2175 ;
  assign y43 = ~n2008 ;
  assign y44 = n1739 ;
  assign y45 = ~n1572 ;
  assign y46 = n1427 ;
  assign y47 = ~n1290 ;
  assign y48 = ~n1136 ;
  assign y49 = ~n1034 ;
  assign y50 = ~n892 ;
  assign y51 = ~n786 ;
  assign y52 = ~n696 ;
  assign y53 = n609 ;
  assign y54 = ~n534 ;
  assign y55 = n457 ;
  assign y56 = ~n401 ;
  assign y57 = ~n341 ;
  assign y58 = n291 ;
  assign y59 = ~n245 ;
  assign y60 = ~n188 ;
  assign y61 = ~n157 ;
  assign y62 = ~n138 ;
  assign y63 = n183 ;
endmodule
