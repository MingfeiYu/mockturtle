module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n757 , n758 , n759 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n933 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n954 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n985 , n986 , n987 , n988 , n991 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1006 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1086 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1163 , n1164 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1310 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1350 , n1351 , n1352 , n1353 , n1356 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1390 , n1395 , n1396 , n1397 , n1398 , n1399 , n1402 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1414 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1443 , n1444 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1474 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1490 , n1491 , n1492 , n1493 , n1494 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1519 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1533 , n1534 , n1535 , n1536 , n1537 , n1539 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1549 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1563 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1598 , n1599 , n1600 , n1601 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1690 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1703 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1730 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1764 , n1766 , n1767 , n1768 , n1769 , n1770 , n1773 , n1775 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1794 , n1801 , n1802 , n1816 , n1817 , n1818 , n1819 , n1820 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1835 , n1840 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2051 , n2052 , n2053 , n2054 , n2055 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2096 , n2097 , n2098 , n2099 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2337 , n2338 , n2339 , n2340 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2839 , n2840 , n2841 , n2842 , n2844 , n2845 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2880 , n2881 , n2882 , n2883 , n2884 , n2887 , n2888 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2945 , n2946 , n2947 , n2948 , n2949 , n2952 , n2953 , n2955 , n2956 , n2957 , n2958 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3103 , n3104 , n3105 , n3108 , n3109 , n3110 , n3111 , n3112 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3435 , n3436 , n3437 , n3438 , n3439 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3475 , n3476 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3694 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3811 , n3814 , n3815 , n3816 , n3818 , n3819 , n3820 , n3821 , n3823 , n3825 , n3826 , n3827 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3969 , n3970 , n3972 , n3973 , n3974 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3989 , n3991 , n3993 , n3994 , n3995 , n3996 , n3997 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4091 , n4094 , n4095 , n4096 , n4098 , n4099 , n4100 , n4101 , n4103 , n4105 , n4106 , n4107 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4174 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4497 , n4498 , n4499 , n4500 , n4501 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4729 , n4730 , n4731 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4770 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4854 , n4855 , n4856 , n4857 , n4858 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5268 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5346 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5484 , n5486 , n5487 , n5488 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5734 , n5735 , n5736 , n5737 , n5738 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5865 , n5866 , n5867 , n5868 , n5869 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5994 , n5995 , n5996 , n5997 , n5998 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 ;
  assign n43 = ~x16 & x17 ;
  assign n44 = n43 ^ x16 ;
  assign n89 = n44 ^ x17 ;
  assign n45 = x18 & ~x19 ;
  assign n91 = x22 & n45 ;
  assign n138 = n89 & n91 ;
  assign n25 = ~x12 & ~x13 ;
  assign n26 = ~x6 & ~x7 ;
  assign n27 = x2 ^ x1 ;
  assign n28 = ~x0 & x1 ;
  assign n29 = n28 ^ x0 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = ~x3 & n30 ;
  assign n32 = ~x4 & n31 ;
  assign n33 = ~x5 & n32 ;
  assign n34 = n26 & n33 ;
  assign n35 = ~x8 & n34 ;
  assign n36 = ~x9 & n35 ;
  assign n37 = ~x10 & n36 ;
  assign n38 = ~x11 & n37 ;
  assign n39 = ~x14 & n38 ;
  assign n40 = n25 & n39 ;
  assign n50 = ~x15 & n40 ;
  assign n80 = n50 ^ x16 ;
  assign n81 = ~x17 & ~n80 ;
  assign n82 = n81 ^ n80 ;
  assign n65 = x19 & ~x22 ;
  assign n84 = ~x18 & n65 ;
  assign n137 = ~n82 & n84 ;
  assign n139 = n138 ^ n137 ;
  assign n41 = ~x22 & ~n40 ;
  assign n42 = n41 ^ x15 ;
  assign n46 = n45 ^ x18 ;
  assign n47 = n46 ^ x19 ;
  assign n48 = n47 ^ x18 ;
  assign n49 = ~n44 & ~n48 ;
  assign n51 = ~x22 & ~n50 ;
  assign n52 = n49 & ~n51 ;
  assign n53 = ~x22 & ~n52 ;
  assign n54 = n53 ^ x20 ;
  assign n57 = x22 ^ x21 ;
  assign n58 = n54 & ~n57 ;
  assign n59 = ~n42 & ~n58 ;
  assign n60 = n59 ^ n42 ;
  assign n564 = n139 ^ n60 ;
  assign n454 = n58 & n139 ;
  assign n61 = n60 ^ n58 ;
  assign n398 = ~n61 & n139 ;
  assign n455 = n454 ^ n398 ;
  assign n565 = n564 ^ n455 ;
  assign n85 = n84 ^ n47 ;
  assign n83 = n65 ^ x19 ;
  assign n86 = n85 ^ n83 ;
  assign n173 = n43 & n86 ;
  assign n92 = n91 ^ n45 ;
  assign n90 = n65 ^ x22 ;
  assign n93 = n92 ^ n90 ;
  assign n67 = x17 ^ x16 ;
  assign n68 = n50 ^ x17 ;
  assign n69 = ~n67 & n68 ;
  assign n141 = n80 ^ n69 ;
  assign n172 = ~n93 & n141 ;
  assign n174 = n173 ^ n172 ;
  assign n151 = ~n44 & n91 ;
  assign n66 = n50 ^ x18 ;
  assign n70 = ~x22 & n69 ;
  assign n71 = ~n66 & n70 ;
  assign n150 = x19 & n71 ;
  assign n152 = n151 ^ n150 ;
  assign n571 = n174 ^ n152 ;
  assign n99 = x21 ^ x20 ;
  assign n100 = n53 ^ x21 ;
  assign n101 = n99 & n100 ;
  assign n87 = n86 ^ n46 ;
  assign n114 = n89 ^ x16 ;
  assign n130 = ~n50 & n114 ;
  assign n131 = n87 & n130 ;
  assign n132 = n131 ^ n52 ;
  assign n94 = n93 ^ n48 ;
  assign n95 = n89 & n94 ;
  assign n88 = ~n82 & n87 ;
  assign n96 = n95 ^ n88 ;
  assign n566 = n132 ^ n96 ;
  assign n168 = n94 & n114 ;
  assign n167 = n81 & n87 ;
  assign n169 = n168 ^ n167 ;
  assign n143 = n43 & n94 ;
  assign n142 = n87 & n141 ;
  assign n144 = n143 ^ n142 ;
  assign n332 = n169 ^ n144 ;
  assign n567 = n566 ^ n332 ;
  assign n568 = n101 & n567 ;
  assign n569 = n568 ^ n101 ;
  assign n111 = n57 & ~n99 ;
  assign n112 = ~n42 & n111 ;
  assign n210 = n86 & n114 ;
  assign n209 = n81 & ~n93 ;
  assign n211 = n210 ^ n209 ;
  assign n106 = n86 & n89 ;
  assign n105 = ~n82 & ~n93 ;
  assign n107 = n106 ^ n105 ;
  assign n257 = n211 ^ n107 ;
  assign n258 = n257 ^ n174 ;
  assign n270 = n112 & ~n258 ;
  assign n570 = n569 ^ n270 ;
  assign n572 = n571 ^ n570 ;
  assign n573 = ~n565 & n572 ;
  assign n494 = ~n61 & n169 ;
  assign n245 = n58 & n169 ;
  assign n583 = n494 ^ n245 ;
  assign n241 = n43 & n85 ;
  assign n240 = n92 & n141 ;
  assign n242 = n241 ^ n240 ;
  assign n247 = ~n60 & n242 ;
  assign n115 = n85 & n114 ;
  assign n113 = n81 & n92 ;
  assign n116 = n115 ^ n113 ;
  assign n120 = ~n42 & n116 ;
  assign n119 = n59 & n116 ;
  assign n121 = n120 ^ n119 ;
  assign n248 = n247 ^ n121 ;
  assign n584 = n583 ^ n248 ;
  assign n402 = ~n61 & n144 ;
  assign n118 = n58 & n116 ;
  assign n122 = n121 ^ n118 ;
  assign n580 = n402 ^ n122 ;
  assign n579 = ~n61 & n152 ;
  assign n581 = n580 ^ n579 ;
  assign n187 = n91 & n114 ;
  assign n186 = n81 & n84 ;
  assign n188 = n187 ^ n186 ;
  assign n574 = n188 ^ n174 ;
  assign n97 = n42 & ~n57 ;
  assign n98 = n97 ^ n61 ;
  assign n102 = n101 ^ n98 ;
  assign n575 = n574 ^ n102 ;
  assign n145 = n112 ^ n111 ;
  assign n289 = ~n139 & ~n145 ;
  assign n200 = n43 & n91 ;
  assign n199 = n84 & n141 ;
  assign n201 = n200 ^ n199 ;
  assign n576 = n289 ^ n201 ;
  assign n406 = n145 & n201 ;
  assign n577 = n576 ^ n406 ;
  assign n578 = ~n575 & ~n577 ;
  assign n582 = n581 ^ n578 ;
  assign n585 = n584 ^ n582 ;
  assign n586 = ~n573 & ~n585 ;
  assign n547 = ~n42 & ~n242 ;
  assign n225 = ~n42 & n201 ;
  assign n548 = n547 ^ n225 ;
  assign n324 = ~n61 & n96 ;
  assign n552 = n324 ^ n102 ;
  assign n63 = n58 ^ n54 ;
  assign n55 = n42 & ~n54 ;
  assign n56 = n55 ^ n42 ;
  assign n62 = n61 ^ n56 ;
  assign n64 = n63 ^ n62 ;
  assign n463 = n98 ^ n64 ;
  assign n549 = n242 ^ n139 ;
  assign n550 = ~n547 & n549 ;
  assign n551 = n463 & n550 ;
  assign n553 = n552 ^ n551 ;
  assign n554 = ~n548 & ~n553 ;
  assign n385 = n56 & n96 ;
  assign n386 = n385 ^ n324 ;
  assign n146 = n144 & n145 ;
  assign n545 = n386 ^ n146 ;
  assign n76 = ~n44 & n46 ;
  assign n77 = n76 ^ n71 ;
  assign n78 = ~n65 & n77 ;
  assign n369 = n145 ^ n78 ;
  assign n368 = ~n78 & ~n145 ;
  assign n370 = n369 ^ n368 ;
  assign n292 = n101 & n169 ;
  assign n291 = ~n98 & n169 ;
  assign n293 = n292 ^ n291 ;
  assign n543 = n370 ^ n293 ;
  assign n464 = n174 & ~n463 ;
  assign n544 = n543 ^ n464 ;
  assign n546 = n545 ^ n544 ;
  assign n555 = n554 ^ n546 ;
  assign n556 = n555 ^ n64 ;
  assign n263 = ~n61 & n132 ;
  assign n561 = n263 ^ n132 ;
  assign n559 = n188 ^ n61 ;
  assign n557 = ~n98 & n188 ;
  assign n483 = n97 & n188 ;
  assign n558 = n557 ^ n483 ;
  assign n560 = n559 ^ n558 ;
  assign n562 = n561 ^ n560 ;
  assign n563 = n556 & ~n562 ;
  assign n587 = n586 ^ n563 ;
  assign n441 = n58 & n211 ;
  assign n376 = ~n61 & n211 ;
  assign n442 = n441 ^ n376 ;
  assign n522 = n442 ^ n121 ;
  assign n450 = n111 & n188 ;
  assign n374 = n188 ^ n112 ;
  assign n230 = ~n112 & ~n188 ;
  assign n375 = n374 ^ n230 ;
  assign n451 = n450 ^ n375 ;
  assign n523 = n522 ^ n451 ;
  assign n520 = n201 ^ n188 ;
  assign n521 = ~n62 & n520 ;
  assign n524 = n523 ^ n521 ;
  assign n515 = n42 & n144 ;
  assign n516 = n101 & n515 ;
  assign n157 = n85 & n89 ;
  assign n156 = ~n82 & n92 ;
  assign n158 = n157 ^ n156 ;
  assign n160 = ~n42 & n158 ;
  assign n514 = n63 & n160 ;
  assign n517 = n516 ^ n514 ;
  assign n286 = ~n61 & n107 ;
  assign n518 = n517 ^ n286 ;
  assign n509 = n102 ^ n62 ;
  assign n510 = n211 & n509 ;
  assign n234 = ~n62 & n211 ;
  assign n511 = n510 ^ n234 ;
  assign n262 = ~n60 & n132 ;
  assign n512 = n511 ^ n262 ;
  assign n507 = n78 ^ n60 ;
  assign n505 = n61 & ~n78 ;
  assign n506 = n505 ^ n58 ;
  assign n508 = n507 ^ n506 ;
  assign n513 = n512 ^ n508 ;
  assign n519 = n518 ^ n513 ;
  assign n525 = n524 ^ n519 ;
  assign n212 = ~n98 & n211 ;
  assign n134 = n98 & ~n132 ;
  assign n133 = n132 ^ n98 ;
  assign n135 = n134 ^ n133 ;
  assign n2654 = n212 ^ n135 ;
  assign n428 = ~n62 & n144 ;
  assign n2652 = n455 ^ n428 ;
  assign n389 = ~n98 & n201 ;
  assign n2653 = n2652 ^ n389 ;
  assign n2655 = n2654 ^ n2653 ;
  assign n313 = ~n42 & ~n169 ;
  assign n314 = ~n63 & n313 ;
  assign n315 = n314 ^ n313 ;
  assign n316 = n315 ^ n64 ;
  assign n312 = ~n102 & n242 ;
  assign n317 = n316 ^ n312 ;
  assign n208 = ~n61 & n201 ;
  assign n318 = n317 ^ n208 ;
  assign n205 = n111 & n169 ;
  assign n170 = n112 & n169 ;
  assign n206 = n205 ^ n170 ;
  assign n2326 = n318 ^ n206 ;
  assign n4187 = n2655 ^ n2326 ;
  assign n381 = n101 & n160 ;
  assign n109 = ~n98 & n107 ;
  assign n2463 = n381 ^ n109 ;
  assign n435 = ~n102 & n174 ;
  assign n4184 = n2463 ^ n435 ;
  assign n140 = ~n64 & n139 ;
  assign n147 = n146 ^ n140 ;
  assign n4185 = n4184 ^ n147 ;
  assign n540 = ~n64 & n242 ;
  assign n232 = n230 ^ n62 ;
  assign n231 = n62 & n230 ;
  assign n233 = n232 ^ n231 ;
  assign n3936 = n540 ^ n233 ;
  assign n154 = n112 & n144 ;
  assign n3937 = n3936 ^ n154 ;
  assign n1112 = n132 & n145 ;
  assign n4183 = n3937 ^ n1112 ;
  assign n4186 = n4185 ^ n4183 ;
  assign n4188 = n4187 ^ n4186 ;
  assign n4189 = n525 & ~n4188 ;
  assign n476 = n58 & n225 ;
  assign n161 = n58 & n160 ;
  assign n618 = n476 ^ n161 ;
  assign n124 = n112 ^ n56 ;
  assign n125 = n116 & n124 ;
  assign n117 = n112 & n116 ;
  assign n123 = n122 ^ n117 ;
  assign n126 = n125 ^ n123 ;
  assign n2370 = n618 ^ n126 ;
  assign n475 = ~n64 & n211 ;
  assign n2371 = n2370 ^ n475 ;
  assign n193 = n92 & n130 ;
  assign n191 = ~n44 & ~n51 ;
  assign n192 = n47 & n191 ;
  assign n194 = n193 ^ n192 ;
  assign n309 = n112 & n194 ;
  assign n307 = n112 ^ n60 ;
  assign n308 = n194 & ~n307 ;
  assign n310 = n309 ^ n308 ;
  assign n305 = ~n102 & n132 ;
  assign n304 = n107 & n112 ;
  assign n306 = n305 ^ n304 ;
  assign n311 = n310 ^ n306 ;
  assign n2372 = n2371 ^ n311 ;
  assign n338 = n112 & n242 ;
  assign n243 = ~n61 & n242 ;
  assign n2367 = n338 ^ n243 ;
  assign n1068 = n242 ^ n174 ;
  assign n1069 = n1068 ^ n61 ;
  assign n1070 = ~n134 & ~n1069 ;
  assign n2368 = n2367 ^ n1070 ;
  assign n380 = n145 & n158 ;
  assign n166 = n96 & ~n98 ;
  assign n1276 = n380 ^ n166 ;
  assign n153 = n112 & n152 ;
  assign n1277 = n1276 ^ n153 ;
  assign n2369 = n2368 ^ n1277 ;
  assign n2373 = n2372 ^ n2369 ;
  assign n432 = ~n98 & n116 ;
  assign n433 = n432 ^ n126 ;
  assign n181 = n119 ^ n117 ;
  assign n180 = ~n102 & n116 ;
  assign n182 = n181 ^ n180 ;
  assign n434 = n433 ^ n182 ;
  assign n436 = n435 ^ n434 ;
  assign n426 = n96 & n112 ;
  assign n178 = n96 & n111 ;
  assign n427 = n426 ^ n178 ;
  assign n429 = n428 ^ n427 ;
  assign n430 = n429 ^ n234 ;
  assign n424 = n304 ^ n170 ;
  assign n219 = n78 & ~n102 ;
  assign n425 = n424 ^ n219 ;
  assign n431 = n430 ^ n425 ;
  assign n437 = n436 ^ n431 ;
  assign n421 = ~n64 & n144 ;
  assign n297 = n112 ^ n102 ;
  assign n298 = n139 & ~n297 ;
  assign n422 = n421 ^ n298 ;
  assign n103 = n96 & ~n102 ;
  assign n420 = n370 ^ n103 ;
  assign n423 = n422 ^ n420 ;
  assign n438 = n437 ^ n423 ;
  assign n1088 = ~n368 & n438 ;
  assign n1089 = n1088 ^ n152 ;
  assign n1090 = n102 & n1089 ;
  assign n1086 = n368 ^ n152 ;
  assign n1091 = n1090 ^ n1086 ;
  assign n2374 = n2373 ^ n1091 ;
  assign n4190 = n4189 ^ n2374 ;
  assign n4191 = n587 & ~n4190 ;
  assign n1193 = n568 ^ n64 ;
  assign n2642 = n194 ^ n144 ;
  assign n2643 = ~n1193 & n2642 ;
  assign n280 = n145 & n211 ;
  assign n279 = n111 & n211 ;
  assign n281 = n280 ^ n279 ;
  assign n595 = n304 ^ n281 ;
  assign n271 = n270 ^ n112 ;
  assign n596 = n595 ^ n271 ;
  assign n295 = n112 & n139 ;
  assign n2375 = n596 ^ n295 ;
  assign n2636 = n2375 ^ n126 ;
  assign n2637 = n2636 ^ n435 ;
  assign n2638 = n2637 ^ n305 ;
  assign n384 = ~n64 & n96 ;
  assign n2634 = n384 ^ n370 ;
  assign n2635 = n2634 ^ n262 ;
  assign n2639 = n2638 ^ n2635 ;
  assign n184 = n58 & n107 ;
  assign n497 = n286 ^ n184 ;
  assign n327 = ~n98 & n194 ;
  assign n498 = n497 ^ n327 ;
  assign n159 = n58 & n158 ;
  assign n162 = n161 ^ n159 ;
  assign n495 = n494 ^ n162 ;
  assign n447 = n145 & n194 ;
  assign n496 = n495 ^ n447 ;
  assign n499 = n498 ^ n496 ;
  assign n2640 = n2639 ^ n499 ;
  assign n1180 = n242 ^ n152 ;
  assign n2632 = ~n98 & n1180 ;
  assign n2630 = n442 ^ n324 ;
  assign n2631 = n2630 ^ n182 ;
  assign n2633 = n2632 ^ n2631 ;
  assign n2641 = n2640 ^ n2633 ;
  assign n2644 = n2643 ^ n2641 ;
  assign n226 = n63 & n225 ;
  assign n831 = n514 ^ n226 ;
  assign n625 = n145 & n174 ;
  assign n832 = n831 ^ n625 ;
  assign n833 = n832 ^ n308 ;
  assign n834 = n833 ^ n386 ;
  assign n2645 = n2644 ^ n834 ;
  assign n2649 = n208 ^ n122 ;
  assign n238 = n78 & ~n98 ;
  assign n2650 = n2649 ^ n238 ;
  assign n228 = ~n62 & n139 ;
  assign n2482 = n286 ^ n228 ;
  assign n365 = n107 & n145 ;
  assign n1262 = n365 ^ n247 ;
  assign n2647 = n2482 ^ n1262 ;
  assign n624 = n174 ^ n145 ;
  assign n626 = n625 ^ n624 ;
  assign n627 = ~n560 & n626 ;
  assign n372 = n112 & n201 ;
  assign n285 = n56 & n107 ;
  assign n287 = n286 ^ n285 ;
  assign n461 = n372 ^ n287 ;
  assign n2646 = n627 ^ n461 ;
  assign n2648 = n2647 ^ n2646 ;
  assign n2651 = n2650 ^ n2648 ;
  assign n2656 = n2655 ^ n2651 ;
  assign n388 = n101 & n201 ;
  assign n390 = n389 ^ n388 ;
  assign n856 = n390 ^ n219 ;
  assign n857 = n856 ^ n312 ;
  assign n415 = ~n62 & n194 ;
  assign n414 = n56 & n194 ;
  assign n416 = n415 ^ n414 ;
  assign n223 = ~n60 & n188 ;
  assign n528 = n416 ^ n223 ;
  assign n529 = n528 ^ n375 ;
  assign n858 = n857 ^ n529 ;
  assign n203 = n62 & ~n201 ;
  assign n446 = n194 ^ n145 ;
  assign n448 = n447 ^ n446 ;
  assign n449 = ~n203 & n448 ;
  assign n853 = n449 ^ n304 ;
  assign n850 = n112 & n158 ;
  assign n851 = n850 ^ n140 ;
  assign n852 = n851 ^ n583 ;
  assign n854 = n853 ^ n852 ;
  assign n288 = n145 ^ n139 ;
  assign n290 = n289 ^ n288 ;
  assign n848 = n290 ^ n234 ;
  assign n322 = ~n98 & n174 ;
  assign n462 = n322 ^ n174 ;
  assign n465 = n464 ^ n462 ;
  assign n328 = n101 & n194 ;
  assign n329 = n328 ^ n327 ;
  assign n466 = n465 ^ n329 ;
  assign n350 = ~n98 & n152 ;
  assign n348 = n145 & n152 ;
  assign n346 = n152 ^ n101 ;
  assign n345 = ~n101 & ~n152 ;
  assign n347 = n346 ^ n345 ;
  assign n349 = n348 ^ n347 ;
  assign n351 = n350 ^ n349 ;
  assign n847 = n466 ^ n351 ;
  assign n849 = n848 ^ n847 ;
  assign n855 = n854 ^ n849 ;
  assign n859 = n858 ^ n855 ;
  assign n2657 = n2656 ^ n859 ;
  assign n2658 = n2645 & n2657 ;
  assign n325 = n324 ^ n263 ;
  assign n321 = ~n61 & n174 ;
  assign n323 = n322 ^ n321 ;
  assign n326 = n325 ^ n323 ;
  assign n330 = n329 ^ n326 ;
  assign n319 = n318 ^ n311 ;
  assign n296 = n295 ^ n290 ;
  assign n299 = n298 ^ n296 ;
  assign n294 = n293 ^ n290 ;
  assign n300 = n299 ^ n294 ;
  assign n301 = n300 ^ n219 ;
  assign n302 = n301 ^ n287 ;
  assign n283 = ~n62 & n169 ;
  assign n108 = n101 & n107 ;
  assign n110 = n109 ^ n108 ;
  assign n282 = n281 ^ n110 ;
  assign n284 = n283 ^ n282 ;
  assign n303 = n302 ^ n284 ;
  assign n320 = n319 ^ n303 ;
  assign n331 = n330 ^ n320 ;
  assign n361 = n290 ^ n161 ;
  assign n202 = n201 ^ n62 ;
  assign n204 = n203 ^ n202 ;
  assign n362 = n361 ^ n204 ;
  assign n357 = n145 & n242 ;
  assign n356 = ~n62 & n158 ;
  assign n358 = n357 ^ n356 ;
  assign n221 = n56 ^ n54 ;
  assign n353 = n194 & n221 ;
  assign n354 = n353 ^ n310 ;
  assign n355 = n354 ^ n295 ;
  assign n359 = n358 ^ n355 ;
  assign n343 = ~n102 & n188 ;
  assign n79 = ~n64 & n78 ;
  assign n344 = n343 ^ n79 ;
  assign n352 = n351 ^ n344 ;
  assign n360 = n359 ^ n352 ;
  assign n363 = n362 ^ n360 ;
  assign n340 = n162 ^ n122 ;
  assign n337 = n234 ^ n180 ;
  assign n339 = n338 ^ n337 ;
  assign n341 = n340 ^ n339 ;
  assign n334 = n107 ^ n78 ;
  assign n333 = n332 ^ n152 ;
  assign n335 = n334 ^ n333 ;
  assign n336 = ~n60 & n335 ;
  assign n342 = n341 ^ n336 ;
  assign n364 = n363 ^ n342 ;
  assign n404 = ~n102 & n144 ;
  assign n401 = n58 & n144 ;
  assign n403 = n402 ^ n401 ;
  assign n405 = n404 ^ n403 ;
  assign n407 = n406 ^ n405 ;
  assign n399 = n398 ^ n243 ;
  assign n396 = n212 ^ n103 ;
  assign n397 = n396 ^ n280 ;
  assign n400 = n399 ^ n397 ;
  assign n408 = n407 ^ n400 ;
  assign n392 = ~n62 & n174 ;
  assign n393 = n392 ^ n140 ;
  assign n387 = n386 ^ n384 ;
  assign n391 = n390 ^ n387 ;
  assign n394 = n393 ^ n391 ;
  assign n382 = n381 ^ n380 ;
  assign n377 = n376 ^ n375 ;
  assign n373 = n372 ^ n182 ;
  assign n378 = n377 ^ n373 ;
  assign n366 = n219 ^ n110 ;
  assign n367 = n366 ^ n365 ;
  assign n371 = n370 ^ n367 ;
  assign n379 = n378 ^ n371 ;
  assign n383 = n382 ^ n379 ;
  assign n395 = n394 ^ n383 ;
  assign n409 = n408 ^ n395 ;
  assign n410 = ~n364 & ~n409 ;
  assign n411 = n331 & n410 ;
  assign n912 = n475 ^ n312 ;
  assign n2544 = n912 ^ n627 ;
  assign n620 = n322 ^ n248 ;
  assign n619 = n618 ^ n393 ;
  assign n621 = n620 ^ n619 ;
  assign n2542 = n174 & n621 ;
  assign n2537 = n2367 ^ n281 ;
  assign n2538 = n2537 ^ n404 ;
  assign n2459 = n596 ^ n348 ;
  assign n2460 = n2459 ^ n380 ;
  assign n2536 = n2460 ^ n180 ;
  assign n2539 = n2538 ^ n2536 ;
  assign n265 = ~n58 & n132 ;
  assign n266 = ~n221 & n265 ;
  assign n267 = n266 ^ n132 ;
  assign n264 = n263 ^ n262 ;
  assign n268 = n267 ^ n264 ;
  assign n222 = n188 & n221 ;
  assign n224 = n223 ^ n222 ;
  assign n1255 = n268 ^ n224 ;
  assign n635 = ~n64 & n152 ;
  assign n1254 = n635 ^ n421 ;
  assign n1256 = n1255 ^ n1254 ;
  assign n527 = n291 ^ n228 ;
  assign n1257 = n1256 ^ n527 ;
  assign n2540 = n2539 ^ n1257 ;
  assign n643 = n435 ^ n309 ;
  assign n644 = n643 ^ n551 ;
  assign n2541 = n2540 ^ n644 ;
  assign n2543 = n2542 ^ n2541 ;
  assign n2545 = n2544 ^ n2543 ;
  assign n1124 = n112 & n132 ;
  assign n841 = ~n98 & n158 ;
  assign n1125 = n1124 ^ n841 ;
  assign n2472 = n1125 ^ n403 ;
  assign n1105 = n194 ^ n169 ;
  assign n1106 = ~n64 & n1105 ;
  assign n175 = ~n60 & n174 ;
  assign n1102 = n402 ^ n175 ;
  assign n1103 = n1102 ^ n510 ;
  assign n1100 = n557 ^ n398 ;
  assign n1101 = n1100 ^ n389 ;
  assign n1104 = n1103 ^ n1101 ;
  assign n1107 = n1106 ^ n1104 ;
  assign n2473 = n2472 ^ n1107 ;
  assign n1214 = n483 ^ n78 ;
  assign n1215 = n54 & n1214 ;
  assign n1212 = n415 ^ n204 ;
  assign n671 = n116 & n145 ;
  assign n885 = n671 ^ n381 ;
  assign n1210 = n885 ^ n347 ;
  assign n896 = n516 ^ n290 ;
  assign n1211 = n1210 ^ n896 ;
  assign n1213 = n1212 ^ n1211 ;
  assign n1216 = n1215 ^ n1213 ;
  assign n2595 = n2473 ^ n1216 ;
  assign n2605 = n1112 ^ n247 ;
  assign n2556 = n520 ^ n139 ;
  assign n2557 = ~n102 & n2556 ;
  assign n2558 = n2557 ^ n212 ;
  assign n2606 = n2605 ^ n2558 ;
  assign n2492 = n455 ^ n162 ;
  assign n2604 = n2492 ^ n543 ;
  assign n2607 = n2606 ^ n2604 ;
  assign n2600 = n426 ^ n329 ;
  assign n2601 = n2600 ^ n295 ;
  assign n2602 = n2601 ^ n117 ;
  assign n2598 = ~n60 & n1105 ;
  assign n2596 = n508 ^ n384 ;
  assign n2597 = n2596 ^ n327 ;
  assign n2599 = n2598 ^ n2597 ;
  assign n2603 = n2602 ^ n2599 ;
  assign n2608 = n2607 ^ n2603 ;
  assign n2609 = ~n2595 & n2608 ;
  assign n2610 = ~n2545 & n2609 ;
  assign n714 = n212 ^ n58 ;
  assign n716 = n188 ^ n116 ;
  assign n717 = n716 ^ n242 ;
  assign n718 = n101 & n717 ;
  assign n195 = n194 ^ n158 ;
  assign n196 = n101 & n195 ;
  assign n189 = n188 ^ n152 ;
  assign n190 = n58 & n189 ;
  assign n197 = n196 ^ n190 ;
  assign n715 = n389 ^ n197 ;
  assign n719 = n718 ^ n715 ;
  assign n531 = ~n78 & ~n101 ;
  assign n721 = n531 ^ n122 ;
  assign n722 = n174 ^ n58 ;
  assign n723 = n722 ^ n511 ;
  assign n724 = ~n721 & n723 ;
  assign n239 = n238 ^ n109 ;
  assign n244 = n243 ^ n239 ;
  assign n246 = n245 ^ n244 ;
  assign n249 = n248 ^ n246 ;
  assign n720 = n366 ^ n249 ;
  assign n725 = n724 ^ n720 ;
  assign n726 = ~n719 & ~n725 ;
  assign n727 = ~n714 & n726 ;
  assign n750 = ~x22 & ~n38 ;
  assign n751 = n750 ^ x12 ;
  assign n699 = n158 ^ n116 ;
  assign n700 = n699 ^ n242 ;
  assign n701 = n111 & n700 ;
  assign n653 = n78 & n112 ;
  assign n697 = n653 ^ n447 ;
  assign n251 = n62 & ~n152 ;
  assign n252 = n251 ^ n139 ;
  assign n253 = n252 ^ n228 ;
  assign n254 = ~n134 & ~n253 ;
  assign n273 = n152 ^ n139 ;
  assign n274 = n101 & n273 ;
  assign n255 = n174 ^ n78 ;
  assign n256 = n42 & n255 ;
  assign n259 = n145 & ~n258 ;
  assign n260 = ~n256 & n259 ;
  assign n261 = n260 ^ n145 ;
  assign n269 = n268 ^ n261 ;
  assign n272 = n271 ^ n269 ;
  assign n275 = n274 ^ n272 ;
  assign n276 = ~n254 & ~n275 ;
  assign n698 = n697 ^ n276 ;
  assign n702 = n701 ^ n698 ;
  assign n710 = n465 ^ n234 ;
  assign n709 = ~n62 & n242 ;
  assign n711 = n710 ^ n709 ;
  assign n708 = ~n102 & n567 ;
  assign n712 = n711 ^ n708 ;
  assign n703 = n116 ^ n107 ;
  assign n704 = n703 ^ n256 ;
  assign n705 = n63 & n704 ;
  assign n706 = n705 ^ n475 ;
  assign n707 = n706 ^ n79 ;
  assign n713 = n712 ^ n707 ;
  assign n728 = n101 & n727 ;
  assign n729 = ~n713 & n728 ;
  assign n730 = n729 ^ n713 ;
  assign n731 = n702 & ~n730 ;
  assign n740 = ~n63 & n731 ;
  assign n947 = n740 ^ n730 ;
  assign n948 = n751 & ~n947 ;
  assign n752 = ~x22 & ~n37 ;
  assign n753 = n752 ^ x11 ;
  assign n657 = n432 ^ n310 ;
  assign n658 = n657 ^ n350 ;
  assign n654 = n653 ^ n234 ;
  assign n655 = n654 ^ n208 ;
  assign n656 = n655 ^ n291 ;
  assign n659 = n658 ^ n656 ;
  assign n648 = n152 ^ n62 ;
  assign n649 = n648 ^ n251 ;
  assign n650 = n649 ^ n354 ;
  assign n646 = n514 ^ n442 ;
  assign n647 = n646 ^ n357 ;
  assign n651 = n650 ^ n647 ;
  assign n645 = n644 ^ n302 ;
  assign n652 = n651 ^ n645 ;
  assign n660 = n659 ^ n652 ;
  assign n600 = ~n58 & ~n201 ;
  assign n629 = n450 ^ n230 ;
  assign n630 = n629 ^ n111 ;
  assign n631 = n630 ^ n162 ;
  assign n632 = ~n600 & ~n631 ;
  assign n622 = n497 ^ n465 ;
  assign n623 = n622 ^ n621 ;
  assign n628 = n627 ^ n623 ;
  assign n633 = n632 ^ n628 ;
  assign n638 = n475 ^ n375 ;
  assign n639 = n638 ^ n170 ;
  assign n634 = n465 ^ n238 ;
  assign n636 = n635 ^ n634 ;
  assign n637 = n636 ^ n414 ;
  assign n640 = n639 ^ n637 ;
  assign n641 = n640 ^ n268 ;
  assign n642 = ~n633 & n641 ;
  assign n661 = n660 ^ n642 ;
  assign n685 = n225 ^ n107 ;
  assign n686 = n101 & n685 ;
  assign n681 = n356 ^ n286 ;
  assign n440 = ~n60 & n78 ;
  assign n682 = n681 ^ n440 ;
  assign n678 = n350 ^ n180 ;
  assign n679 = n678 ^ n347 ;
  assign n675 = ~n62 & n132 ;
  assign n676 = n675 ^ n508 ;
  assign n677 = n676 ^ n117 ;
  assign n680 = n679 ^ n677 ;
  assign n683 = n682 ^ n680 ;
  assign n672 = n671 ^ n281 ;
  assign n669 = n454 ^ n372 ;
  assign n670 = n669 ^ n146 ;
  assign n673 = n672 ^ n670 ;
  assign n666 = n283 ^ n280 ;
  assign n667 = n666 ^ n206 ;
  assign n663 = n376 ^ n122 ;
  assign n664 = n663 ^ n243 ;
  assign n662 = n175 ^ n154 ;
  assign n665 = n664 ^ n662 ;
  assign n668 = n667 ^ n665 ;
  assign n674 = n673 ^ n668 ;
  assign n684 = n683 ^ n674 ;
  assign n687 = n686 ^ n684 ;
  assign n688 = n661 & n687 ;
  assign n502 = n497 ^ n166 ;
  assign n503 = n502 ^ n494 ;
  assign n504 = n503 ^ n408 ;
  assign n526 = n525 ^ n275 ;
  assign n532 = n132 ^ n60 ;
  assign n533 = n532 ^ n262 ;
  assign n534 = ~n531 & ~n533 ;
  assign n535 = n534 ^ n304 ;
  assign n530 = n529 ^ n527 ;
  assign n536 = n535 ^ n530 ;
  assign n537 = n526 & n536 ;
  assign n538 = ~n504 & n537 ;
  assign n541 = n540 ^ n376 ;
  assign n539 = n309 ^ n233 ;
  assign n542 = n541 ^ n539 ;
  assign n588 = n587 ^ n542 ;
  assign n611 = n188 ^ n132 ;
  assign n612 = n58 & n611 ;
  assign n608 = n262 ^ n223 ;
  assign n609 = n608 ^ n455 ;
  assign n610 = n609 ^ n356 ;
  assign n613 = n612 ^ n610 ;
  assign n605 = n448 ^ n132 ;
  assign n606 = ~n251 & n605 ;
  assign n597 = n596 ^ n225 ;
  assign n602 = n201 ^ n158 ;
  assign n598 = n158 ^ n58 ;
  assign n599 = n598 ^ n159 ;
  assign n601 = n600 ^ n599 ;
  assign n603 = n602 ^ n601 ;
  assign n604 = ~n597 & n603 ;
  assign n607 = n606 ^ n604 ;
  assign n614 = n613 ^ n607 ;
  assign n218 = ~n60 & n96 ;
  assign n592 = n353 ^ n218 ;
  assign n591 = n290 ^ n135 ;
  assign n593 = n592 ^ n591 ;
  assign n589 = n543 ^ n153 ;
  assign n590 = n589 ^ n350 ;
  assign n594 = n593 ^ n590 ;
  assign n615 = n614 ^ n594 ;
  assign n616 = ~n588 & n615 ;
  assign n617 = n538 & n616 ;
  assign n689 = n688 ^ n617 ;
  assign n690 = ~x12 & ~x22 ;
  assign n691 = n38 & n690 ;
  assign n692 = n691 ^ x22 ;
  assign n738 = n692 ^ x13 ;
  assign n930 = n738 ^ n688 ;
  assign n933 = n731 ^ n688 ;
  assign n936 = ~n930 & n933 ;
  assign n695 = n692 ^ x14 ;
  assign n693 = x13 & ~x22 ;
  assign n694 = n692 & n693 ;
  assign n696 = n695 ^ n694 ;
  assign n732 = n731 ^ n696 ;
  assign n937 = n936 ^ n732 ;
  assign n938 = ~n689 & n937 ;
  assign n939 = n938 ^ n732 ;
  assign n942 = n939 ^ n727 ;
  assign n943 = n942 ^ n730 ;
  assign n944 = n943 ^ n939 ;
  assign n945 = n753 & ~n944 ;
  assign n946 = n945 ^ n942 ;
  assign n949 = n948 ^ n946 ;
  assign n826 = ~x22 & ~n35 ;
  assign n827 = n826 ^ x9 ;
  assign n961 = ~n727 & ~n827 ;
  assign n962 = n961 ^ n727 ;
  assign n950 = n731 ^ n617 ;
  assign n954 = n751 ^ n731 ;
  assign n957 = n950 & ~n954 ;
  assign n951 = n738 ^ n731 ;
  assign n958 = n957 ^ n951 ;
  assign n959 = ~n689 & n958 ;
  assign n960 = n959 ^ n951 ;
  assign n963 = n962 ^ n960 ;
  assign n913 = n912 ^ n405 ;
  assign n910 = n596 ^ n243 ;
  assign n911 = n910 ^ n654 ;
  assign n914 = n913 ^ n911 ;
  assign n907 = n380 ^ n322 ;
  assign n906 = n682 ^ n110 ;
  assign n908 = n907 ^ n906 ;
  assign n902 = n505 ^ n316 ;
  assign n909 = n908 ^ n902 ;
  assign n915 = n914 ^ n909 ;
  assign n903 = n169 ^ n158 ;
  assign n904 = ~n463 & ~n903 ;
  assign n905 = n902 & n904 ;
  assign n916 = n915 ^ n905 ;
  assign n897 = n896 ^ n338 ;
  assign n171 = n170 ^ n166 ;
  assign n898 = n897 ^ n171 ;
  assign n895 = n426 ^ n393 ;
  assign n899 = n898 ^ n895 ;
  assign n835 = n188 ^ n78 ;
  assign n836 = n835 ^ n144 ;
  assign n837 = ~n62 & n836 ;
  assign n900 = n899 ^ n837 ;
  assign n891 = n365 ^ n206 ;
  assign n129 = ~n64 & n107 ;
  assign n890 = n435 ^ n129 ;
  assign n892 = n891 ^ n890 ;
  assign n888 = n441 ^ n109 ;
  assign n889 = n888 ^ n649 ;
  assign n893 = n892 ^ n889 ;
  assign n884 = n841 ^ n498 ;
  assign n886 = n885 ^ n884 ;
  assign n882 = n427 ^ n421 ;
  assign n883 = n882 ^ n676 ;
  assign n887 = n886 ^ n883 ;
  assign n894 = n893 ^ n887 ;
  assign n901 = n900 ^ n894 ;
  assign n917 = n916 ^ n901 ;
  assign n918 = ~n588 & n917 ;
  assign n844 = n596 ^ n427 ;
  assign n842 = n841 ^ n432 ;
  assign n843 = n842 ^ n540 ;
  assign n845 = n844 ^ n843 ;
  assign n838 = n837 ^ n161 ;
  assign n458 = n254 ^ n146 ;
  assign n839 = n838 ^ n458 ;
  assign n840 = n839 ^ n834 ;
  assign n846 = n845 ^ n840 ;
  assign n867 = n579 ^ n140 ;
  assign n864 = ~n60 & n152 ;
  assign n865 = n864 ^ n218 ;
  assign n866 = n865 ^ n263 ;
  assign n868 = n867 ^ n866 ;
  assign n207 = n206 ^ n204 ;
  assign n869 = n868 ^ n207 ;
  assign n861 = n109 ^ n103 ;
  assign n860 = n515 ^ n174 ;
  assign n862 = n861 ^ n860 ;
  assign n863 = n101 & n862 ;
  assign n870 = n869 ^ n863 ;
  assign n875 = n145 ^ n60 ;
  assign n876 = n566 & ~n875 ;
  assign n873 = n635 ^ n494 ;
  assign n871 = n653 ^ n338 ;
  assign n872 = n871 ^ n129 ;
  assign n874 = n873 ^ n872 ;
  assign n877 = n876 ^ n874 ;
  assign n486 = n112 ^ n63 ;
  assign n485 = ~n63 & ~n112 ;
  assign n487 = n486 ^ n485 ;
  assign n488 = n487 ^ n316 ;
  assign n489 = n488 ^ n117 ;
  assign n482 = n280 ^ n126 ;
  assign n484 = n483 ^ n482 ;
  assign n490 = n489 ^ n484 ;
  assign n878 = n877 ^ n490 ;
  assign n879 = ~n870 & ~n878 ;
  assign n880 = n859 & n879 ;
  assign n881 = ~n846 & n880 ;
  assign n920 = n918 ^ n881 ;
  assign n964 = n918 ^ n688 ;
  assign n965 = n918 ^ n696 ;
  assign n966 = n964 & n965 ;
  assign n967 = n966 ^ n918 ;
  assign n968 = ~n920 & ~n967 ;
  assign n969 = n968 ^ n688 ;
  assign n970 = n969 ^ n960 ;
  assign n971 = n963 & n970 ;
  assign n972 = n971 ^ n962 ;
  assign n973 = n972 ^ n939 ;
  assign n974 = ~n949 & n973 ;
  assign n779 = ~n738 & ~n740 ;
  assign n759 = n751 ^ n740 ;
  assign n780 = n779 ^ n759 ;
  assign n828 = ~x22 & ~n36 ;
  assign n829 = n828 ^ x10 ;
  assign n1143 = n829 ^ n727 ;
  assign n991 = n829 ^ n730 ;
  assign n1144 = n1143 ^ n991 ;
  assign n781 = n780 & n1144 ;
  assign n782 = n781 ^ n759 ;
  assign n733 = n696 ^ n617 ;
  assign n734 = n732 & n733 ;
  assign n735 = n734 ^ n696 ;
  assign n736 = ~n689 & ~n735 ;
  assign n737 = n736 ^ n731 ;
  assign n825 = n782 ^ n737 ;
  assign n940 = n939 ^ n825 ;
  assign n830 = n829 ^ n827 ;
  assign n919 = n881 & n918 ;
  assign n921 = n920 ^ n919 ;
  assign n923 = n688 & ~n921 ;
  assign n922 = n921 ^ n688 ;
  assign n924 = n923 ^ n922 ;
  assign n925 = n924 ^ n827 ;
  assign n926 = n830 & n925 ;
  assign n927 = n926 ^ n829 ;
  assign n928 = n927 ^ n753 ;
  assign n929 = ~n727 & n928 ;
  assign n941 = n940 ^ n929 ;
  assign n975 = n974 ^ n941 ;
  assign n977 = n975 ^ n927 ;
  assign n978 = n825 ^ n727 ;
  assign n979 = n978 ^ n975 ;
  assign n980 = n979 ^ n753 ;
  assign n981 = ~n977 & ~n980 ;
  assign n976 = ~n825 & ~n975 ;
  assign n982 = n981 ^ n976 ;
  assign n985 = ~n727 & n982 ;
  assign n986 = n985 ^ n976 ;
  assign n987 = n986 ^ n975 ;
  assign n754 = n753 ^ n751 ;
  assign n755 = ~n727 & n754 ;
  assign n747 = ~n688 & ~n731 ;
  assign n748 = ~n617 & n747 ;
  assign n749 = n748 ^ n731 ;
  assign n757 = n755 ^ n749 ;
  assign n743 = n740 ^ n727 ;
  assign n744 = n738 & n743 ;
  assign n739 = n738 ^ n696 ;
  assign n742 = n739 & ~n947 ;
  assign n745 = n744 ^ n742 ;
  assign n746 = n745 ^ n740 ;
  assign n758 = n757 ^ n746 ;
  assign n783 = ~n758 & ~n782 ;
  assign n784 = n737 & n783 ;
  assign n809 = n784 ^ n782 ;
  assign n804 = n727 & n758 ;
  assign n805 = n782 & ~n804 ;
  assign n810 = n809 ^ n805 ;
  assign n785 = n746 & ~n757 ;
  assign n806 = n785 ^ n758 ;
  assign n807 = ~n753 & n806 ;
  assign n808 = n805 & n807 ;
  assign n811 = n810 ^ n808 ;
  assign n790 = n738 & ~n757 ;
  assign n787 = n746 & ~n782 ;
  assign n791 = n790 ^ n787 ;
  assign n792 = n737 & n791 ;
  assign n793 = n792 ^ n787 ;
  assign n794 = ~n727 & n793 ;
  assign n812 = ~n737 & ~n794 ;
  assign n820 = ~n804 & n812 ;
  assign n821 = ~n785 & n820 ;
  assign n822 = n821 ^ n785 ;
  assign n813 = n812 ^ n794 ;
  assign n814 = n813 ^ n785 ;
  assign n823 = n822 ^ n814 ;
  assign n824 = ~n811 & ~n823 ;
  assign n988 = n987 ^ n824 ;
  assign n1152 = n969 ^ n963 ;
  assign n1145 = n727 & n753 ;
  assign n1146 = n1145 ^ n991 ;
  assign n1147 = n1144 & ~n1146 ;
  assign n1148 = n1147 ^ n991 ;
  assign n1149 = n743 & ~n1148 ;
  assign n1019 = ~x6 & ~x22 ;
  assign n1020 = n33 & n1019 ;
  assign n1018 = x22 ^ x7 ;
  assign n1021 = n1020 ^ n1018 ;
  assign n1016 = ~x22 & ~n34 ;
  assign n1017 = n1016 ^ x8 ;
  assign n1022 = n1021 ^ n1017 ;
  assign n1063 = n376 ^ n110 ;
  assign n1062 = n865 ^ n416 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1059 = n435 ^ n380 ;
  assign n213 = n212 ^ n208 ;
  assign n1060 = n1059 ^ n213 ;
  assign n1056 = n403 ^ n103 ;
  assign n1057 = n1056 ^ n675 ;
  assign n1058 = n1057 ^ n129 ;
  assign n1061 = n1060 ^ n1058 ;
  assign n1065 = n1064 ^ n1061 ;
  assign n443 = n442 ^ n440 ;
  assign n444 = n443 ^ n175 ;
  assign n1053 = n444 ^ n285 ;
  assign n1054 = n1053 ^ n375 ;
  assign n1049 = n850 ^ n404 ;
  assign n1050 = n1049 ^ n447 ;
  assign n1051 = n1050 ^ n475 ;
  assign n1048 = n508 ^ n308 ;
  assign n1052 = n1051 ^ n1048 ;
  assign n1055 = n1054 ^ n1052 ;
  assign n1066 = n1065 ^ n1055 ;
  assign n1028 = n350 ^ n204 ;
  assign n1029 = n1028 ^ n119 ;
  assign n1025 = n618 ^ n514 ;
  assign n1023 = n281 ^ n268 ;
  assign n1024 = n1023 ^ n381 ;
  assign n1026 = n1025 ^ n1024 ;
  assign n1027 = n1026 ^ n582 ;
  assign n1030 = n1029 ^ n1027 ;
  assign n1043 = n343 ^ n135 ;
  assign n1042 = n338 ^ n322 ;
  assign n1044 = n1043 ^ n1042 ;
  assign n1039 = n357 ^ n280 ;
  assign n1040 = n1039 ^ n497 ;
  assign n1038 = n329 ^ n316 ;
  assign n1041 = n1040 ^ n1038 ;
  assign n1045 = n1044 ^ n1041 ;
  assign n1036 = ~n62 & n699 ;
  assign n1032 = ~n64 & n189 ;
  assign n1033 = n1032 ^ n283 ;
  assign n1034 = n1033 ^ n291 ;
  assign n1031 = n857 ^ n321 ;
  assign n1035 = n1034 ^ n1031 ;
  assign n1037 = n1036 ^ n1035 ;
  assign n1046 = n1045 ^ n1037 ;
  assign n1047 = ~n1030 & n1046 ;
  assign n1067 = n1066 ^ n1047 ;
  assign n1071 = n1051 ^ n667 ;
  assign n1078 = n494 ^ n160 ;
  assign n1077 = n286 ^ n140 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1080 = n1079 ^ n343 ;
  assign n1075 = n281 ^ n170 ;
  assign n1073 = n328 ^ n243 ;
  assign n1072 = n558 ^ n540 ;
  assign n1074 = n1073 ^ n1072 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1081 = n1080 ^ n1076 ;
  assign n1082 = ~n1071 & ~n1081 ;
  assign n1083 = n1082 ^ n1070 ;
  assign n1092 = n1091 ^ n1083 ;
  assign n1130 = n154 ^ n98 ;
  assign n1131 = n152 ^ n116 ;
  assign n1132 = n1131 ^ n144 ;
  assign n1133 = ~n1130 & n1132 ;
  assign n1126 = n1125 ^ n426 ;
  assign n1122 = n625 ^ n376 ;
  assign n1123 = n1122 ^ n182 ;
  assign n1127 = n1126 ^ n1123 ;
  assign n1118 = n579 ^ n321 ;
  assign n1119 = n1118 ^ n309 ;
  assign n1117 = n649 ^ n384 ;
  assign n1120 = n1119 ^ n1117 ;
  assign n1121 = n1120 ^ n213 ;
  assign n1128 = n1127 ^ n1121 ;
  assign n1109 = n653 ^ n180 ;
  assign n1110 = n1109 ^ n386 ;
  assign n1113 = n1112 ^ n218 ;
  assign n1111 = n653 ^ n312 ;
  assign n1114 = n1113 ^ n1111 ;
  assign n1115 = ~n1110 & ~n1114 ;
  assign n1097 = n671 ^ n524 ;
  assign n1096 = n238 ^ n79 ;
  assign n1098 = n1097 ^ n1096 ;
  assign n1093 = n375 ^ n146 ;
  assign n136 = n135 ^ n129 ;
  assign n1094 = n1093 ^ n136 ;
  assign n1095 = n1094 ^ n622 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1108 = n1107 ^ n1099 ;
  assign n1116 = n1115 ^ n1108 ;
  assign n1129 = n1128 ^ n1116 ;
  assign n1134 = n1133 ^ n1129 ;
  assign n1135 = ~n1092 & n1134 ;
  assign n1136 = ~n881 & ~n1135 ;
  assign n1137 = n1067 & n1136 ;
  assign n1138 = n1137 ^ n881 ;
  assign n1139 = n1138 ^ n1021 ;
  assign n1140 = ~n1022 & ~n1139 ;
  assign n1141 = n1140 ^ n1021 ;
  assign n1142 = ~n727 & ~n1141 ;
  assign n1150 = n1149 ^ n1142 ;
  assign n999 = n696 ^ n688 ;
  assign n1000 = n920 & n999 ;
  assign n996 = ~n688 & n919 ;
  assign n997 = n996 ^ n923 ;
  assign n998 = n930 & n997 ;
  assign n1001 = n1000 ^ n998 ;
  assign n1002 = n1001 ^ n961 ;
  assign n993 = n730 & n830 ;
  assign n994 = n993 ^ n829 ;
  assign n995 = ~n740 & n994 ;
  assign n1003 = n1002 ^ n995 ;
  assign n1006 = n753 ^ n731 ;
  assign n1009 = n933 & ~n1006 ;
  assign n1010 = n1009 ^ n954 ;
  assign n1011 = ~n689 & ~n1010 ;
  assign n1012 = n1011 ^ n954 ;
  assign n1013 = n1012 ^ n1001 ;
  assign n1014 = n1003 & ~n1013 ;
  assign n1015 = n1014 ^ n1001 ;
  assign n1151 = n1150 ^ n1015 ;
  assign n1153 = n1152 ^ n1151 ;
  assign n1174 = ~n727 & ~n1022 ;
  assign n1158 = ~n727 & ~n1021 ;
  assign n1156 = n920 & n930 ;
  assign n1154 = n751 ^ n688 ;
  assign n1155 = n997 & ~n1154 ;
  assign n1157 = n1156 ^ n1155 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1160 = n1135 ^ n1067 ;
  assign n1163 = n1067 ^ n881 ;
  assign n1164 = n881 ^ n696 ;
  assign n1167 = ~n1163 & ~n1164 ;
  assign n1168 = n1167 ^ n1067 ;
  assign n1169 = n1160 & n1168 ;
  assign n1161 = n1158 ^ n881 ;
  assign n1170 = n1169 ^ n1161 ;
  assign n1171 = ~n1159 & n1170 ;
  assign n1172 = n1171 ^ n1158 ;
  assign n1173 = n1172 ^ n1138 ;
  assign n1175 = n1174 ^ n1173 ;
  assign n1294 = n829 ^ n688 ;
  assign n1295 = n1294 ^ n1006 ;
  assign n1296 = n1295 ^ n1006 ;
  assign n1297 = n829 ^ n731 ;
  assign n1300 = n1296 & ~n1297 ;
  assign n1301 = n1300 ^ n1006 ;
  assign n1302 = ~n689 & ~n1301 ;
  assign n1303 = n1302 ^ n1006 ;
  assign n1176 = ~x22 & ~n33 ;
  assign n1177 = n1176 ^ x6 ;
  assign n1178 = ~n727 & n1177 ;
  assign n1194 = n144 & ~n1193 ;
  assign n1190 = n1112 ^ n447 ;
  assign n1189 = n263 ^ n233 ;
  assign n1191 = n1190 ^ n1189 ;
  assign n1192 = n1191 ^ n286 ;
  assign n1195 = n1194 ^ n1192 ;
  assign n1196 = n476 ^ n380 ;
  assign n1197 = n1196 ^ n515 ;
  assign n1198 = n1197 ^ n219 ;
  assign n1199 = n1198 ^ n673 ;
  assign n1200 = n1199 ^ n1094 ;
  assign n1201 = n1195 & n1200 ;
  assign n1179 = n554 ^ n63 ;
  assign n1185 = ~n221 & n1180 ;
  assign n1186 = n1185 ^ n116 ;
  assign n1187 = n1179 & n1186 ;
  assign n1188 = n1187 ^ n625 ;
  assign n1202 = n1201 ^ n1188 ;
  assign n1205 = n174 ^ n169 ;
  assign n1206 = n1205 ^ n195 ;
  assign n1207 = ~n98 & n1206 ;
  assign n1203 = n583 ^ n579 ;
  assign n1204 = n1203 ^ n153 ;
  assign n1208 = n1207 ^ n1204 ;
  assign n1209 = ~n1125 & ~n1208 ;
  assign n1217 = n1216 ^ n1209 ;
  assign n1224 = n647 ^ n394 ;
  assign n1225 = n1224 ^ n1064 ;
  assign n1220 = n435 ^ n293 ;
  assign n1221 = n1220 ^ n154 ;
  assign n1222 = n1221 ^ n234 ;
  assign n1218 = n508 ^ n304 ;
  assign n1219 = n1218 ^ n1043 ;
  assign n1223 = n1222 ^ n1219 ;
  assign n1226 = n1225 ^ n1223 ;
  assign n1227 = n1217 & ~n1226 ;
  assign n1228 = n1202 & n1227 ;
  assign n1229 = n1135 & n1228 ;
  assign n1230 = ~n1178 & ~n1229 ;
  assign n235 = n234 ^ n233 ;
  assign n1231 = n334 ^ n235 ;
  assign n1246 = n1131 ^ n611 ;
  assign n1248 = n145 & ~n1246 ;
  assign n1243 = ~n102 & n602 ;
  assign n1240 = n427 ^ n325 ;
  assign n1241 = n1240 ^ n512 ;
  assign n1242 = n1241 ^ n1109 ;
  assign n1244 = n1243 ^ n1242 ;
  assign n1237 = n289 & ~n1131 ;
  assign n1238 = n55 & ~n1237 ;
  assign n1234 = n1124 ^ n426 ;
  assign n1232 = n328 ^ n108 ;
  assign n1233 = n1232 ^ n375 ;
  assign n1235 = n1234 ^ n1233 ;
  assign n1236 = n1235 ^ n1042 ;
  assign n1239 = n1238 ^ n1236 ;
  assign n1245 = n1244 ^ n1239 ;
  assign n1249 = n1248 ^ n1245 ;
  assign n1259 = ~n60 & ~n1237 ;
  assign n1250 = n540 ^ n465 ;
  assign n1251 = n1250 ^ n384 ;
  assign n1252 = n1251 ^ n618 ;
  assign n1253 = n1252 ^ n494 ;
  assign n1258 = n1257 ^ n1253 ;
  assign n1260 = n1259 ^ n1258 ;
  assign n1261 = n1249 & ~n1260 ;
  assign n1283 = ~n485 & n1261 ;
  assign n1284 = ~n1231 & n1283 ;
  assign n1268 = n1100 ^ n441 ;
  assign n1269 = n1268 ^ n175 ;
  assign n1266 = n305 ^ n295 ;
  assign n1265 = n356 ^ n316 ;
  assign n1267 = n1266 ^ n1265 ;
  assign n1270 = n1269 ^ n1267 ;
  assign n1263 = n1119 ^ n528 ;
  assign n1264 = n1263 ^ n1262 ;
  assign n1271 = n1270 ^ n1264 ;
  assign n1274 = n841 ^ n516 ;
  assign n1272 = n376 ^ n208 ;
  assign n1273 = n1272 ^ n508 ;
  assign n1275 = n1274 ^ n1273 ;
  assign n1278 = n1277 ^ n1275 ;
  assign n1279 = n1271 & ~n1278 ;
  assign n1280 = n1279 ^ n1188 ;
  assign n1281 = n1280 ^ n1261 ;
  assign n1285 = n1284 ^ n1281 ;
  assign n1290 = ~n1135 & ~n1285 ;
  assign n1287 = n1285 ^ n1228 ;
  assign n1286 = ~n1228 & n1285 ;
  assign n1288 = n1287 ^ n1286 ;
  assign n1289 = ~n1135 & n1288 ;
  assign n1291 = n1290 ^ n1289 ;
  assign n1292 = n1230 & ~n1291 ;
  assign n1293 = n1292 ^ n1291 ;
  assign n1304 = n1303 ^ n1293 ;
  assign n1305 = n1017 ^ n740 ;
  assign n1316 = n1305 ^ n1293 ;
  assign n1306 = n1305 ^ n1144 ;
  assign n1307 = n1306 ^ n1017 ;
  assign n1313 = ~n827 & n1307 ;
  assign n1314 = n1313 ^ n1017 ;
  assign n1315 = n1144 & ~n1314 ;
  assign n1317 = n1316 ^ n1315 ;
  assign n1318 = n1304 & n1317 ;
  assign n1319 = n1318 ^ n1303 ;
  assign n1320 = n1319 ^ n1172 ;
  assign n1321 = ~n1175 & n1320 ;
  assign n1322 = n1321 ^ n1172 ;
  assign n1323 = n1322 ^ n1151 ;
  assign n1324 = ~n1153 & ~n1323 ;
  assign n1325 = n1324 ^ n1151 ;
  assign n1326 = n972 ^ n949 ;
  assign n1327 = n1142 ^ n1015 ;
  assign n1328 = ~n1150 & n1327 ;
  assign n1329 = n1328 ^ n1015 ;
  assign n1330 = n1329 ^ n1326 ;
  assign n1331 = ~n727 & n830 ;
  assign n1332 = n1331 ^ n924 ;
  assign n1333 = n1332 ^ n1329 ;
  assign n1334 = ~n1330 & n1333 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1336 = ~n1326 & n1335 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1338 = ~n1325 & n1337 ;
  assign n1339 = n1334 ^ n1326 ;
  assign n1340 = ~n1325 & ~n1336 ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1344 = n1317 ^ n1303 ;
  assign n1343 = n1170 ^ n1157 ;
  assign n1345 = n1344 ^ n1343 ;
  assign n1353 = n1135 ^ n881 ;
  assign n1356 = n881 ^ n738 ;
  assign n1359 = n1353 & n1356 ;
  assign n1360 = n1359 ^ n1164 ;
  assign n1361 = n1160 & n1360 ;
  assign n1362 = n1361 ^ n1164 ;
  assign n1346 = n1021 ^ n730 ;
  assign n1347 = n1346 ^ n1017 ;
  assign n1350 = ~n1144 & n1347 ;
  assign n1351 = n1350 ^ n1017 ;
  assign n1352 = n743 & n1351 ;
  assign n1363 = n1362 ^ n1352 ;
  assign n1364 = n827 ^ n731 ;
  assign n1369 = n950 & ~n1364 ;
  assign n1370 = n1369 ^ n1297 ;
  assign n1371 = ~n689 & ~n1370 ;
  assign n1372 = n1371 ^ n1297 ;
  assign n1373 = n1372 ^ n1362 ;
  assign n1374 = n1363 & ~n1373 ;
  assign n1375 = n1374 ^ n1362 ;
  assign n1376 = n1375 ^ n1343 ;
  assign n1377 = n1345 & ~n1376 ;
  assign n1378 = n1377 ^ n1344 ;
  assign n1342 = n1012 ^ n1003 ;
  assign n1380 = n1378 ^ n1342 ;
  assign n1379 = n1342 & ~n1378 ;
  assign n1381 = n1380 ^ n1379 ;
  assign n2227 = n1319 ^ n1175 ;
  assign n2198 = n1375 ^ n1345 ;
  assign n2182 = n920 & ~n1154 ;
  assign n2087 = n753 ^ n688 ;
  assign n2181 = n997 & ~n2087 ;
  assign n2183 = n2182 ^ n2181 ;
  assign n2184 = n2183 ^ n1178 ;
  assign n1530 = n1291 ^ n1229 ;
  assign n1528 = n1228 ^ n1135 ;
  assign n1529 = n1528 ^ n1286 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n2112 = n1531 ^ n1288 ;
  assign n2113 = ~n696 & ~n2112 ;
  assign n1580 = ~x22 & ~n32 ;
  assign n1581 = n1580 ^ x5 ;
  assign n2109 = n1581 ^ n727 ;
  assign n2001 = n727 & ~n1581 ;
  assign n2110 = n2109 ^ n2001 ;
  assign n2191 = ~n1530 & n2110 ;
  assign n2192 = n2191 ^ n1228 ;
  assign n2193 = ~n2113 & ~n2192 ;
  assign n2185 = n1229 ^ n1228 ;
  assign n2194 = n2193 ^ n2185 ;
  assign n2195 = n2194 ^ n2183 ;
  assign n2196 = ~n2184 & n2195 ;
  assign n2197 = n2196 ^ n1293 ;
  assign n2199 = n2198 ^ n2197 ;
  assign n2044 = n881 ^ n751 ;
  assign n2096 = n1353 & ~n2044 ;
  assign n2097 = n2096 ^ n1356 ;
  assign n2098 = n1160 & n2097 ;
  assign n2088 = n920 & ~n2087 ;
  assign n2086 = n997 & ~n1294 ;
  assign n2089 = n2088 ^ n2086 ;
  assign n2090 = n2089 ^ n1356 ;
  assign n2099 = n2098 ^ n2090 ;
  assign n2055 = n1017 ^ n731 ;
  assign n2104 = n950 & ~n2055 ;
  assign n2105 = n2104 ^ n1364 ;
  assign n2106 = ~n689 & ~n2105 ;
  assign n2107 = n2106 ^ n1364 ;
  assign n2167 = n2107 ^ n2089 ;
  assign n2168 = n2099 & ~n2167 ;
  assign n2169 = n2168 ^ n2089 ;
  assign n2166 = n1372 ^ n1363 ;
  assign n2170 = n2169 ^ n2166 ;
  assign n1387 = n881 ^ n753 ;
  assign n2051 = n1353 & ~n1387 ;
  assign n2052 = n2051 ^ n2044 ;
  assign n2053 = n1160 & ~n2052 ;
  assign n2042 = n920 & ~n1294 ;
  assign n1384 = n827 ^ n688 ;
  assign n2041 = n997 & ~n1384 ;
  assign n2043 = n2042 ^ n2041 ;
  assign n2045 = n2044 ^ n2043 ;
  assign n2054 = n2053 ^ n2045 ;
  assign n2118 = ~n947 & ~n1021 ;
  assign n2117 = ~n1144 & n1177 ;
  assign n2119 = n2118 ^ n2117 ;
  assign n2120 = n2119 ^ n727 ;
  assign n2122 = n2120 ^ n2043 ;
  assign n1620 = n1021 ^ n688 ;
  assign n2060 = n950 & ~n1620 ;
  assign n2061 = n2060 ^ n2055 ;
  assign n2062 = ~n689 & ~n2061 ;
  assign n2063 = n2062 ^ n2055 ;
  assign n2121 = n2120 ^ n2063 ;
  assign n2123 = n2122 ^ n2121 ;
  assign n2124 = n2054 & ~n2123 ;
  assign n2125 = n2124 ^ n2121 ;
  assign n1482 = ~x22 & ~n31 ;
  assign n1483 = n1482 ^ x4 ;
  assign n1999 = ~n727 & ~n1483 ;
  assign n2039 = n1999 ^ n727 ;
  assign n2126 = n2039 ^ n1228 ;
  assign n1572 = n1228 ^ n738 ;
  assign n1414 = n1285 ^ n1135 ;
  assign n2127 = n1287 & ~n1414 ;
  assign n2128 = ~n1572 & n2127 ;
  assign n2129 = n2128 ^ n1228 ;
  assign n2130 = n2129 ^ n2039 ;
  assign n2032 = n1528 ^ n696 ;
  assign n2033 = n2032 ^ n1285 ;
  assign n2034 = n2033 ^ n739 ;
  assign n2035 = ~n1528 & ~n2034 ;
  assign n2036 = n2035 ^ n739 ;
  assign n2037 = n1287 & n2036 ;
  assign n2038 = n2037 ^ n2032 ;
  assign n2040 = n2039 ^ n2038 ;
  assign n2131 = n2129 ^ n1285 ;
  assign n2134 = ~n2040 & ~n2131 ;
  assign n2135 = n2130 & n2134 ;
  assign n2136 = n2135 ^ n2130 ;
  assign n2137 = n2136 ^ n2039 ;
  assign n2138 = n2126 & ~n2137 ;
  assign n2139 = n2138 ^ n1228 ;
  assign n2171 = n2139 ^ n2120 ;
  assign n2172 = n2125 & n2171 ;
  assign n2173 = n2172 ^ n2120 ;
  assign n2178 = n2173 ^ n2169 ;
  assign n2179 = n2170 & ~n2178 ;
  assign n2180 = n2179 ^ n2173 ;
  assign n2224 = n2197 ^ n2180 ;
  assign n2225 = n2199 & ~n2224 ;
  assign n2226 = n2225 ^ n2197 ;
  assign n2228 = n2227 ^ n2226 ;
  assign n2174 = n2173 ^ n2170 ;
  assign n2140 = n2139 ^ n2125 ;
  assign n2114 = ~n1530 & ~n2113 ;
  assign n2108 = n2107 ^ n2099 ;
  assign n2111 = n2110 ^ n2108 ;
  assign n2115 = n2114 ^ n2111 ;
  assign n2076 = ~n947 & n1177 ;
  assign n2075 = ~n1144 & n1581 ;
  assign n2077 = n2076 ^ n2075 ;
  assign n2078 = n2077 ^ n727 ;
  assign n1390 = n881 ^ n829 ;
  assign n1395 = n1353 & ~n1390 ;
  assign n1396 = n1395 ^ n1387 ;
  assign n1397 = n1160 & ~n1396 ;
  assign n1385 = n920 & ~n1384 ;
  assign n1382 = n1017 ^ n688 ;
  assign n1383 = n997 & ~n1382 ;
  assign n1386 = n1385 ^ n1383 ;
  assign n1388 = n1387 ^ n1386 ;
  assign n1398 = n1397 ^ n1388 ;
  assign n1402 = n1177 ^ n688 ;
  assign n1405 = n933 & n1402 ;
  assign n1399 = n1021 ^ n731 ;
  assign n1406 = n1405 ^ n1399 ;
  assign n1407 = ~n689 & n1406 ;
  assign n1408 = n1407 ^ n1399 ;
  assign n2072 = n1408 ^ n1386 ;
  assign n2073 = n1398 & n2072 ;
  assign n2074 = n2073 ^ n1408 ;
  assign n2079 = n2078 ^ n2074 ;
  assign n473 = n166 ^ n154 ;
  assign n1430 = n1274 ^ n473 ;
  assign n1429 = n398 ^ n337 ;
  assign n1431 = n1430 ^ n1429 ;
  assign n1432 = n1431 ^ n639 ;
  assign n1425 = n514 ^ n291 ;
  assign n1426 = n1425 ^ n540 ;
  assign n1424 = n145 & n835 ;
  assign n1427 = n1426 ^ n1424 ;
  assign n1422 = n485 ^ n98 ;
  assign n1423 = n132 & n1422 ;
  assign n1428 = n1427 ^ n1423 ;
  assign n1433 = n1432 ^ n1428 ;
  assign n1451 = n649 ^ n228 ;
  assign n1452 = n1451 ^ n596 ;
  assign n1453 = n1452 ^ n249 ;
  assign n1434 = n139 ^ n78 ;
  assign n1443 = ~n42 & ~n1434 ;
  assign n1435 = n1434 ^ n152 ;
  assign n1437 = n1435 ^ n111 ;
  assign n1436 = n1435 ^ n42 ;
  assign n1438 = n1437 ^ n1436 ;
  assign n1444 = n1443 ^ n1438 ;
  assign n1447 = n1443 ^ n42 ;
  assign n1448 = ~n58 & ~n1447 ;
  assign n1449 = n1448 ^ n1435 ;
  assign n1450 = ~n1444 & n1449 ;
  assign n1454 = n1453 ^ n1450 ;
  assign n1455 = n1433 & ~n1454 ;
  assign n1421 = n426 ^ n331 ;
  assign n1456 = n1455 ^ n1421 ;
  assign n1457 = ~n696 & ~n1228 ;
  assign n1458 = ~n1456 & n1457 ;
  assign n1459 = n1458 ^ n1228 ;
  assign n2082 = n2078 ^ n1459 ;
  assign n1460 = x22 ^ x2 ;
  assign n1461 = ~x1 & n1460 ;
  assign n1462 = ~x22 & n1461 ;
  assign n1463 = n1462 ^ n1460 ;
  assign n1466 = n1463 ^ x22 ;
  assign n1464 = n29 & n1463 ;
  assign n1465 = n1464 ^ n30 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1468 = n1467 ^ x3 ;
  assign n1469 = ~n727 & ~n1468 ;
  assign n1470 = n1469 ^ n1459 ;
  assign n1410 = n1135 ^ n751 ;
  assign n1417 = ~n1410 & ~n1414 ;
  assign n1411 = n1135 ^ n738 ;
  assign n1418 = n1417 ^ n1411 ;
  assign n1419 = n1287 & n1418 ;
  assign n1420 = n1419 ^ n1411 ;
  assign n2080 = n1459 ^ n1420 ;
  assign n2081 = ~n1470 & ~n2080 ;
  assign n2083 = n2082 ^ n2081 ;
  assign n2084 = ~n2079 & n2083 ;
  assign n2085 = n2084 ^ n2078 ;
  assign n2116 = n2115 ^ n2085 ;
  assign n2141 = n2140 ^ n2116 ;
  assign n2064 = n2063 ^ n2054 ;
  assign n2065 = n2064 ^ n2040 ;
  assign n1476 = ~n738 & ~n1228 ;
  assign n1477 = n1476 ^ n696 ;
  assign n1478 = ~n1456 & ~n1477 ;
  assign n1474 = n1228 ^ n696 ;
  assign n1479 = n1478 ^ n1474 ;
  assign n2007 = ~n727 & n1479 ;
  assign n2000 = n1999 ^ n740 ;
  assign n2002 = n2001 ^ n1483 ;
  assign n2004 = ~n730 & ~n2002 ;
  assign n2005 = n2004 ^ n1483 ;
  assign n2006 = ~n2000 & n2005 ;
  assign n2008 = n2007 ^ n2006 ;
  assign n1970 = n920 & ~n1382 ;
  assign n1969 = n997 & n1620 ;
  assign n1971 = n1970 ^ n1969 ;
  assign n1972 = n1971 ^ n1390 ;
  assign n1623 = n881 ^ n827 ;
  assign n1966 = n1353 & ~n1623 ;
  assign n1967 = n1966 ^ n1390 ;
  assign n1968 = n1160 & ~n1967 ;
  assign n1973 = n1972 ^ n1968 ;
  assign n1582 = n1581 ^ n731 ;
  assign n1979 = n950 & ~n1582 ;
  assign n1974 = n1177 ^ n731 ;
  assign n1980 = n1979 ^ n1974 ;
  assign n1981 = ~n689 & ~n1980 ;
  assign n1982 = n1981 ^ n1974 ;
  assign n1996 = n1982 ^ n1971 ;
  assign n1997 = n1973 & ~n1996 ;
  assign n1998 = n1997 ^ n1982 ;
  assign n2066 = n2007 ^ n1998 ;
  assign n2067 = n2008 & ~n2066 ;
  assign n2068 = n2067 ^ n2007 ;
  assign n2069 = n2068 ^ n2040 ;
  assign n2070 = n2065 & ~n2069 ;
  assign n2071 = n2070 ^ n2064 ;
  assign n2142 = n2141 ^ n2071 ;
  assign n1471 = n1470 ^ n1420 ;
  assign n1409 = n1408 ^ n1398 ;
  assign n1472 = n1471 ^ n1409 ;
  assign n1484 = n1483 ^ n1468 ;
  assign n1490 = ~n1144 & n1484 ;
  assign n1485 = n1483 ^ n730 ;
  assign n1491 = n1490 ^ n1485 ;
  assign n1492 = n743 & n1491 ;
  assign n1480 = n1479 ^ n727 ;
  assign n1493 = n1492 ^ n1480 ;
  assign n1494 = n1135 ^ n753 ;
  assign n1499 = ~n1414 & ~n1494 ;
  assign n1500 = n1499 ^ n1410 ;
  assign n1501 = n1287 & ~n1500 ;
  assign n1502 = n1501 ^ n1410 ;
  assign n1503 = n1502 ^ n1480 ;
  assign n1504 = ~n1493 & n1503 ;
  assign n1481 = n1480 ^ n1471 ;
  assign n1505 = n1504 ^ n1481 ;
  assign n1506 = n1472 & n1505 ;
  assign n1507 = n1506 ^ n1471 ;
  assign n1614 = n920 & ~n1402 ;
  assign n1612 = n1581 ^ n688 ;
  assign n1613 = n997 & ~n1612 ;
  assign n1615 = n1614 ^ n1613 ;
  assign n1546 = n1021 ^ n881 ;
  assign n1606 = n1353 & n1546 ;
  assign n1601 = n1017 ^ n881 ;
  assign n1607 = n1606 ^ n1601 ;
  assign n1608 = n1160 & ~n1607 ;
  assign n1609 = n1608 ^ n1601 ;
  assign n1563 = n1135 ^ n829 ;
  assign n1610 = n1609 ^ n1563 ;
  assign n1534 = n1135 ^ n827 ;
  assign n1598 = ~n1414 & ~n1534 ;
  assign n1599 = n1598 ^ n1563 ;
  assign n1600 = n1287 & ~n1599 ;
  assign n1611 = n1610 ^ n1600 ;
  assign n1907 = n1615 ^ n1611 ;
  assign n1657 = n1483 ^ n688 ;
  assign n1678 = n920 & ~n1657 ;
  assign n1677 = n997 & ~n1468 ;
  assign n1679 = n1678 ^ n1677 ;
  assign n1680 = n1679 ^ n996 ;
  assign n1527 = n1135 ^ n1017 ;
  assign n1673 = ~n1287 & ~n1527 ;
  assign n1671 = n1135 ^ n1021 ;
  assign n1672 = n1671 & n2127 ;
  assign n1674 = n1673 ^ n1672 ;
  assign n1549 = n1177 ^ n881 ;
  assign n1675 = n1674 ^ n1549 ;
  assign n1663 = n1581 ^ n881 ;
  assign n1668 = n1353 & ~n1663 ;
  assign n1669 = n1668 ^ n1549 ;
  assign n1670 = n1160 & ~n1669 ;
  assign n1676 = n1675 ^ n1670 ;
  assign n1685 = n1680 ^ n1676 ;
  assign n1651 = n827 & ~n1228 ;
  assign n1652 = n1651 ^ n829 ;
  assign n1653 = ~n1456 & n1652 ;
  assign n1649 = n1228 ^ n829 ;
  assign n1654 = n1653 ^ n1649 ;
  assign n1646 = n924 & ~n996 ;
  assign n1647 = n1468 & n1646 ;
  assign n1648 = n1647 ^ n996 ;
  assign n1686 = n1654 ^ n1648 ;
  assign n1687 = ~n1685 & ~n1686 ;
  assign n1681 = n1680 ^ n1674 ;
  assign n1682 = ~n1676 & n1681 ;
  assign n1683 = n1682 ^ n1674 ;
  assign n1659 = n920 & ~n1612 ;
  assign n1658 = n997 & ~n1657 ;
  assign n1660 = n1659 ^ n1658 ;
  assign n1516 = n689 & ~n1468 ;
  assign n1661 = n1660 ^ n1516 ;
  assign n1655 = n1648 & ~n1654 ;
  assign n1552 = n1353 & ~n1549 ;
  assign n1553 = n1552 ^ n1546 ;
  assign n1554 = n1160 & n1553 ;
  assign n1555 = n1554 ^ n1546 ;
  assign n1541 = n829 & ~n1228 ;
  assign n1542 = n1541 ^ n753 ;
  assign n1543 = ~n1456 & n1542 ;
  assign n1539 = n1228 ^ n753 ;
  assign n1544 = n1543 ^ n1539 ;
  assign n1535 = ~n1287 & ~n1534 ;
  assign n1533 = ~n1527 & n2127 ;
  assign n1536 = n1535 ^ n1533 ;
  assign n1545 = n1544 ^ n1536 ;
  assign n1645 = n1555 ^ n1545 ;
  assign n1656 = n1655 ^ n1645 ;
  assign n1662 = n1661 ^ n1656 ;
  assign n1684 = n1683 ^ n1662 ;
  assign n1688 = n1687 ^ n1684 ;
  assign n1698 = ~n1287 & n1671 ;
  assign n1696 = n1177 ^ n1135 ;
  assign n1697 = ~n1696 & n2127 ;
  assign n1699 = n1698 ^ n1697 ;
  assign n1692 = n1017 & ~n1228 ;
  assign n1693 = n1692 ^ n827 ;
  assign n1694 = ~n1456 & n1693 ;
  assign n1690 = n1228 ^ n827 ;
  assign n1695 = n1694 ^ n1690 ;
  assign n1700 = n1699 ^ n1695 ;
  assign n1703 = n1483 ^ n881 ;
  assign n1708 = n1353 & ~n1703 ;
  assign n1709 = n1708 ^ n1663 ;
  assign n1710 = n1160 & ~n1709 ;
  assign n1701 = n1699 ^ n1663 ;
  assign n1711 = n1710 ^ n1701 ;
  assign n1712 = ~n1700 & ~n1711 ;
  assign n1713 = n1712 ^ n1699 ;
  assign n1752 = n1713 ^ n1684 ;
  assign n1718 = ~n1160 & ~n1468 ;
  assign n1719 = ~n1138 & ~n1718 ;
  assign n1720 = n1483 ^ n1067 ;
  assign n1721 = n1720 ^ n1484 ;
  assign n1722 = n1703 ^ n1484 ;
  assign n1723 = ~n1721 & n1722 ;
  assign n1724 = n1723 ^ n1484 ;
  assign n1725 = n1160 & ~n1724 ;
  assign n1726 = n1725 ^ n1703 ;
  assign n1727 = ~n1719 & n1726 ;
  assign n1716 = ~n1287 & ~n1696 ;
  assign n1714 = n1581 ^ n1135 ;
  assign n1715 = ~n1714 & n2127 ;
  assign n1717 = n1716 ^ n1715 ;
  assign n1728 = n1727 ^ n1717 ;
  assign n1732 = ~n1021 & ~n1228 ;
  assign n1733 = n1732 ^ n1017 ;
  assign n1734 = ~n1456 & n1733 ;
  assign n1730 = n1228 ^ n1017 ;
  assign n1735 = n1734 ^ n1730 ;
  assign n1736 = n1735 ^ n1717 ;
  assign n1737 = ~n1728 & n1736 ;
  assign n1738 = n1737 ^ n1727 ;
  assign n1741 = n920 & ~n1468 ;
  assign n1742 = n1726 ^ n1719 ;
  assign n1743 = n1742 ^ n1727 ;
  assign n1744 = n1717 & ~n1735 ;
  assign n1745 = n1744 ^ n1738 ;
  assign n1746 = n1745 ^ n1741 ;
  assign n1747 = ~n1743 & n1746 ;
  assign n1748 = n1747 ^ n1744 ;
  assign n1749 = ~n1741 & ~n1748 ;
  assign n1750 = ~n1738 & n1749 ;
  assign n1739 = n1738 ^ n1713 ;
  assign n1751 = n1750 ^ n1739 ;
  assign n1753 = n1752 ^ n1751 ;
  assign n1754 = n1753 ^ n1752 ;
  assign n1755 = n1711 ^ n1695 ;
  assign n1756 = n1755 ^ n1748 ;
  assign n1757 = n1742 ^ n1736 ;
  assign n1766 = n1177 & ~n1228 ;
  assign n1767 = n1766 ^ n1021 ;
  assign n1768 = ~n1456 & ~n1767 ;
  assign n1764 = n1228 ^ n1021 ;
  assign n1769 = n1768 ^ n1764 ;
  assign n1760 = ~n1287 & ~n1714 ;
  assign n1758 = n1483 ^ n1135 ;
  assign n1759 = ~n1758 & n2127 ;
  assign n1761 = n1760 ^ n1759 ;
  assign n1770 = n1769 ^ n1761 ;
  assign n1777 = ~n1228 & n1581 ;
  assign n1778 = n1777 ^ n1177 ;
  assign n1779 = ~n1456 & n1778 ;
  assign n1775 = n1228 ^ n1177 ;
  assign n1780 = n1779 ^ n1775 ;
  assign n1781 = n1468 ^ n1228 ;
  assign n1782 = ~n1287 & n1781 ;
  assign n1783 = n1782 ^ n1228 ;
  assign n1784 = ~n1135 & n1783 ;
  assign n1785 = ~n1780 & n1784 ;
  assign n1786 = n1785 ^ n1769 ;
  assign n1787 = n1770 & n1786 ;
  assign n1788 = n1787 ^ n1769 ;
  assign n1789 = n1757 & n1788 ;
  assign n1791 = n1285 & ~n1468 ;
  assign n1790 = n1456 & n1581 ;
  assign n1792 = n1791 ^ n1790 ;
  assign n1840 = n1483 ^ n1228 ;
  assign n1801 = n1840 ^ n1456 ;
  assign n1825 = ~n1483 & n1801 ;
  assign n1818 = n1456 ^ n1228 ;
  assign n1835 = n1581 ^ n1483 ;
  assign n1816 = n1835 ^ n1456 ;
  assign n1817 = n1816 ^ n1468 ;
  assign n1819 = n1818 ^ n1817 ;
  assign n1820 = ~n1781 & n1819 ;
  assign n1826 = n1825 ^ n1820 ;
  assign n1827 = n1826 ^ n1818 ;
  assign n1828 = n1825 ^ n1816 ;
  assign n1829 = n1828 ^ n1818 ;
  assign n1830 = ~n1827 & n1829 ;
  assign n1831 = n1456 & n1830 ;
  assign n1832 = n1831 ^ n1825 ;
  assign n1844 = n1832 ^ n1801 ;
  assign n1794 = n1581 ^ n1456 ;
  assign n1845 = n1844 ^ n1794 ;
  assign n1802 = n1581 ^ n1228 ;
  assign n1846 = n1845 ^ n1802 ;
  assign n1847 = ~n1792 & ~n1846 ;
  assign n1848 = n1758 ^ n1468 ;
  assign n1849 = n1848 ^ n1285 ;
  assign n1850 = n1849 ^ n1758 ;
  assign n1851 = n1758 ^ n1484 ;
  assign n1852 = n1850 & n1851 ;
  assign n1853 = n1852 ^ n1758 ;
  assign n1854 = n1287 & ~n1853 ;
  assign n1855 = n1854 ^ n1758 ;
  assign n1862 = n1855 ^ n1770 ;
  assign n1856 = n1770 & ~n1855 ;
  assign n1863 = n1862 ^ n1856 ;
  assign n1864 = ~n1784 & n1863 ;
  assign n1858 = ~n1718 & ~n1784 ;
  assign n1859 = n1858 ^ n1770 ;
  assign n1860 = n1780 & ~n1859 ;
  assign n1857 = ~n1718 & ~n1856 ;
  assign n1861 = n1860 ^ n1857 ;
  assign n1865 = n1864 ^ n1861 ;
  assign n1866 = ~n1847 & n1865 ;
  assign n1867 = n1858 ^ n1757 ;
  assign n1868 = ~n1770 & ~n1867 ;
  assign n1869 = n1868 ^ n1757 ;
  assign n1870 = n1780 & n1869 ;
  assign n1878 = ~n1857 & n1870 ;
  assign n1879 = ~n1863 & n1878 ;
  assign n1880 = n1879 ^ n1863 ;
  assign n1871 = n1870 ^ n1869 ;
  assign n1872 = n1871 ^ n1863 ;
  assign n1881 = n1880 ^ n1872 ;
  assign n1882 = ~n1866 & n1881 ;
  assign n1883 = ~n1789 & n1882 ;
  assign n1886 = n1883 ^ n1755 ;
  assign n1887 = n1886 ^ n1789 ;
  assign n1884 = ~n1769 & n1868 ;
  assign n1885 = n1883 & n1884 ;
  assign n1888 = n1887 ^ n1885 ;
  assign n1889 = ~n1756 & n1888 ;
  assign n1890 = n1889 ^ n1755 ;
  assign n1891 = n1890 ^ n1684 ;
  assign n1892 = n1891 ^ n1752 ;
  assign n1893 = ~n1754 & n1892 ;
  assign n1894 = n1893 ^ n1752 ;
  assign n1895 = ~n1688 & n1894 ;
  assign n1896 = n1895 ^ n1687 ;
  assign n1897 = n1686 ^ n1685 ;
  assign n1898 = n1897 ^ n1687 ;
  assign n1899 = n1890 ^ n1751 ;
  assign n1900 = n1898 & ~n1899 ;
  assign n1903 = n1713 & n1890 ;
  assign n1904 = n1903 ^ n1684 ;
  assign n1905 = n1900 & ~n1904 ;
  assign n1906 = ~n1896 & ~n1905 ;
  assign n1909 = n1907 ^ n1906 ;
  assign n1908 = n1906 & ~n1907 ;
  assign n1910 = n1909 ^ n1908 ;
  assign n1636 = ~n947 & ~n1468 ;
  assign n1517 = ~n749 & ~n1516 ;
  assign n1521 = n753 & ~n1228 ;
  assign n1522 = n1521 ^ n751 ;
  assign n1523 = ~n1456 & n1522 ;
  assign n1519 = n1228 ^ n751 ;
  assign n1524 = n1523 ^ n1519 ;
  assign n1634 = n1517 & ~n1524 ;
  assign n1630 = n1353 & ~n1601 ;
  assign n1631 = n1630 ^ n1623 ;
  assign n1632 = n1160 & ~n1631 ;
  assign n1621 = n920 & n1620 ;
  assign n1619 = n997 & ~n1402 ;
  assign n1622 = n1621 ^ n1619 ;
  assign n1624 = n1623 ^ n1622 ;
  assign n1633 = n1632 ^ n1624 ;
  assign n1635 = n1634 ^ n1633 ;
  assign n1637 = n1636 ^ n1635 ;
  assign n1616 = n1615 ^ n1609 ;
  assign n1617 = n1611 & ~n1616 ;
  assign n1618 = n1617 ^ n1609 ;
  assign n1638 = n1637 ^ n1618 ;
  assign n1508 = n1483 ^ n731 ;
  assign n1587 = n950 & ~n1508 ;
  assign n1588 = n1587 ^ n1582 ;
  assign n1589 = ~n689 & ~n1588 ;
  assign n1590 = n1589 ^ n1582 ;
  assign n1576 = n751 & ~n1228 ;
  assign n1577 = n1576 ^ n738 ;
  assign n1578 = ~n1456 & ~n1577 ;
  assign n1568 = ~n1414 & ~n1563 ;
  assign n1569 = n1568 ^ n1494 ;
  assign n1570 = n1287 & ~n1569 ;
  assign n1571 = n1570 ^ n1494 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1579 = n1578 ^ n1573 ;
  assign n1591 = n1590 ^ n1579 ;
  assign n1509 = n1508 ^ n1484 ;
  assign n1512 = n950 & n1509 ;
  assign n1513 = n1512 ^ n1508 ;
  assign n1514 = ~n689 & ~n1513 ;
  assign n1515 = n1514 ^ n1508 ;
  assign n1592 = n1591 ^ n1515 ;
  assign n1525 = n1524 ^ n1517 ;
  assign n1526 = n1525 ^ n1515 ;
  assign n1556 = n1555 ^ n1544 ;
  assign n1557 = n1545 & ~n1556 ;
  assign n1558 = n1557 ^ n1555 ;
  assign n1559 = n1558 ^ n1515 ;
  assign n1560 = n1526 & ~n1559 ;
  assign n1593 = n1592 ^ n1560 ;
  assign n1644 = n1638 ^ n1593 ;
  assign n1911 = n1910 ^ n1644 ;
  assign n1927 = n1558 ^ n1526 ;
  assign n1912 = n1516 & n1660 ;
  assign n1915 = n1655 & n1912 ;
  assign n1916 = n1915 ^ n1661 ;
  assign n1913 = n1912 ^ n1661 ;
  assign n1914 = ~n1655 & ~n1913 ;
  assign n1917 = n1916 ^ n1914 ;
  assign n1918 = n1917 ^ n1655 ;
  assign n1919 = n1915 ^ n1645 ;
  assign n1920 = n1683 ^ n1645 ;
  assign n1921 = ~n1919 & n1920 ;
  assign n1922 = n1921 ^ n1915 ;
  assign n1923 = n1921 & n1922 ;
  assign n1924 = n1918 & n1923 ;
  assign n1925 = n1924 ^ n1922 ;
  assign n1930 = n1914 ^ n1645 ;
  assign n1931 = n1920 & n1930 ;
  assign n1932 = n1931 ^ n1914 ;
  assign n1933 = ~n1918 & n1932 ;
  assign n1934 = n1931 & n1933 ;
  assign n1935 = n1934 ^ n1932 ;
  assign n1940 = ~n1925 & ~n1935 ;
  assign n1941 = n1927 & n1940 ;
  assign n1942 = n1941 ^ n1927 ;
  assign n1926 = n1925 ^ n1644 ;
  assign n1928 = n1927 ^ n1926 ;
  assign n1943 = n1942 ^ n1928 ;
  assign n1944 = ~n1911 & n1943 ;
  assign n1945 = n1944 ^ n1910 ;
  assign n1946 = n1935 ^ n1925 ;
  assign n1947 = ~n1644 & n1946 ;
  assign n1948 = n1947 ^ n1925 ;
  assign n1949 = n1927 ^ n1644 ;
  assign n1950 = n1949 ^ n1908 ;
  assign n1951 = n1948 & ~n1950 ;
  assign n1952 = n1951 ^ n1644 ;
  assign n1953 = ~n1908 & ~n1952 ;
  assign n1954 = ~n1945 & ~n1953 ;
  assign n1642 = n1502 ^ n1493 ;
  assign n1639 = n1638 ^ n1591 ;
  assign n1640 = n1593 & n1639 ;
  assign n1641 = n1640 ^ n1638 ;
  assign n1643 = n1642 ^ n1641 ;
  assign n1955 = n1954 ^ n1643 ;
  assign n1986 = n1635 ^ n1618 ;
  assign n1987 = ~n1637 & n1986 ;
  assign n1988 = n1987 ^ n1635 ;
  assign n1983 = n1982 ^ n1973 ;
  assign n1959 = n1634 ^ n1622 ;
  assign n1960 = n1633 & n1959 ;
  assign n1961 = n1960 ^ n1634 ;
  assign n1984 = n1983 ^ n1961 ;
  assign n1956 = n1590 ^ n1571 ;
  assign n1957 = ~n1579 & n1956 ;
  assign n1958 = n1957 ^ n1571 ;
  assign n1985 = n1984 ^ n1958 ;
  assign n1990 = n1988 ^ n1985 ;
  assign n1989 = ~n1985 & ~n1988 ;
  assign n1991 = n1990 ^ n1989 ;
  assign n2009 = n2008 ^ n1998 ;
  assign n1995 = n1505 ^ n1409 ;
  assign n2010 = n2009 ^ n1995 ;
  assign n1992 = n1961 ^ n1958 ;
  assign n1993 = ~n1984 & ~n1992 ;
  assign n1994 = n1993 ^ n1958 ;
  assign n2011 = n2010 ^ n1994 ;
  assign n2012 = n2011 ^ n1641 ;
  assign n2013 = n2012 ^ n2011 ;
  assign n2014 = n2011 ^ n1642 ;
  assign n2015 = n2014 ^ n2011 ;
  assign n2016 = n2013 & n2015 ;
  assign n2017 = n2016 ^ n2011 ;
  assign n2018 = n1991 & ~n2017 ;
  assign n2019 = ~n1955 & n2018 ;
  assign n2020 = n2011 ^ n1989 ;
  assign n2021 = n1954 ^ n1641 ;
  assign n2022 = ~n1643 & n2021 ;
  assign n2023 = n2022 ^ n1643 ;
  assign n2024 = n2023 ^ n1954 ;
  assign n2025 = n2024 ^ n2011 ;
  assign n2026 = ~n2020 & ~n2025 ;
  assign n2027 = n2026 ^ n2011 ;
  assign n2028 = ~n2019 & n2027 ;
  assign n2029 = n1507 & n2028 ;
  assign n2143 = n2142 ^ n2029 ;
  assign n2145 = n2083 ^ n2074 ;
  assign n2144 = n2068 ^ n2065 ;
  assign n2146 = n2145 ^ n2144 ;
  assign n2148 = n2009 ^ n1994 ;
  assign n2149 = n2010 & n2148 ;
  assign n2150 = n2149 ^ n2009 ;
  assign n2152 = n2150 ^ n2144 ;
  assign n2153 = ~n2146 & n2152 ;
  assign n2147 = n2146 ^ n2029 ;
  assign n2151 = n2150 ^ n2147 ;
  assign n2154 = n2153 ^ n2151 ;
  assign n2155 = n2143 & n2154 ;
  assign n2156 = n2155 ^ n2142 ;
  assign n2157 = n2028 ^ n1507 ;
  assign n2158 = n2157 ^ n2029 ;
  assign n2159 = n2144 ^ n2142 ;
  assign n2162 = n2153 & ~n2159 ;
  assign n2163 = n2162 ^ n2142 ;
  assign n2164 = n2158 & n2163 ;
  assign n2165 = ~n2156 & ~n2164 ;
  assign n2176 = n2174 ^ n2165 ;
  assign n2175 = ~n2165 & ~n2174 ;
  assign n2177 = n2176 ^ n2175 ;
  assign n2204 = n2194 ^ n2184 ;
  assign n2201 = n2108 ^ n2085 ;
  assign n2202 = ~n2115 & n2201 ;
  assign n2203 = n2202 ^ n2108 ;
  assign n2205 = n2204 ^ n2203 ;
  assign n2206 = n2116 ^ n2071 ;
  assign n2207 = ~n2141 & n2206 ;
  assign n2208 = n2207 ^ n2116 ;
  assign n2209 = n2208 ^ n2203 ;
  assign n2210 = n2205 & ~n2209 ;
  assign n2211 = n2210 ^ n2205 ;
  assign n2200 = n2199 ^ n2180 ;
  assign n2214 = n2203 ^ n2200 ;
  assign n2215 = n2211 & n2214 ;
  assign n2216 = n2215 ^ n2200 ;
  assign n2217 = n2177 & n2216 ;
  assign n2218 = n2200 ^ n2175 ;
  assign n2219 = n2210 ^ n2208 ;
  assign n2220 = n2219 ^ n2200 ;
  assign n2221 = n2218 & ~n2220 ;
  assign n2222 = n2221 ^ n2200 ;
  assign n2223 = ~n2217 & ~n2222 ;
  assign n2229 = n2228 ^ n2223 ;
  assign n2230 = ~n1381 & ~n2229 ;
  assign n2232 = n1322 ^ n1153 ;
  assign n2231 = ~n2227 & ~n2228 ;
  assign n2233 = n2232 ^ n2231 ;
  assign n2234 = n2232 ^ n1379 ;
  assign n2235 = n2232 ^ n2227 ;
  assign n2236 = n2235 ^ n2223 ;
  assign n2237 = n2236 ^ n2226 ;
  assign n2238 = n2237 ^ n2235 ;
  assign n2239 = n2232 ^ n2223 ;
  assign n2240 = n2239 ^ n2235 ;
  assign n2241 = ~n2238 & n2240 ;
  assign n2242 = n2241 ^ n2235 ;
  assign n2243 = ~n2234 & ~n2242 ;
  assign n2244 = n2243 ^ n1379 ;
  assign n2245 = ~n2233 & ~n2244 ;
  assign n2246 = n2230 & n2245 ;
  assign n2247 = n2246 ^ n2244 ;
  assign n2250 = n1332 ^ n1330 ;
  assign n2251 = n2250 ^ n1325 ;
  assign n2252 = n2251 ^ n1341 ;
  assign n2253 = n2252 ^ n1338 ;
  assign n2248 = n1336 ^ n1325 ;
  assign n2249 = n2248 ^ n1340 ;
  assign n2254 = n2253 ^ n2249 ;
  assign n2255 = n2254 ^ n2253 ;
  assign n2256 = n975 & n2255 ;
  assign n2257 = n2256 ^ n2253 ;
  assign n2258 = n2247 & ~n2257 ;
  assign n2259 = ~n1341 & ~n2258 ;
  assign n2260 = n975 & n2259 ;
  assign n2261 = ~n1338 & n2260 ;
  assign n2262 = n2261 ^ n2259 ;
  assign n2263 = n2262 ^ n2258 ;
  assign n2264 = n2263 ^ n987 ;
  assign n2265 = n988 & n2264 ;
  assign n2266 = n2265 ^ n987 ;
  assign n799 = n751 & n753 ;
  assign n800 = n799 ^ n754 ;
  assign n801 = n800 ^ n739 ;
  assign n802 = ~n727 & ~n801 ;
  assign n796 = ~n696 & ~n730 ;
  assign n797 = n796 ^ n696 ;
  assign n786 = n785 ^ n784 ;
  assign n795 = ~n786 & ~n794 ;
  assign n798 = n797 ^ n795 ;
  assign n803 = n802 ^ n798 ;
  assign n2267 = n2266 ^ n803 ;
  assign n467 = n466 ^ n322 ;
  assign n468 = n467 ^ n228 ;
  assign n469 = n468 ^ n461 ;
  assign n164 = ~n62 & n78 ;
  assign n456 = n455 ^ n164 ;
  assign n457 = n456 ^ n267 ;
  assign n459 = n458 ^ n457 ;
  assign n452 = n451 ^ n449 ;
  assign n445 = n444 ^ n391 ;
  assign n453 = n452 ^ n445 ;
  assign n460 = n459 ^ n453 ;
  assign n470 = n469 ^ n460 ;
  assign n417 = n416 ^ n403 ;
  assign n418 = n417 ^ n233 ;
  assign n412 = n343 ^ n281 ;
  assign n413 = n412 ^ n351 ;
  assign n419 = n418 ^ n413 ;
  assign n439 = n438 ^ n419 ;
  assign n471 = n470 ^ n439 ;
  assign n492 = n389 ^ n248 ;
  assign n479 = n382 ^ n140 ;
  assign n477 = n476 ^ n475 ;
  assign n478 = n477 ^ n224 ;
  assign n480 = n479 ^ n478 ;
  assign n472 = n356 ^ n238 ;
  assign n474 = n473 ^ n472 ;
  assign n481 = n480 ^ n474 ;
  assign n491 = n490 ^ n481 ;
  assign n493 = n492 ^ n491 ;
  assign n500 = n499 ^ n493 ;
  assign n501 = ~n471 & ~n500 ;
  assign n2268 = n2267 ^ n501 ;
  assign n2285 = n2263 ^ n988 ;
  assign n2283 = n78 & ~n485 ;
  assign n2281 = n1037 ^ n286 ;
  assign n2276 = n882 ^ n622 ;
  assign n2277 = n2276 ^ n843 ;
  assign n2278 = n2277 ^ n607 ;
  assign n2273 = n1102 ^ n166 ;
  assign n2271 = n389 ^ n206 ;
  assign n2272 = n2271 ^ n268 ;
  assign n2274 = n2273 ^ n2272 ;
  assign n2269 = n625 ^ n117 ;
  assign n2270 = n2269 ^ n512 ;
  assign n2275 = n2274 ^ n2270 ;
  assign n2279 = n2278 ^ n2275 ;
  assign n2280 = n2279 ^ n1226 ;
  assign n2282 = n2281 ^ n2280 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2286 = n2285 ^ n2284 ;
  assign n2304 = n1122 ^ n403 ;
  assign n2303 = n516 ^ n512 ;
  assign n2305 = n2304 ^ n2303 ;
  assign n2299 = n283 ^ n212 ;
  assign n2297 = n428 ^ n109 ;
  assign n2298 = n2297 ^ n496 ;
  assign n2300 = n2299 ^ n2298 ;
  assign n2301 = n2300 ^ n644 ;
  assign n2295 = n468 ^ n398 ;
  assign n2296 = n2295 ^ n299 ;
  assign n2302 = n2301 ^ n2296 ;
  assign n2306 = n2305 ^ n2302 ;
  assign n148 = n147 ^ n136 ;
  assign n127 = n126 ^ n110 ;
  assign n104 = n103 ^ n79 ;
  assign n128 = n127 ^ n104 ;
  assign n149 = n148 ^ n128 ;
  assign n2311 = n613 ^ n149 ;
  assign n2308 = n427 ^ n122 ;
  assign n2307 = n841 ^ n650 ;
  assign n2309 = n2308 ^ n2307 ;
  assign n2310 = n2309 ^ n647 ;
  assign n2312 = n2311 ^ n2310 ;
  assign n2318 = n850 ^ n204 ;
  assign n2319 = n2318 ^ n557 ;
  assign n2315 = n372 ^ n327 ;
  assign n2316 = n2315 ^ n226 ;
  assign n2314 = n627 ^ n402 ;
  assign n2317 = n2316 ^ n2314 ;
  assign n2320 = n2319 ^ n2317 ;
  assign n2313 = n535 ^ n261 ;
  assign n2321 = n2320 ^ n2313 ;
  assign n2322 = n2321 ^ n659 ;
  assign n2323 = ~n2312 & ~n2322 ;
  assign n2324 = n2306 & n2323 ;
  assign n2290 = n1332 ^ n1326 ;
  assign n2287 = n2247 ^ n1325 ;
  assign n2291 = n2287 ^ n1333 ;
  assign n2292 = ~n2290 & n2291 ;
  assign n2293 = n2292 ^ n975 ;
  assign n2288 = n1329 ^ n1325 ;
  assign n2289 = n2287 & ~n2288 ;
  assign n2294 = n2293 ^ n2289 ;
  assign n2325 = n2324 ^ n2294 ;
  assign n2358 = n375 ^ n126 ;
  assign n2359 = n2358 ^ n98 ;
  assign n2360 = n716 & n2359 ;
  assign n2356 = n2251 ^ n2247 ;
  assign n2352 = n671 ^ n348 ;
  assign n2353 = n2352 ^ n121 ;
  assign n2354 = n2353 ^ n2306 ;
  assign n2346 = n180 ^ n60 ;
  assign n2347 = n2346 ^ n279 ;
  assign n2340 = n1206 ^ n62 ;
  assign n2343 = ~n78 & n2340 ;
  assign n2344 = n2343 ^ n62 ;
  assign n2345 = ~n507 & ~n2344 ;
  assign n2348 = n2347 ^ n2345 ;
  assign n2331 = n153 ^ n63 ;
  assign n2332 = n152 ^ n96 ;
  assign n2337 = ~n42 & n2332 ;
  assign n2338 = n2337 ^ n685 ;
  assign n2339 = n2331 & n2338 ;
  assign n2349 = n2348 ^ n2339 ;
  assign n2350 = n2349 ^ n481 ;
  assign n2328 = n1125 ^ n286 ;
  assign n2327 = n2326 ^ n292 ;
  assign n2329 = n2328 ^ n2327 ;
  assign n2330 = n2329 ^ n865 ;
  assign n2351 = n2350 ^ n2330 ;
  assign n2355 = n2354 ^ n2351 ;
  assign n2357 = n2356 ^ n2355 ;
  assign n2361 = n2360 ^ n2357 ;
  assign n2392 = n507 ^ n194 ;
  assign n2393 = ~n251 & ~n2392 ;
  assign n2388 = n55 & n549 ;
  assign n2387 = n416 ^ n392 ;
  assign n2389 = n2388 ^ n2387 ;
  assign n2383 = n841 ^ n125 ;
  assign n2384 = n2383 ^ n222 ;
  assign n2381 = n540 ^ n283 ;
  assign n2382 = n2381 ^ n675 ;
  assign n2385 = n2384 ^ n2382 ;
  assign n2378 = n494 ^ n403 ;
  assign n2379 = n2378 ^ n324 ;
  assign n2376 = n850 ^ n287 ;
  assign n2377 = n2376 ^ n2375 ;
  assign n2380 = n2379 ^ n2377 ;
  assign n2386 = n2385 ^ n2380 ;
  assign n2390 = n2389 ^ n2386 ;
  assign n2391 = n2390 ^ n1116 ;
  assign n2394 = n2393 ^ n2391 ;
  assign n2395 = n2374 & n2394 ;
  assign n2364 = n2228 ^ n1380 ;
  assign n2365 = n2229 & ~n2364 ;
  assign n2362 = n2232 ^ n1381 ;
  assign n2363 = n2362 ^ n2231 ;
  assign n2366 = n2365 ^ n2363 ;
  assign n2396 = n2395 ^ n2366 ;
  assign n2398 = n555 & ~n1065 ;
  assign n2404 = n223 ^ n121 ;
  assign n2405 = n2404 ^ n1100 ;
  assign n2406 = n2405 ^ n649 ;
  assign n2407 = n2406 ^ n1076 ;
  assign n2408 = n2407 ^ n1053 ;
  assign n2399 = n1112 ^ n427 ;
  assign n2400 = n2399 ^ n305 ;
  assign n227 = n226 ^ n224 ;
  assign n229 = n228 ^ n227 ;
  assign n2401 = n2400 ^ n229 ;
  assign n2402 = n2401 ^ n1051 ;
  assign n2403 = n2402 ^ n363 ;
  assign n2409 = n2408 ^ n2403 ;
  assign n2410 = n2398 & ~n2409 ;
  assign n2397 = n2364 ^ n2223 ;
  assign n2411 = n2410 ^ n2397 ;
  assign n2561 = n324 ^ n206 ;
  assign n2562 = n2561 ^ n514 ;
  assign n2559 = n2558 ^ n350 ;
  assign n2560 = n2559 ^ n583 ;
  assign n2563 = n2562 ^ n2560 ;
  assign n2431 = n671 ^ n287 ;
  assign n2432 = n2431 ^ n372 ;
  assign n2564 = n2563 ^ n2432 ;
  assign n2565 = n2564 ^ n1095 ;
  assign n2552 = n441 ^ n398 ;
  assign n2553 = n2552 ^ n434 ;
  assign n2554 = n2553 ^ n853 ;
  assign n2550 = n709 ^ n618 ;
  assign n2548 = n557 ^ n110 ;
  assign n2546 = n625 ^ n511 ;
  assign n2547 = n2546 ^ n154 ;
  assign n2549 = n2548 ^ n2547 ;
  assign n2551 = n2550 ^ n2549 ;
  assign n2555 = n2554 ^ n2551 ;
  assign n2566 = n2565 ^ n2555 ;
  assign n2567 = ~n2545 & n2566 ;
  assign n2440 = n382 ^ n136 ;
  assign n2441 = n2440 ^ n2319 ;
  assign n2438 = n664 ^ n208 ;
  assign n2436 = n864 ^ n223 ;
  assign n2437 = n2436 ^ n355 ;
  assign n2439 = n2438 ^ n2437 ;
  assign n2442 = n2441 ^ n2439 ;
  assign n2427 = n55 & n78 ;
  assign n2424 = n596 ^ n435 ;
  assign n2425 = n2424 ^ n444 ;
  assign n2419 = n132 ^ n102 ;
  assign n2420 = n565 ^ n152 ;
  assign n2421 = n2420 ^ n864 ;
  assign n2422 = ~n2419 & ~n2421 ;
  assign n2415 = n291 ^ n212 ;
  assign n2414 = n709 ^ n649 ;
  assign n2416 = n2415 ^ n2414 ;
  assign n2417 = n2416 ^ n281 ;
  assign n2418 = n2417 ^ n415 ;
  assign n2423 = n2422 ^ n2418 ;
  assign n2426 = n2425 ^ n2423 ;
  assign n2428 = n2427 ^ n2426 ;
  assign n2430 = n895 ^ n327 ;
  assign n2433 = n2432 ^ n2430 ;
  assign n2429 = n124 & n1105 ;
  assign n2434 = n2433 ^ n2429 ;
  assign n2435 = ~n2428 & ~n2434 ;
  assign n2443 = n2442 ^ n2435 ;
  assign n2444 = ~n846 & n2443 ;
  assign n2412 = n2208 ^ n2205 ;
  assign n2413 = n2412 ^ n2176 ;
  assign n2445 = n2444 ^ n2413 ;
  assign n2461 = n2460 ^ n2402 ;
  assign n2456 = n365 ^ n79 ;
  assign n155 = n154 ^ n153 ;
  assign n2455 = n384 ^ n155 ;
  assign n2457 = n2456 ^ n2455 ;
  assign n2453 = n2431 ^ n2358 ;
  assign n2450 = n1039 ^ n206 ;
  assign n2451 = n2450 ^ n304 ;
  assign n2452 = n2451 ^ n1254 ;
  assign n2454 = n2453 ^ n2452 ;
  assign n2458 = n2457 ^ n2454 ;
  assign n2462 = n2461 ^ n2458 ;
  assign n2474 = n2473 ^ n633 ;
  assign n2468 = n539 ^ n180 ;
  assign n2465 = n329 ^ n146 ;
  assign n2466 = n2465 ^ n310 ;
  assign n2467 = n2466 ^ n263 ;
  assign n2469 = n2468 ^ n2467 ;
  assign n2464 = n2463 ^ n1064 ;
  assign n2470 = n2469 ^ n2464 ;
  assign n2471 = n2470 ^ n2423 ;
  assign n2475 = n2474 ^ n2471 ;
  assign n2476 = n2462 & n2475 ;
  assign n2446 = n2150 ^ n2146 ;
  assign n2447 = n2446 ^ n1507 ;
  assign n2448 = ~n2157 & n2447 ;
  assign n2160 = n2153 ^ n2142 ;
  assign n2449 = n2448 ^ n2160 ;
  assign n2477 = n2476 ^ n2449 ;
  assign n2498 = n242 ^ n211 ;
  assign n2499 = ~n98 & n2498 ;
  assign n2500 = n2499 ^ n841 ;
  assign n2501 = n2500 ^ n709 ;
  assign n2502 = n2501 ^ n892 ;
  assign n2495 = n310 ^ n103 ;
  assign n2496 = n2495 ^ n2431 ;
  assign n2493 = n2492 ^ n625 ;
  assign n2491 = n1255 ^ n850 ;
  assign n2494 = n2493 ^ n2491 ;
  assign n2497 = n2496 ^ n2494 ;
  assign n2503 = n2502 ^ n2497 ;
  assign n2487 = n96 ^ n42 ;
  assign n2488 = ~n314 & ~n345 ;
  assign n2489 = ~n2487 & n2488 ;
  assign n2483 = n511 ^ n404 ;
  assign n2484 = n2483 ^ n406 ;
  assign n2485 = n2484 ^ n2482 ;
  assign n2479 = n2315 ^ n477 ;
  assign n2480 = n2479 ^ n118 ;
  assign n2481 = n2480 ^ n450 ;
  assign n2486 = n2485 ^ n2481 ;
  assign n2490 = n2489 ^ n2486 ;
  assign n2504 = n2503 ^ n2490 ;
  assign n2505 = n2504 ^ n363 ;
  assign n2478 = n2446 ^ n2157 ;
  assign n2506 = n2505 ^ n2478 ;
  assign n2507 = n463 & ~n1202 ;
  assign n2515 = n111 & n152 ;
  assign n2513 = n292 ^ n180 ;
  assign n2514 = n2513 ^ n108 ;
  assign n2516 = n2515 ^ n2514 ;
  assign n2517 = ~n861 & ~n2516 ;
  assign n2508 = n1114 ^ n845 ;
  assign n2509 = n2508 ^ n517 ;
  assign n2510 = n2509 ^ n1218 ;
  assign n2511 = n2510 ^ n2442 ;
  assign n2512 = n2511 ^ n470 ;
  assign n2518 = n2517 ^ n2512 ;
  assign n2519 = n2507 & ~n2518 ;
  assign n2520 = n2519 ^ n2518 ;
  assign n2522 = n2024 ^ n2022 ;
  assign n2523 = n2522 ^ n1988 ;
  assign n2524 = ~n1990 & n2523 ;
  assign n2521 = n2022 ^ n2011 ;
  assign n2525 = n2524 ^ n2521 ;
  assign n2526 = ~n2520 & n2525 ;
  assign n2527 = n2526 ^ n2478 ;
  assign n2528 = n2506 & n2527 ;
  assign n2529 = n2528 ^ n2505 ;
  assign n2530 = n2529 ^ n2449 ;
  assign n2531 = n2477 & ~n2530 ;
  assign n2532 = n2531 ^ n2449 ;
  assign n2533 = n2532 ^ n2413 ;
  assign n2534 = ~n2445 & ~n2533 ;
  assign n2535 = n2534 ^ n2413 ;
  assign n2568 = n2567 ^ n2535 ;
  assign n2212 = n2211 ^ n2200 ;
  assign n2572 = n2567 ^ n2212 ;
  assign n2569 = n2205 ^ n2174 ;
  assign n2570 = n2569 ^ n2208 ;
  assign n2571 = ~n2176 & ~n2570 ;
  assign n2573 = n2572 ^ n2571 ;
  assign n2574 = ~n2568 & n2573 ;
  assign n2575 = n2574 ^ n2567 ;
  assign n2576 = n2575 ^ n2397 ;
  assign n2577 = ~n2411 & ~n2576 ;
  assign n2578 = n2577 ^ n2397 ;
  assign n2579 = n2578 ^ n2366 ;
  assign n2580 = n2396 & n2579 ;
  assign n2581 = n2580 ^ n2578 ;
  assign n2582 = n2581 ^ n2356 ;
  assign n2583 = ~n2361 & n2582 ;
  assign n2584 = n2583 ^ n2356 ;
  assign n2587 = n2584 ^ n2294 ;
  assign n2588 = n2325 & n2587 ;
  assign n2585 = n2584 ^ n2285 ;
  assign n2589 = n2588 ^ n2585 ;
  assign n2590 = ~n2286 & n2589 ;
  assign n2591 = n2590 ^ n2285 ;
  assign n2592 = n2591 ^ n2267 ;
  assign n2593 = ~n2268 & n2592 ;
  assign n2594 = n2593 ^ n2267 ;
  assign n2611 = n2610 ^ n2594 ;
  assign n2624 = n2610 ^ n2266 ;
  assign n2612 = ~n738 & ~n800 ;
  assign n2615 = n2612 ^ n800 ;
  assign n2616 = ~n696 & n2615 ;
  assign n2617 = ~n727 & n2616 ;
  assign n2618 = n2617 ^ n797 ;
  assign n2619 = n795 & ~n2266 ;
  assign n2620 = ~n2618 & n2619 ;
  assign n2621 = n2620 ^ n2266 ;
  assign n2625 = n2624 ^ n2621 ;
  assign n5689 = ~n738 & n800 ;
  assign n2614 = ~n727 & n5689 ;
  assign n2622 = n796 & ~n2621 ;
  assign n2623 = n2614 & n2622 ;
  assign n2626 = n2625 ^ n2623 ;
  assign n2627 = ~n2611 & n2626 ;
  assign n2628 = n2627 ^ n2610 ;
  assign n2629 = n411 & n2628 ;
  assign n2659 = n2658 ^ n2629 ;
  assign n2771 = x22 & n28 ;
  assign n2772 = n2771 ^ n27 ;
  assign n4566 = ~n28 & n2772 ;
  assign n4573 = n4566 ^ n2772 ;
  assign n3502 = n30 ^ n29 ;
  assign n2774 = x0 & x2 ;
  assign n2761 = x0 & ~x22 ;
  assign n2775 = n2774 ^ n2761 ;
  assign n3737 = n3502 ^ n2775 ;
  assign n4574 = n4573 ^ n3737 ;
  assign n2780 = ~n1468 & n4574 ;
  assign n2781 = ~n4574 ^ n2780 ;
  assign n2792 = ~n1483 & ~n2781 ;
  assign n2805 = ~n1581 & n2792 ;
  assign n2795 = n2792 ^ n2781 ;
  assign n2789 = ~n4574 ^ n1468 ;
  assign n2790 = ~n1483 & ~n2789 ;
  assign n2791 = n2790 ^ n1483 ;
  assign n2793 = n2792 ^ n2791 ;
  assign n2796 = n2795 ^ n2793 ;
  assign n4167 = n2805 ^ n2796 ;
  assign n4168 = ~n2659 & n4167 ;
  assign n3229 = n1581 & ~n2789 ;
  assign n3189 = n3229 ^ n2789 ;
  assign n4165 = n3189 ^ n1581 ;
  assign n2801 = n1581 & n2789 ;
  assign n2800 = n1581 & ~n2796 ;
  assign n2802 = n2801 ^ n2800 ;
  assign n2798 = n2792 ^ n1581 ;
  assign n2797 = n2796 ^ n2789 ;
  assign n2799 = n2798 ^ n2797 ;
  assign n2803 = n2802 ^ n2799 ;
  assign n2804 = n2803 ^ n2792 ;
  assign n2806 = n2805 ^ n2804 ;
  assign n4166 = n4165 ^ n2806 ;
  assign n4169 = n4168 ^ n4166 ;
  assign n2820 = n2628 ^ n411 ;
  assign n4174 = n2803 & n2820 ;
  assign n4176 = n4174 ^ n2805 ;
  assign n4170 = n2805 ^ n2792 ;
  assign n4177 = n4176 ^ n4170 ;
  assign n4178 = ~n4169 & ~n4177 ;
  assign n2660 = ~n2629 & ~n2658 ;
  assign n2661 = n2660 ^ n2659 ;
  assign n214 = n213 ^ n207 ;
  assign n179 = n178 ^ n132 ;
  assign n183 = n182 ^ n179 ;
  assign n185 = n184 ^ n183 ;
  assign n198 = n197 ^ n185 ;
  assign n215 = n214 ^ n198 ;
  assign n176 = n175 ^ n171 ;
  assign n163 = n162 ^ n155 ;
  assign n165 = n164 ^ n163 ;
  assign n177 = n176 ^ n165 ;
  assign n216 = n215 ^ n177 ;
  assign n217 = ~n149 & ~n216 ;
  assign n236 = n235 ^ n229 ;
  assign n220 = n219 ^ n218 ;
  assign n237 = n236 ^ n220 ;
  assign n250 = n249 ^ n237 ;
  assign n277 = n276 ^ n250 ;
  assign n278 = n217 & ~n277 ;
  assign n2662 = n2661 ^ n278 ;
  assign n4158 = n2662 ^ n1581 ;
  assign n4157 = n2662 ^ n1483 ;
  assign n4159 = n4158 ^ n4157 ;
  assign n2735 = n2658 ^ n411 ;
  assign n2696 = ~n2614 & n2618 ;
  assign n2697 = n2696 ^ n2266 ;
  assign n2698 = n803 & ~n2697 ;
  assign n2691 = ~n2594 & n2610 ;
  assign n2727 = n2691 ^ n2611 ;
  assign n2728 = ~n2698 & n2727 ;
  assign n2699 = n2691 & n2698 ;
  assign n2736 = n2728 ^ n2699 ;
  assign n2737 = n2736 ^ n2628 ;
  assign n2721 = n2591 ^ n2268 ;
  assign n2719 = n2589 ^ n2284 ;
  assign n2700 = n2584 ^ n2325 ;
  assign n2701 = n2581 ^ n2361 ;
  assign n2702 = n2578 ^ n2396 ;
  assign n2703 = n2575 ^ n2411 ;
  assign n2704 = n2573 ^ n2535 ;
  assign n2705 = n2532 ^ n2445 ;
  assign n2706 = n2529 ^ n2477 ;
  assign n2710 = n2526 ^ n2506 ;
  assign n2738 = n2706 & ~n2710 ;
  assign n2739 = ~n2705 & ~n2738 ;
  assign n2740 = n2704 & ~n2739 ;
  assign n2741 = ~n2703 & ~n2740 ;
  assign n2742 = ~n2702 & ~n2741 ;
  assign n2743 = n2701 & ~n2742 ;
  assign n2744 = ~n2700 & ~n2743 ;
  assign n2745 = n2719 & ~n2744 ;
  assign n2746 = ~n2721 & ~n2745 ;
  assign n2747 = ~n2737 & ~n2746 ;
  assign n2748 = n2747 ^ n2658 ;
  assign n2749 = n2735 & n2748 ;
  assign n2750 = n2747 ^ n2628 ;
  assign n2751 = n2749 & ~n2750 ;
  assign n2752 = n2751 ^ n2658 ;
  assign n2707 = n2525 ^ n2520 ;
  assign n2708 = n2506 & ~n2707 ;
  assign n2709 = n2708 ^ n2707 ;
  assign n2711 = n2710 ^ n2709 ;
  assign n2712 = ~n2706 & ~n2711 ;
  assign n2713 = n2705 & ~n2712 ;
  assign n2714 = ~n2704 & ~n2713 ;
  assign n2715 = n2703 & ~n2714 ;
  assign n2716 = n2702 & ~n2715 ;
  assign n2717 = ~n2701 & ~n2716 ;
  assign n2718 = n2700 & ~n2717 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2722 = ~n2720 & n2721 ;
  assign n2729 = ~n2722 & n2728 ;
  assign n2723 = ~n2699 & n2722 ;
  assign n2724 = n2628 & n2723 ;
  assign n2725 = n2724 ^ n2699 ;
  assign n2726 = n2725 ^ n2628 ;
  assign n2730 = n2729 ^ n2726 ;
  assign n2731 = n411 & ~n2730 ;
  assign n2732 = n2731 ^ n2725 ;
  assign n2733 = n2660 & ~n2732 ;
  assign n3688 = n2752 ^ n2733 ;
  assign n4160 = n4157 ^ n3688 ;
  assign n4161 = n4160 ^ n4157 ;
  assign n4162 = n4159 & n4161 ;
  assign n4163 = n4162 ^ n4157 ;
  assign n4164 = ~n2789 & ~n4163 ;
  assign n4179 = n4178 ^ n4164 ;
  assign n2868 = n1581 ^ n1021 ;
  assign n1773 = n1581 ^ n1177 ;
  assign n2869 = n1177 ^ n1017 ;
  assign n2870 = ~n1773 & n2869 ;
  assign n2871 = n2868 & n2870 ;
  assign n3184 = n2744 ^ n2718 ;
  assign n3182 = n2745 ^ n2744 ;
  assign n3183 = n3182 ^ n2720 ;
  assign n3185 = n3184 ^ n3183 ;
  assign n3186 = n3185 ^ n2718 ;
  assign n3866 = n3186 ^ n2700 ;
  assign n3867 = n2871 & n3866 ;
  assign n3863 = n1773 & ~n2721 ;
  assign n2864 = n1021 & ~n1773 ;
  assign n2862 = n1177 & n1581 ;
  assign n2863 = n2862 ^ n1773 ;
  assign n2865 = n2864 ^ n2863 ;
  assign n2989 = n2865 ^ n1017 ;
  assign n3860 = ~n1017 & ~n3186 ;
  assign n3861 = n2989 & n3860 ;
  assign n3858 = n2989 ^ n2719 ;
  assign n3862 = n3861 ^ n3858 ;
  assign n3864 = n3863 ^ n3862 ;
  assign n3853 = n2719 ^ n1021 ;
  assign n3854 = n3853 ^ n2719 ;
  assign n3855 = ~n3186 & n3854 ;
  assign n3856 = n3855 ^ n2719 ;
  assign n3857 = n2865 & n3856 ;
  assign n3865 = n3864 ^ n3857 ;
  assign n3868 = n3867 ^ n3865 ;
  assign n3808 = n2701 ^ n829 ;
  assign n1310 = n1017 ^ n827 ;
  assign n2855 = n2743 ^ n2717 ;
  assign n2856 = n2855 ^ n2716 ;
  assign n3804 = n1310 & n2856 ;
  assign n2896 = n829 & n1310 ;
  assign n2905 = ~n753 & n2896 ;
  assign n1537 = n829 ^ n753 ;
  assign n2899 = n827 & n1017 ;
  assign n2900 = n2899 ^ n1310 ;
  assign n2903 = n2900 ^ n753 ;
  assign n2904 = n1537 & n2903 ;
  assign n2906 = n2905 ^ n2904 ;
  assign n3800 = n2703 & n2906 ;
  assign n2897 = n2896 ^ n1310 ;
  assign n2898 = n2897 ^ n829 ;
  assign n2901 = n2900 ^ n2898 ;
  assign n3799 = ~n2702 & n2901 ;
  assign n3801 = n3800 ^ n3799 ;
  assign n3802 = n3801 ^ n753 ;
  assign n2859 = n2742 ^ n2716 ;
  assign n3797 = n1310 & ~n2859 ;
  assign n3803 = n3802 ^ n3797 ;
  assign n3805 = n3804 ^ n3803 ;
  assign n3844 = n3808 ^ n3805 ;
  assign n3845 = n3844 ^ n3804 ;
  assign n3846 = n3845 ^ n3801 ;
  assign n3838 = n3805 ^ n3797 ;
  assign n3798 = n3797 ^ n753 ;
  assign n3806 = n3805 ^ n3798 ;
  assign n3807 = n3806 ^ n3801 ;
  assign n3811 = n3808 ^ n3807 ;
  assign n3839 = n3838 ^ n3811 ;
  assign n3835 = n3804 ^ n3798 ;
  assign n3836 = n3835 ^ n3805 ;
  assign n3837 = n3836 ^ n3811 ;
  assign n3840 = n3839 ^ n3837 ;
  assign n3841 = n3840 ^ n3811 ;
  assign n3814 = n3804 ^ n753 ;
  assign n3815 = n3814 ^ n3801 ;
  assign n3816 = n3815 ^ n3805 ;
  assign n3809 = n3808 ^ n3804 ;
  assign n3818 = n3816 ^ n3809 ;
  assign n3819 = n3818 ^ n3801 ;
  assign n3820 = n3819 ^ n3808 ;
  assign n3823 = n3809 & ~n3815 ;
  assign n3821 = n3809 ^ n3808 ;
  assign n3825 = n3823 ^ n3821 ;
  assign n3826 = n3820 & n3825 ;
  assign n3831 = n3826 ^ n3823 ;
  assign n3827 = n3826 ^ n3808 ;
  assign n3829 = n3816 ^ n3815 ;
  assign n3830 = n3827 & ~n3829 ;
  assign n3832 = n3831 ^ n3830 ;
  assign n3833 = n3832 ^ n3815 ;
  assign n3834 = n3833 ^ n3821 ;
  assign n3842 = n3841 ^ n3834 ;
  assign n3843 = n3842 ^ n3808 ;
  assign n3847 = n3846 ^ n3843 ;
  assign n3848 = n3847 ^ n3808 ;
  assign n3146 = ~n696 & n799 ;
  assign n3147 = n3146 ^ n799 ;
  assign n3144 = n696 & ~n800 ;
  assign n3145 = n3144 ^ n800 ;
  assign n3148 = n3147 ^ n3145 ;
  assign n3149 = n739 & ~n3148 ;
  assign n3788 = n2706 & n3149 ;
  assign n3141 = n738 & n799 ;
  assign n3142 = n3141 ^ n2612 ;
  assign n3787 = n2705 & n3142 ;
  assign n3789 = n3788 ^ n3787 ;
  assign n2942 = n2739 ^ n2713 ;
  assign n3004 = n2942 ^ n2704 ;
  assign n3781 = n3004 ^ n2704 ;
  assign n3782 = n2704 ^ n739 ;
  assign n3783 = n3782 ^ n2704 ;
  assign n3784 = ~n3781 & n3783 ;
  assign n3785 = n3784 ^ n2704 ;
  assign n3786 = n754 & n3785 ;
  assign n3790 = n3789 ^ n3786 ;
  assign n3791 = n3790 ^ n2710 ;
  assign n3150 = n2707 & n3149 ;
  assign n3143 = ~n2710 & n3142 ;
  assign n3151 = n3150 ^ n3143 ;
  assign n3136 = n2706 ^ n739 ;
  assign n3137 = n3136 ^ n2706 ;
  assign n3138 = ~n2709 & n3137 ;
  assign n3139 = n3138 ^ n2706 ;
  assign n3140 = n754 & n3139 ;
  assign n3152 = n3151 ^ n3140 ;
  assign n3154 = n3145 ^ n799 ;
  assign n3155 = n799 ^ n738 ;
  assign n3156 = n2707 & ~n3155 ;
  assign n3157 = n3156 ^ n799 ;
  assign n3158 = ~n3154 & ~n3157 ;
  assign n3159 = n3158 ^ n799 ;
  assign n3160 = ~n2708 & ~n3159 ;
  assign n3412 = ~n3152 & ~n3160 ;
  assign n2921 = n2738 ^ n2712 ;
  assign n3414 = n2705 ^ n739 ;
  assign n3415 = n3414 ^ n2705 ;
  assign n3416 = ~n2921 & n3415 ;
  assign n3417 = n3416 ^ n2705 ;
  assign n3418 = n754 & ~n3417 ;
  assign n3428 = n3418 ^ n800 ;
  assign n5847 = n738 & ~n3145 ;
  assign n3427 = ~n2710 & n5847 ;
  assign n3429 = n3428 ^ n3427 ;
  assign n3419 = n3418 ^ n799 ;
  assign n3420 = n3419 ^ n3418 ;
  assign n3421 = ~n696 & n738 ;
  assign n3422 = n3421 ^ n739 ;
  assign n3423 = ~n2710 & n3422 ;
  assign n3424 = n3420 & n3423 ;
  assign n3425 = n3424 ^ n3419 ;
  assign n3430 = n3429 ^ n3425 ;
  assign n3431 = n3425 ^ n3418 ;
  assign n3432 = n3431 ^ n738 ;
  assign n3435 = ~n2706 & ~n3432 ;
  assign n3436 = n3435 ^ n738 ;
  assign n3437 = ~n3430 & ~n3436 ;
  assign n3438 = n3437 ^ n3429 ;
  assign n3775 = ~n3412 & ~n3438 ;
  assign n3776 = ~n696 & n3775 ;
  assign n3777 = n2707 & n3776 ;
  assign n3778 = n3777 ^ n3775 ;
  assign n3779 = n3778 ^ n3438 ;
  assign n3792 = n3791 ^ n3779 ;
  assign n3793 = n3792 ^ n3790 ;
  assign n3794 = n696 & n3779 ;
  assign n3795 = ~n3793 & n3794 ;
  assign n3796 = n3795 ^ n3792 ;
  assign n3849 = n3848 ^ n3796 ;
  assign n3413 = n3412 ^ n2707 ;
  assign n3439 = n3438 ^ n696 ;
  assign n3442 = n3412 & n3439 ;
  assign n3443 = n3442 ^ n696 ;
  assign n3444 = ~n3413 & ~n3443 ;
  assign n3445 = n3444 ^ n3438 ;
  assign n3066 = n2741 ^ n2715 ;
  assign n3408 = n1310 & ~n3066 ;
  assign n3409 = n2702 ^ n829 ;
  assign n3410 = n3408 & n3409 ;
  assign n3398 = n2704 & n2906 ;
  assign n3397 = n2703 & n2901 ;
  assign n3399 = n3398 ^ n3397 ;
  assign n3400 = n3399 ^ n753 ;
  assign n3403 = n3400 ^ n2702 ;
  assign n3404 = ~n3066 & n3403 ;
  assign n3405 = n3404 ^ n2702 ;
  assign n3406 = n1310 & ~n3405 ;
  assign n3407 = n3406 ^ n3400 ;
  assign n3411 = n3410 ^ n3407 ;
  assign n3446 = n3445 ^ n3411 ;
  assign n3161 = ~n696 & n3160 ;
  assign n2979 = n2740 ^ n2714 ;
  assign n3104 = n2705 & n2906 ;
  assign n3103 = n2704 & n2901 ;
  assign n3105 = n3104 ^ n3103 ;
  assign n3108 = ~n2979 & ~n3105 ;
  assign n3109 = n3108 ^ n1310 ;
  assign n3110 = ~n753 & n3109 ;
  assign n3111 = n3110 ^ n1310 ;
  assign n3118 = ~n829 & ~n2979 ;
  assign n3119 = n3118 ^ n2703 ;
  assign n3120 = n3111 & n3119 ;
  assign n3122 = ~n2703 & n2897 ;
  assign n3123 = ~n2979 & n3122 ;
  assign n3121 = n3066 ^ n2714 ;
  assign n3124 = n3123 ^ n3121 ;
  assign n3125 = n3124 ^ n3123 ;
  assign n3126 = n3123 ^ n1310 ;
  assign n3127 = n3126 ^ n3123 ;
  assign n3128 = n3125 & n3127 ;
  assign n3129 = n3128 ^ n3123 ;
  assign n3130 = n3105 ^ n753 ;
  assign n3131 = n3130 ^ n3105 ;
  assign n3132 = n3131 ^ n3123 ;
  assign n3133 = n3129 & ~n3132 ;
  assign n3134 = n3133 ^ n3130 ;
  assign n3135 = ~n3120 & n3134 ;
  assign n3153 = n3152 ^ n3135 ;
  assign n3162 = n3161 ^ n3153 ;
  assign n2967 = n2710 ^ n2707 ;
  assign n2968 = n2967 ^ n2710 ;
  assign n2969 = n2710 ^ n751 ;
  assign n2970 = n2969 ^ n2710 ;
  assign n2971 = n2968 & n2970 ;
  assign n2972 = n2971 ^ n2710 ;
  assign n2973 = ~n754 & ~n2972 ;
  assign n2974 = n2973 ^ n2710 ;
  assign n2966 = ~n738 & n2707 ;
  assign n2975 = n2974 ^ n2966 ;
  assign n2938 = n2706 & n2906 ;
  assign n2937 = n2705 & n2901 ;
  assign n2939 = n2938 ^ n2937 ;
  assign n2936 = n1310 & n2704 ;
  assign n2940 = n2939 ^ n2936 ;
  assign n2941 = n2940 ^ n2939 ;
  assign n2945 = n2941 & n2942 ;
  assign n2946 = n2945 ^ n2939 ;
  assign n2947 = ~n753 & n2946 ;
  assign n2949 = n2939 ^ n753 ;
  assign n2952 = n2949 ^ n2936 ;
  assign n2955 = n2952 ^ n2942 ;
  assign n2956 = n2955 ^ n2952 ;
  assign n2948 = n2704 ^ n829 ;
  assign n2953 = n2952 ^ n2948 ;
  assign n2957 = n2952 ^ n1310 ;
  assign n2958 = n2957 ^ n2952 ;
  assign n2961 = n2953 & n2958 ;
  assign n2962 = ~n2956 & n2961 ;
  assign n2963 = n2962 ^ n2956 ;
  assign n2964 = n2963 ^ n2955 ;
  assign n2965 = ~n2947 & ~n2964 ;
  assign n2976 = n2975 ^ n2965 ;
  assign n2888 = n754 & n2707 ;
  assign n2907 = n2707 & n2906 ;
  assign n2902 = ~n2710 & n2901 ;
  assign n2908 = n2907 ^ n2902 ;
  assign n2891 = n2706 ^ n1537 ;
  assign n2892 = n2891 ^ n2706 ;
  assign n2893 = ~n2709 & n2892 ;
  assign n2894 = n2893 ^ n2706 ;
  assign n2895 = n1310 & n2894 ;
  assign n2909 = n2908 ^ n2895 ;
  assign n2910 = n2506 ^ n830 ;
  assign n2911 = n1310 & n2910 ;
  assign n2912 = n2911 ^ n830 ;
  assign n2913 = n2707 ^ n1310 ;
  assign n2914 = n2913 ^ n753 ;
  assign n2915 = n2912 & ~n2914 ;
  assign n2916 = n2915 ^ n1310 ;
  assign n2917 = n753 & n2916 ;
  assign n2918 = n2917 ^ n753 ;
  assign n2919 = ~n2909 & n2918 ;
  assign n2920 = ~n2888 & ~n2919 ;
  assign n2930 = ~n2710 & n2906 ;
  assign n2929 = n2706 & n2901 ;
  assign n2931 = n2930 ^ n2929 ;
  assign n2932 = n2931 ^ n753 ;
  assign n2924 = n2705 ^ n1537 ;
  assign n2925 = n2924 ^ n2705 ;
  assign n2926 = ~n2921 & n2925 ;
  assign n2927 = n2926 ^ n2705 ;
  assign n2928 = n1310 & n2927 ;
  assign n2933 = n2932 ^ n2928 ;
  assign n2934 = n2920 & n2933 ;
  assign n2935 = n2934 ^ n2933 ;
  assign n3163 = n2975 ^ n2935 ;
  assign n3164 = n2976 & ~n3163 ;
  assign n3165 = n3164 ^ n2975 ;
  assign n3394 = n3165 ^ n3135 ;
  assign n3395 = n3162 & ~n3394 ;
  assign n3396 = n3395 ^ n3135 ;
  assign n3772 = n3411 ^ n3396 ;
  assign n3773 = n3446 & ~n3772 ;
  assign n3774 = n3773 ^ n3445 ;
  assign n3850 = n3849 ^ n3774 ;
  assign n3869 = n3868 ^ n3850 ;
  assign n3465 = n1773 & ~n2719 ;
  assign n3461 = n1021 & ~n3184 ;
  assign n3462 = n3461 ^ n2744 ;
  assign n3463 = n2865 & n3462 ;
  assign n3448 = n3184 ^ n2871 ;
  assign n3450 = n3184 ^ n2701 ;
  assign n3454 = ~n3448 & n3450 ;
  assign n3449 = n3448 ^ n2871 ;
  assign n3451 = n3450 ^ n1017 ;
  assign n3452 = n2865 & ~n3451 ;
  assign n3453 = ~n3449 & n3452 ;
  assign n3455 = n3454 ^ n3453 ;
  assign n3456 = n3455 ^ n1017 ;
  assign n3457 = n3456 ^ n2744 ;
  assign n3447 = n3446 ^ n3396 ;
  assign n3458 = n3457 ^ n3447 ;
  assign n3464 = n3463 ^ n3458 ;
  assign n3466 = n3465 ^ n3464 ;
  assign n3167 = ~n2855 & n2865 ;
  assign n3176 = n2989 & ~n3167 ;
  assign n3174 = n1773 & ~n2700 ;
  assign n3169 = n2855 ^ n2702 ;
  assign n3170 = n2871 & n3169 ;
  assign n3171 = n3170 ^ n2865 ;
  assign n3168 = n1021 & n3167 ;
  assign n3172 = n3171 ^ n3168 ;
  assign n3166 = n3165 ^ n3162 ;
  assign n3173 = n3172 ^ n3166 ;
  assign n3175 = n3174 ^ n3173 ;
  assign n3177 = n3176 ^ n3175 ;
  assign n3100 = ~n2701 & ~n2865 ;
  assign n3178 = n3177 ^ n3100 ;
  assign n2977 = n2976 ^ n2935 ;
  assign n2860 = n1773 & ~n2859 ;
  assign n2874 = n2701 ^ n1021 ;
  assign n2857 = n1773 & n2856 ;
  assign n2875 = n2874 ^ n2857 ;
  assign n2876 = ~n2860 & ~n2875 ;
  assign n2883 = n2876 ^ n2857 ;
  assign n2872 = n2703 & n2871 ;
  assign n2866 = ~n2702 & ~n2865 ;
  assign n2858 = n2857 ^ n1017 ;
  assign n2861 = n2860 ^ n2858 ;
  assign n2867 = n2866 ^ n2861 ;
  assign n2873 = n2872 ^ n2867 ;
  assign n2877 = n2876 ^ n2875 ;
  assign n2878 = n2877 ^ n2857 ;
  assign n2880 = ~n1017 & ~n2878 ;
  assign n2881 = n2880 ^ n2857 ;
  assign n2882 = n2873 & ~n2881 ;
  assign n2884 = n2883 ^ n2882 ;
  assign n2887 = n2884 ^ n2874 ;
  assign n2978 = n2977 ^ n2887 ;
  assign n3083 = n1773 & ~n2702 ;
  assign n3077 = n3066 ^ n2989 ;
  assign n3080 = ~n1017 & ~n3066 ;
  assign n3081 = n3077 & n3080 ;
  assign n3076 = n2704 ^ n2703 ;
  assign n3078 = n3077 ^ n3076 ;
  assign n3082 = n3081 ^ n3078 ;
  assign n3084 = n3083 ^ n3082 ;
  assign n3069 = n3066 ^ n2703 ;
  assign n3070 = n3069 ^ n2703 ;
  assign n3071 = n2703 ^ n1021 ;
  assign n3072 = n3071 ^ n2703 ;
  assign n3073 = ~n3070 & n3072 ;
  assign n3074 = n3073 ^ n2703 ;
  assign n3075 = n2865 & ~n3074 ;
  assign n3085 = n3084 ^ n3075 ;
  assign n3067 = n3066 ^ n2704 ;
  assign n3068 = ~n2871 & ~n3067 ;
  assign n3086 = n3085 ^ n3068 ;
  assign n3002 = n2917 ^ n2909 ;
  assign n2998 = n1773 & n2703 ;
  assign n2992 = n2705 ^ n2704 ;
  assign n2990 = n2989 ^ n2740 ;
  assign n2991 = n2990 ^ n2714 ;
  assign n2993 = n2992 ^ n2991 ;
  assign n2994 = n2993 ^ n2992 ;
  assign n2995 = n1017 & ~n2979 ;
  assign n2996 = ~n2994 & n2995 ;
  assign n2997 = n2996 ^ n2993 ;
  assign n2999 = n2998 ^ n2997 ;
  assign n2984 = n2704 ^ n1021 ;
  assign n2985 = n2984 ^ n2704 ;
  assign n2986 = ~n2979 & ~n2985 ;
  assign n2987 = n2986 ^ n2704 ;
  assign n2988 = n2865 & ~n2987 ;
  assign n3000 = n2999 ^ n2988 ;
  assign n2980 = n2979 ^ n2705 ;
  assign n2981 = ~n2871 & ~n2980 ;
  assign n3001 = n3000 ^ n2981 ;
  assign n3003 = n3002 ^ n3001 ;
  assign n3022 = n829 & n2707 ;
  assign n3018 = n827 & n2968 ;
  assign n3019 = n3018 ^ n2710 ;
  assign n3020 = ~n1310 & ~n3019 ;
  assign n3021 = n3020 ^ n2710 ;
  assign n3023 = n3022 ^ n3021 ;
  assign n3062 = n3023 ^ n3002 ;
  assign n3013 = n2706 & n2871 ;
  assign n3012 = n2705 & ~n2865 ;
  assign n3014 = n3013 ^ n3012 ;
  assign n3006 = n2984 ^ n1017 ;
  assign n3007 = n3006 ^ n2704 ;
  assign n3008 = ~n2942 & ~n3007 ;
  assign n3009 = n3008 ^ n2704 ;
  assign n3010 = n1773 & n3009 ;
  assign n3011 = n3010 ^ n1017 ;
  assign n3015 = n3014 ^ n3011 ;
  assign n3024 = n3023 ^ n3015 ;
  assign n3042 = n1310 & n2707 ;
  assign n3025 = n1773 & ~n2710 ;
  assign n3026 = n2864 ^ n2862 ;
  assign n3027 = n1017 & ~n3026 ;
  assign n3028 = ~n2707 & n3027 ;
  assign n3029 = ~n3025 & n3028 ;
  assign n3030 = n3029 ^ n3027 ;
  assign n3031 = n3030 ^ n1017 ;
  assign n3038 = n2707 & n2871 ;
  assign n3037 = ~n2710 & ~n2865 ;
  assign n3039 = n3038 ^ n3037 ;
  assign n3032 = n2706 ^ n1022 ;
  assign n3033 = n3032 ^ n2706 ;
  assign n3034 = ~n2709 & ~n3033 ;
  assign n3035 = n3034 ^ n2706 ;
  assign n3036 = n1773 & n3035 ;
  assign n3040 = n3039 ^ n3036 ;
  assign n3041 = n3031 & ~n3040 ;
  assign n3044 = n3042 ^ n3041 ;
  assign n3043 = n3041 & n3042 ;
  assign n3045 = n3044 ^ n3043 ;
  assign n3057 = n1773 & n2705 ;
  assign n3048 = n2865 & ~n2921 ;
  assign n3054 = n2921 ^ n1017 ;
  assign n3055 = ~n3048 & ~n3054 ;
  assign n3052 = n2706 & ~n2865 ;
  assign n3049 = n1021 & n3048 ;
  assign n3046 = n2921 ^ n2710 ;
  assign n3047 = ~n2871 & n3046 ;
  assign n3050 = n3049 ^ n3047 ;
  assign n3051 = n3050 ^ n2710 ;
  assign n3053 = n3052 ^ n3051 ;
  assign n3056 = n3055 ^ n3053 ;
  assign n3058 = n3057 ^ n3056 ;
  assign n3059 = n3045 & ~n3058 ;
  assign n3060 = n3059 ^ n3023 ;
  assign n3061 = ~n3024 & ~n3060 ;
  assign n3063 = n3062 ^ n3061 ;
  assign n3064 = ~n3003 & ~n3063 ;
  assign n3065 = n3064 ^ n3002 ;
  assign n3087 = n3086 ^ n3065 ;
  assign n3088 = n2919 ^ n2888 ;
  assign n3089 = n3088 ^ n2933 ;
  assign n3092 = n2919 & ~n2933 ;
  assign n3093 = ~n3089 & n3092 ;
  assign n3090 = n3089 ^ n3086 ;
  assign n3094 = n3093 ^ n3090 ;
  assign n3095 = ~n3087 & ~n3094 ;
  assign n3096 = n3095 ^ n3086 ;
  assign n3097 = n3096 ^ n2887 ;
  assign n3098 = ~n2978 & n3097 ;
  assign n3099 = n3098 ^ n2887 ;
  assign n3467 = n3166 ^ n3099 ;
  assign n3468 = ~n3178 & n3467 ;
  assign n3469 = n3468 ^ n3166 ;
  assign n3769 = n3469 ^ n3447 ;
  assign n3770 = n3466 & ~n3769 ;
  assign n3771 = n3770 ^ n3447 ;
  assign n3870 = n3869 ^ n3771 ;
  assign n3758 = n2796 & n2820 ;
  assign n3753 = n3688 ^ n2732 ;
  assign n3754 = n3753 ^ n2737 ;
  assign n3755 = ~n3189 & n3754 ;
  assign n3751 = n2796 ^ n1581 ;
  assign n3752 = n3751 ^ n2737 ;
  assign n3756 = n3755 ^ n3752 ;
  assign n3748 = ~n1581 & ~n2796 ;
  assign n3749 = n3748 ^ n2792 ;
  assign n3750 = n2737 & ~n3749 ;
  assign n3757 = n3756 ^ n3750 ;
  assign n3759 = n3758 ^ n3757 ;
  assign n3760 = n2659 ^ n1483 ;
  assign n2811 = n2746 ^ n2730 ;
  assign n2812 = n2811 ^ n2747 ;
  assign n2813 = n2812 ^ n2746 ;
  assign n2814 = n2736 ^ n411 ;
  assign n2815 = n2813 & ~n2814 ;
  assign n3761 = n3760 ^ n2815 ;
  assign n3762 = n3761 ^ n3760 ;
  assign n3763 = n1581 & ~n2659 ;
  assign n3764 = n3763 ^ n3760 ;
  assign n3765 = ~n3762 & n3764 ;
  assign n3766 = n3765 ^ n3760 ;
  assign n3767 = ~n2789 & n3766 ;
  assign n3768 = n3759 & ~n3767 ;
  assign n3871 = n3870 ^ n3768 ;
  assign n4145 = n3848 ^ n3774 ;
  assign n4146 = n3796 ^ n3774 ;
  assign n4147 = n4145 & n4146 ;
  assign n4148 = n4147 ^ n3848 ;
  assign n4140 = n2705 & n3149 ;
  assign n4139 = n2704 & n3142 ;
  assign n4141 = n4140 ^ n4139 ;
  assign n4136 = n739 & ~n2979 ;
  assign n4137 = n4136 ^ n2703 ;
  assign n4138 = n754 & n4137 ;
  assign n4142 = n4141 ^ n4138 ;
  assign n4131 = n2710 ^ n2706 ;
  assign n4129 = n3790 ^ n3779 ;
  assign n4130 = n3791 & ~n4129 ;
  assign n4132 = n4131 ^ n4130 ;
  assign n4133 = ~n696 & n4132 ;
  assign n4143 = n4142 ^ n4133 ;
  assign n4088 = n2700 ^ n829 ;
  assign n3230 = n3184 ^ n2743 ;
  assign n4084 = n1310 & n3230 ;
  assign n4080 = ~n2702 & n2906 ;
  assign n4079 = ~n2701 & n2901 ;
  assign n4081 = n4080 ^ n4079 ;
  assign n4082 = n4081 ^ n753 ;
  assign n4077 = n1310 & ~n2855 ;
  assign n4083 = n4082 ^ n4077 ;
  assign n4085 = n4084 ^ n4083 ;
  assign n4124 = n4088 ^ n4085 ;
  assign n4125 = n4124 ^ n4084 ;
  assign n4126 = n4125 ^ n4081 ;
  assign n4118 = n4085 ^ n4077 ;
  assign n4078 = n4077 ^ n753 ;
  assign n4086 = n4085 ^ n4078 ;
  assign n4087 = n4086 ^ n4081 ;
  assign n4091 = n4088 ^ n4087 ;
  assign n4119 = n4118 ^ n4091 ;
  assign n4115 = n4084 ^ n4078 ;
  assign n4116 = n4115 ^ n4085 ;
  assign n4117 = n4116 ^ n4091 ;
  assign n4120 = n4119 ^ n4117 ;
  assign n4121 = n4120 ^ n4091 ;
  assign n4094 = n4084 ^ n753 ;
  assign n4095 = n4094 ^ n4081 ;
  assign n4096 = n4095 ^ n4085 ;
  assign n4089 = n4088 ^ n4084 ;
  assign n4098 = n4096 ^ n4089 ;
  assign n4099 = n4098 ^ n4081 ;
  assign n4100 = n4099 ^ n4088 ;
  assign n4103 = n4089 & ~n4095 ;
  assign n4101 = n4089 ^ n4088 ;
  assign n4105 = n4103 ^ n4101 ;
  assign n4106 = n4100 & n4105 ;
  assign n4111 = n4106 ^ n4103 ;
  assign n4107 = n4106 ^ n4088 ;
  assign n4109 = n4096 ^ n4095 ;
  assign n4110 = n4107 & ~n4109 ;
  assign n4112 = n4111 ^ n4110 ;
  assign n4113 = n4112 ^ n4095 ;
  assign n4114 = n4113 ^ n4101 ;
  assign n4122 = n4121 ^ n4114 ;
  assign n4123 = n4122 ^ n4088 ;
  assign n4127 = n4126 ^ n4123 ;
  assign n4128 = n4127 ^ n4088 ;
  assign n4144 = n4143 ^ n4128 ;
  assign n4149 = n4148 ^ n4144 ;
  assign n4074 = n3868 ^ n3771 ;
  assign n4075 = n3869 & ~n4074 ;
  assign n4076 = n4075 ^ n3868 ;
  assign n4150 = n4149 ^ n4076 ;
  assign n2836 = n2746 ^ n2722 ;
  assign n4069 = n2836 ^ n2719 ;
  assign n4070 = n2871 & n4069 ;
  assign n4066 = n1773 & n2737 ;
  assign n4061 = n2836 & n2865 ;
  assign n4064 = n4061 ^ n2865 ;
  assign n4065 = ~n1017 & ~n4064 ;
  assign n4067 = n4066 ^ n4065 ;
  assign n4068 = n4067 ^ n2865 ;
  assign n4071 = n4070 ^ n4068 ;
  assign n4062 = ~n1021 & n2865 ;
  assign n4063 = ~n4061 & ~n4062 ;
  assign n4072 = n4071 ^ n4063 ;
  assign n4060 = ~n2721 & ~n2865 ;
  assign n4073 = n4072 ^ n4060 ;
  assign n4151 = n4150 ^ n4073 ;
  assign n4152 = n4151 ^ n3768 ;
  assign n4153 = n4152 ^ n4151 ;
  assign n3470 = n3469 ^ n3466 ;
  assign n3179 = n3178 ^ n3099 ;
  assign n2842 = n2721 ^ n1581 ;
  assign n2844 = n2796 & n2842 ;
  assign n2845 = n2844 ^ n2805 ;
  assign n2851 = n2719 & n2803 ;
  assign n2852 = n2851 ^ n2792 ;
  assign n2853 = ~n2845 & ~n2852 ;
  assign n2782 = n2737 ^ n1483 ;
  assign n2834 = n2782 ^ n1835 ;
  assign n2835 = n2834 ^ n2782 ;
  assign n2839 = n2835 & n2836 ;
  assign n2840 = n2839 ^ n2782 ;
  assign n2841 = ~n2789 & ~n2840 ;
  assign n2854 = n2853 ^ n2841 ;
  assign n3180 = n3179 ^ n2854 ;
  assign n3211 = n3096 ^ n2978 ;
  assign n3190 = n2836 ^ n2720 ;
  assign n3191 = ~n3189 & ~n3190 ;
  assign n3181 = n2721 ^ n1483 ;
  assign n3187 = ~n2789 & ~n3186 ;
  assign n3188 = ~n3181 & n3187 ;
  assign n3192 = n3191 ^ n3188 ;
  assign n3201 = ~n2700 & n2806 ;
  assign n3200 = ~n2719 & ~n2793 ;
  assign n3202 = n3201 ^ n3200 ;
  assign n3203 = n3202 ^ n1581 ;
  assign n3193 = n2719 ^ n1483 ;
  assign n3194 = n3193 ^ n2719 ;
  assign n3195 = n1581 & ~n2700 ;
  assign n3196 = n3195 ^ n2719 ;
  assign n3197 = ~n3194 & ~n3196 ;
  assign n3198 = n3197 ^ n2719 ;
  assign n3199 = ~n2781 & ~n3198 ;
  assign n3204 = n3203 ^ n3199 ;
  assign n3205 = ~n3192 & n3204 ;
  assign n3209 = n3205 ^ n3192 ;
  assign n3206 = n3190 ^ n3186 ;
  assign n3207 = n3206 & n3229 ;
  assign n3208 = n3205 & n3207 ;
  assign n3210 = n3209 ^ n3208 ;
  assign n3212 = n3211 ^ n3210 ;
  assign n3225 = n3094 ^ n3065 ;
  assign n3214 = ~n2701 & n2803 ;
  assign n3213 = ~n2700 & n2796 ;
  assign n3215 = n3214 ^ n3213 ;
  assign n3223 = n3215 ^ n1581 ;
  assign n3218 = n3193 ^ n1581 ;
  assign n3219 = ~n3184 & ~n3218 ;
  assign n3216 = ~n1581 & n3215 ;
  assign n3217 = n3185 & n3216 ;
  assign n3220 = n3219 ^ n3217 ;
  assign n3221 = n3220 ^ n3183 ;
  assign n3222 = ~n2789 & ~n3221 ;
  assign n3224 = n3223 ^ n3222 ;
  assign n3226 = n3225 ^ n3224 ;
  assign n3243 = n3063 ^ n3001 ;
  assign n3232 = ~n2702 & n2803 ;
  assign n3231 = ~n2701 & n2796 ;
  assign n3233 = n3232 ^ n3231 ;
  assign n3239 = n3233 ^ n1581 ;
  assign n3236 = ~n2789 & ~n2855 ;
  assign n3237 = n2700 ^ n1483 ;
  assign n3238 = n3236 & ~n3237 ;
  assign n3240 = n3239 ^ n3238 ;
  assign n3234 = n3230 & ~n3233 ;
  assign n3235 = n3229 & n3234 ;
  assign n3241 = n3240 ^ n3235 ;
  assign n3227 = n3184 ^ n2717 ;
  assign n3228 = ~n3189 & ~n3227 ;
  assign n3242 = n3241 ^ n3228 ;
  assign n3244 = n3243 ^ n3242 ;
  assign n3261 = ~n2789 & ~n2859 ;
  assign n3262 = n2701 ^ n1483 ;
  assign n3263 = n3261 & n3262 ;
  assign n3249 = n2855 ^ n2742 ;
  assign n3250 = n3229 & ~n3249 ;
  assign n3247 = n2703 & n2803 ;
  assign n3246 = ~n2702 & n2796 ;
  assign n3248 = n3247 ^ n3246 ;
  assign n3251 = n3250 ^ n3248 ;
  assign n3252 = ~n2789 & n2856 ;
  assign n3253 = n3252 ^ n3250 ;
  assign n3254 = ~n3251 & n3253 ;
  assign n3255 = n3254 ^ n3250 ;
  assign n3256 = n3250 ^ n1581 ;
  assign n3257 = n3256 ^ n3248 ;
  assign n3258 = n3257 ^ n3250 ;
  assign n3259 = n3255 & ~n3258 ;
  assign n3260 = n3259 ^ n3257 ;
  assign n3264 = n3263 ^ n3260 ;
  assign n3245 = n3060 ^ n3015 ;
  assign n3265 = n3264 ^ n3245 ;
  assign n3293 = n3058 ^ n3045 ;
  assign n3294 = n3293 ^ n3043 ;
  assign n3266 = n2859 ^ n2741 ;
  assign n3268 = n2704 & n2803 ;
  assign n3267 = n2703 & n2796 ;
  assign n3269 = n3268 ^ n3267 ;
  assign n3270 = n3269 ^ n1581 ;
  assign n3271 = n3270 ^ n2801 ;
  assign n3272 = n3271 ^ n3269 ;
  assign n3273 = n3266 & n3272 ;
  assign n3274 = n3273 ^ n3270 ;
  assign n3279 = ~n3066 & ~n3269 ;
  assign n3280 = n3279 ^ n2789 ;
  assign n3281 = n1581 & ~n3280 ;
  assign n3282 = n3281 ^ n2789 ;
  assign n3283 = n2702 ^ n1483 ;
  assign n3284 = n3283 ^ n2702 ;
  assign n3289 = ~n3066 & n3284 ;
  assign n3290 = n3289 ^ n2702 ;
  assign n3291 = ~n3282 & ~n3290 ;
  assign n3292 = ~n3274 & ~n3291 ;
  assign n3295 = n3294 ^ n3292 ;
  assign n3310 = n3040 ^ n3030 ;
  assign n3297 = n2705 & n2803 ;
  assign n3296 = n2704 & n2796 ;
  assign n3298 = n3297 ^ n3296 ;
  assign n3307 = n3121 & n3229 ;
  assign n3308 = ~n3298 & n3307 ;
  assign n3304 = n3066 ^ n2740 ;
  assign n3305 = ~n3189 & ~n3304 ;
  assign n3300 = ~n2789 & ~n2979 ;
  assign n3301 = n2703 ^ n1483 ;
  assign n3302 = n3300 & n3301 ;
  assign n3299 = n3298 ^ n1581 ;
  assign n3303 = n3302 ^ n3299 ;
  assign n3306 = n3305 ^ n3303 ;
  assign n3309 = n3308 ^ n3306 ;
  assign n3311 = n3310 ^ n3309 ;
  assign n3330 = n2862 ^ n1021 ;
  assign n3331 = n2707 & ~n3330 ;
  assign n3332 = n3331 ^ n3025 ;
  assign n3325 = n2705 ^ n1581 ;
  assign n3313 = n2704 ^ n1483 ;
  assign n3312 = n2704 ^ n1581 ;
  assign n3314 = n3313 ^ n3312 ;
  assign n3315 = ~n2942 & n3314 ;
  assign n3316 = n3315 ^ n3312 ;
  assign n3326 = n3325 ^ n3316 ;
  assign n3317 = n2705 ^ n1468 ;
  assign n3318 = n3317 ^ n1581 ;
  assign n3319 = n3318 ^ n2705 ;
  assign n3322 = n2706 & ~n3319 ;
  assign n3323 = n3322 ^ n2705 ;
  assign n3324 = n1484 & n3323 ;
  assign n3327 = n3326 ^ n3324 ;
  assign n3328 = n2789 & n3327 ;
  assign n3329 = n3328 ^ n3316 ;
  assign n3333 = n3332 ^ n3329 ;
  assign n3340 = ~n2710 & n2803 ;
  assign n3339 = n2706 & n2796 ;
  assign n3341 = n3340 ^ n3339 ;
  assign n3334 = n2705 ^ n1835 ;
  assign n3335 = n3334 ^ n2705 ;
  assign n3336 = ~n2921 & n3335 ;
  assign n3337 = n3336 ^ n2705 ;
  assign n3338 = ~n2789 & n3337 ;
  assign n3342 = n3341 ^ n3338 ;
  assign n3343 = n2710 ^ n1835 ;
  assign n3344 = n3343 ^ n2710 ;
  assign n3345 = n2968 & n3344 ;
  assign n3346 = n3345 ^ n2710 ;
  assign n3347 = n1484 & ~n3346 ;
  assign n3348 = n3347 ^ n2710 ;
  assign n3349 = n3348 ^ n2706 ;
  assign n3350 = n3349 ^ n1835 ;
  assign n3351 = n3350 ^ n3349 ;
  assign n3352 = n3349 ^ n2709 ;
  assign n3353 = n3352 ^ n3349 ;
  assign n3354 = n3351 & ~n3353 ;
  assign n3355 = n3354 ^ n3349 ;
  assign n3356 = ~n2789 & ~n3355 ;
  assign n3357 = n3356 ^ n3348 ;
  assign n3358 = n1581 & n3357 ;
  assign n3359 = ~n2708 & ~n2797 ;
  assign n3360 = n3358 & n3359 ;
  assign n3361 = n3360 ^ n3358 ;
  assign n3362 = ~n3342 & ~n3361 ;
  assign n3367 = n3362 ^ n1177 ;
  assign n3368 = n1773 & n2707 ;
  assign n3369 = n3367 & n3368 ;
  assign n3364 = n3342 ^ n1581 ;
  assign n3363 = n3362 ^ n1581 ;
  assign n3365 = n3364 ^ n3363 ;
  assign n3366 = n3365 ^ n3332 ;
  assign n3370 = n3369 ^ n3366 ;
  assign n3371 = n3333 & ~n3370 ;
  assign n3372 = n3371 ^ n3332 ;
  assign n3373 = n3372 ^ n3309 ;
  assign n3374 = n3311 & ~n3373 ;
  assign n3375 = n3374 ^ n3310 ;
  assign n3376 = n3375 ^ n3292 ;
  assign n3377 = n3295 & n3376 ;
  assign n3378 = n3377 ^ n3294 ;
  assign n3379 = n3378 ^ n3245 ;
  assign n3380 = ~n3265 & ~n3379 ;
  assign n3381 = n3380 ^ n3264 ;
  assign n3382 = n3381 ^ n3242 ;
  assign n3383 = n3244 & ~n3382 ;
  assign n3384 = n3383 ^ n3243 ;
  assign n3385 = n3384 ^ n3224 ;
  assign n3386 = ~n3226 & ~n3385 ;
  assign n3387 = n3386 ^ n3225 ;
  assign n3388 = n3387 ^ n3210 ;
  assign n3389 = n3212 & ~n3388 ;
  assign n3390 = n3389 ^ n3210 ;
  assign n3391 = n3390 ^ n2854 ;
  assign n3392 = n3180 & ~n3391 ;
  assign n3393 = n3392 ^ n3179 ;
  assign n3471 = n3470 ^ n3393 ;
  assign n2819 = ~n2789 & ~n2813 ;
  assign n2821 = n2820 ^ n1483 ;
  assign n2807 = ~n2721 & n2806 ;
  assign n2794 = n2737 & ~n2793 ;
  assign n2808 = n2807 ^ n2794 ;
  assign n2783 = n2782 ^ n2737 ;
  assign n2784 = n1581 & ~n2721 ;
  assign n2785 = n2784 ^ n2737 ;
  assign n2786 = ~n2783 & n2785 ;
  assign n2787 = n2786 ^ n2737 ;
  assign n2788 = ~n2781 & n2787 ;
  assign n2809 = n2808 ^ n2788 ;
  assign n2822 = n2809 ^ n1581 ;
  assign n2810 = ~n1581 & ~n2809 ;
  assign n2823 = n2822 ^ n2810 ;
  assign n2824 = n2821 & n2823 ;
  assign n2825 = n2819 & n2824 ;
  assign n2826 = n2825 ^ n2823 ;
  assign n2831 = n2826 ^ n2810 ;
  assign n2816 = n2815 ^ n2747 ;
  assign n2828 = n2816 ^ n2813 ;
  assign n2829 = n2828 & n3229 ;
  assign n2830 = n2826 & n2829 ;
  assign n2832 = n2831 ^ n2830 ;
  assign n2817 = ~n2789 & ~n2816 ;
  assign n2818 = n2810 & n2817 ;
  assign n2833 = n2832 ^ n2818 ;
  assign n3742 = n3393 ^ n2833 ;
  assign n3743 = n3471 & n3742 ;
  assign n3744 = n3743 ^ n2833 ;
  assign n4154 = n4153 ^ n3744 ;
  assign n4155 = n3871 & n4154 ;
  assign n4156 = n4155 ^ n4152 ;
  assign n4180 = n4179 ^ n4156 ;
  assign n2673 = n333 ^ n96 ;
  assign n2674 = n63 & n2673 ;
  assign n2675 = n2674 ^ n276 ;
  assign n2683 = n101 ^ n60 ;
  assign n2684 = n273 ^ n201 ;
  assign n2685 = ~n2683 & n2684 ;
  assign n2679 = n579 ^ n162 ;
  assign n2677 = n1100 ^ n343 ;
  assign n2676 = ~n64 & n255 ;
  assign n2678 = n2677 ^ n2676 ;
  assign n2680 = n2679 ^ n2678 ;
  assign n2681 = n2680 ^ n706 ;
  assign n2682 = n2681 ^ n725 ;
  assign n2686 = n2685 ^ n2682 ;
  assign n2687 = n2675 & ~n2686 ;
  assign n2688 = n278 & ~n2661 ;
  assign n3713 = n2687 & ~n2688 ;
  assign n3716 = n3713 ^ n2687 ;
  assign n3724 = n390 ^ n208 ;
  assign n3725 = n3724 ^ n719 ;
  assign n3723 = n2675 ^ n140 ;
  assign n3726 = n3725 ^ n3723 ;
  assign n3721 = n1105 ^ n139 ;
  assign n3722 = n58 & n3721 ;
  assign n3727 = n3726 ^ n3722 ;
  assign n3717 = n550 ^ n195 ;
  assign n3718 = n3717 ^ n520 ;
  assign n3719 = n63 & n3718 ;
  assign n3720 = ~n2550 & ~n3719 ;
  assign n3728 = n3727 ^ n3720 ;
  assign n3729 = ~n3716 & n3728 ;
  assign n2689 = n2688 ^ n2687 ;
  assign n4048 = n3729 ^ n2689 ;
  assign n4049 = n4048 ^ x2 ;
  assign n4050 = n4049 ^ n4048 ;
  assign n2753 = ~n278 & ~n2752 ;
  assign n3714 = ~n2753 & n3713 ;
  assign n4043 = ~n3714 & n3729 ;
  assign n2734 = n278 & ~n2733 ;
  assign n3710 = n2734 ^ n2688 ;
  assign n3711 = ~n2687 & ~n3710 ;
  assign n3712 = n3711 ^ n2688 ;
  assign n4042 = ~n3712 & ~n3728 ;
  assign n4044 = n4043 ^ n4042 ;
  assign n4045 = n27 & ~n4044 ;
  assign n4032 = n835 ^ n602 ;
  assign n4033 = ~n98 & n4032 ;
  assign n4029 = n205 ^ n146 ;
  assign n4030 = n4029 ^ n357 ;
  assign n4028 = n850 ^ n312 ;
  assign n4031 = n4030 ^ n4028 ;
  assign n4034 = n4033 ^ n4031 ;
  assign n4035 = n1249 & ~n4034 ;
  assign n4036 = n570 ^ n401 ;
  assign n4037 = n4036 ^ n218 ;
  assign n4038 = n4035 & ~n4037 ;
  assign n4039 = n111 & n3718 ;
  assign n4040 = n4038 & n4039 ;
  assign n4041 = n4040 ^ n4038 ;
  assign n4046 = n4045 ^ n4041 ;
  assign n4051 = n4046 ^ n3729 ;
  assign n4052 = n4051 ^ n4046 ;
  assign n4053 = n4052 ^ n4048 ;
  assign n4054 = ~n4050 & ~n4053 ;
  assign n4055 = n4054 ^ n4048 ;
  assign n4056 = ~x1 & ~n4055 ;
  assign n4057 = n4056 ^ n4051 ;
  assign n4058 = ~x0 & ~n4057 ;
  assign n4047 = ~n4574 ^ n4046 ;
  assign n4059 = n4058 ^ n4047 ;
  assign n4181 = n4180 ^ n4059 ;
  assign n3872 = n3871 ^ n3744 ;
  assign n2768 = x0 & n27 ;
  assign n2763 = n2761 ^ x0 ;
  assign n2764 = n2763 ^ x1 ;
  assign n2765 = n2764 ^ n28 ;
  assign n2762 = x2 & n2761 ;
  assign n2766 = n2765 ^ n2762 ;
  assign n2767 = ~n1465 & n2766 ;
  assign n2769 = n2768 ^ n2767 ;
  assign n2770 = n2769 ^ n1465 ;
  assign n3738 = n3737 ^ n2770 ;
  assign n3734 = ~n2662 & ~n3502 ;
  assign n3531 = n2768 ^ x0 ;
  assign n3733 = n3531 & n3729 ;
  assign n3735 = n3734 ^ n3733 ;
  assign n2773 = n2772 ^ n2770 ;
  assign n3736 = n3735 ^ n2773 ;
  assign n3739 = n3738 ^ n3736 ;
  assign n3732 = n28 & ~n2689 ;
  assign n3740 = n3739 ^ n3732 ;
  assign n3715 = n3714 ^ n3712 ;
  assign n3730 = n3729 ^ n3715 ;
  assign n3731 = n2768 & n3730 ;
  assign n3741 = n3740 ^ n3731 ;
  assign n3873 = n3872 ^ n3741 ;
  assign n3472 = n3471 ^ n2833 ;
  assign n2754 = n2753 ^ n2734 ;
  assign n2755 = n27 & n2754 ;
  assign n2672 = x22 ^ x1 ;
  assign n2690 = n2689 ^ n2672 ;
  assign n2756 = n2755 ^ n2690 ;
  assign n2671 = n2662 ^ n1460 ;
  assign n2757 = n2756 ^ n2671 ;
  assign n2663 = n2662 ^ x22 ;
  assign n2664 = n2663 ^ n2659 ;
  assign n2665 = n2664 ^ n2663 ;
  assign n2668 = x2 & ~n2665 ;
  assign n2669 = n2668 ^ n2663 ;
  assign n2670 = ~x1 & ~n2669 ;
  assign n2758 = n2757 ^ n2670 ;
  assign n2759 = ~x0 & ~n2758 ;
  assign n2760 = n2759 ^ n2756 ;
  assign n3473 = n3472 ^ n2760 ;
  assign n3685 = n3390 ^ n3180 ;
  assign n3686 = n3685 ^ n3472 ;
  assign n3668 = n2737 ^ n1460 ;
  assign n3666 = ~n4574 ^ n2820 ;
  assign n3665 = n27 & ~n2813 ;
  assign n3667 = n3666 ^ n3665 ;
  assign n3669 = n3668 ^ n3667 ;
  assign n3657 = n2737 ^ x22 ;
  assign n3658 = n3657 ^ n2721 ;
  assign n3659 = n3658 ^ n3657 ;
  assign n3662 = x2 & ~n3659 ;
  assign n3663 = n3662 ^ n3657 ;
  assign n3664 = ~x1 & ~n3663 ;
  assign n3670 = n3669 ^ n3664 ;
  assign n3671 = ~x0 & n3670 ;
  assign n3672 = n3671 ^ n3667 ;
  assign n3489 = n3381 ^ n3244 ;
  assign n3673 = n3672 ^ n3489 ;
  assign n3503 = ~n2701 & ~n3502 ;
  assign n3491 = n3375 ^ n3295 ;
  assign n3501 = ~n4574 ^ n3491 ;
  assign n3504 = n3503 ^ n3501 ;
  assign n3500 = n28 & ~n2700 ;
  assign n3505 = n3504 ^ n3500 ;
  assign n3497 = n27 & ~n3184 ;
  assign n3498 = n3497 ^ n2719 ;
  assign n3499 = x0 & ~n3498 ;
  assign n3506 = n3505 ^ n3499 ;
  assign n3521 = n2703 & ~n3502 ;
  assign n3519 = n28 & ~n2702 ;
  assign n3517 = n3370 ^ n3329 ;
  assign n3518 = ~n4574 ^ n3517 ;
  assign n3520 = n3519 ^ n3518 ;
  assign n3522 = n3521 ^ n3520 ;
  assign n3510 = n2859 ^ n2701 ;
  assign n3511 = n3510 ^ n2701 ;
  assign n3514 = n27 & ~n3511 ;
  assign n3515 = n3514 ^ n2701 ;
  assign n3516 = x0 & ~n3515 ;
  assign n3523 = n3522 ^ n3516 ;
  assign n3542 = n28 & n2704 ;
  assign n3533 = n3357 ^ n2802 ;
  assign n3534 = n3533 ^ n3357 ;
  assign n3535 = ~n2710 & ~n2789 ;
  assign n3536 = ~n2707 & ~n3535 ;
  assign n3537 = n3534 & n3536 ;
  assign n3538 = n3537 ^ n3533 ;
  assign n3539 = ~n4574 ^ n3538 ;
  assign n3532 = n2703 & n3531 ;
  assign n3540 = n3539 ^ n3532 ;
  assign n3530 = n2705 & ~n3502 ;
  assign n3541 = n3540 ^ n3530 ;
  assign n3543 = n3542 ^ n3541 ;
  assign n3112 = n2979 ^ n2703 ;
  assign n3529 = n2768 & ~n3112 ;
  assign n3544 = n3543 ^ n3529 ;
  assign n3550 = n2780 ^ n1468 ;
  assign n3551 = n3550 ^ n1483 ;
  assign n3552 = n2707 & ~n3551 ;
  assign n3553 = n3552 ^ n3535 ;
  assign n3524 = n3367 ^ n3361 ;
  assign n3525 = n3524 ^ n3364 ;
  assign n3526 = ~n2707 & ~n3525 ;
  assign n3527 = n3526 ^ n3367 ;
  assign n3586 = n3553 ^ n3527 ;
  assign n3557 = n2704 & n3531 ;
  assign n2776 = n2775 ^ n1464 ;
  assign n2777 = n2776 ^ n2773 ;
  assign n2778 = n2777 ^ n2767 ;
  assign n3549 = n2778 ^ x0 ;
  assign n3554 = n3553 ^ n3549 ;
  assign n3320 = n2706 ^ n2705 ;
  assign n3548 = n28 & n3320 ;
  assign n3555 = n3554 ^ n3548 ;
  assign n3546 = n30 ^ x0 ;
  assign n3547 = ~n2706 & ~n3546 ;
  assign n3556 = n3555 ^ n3547 ;
  assign n3558 = n3557 ^ n3556 ;
  assign n3545 = n2768 & ~n3004 ;
  assign n3559 = n3558 ^ n3545 ;
  assign n3571 = n2506 & ~n2706 ;
  assign n3572 = n3571 ^ n1468 ;
  assign n3573 = ~n2707 & n3572 ;
  assign n3574 = n3573 ^ n1468 ;
  assign n3575 = n3574 & ~n4574 ;
  assign n3583 = n3575 ^ n3553 ;
  assign n3566 = ~n2710 & ~n3502 ;
  assign n3565 = n28 & n2706 ;
  assign n3567 = n3566 ^ n3565 ;
  assign n3562 = n27 & ~n2921 ;
  assign n3563 = n3562 ^ n2705 ;
  assign n3564 = x0 & n3563 ;
  assign n3568 = n3567 ^ n3564 ;
  assign n3576 = n3575 ^ n2780 ;
  assign n3577 = n3576 ^ n3575 ;
  assign n3580 = n2707 & n3577 ;
  assign n3581 = n3580 ^ n3575 ;
  assign n3582 = n3568 & n3581 ;
  assign n3584 = n3583 ^ n3582 ;
  assign n3585 = ~n3559 & n3584 ;
  assign n3587 = n3586 ^ n3585 ;
  assign n3588 = n3587 ^ n3527 ;
  assign n3589 = n3588 ^ n3538 ;
  assign n3590 = n3544 & ~n3589 ;
  assign n3591 = n3590 ^ n3587 ;
  assign n3285 = n3066 ^ n2702 ;
  assign n3599 = n2768 & n3285 ;
  assign n3595 = ~n4574 ^ n3527 ;
  assign n3594 = n2704 & ~n3502 ;
  assign n3596 = n3595 ^ n3594 ;
  assign n3593 = ~n2702 & n3531 ;
  assign n3597 = n3596 ^ n3593 ;
  assign n3592 = n28 & n2703 ;
  assign n3598 = n3597 ^ n3592 ;
  assign n3600 = n3599 ^ n3598 ;
  assign n3601 = ~n3591 & ~n3600 ;
  assign n3528 = n3527 ^ n3517 ;
  assign n3602 = n3601 ^ n3528 ;
  assign n3603 = ~n3523 & n3602 ;
  assign n3604 = n3603 ^ n3517 ;
  assign n3621 = n3604 ^ n3491 ;
  assign n3612 = x2 & ~n2702 ;
  assign n3613 = n3612 ^ n2701 ;
  assign n3614 = ~x1 & ~n3613 ;
  assign n3507 = n27 & ~n2855 ;
  assign n3508 = n3507 ^ n2700 ;
  assign n3606 = n3508 ^ n2701 ;
  assign n3615 = n3614 ^ n3606 ;
  assign n3616 = ~x0 & n3615 ;
  assign n3509 = ~n4574 ^ n3508 ;
  assign n3605 = n3604 ^ n3509 ;
  assign n3617 = n3616 ^ n3605 ;
  assign n3618 = n3604 ^ n3372 ;
  assign n3619 = n3618 ^ n3311 ;
  assign n3620 = n3617 & ~n3619 ;
  assign n3622 = n3621 ^ n3620 ;
  assign n3623 = n3506 & ~n3622 ;
  assign n3488 = n3378 ^ n3265 ;
  assign n3492 = n3491 ^ n3488 ;
  assign n3624 = n3623 ^ n3492 ;
  assign n3635 = ~n2700 & ~n3502 ;
  assign n3633 = n28 & ~n2719 ;
  assign n3632 = ~n4574 ^ n3488 ;
  assign n3634 = n3633 ^ n3632 ;
  assign n3636 = n3635 ^ n3634 ;
  assign n3629 = n27 & ~n3186 ;
  assign n3630 = n3629 ^ n2721 ;
  assign n3631 = x0 & ~n3630 ;
  assign n3637 = n3636 ^ n3631 ;
  assign n3638 = n3624 & n3637 ;
  assign n3490 = n3489 ^ n3488 ;
  assign n3639 = n3638 ^ n3490 ;
  assign n3648 = n2721 ^ n2719 ;
  assign n3649 = n3648 ^ n2721 ;
  assign n3650 = x2 & ~n3649 ;
  assign n3651 = n3650 ^ n2721 ;
  assign n3652 = ~x1 & ~n3651 ;
  assign n3641 = n27 & ~n2836 ;
  assign n3642 = n3641 ^ n2737 ;
  assign n3644 = n3642 ^ n2721 ;
  assign n3653 = n3652 ^ n3644 ;
  assign n3654 = ~x0 & ~n3653 ;
  assign n3640 = ~n4574 ^ n3489 ;
  assign n3643 = n3642 ^ n3640 ;
  assign n3655 = n3654 ^ n3643 ;
  assign n3656 = n3639 & n3655 ;
  assign n3674 = n3673 ^ n3656 ;
  assign n3675 = n3672 ^ n3226 ;
  assign n3676 = n3675 ^ n3384 ;
  assign n3677 = ~n3674 & n3676 ;
  assign n3678 = n3677 ^ n3672 ;
  assign n3485 = n28 & ~n2820 ;
  assign n3483 = n2768 & ~n2815 ;
  assign n3478 = n2767 ^ n27 ;
  assign n3479 = n3478 ^ n2659 ;
  assign n3480 = n3479 ^ x1 ;
  assign n3481 = x0 & n3480 ;
  assign n3476 = n2777 ^ x1 ;
  assign n3482 = n3481 ^ n3476 ;
  assign n3484 = n3483 ^ n3482 ;
  assign n3486 = n3485 ^ n3484 ;
  assign n3475 = ~n2737 & ~n3502 ;
  assign n3487 = n3486 ^ n3475 ;
  assign n3679 = n3678 ^ n3487 ;
  assign n3680 = n3487 ^ n3212 ;
  assign n3681 = n3680 ^ n3387 ;
  assign n3682 = n3679 & ~n3681 ;
  assign n3683 = n3682 ^ n3678 ;
  assign n3684 = n3683 ^ n2760 ;
  assign n3687 = n3686 ^ n3684 ;
  assign n3698 = ~x2 & ~n2820 ;
  assign n3694 = n2820 ^ n2659 ;
  assign n3699 = n3698 ^ n3694 ;
  assign n3700 = ~x1 & n3699 ;
  assign n3689 = n27 & ~n3688 ;
  assign n3690 = n3689 ^ n2662 ;
  assign n3692 = n3690 ^ n2659 ;
  assign n3701 = n3700 ^ n3692 ;
  assign n3702 = ~x0 & ~n3701 ;
  assign n3691 = ~n4574 ^ n3690 ;
  assign n3703 = n3702 ^ n3691 ;
  assign n3704 = n3703 ^ n2760 ;
  assign n3705 = n3704 ^ n3686 ;
  assign n3706 = ~n3687 & n3705 ;
  assign n3707 = n3706 ^ n3686 ;
  assign n3708 = ~n3473 & ~n3707 ;
  assign n3709 = n3708 ^ n3472 ;
  assign n4025 = n3741 ^ n3709 ;
  assign n4026 = ~n3873 & n4025 ;
  assign n4027 = n4026 ^ n3741 ;
  assign n4182 = n4181 ^ n4027 ;
  assign n4192 = n4191 ^ n4182 ;
  assign n3887 = n145 & n333 ;
  assign n3883 = n709 ^ n109 ;
  assign n3882 = n416 ^ n122 ;
  assign n3884 = n3883 ^ n3882 ;
  assign n3885 = n3884 ^ n1059 ;
  assign n3880 = n2381 ^ n220 ;
  assign n3876 = n97 & n139 ;
  assign n3877 = n3876 ^ n625 ;
  assign n3878 = n3877 ^ n208 ;
  assign n3879 = n3878 ^ n494 ;
  assign n3881 = n3880 ^ n3879 ;
  assign n3886 = n3885 ^ n3881 ;
  assign n3888 = n3887 ^ n3886 ;
  assign n3889 = n3888 ^ n848 ;
  assign n3875 = n132 & ~n2374 ;
  assign n3890 = n3889 ^ n3875 ;
  assign n3902 = n633 ^ n79 ;
  assign n3899 = n2653 ^ n2600 ;
  assign n3896 = n910 ^ n175 ;
  assign n3897 = n3896 ^ n396 ;
  assign n3898 = n3897 ^ n2307 ;
  assign n3900 = n3899 ^ n3898 ;
  assign n3891 = n583 ^ n238 ;
  assign n3892 = n3891 ^ n432 ;
  assign n3893 = n3892 ^ n129 ;
  assign n3894 = n3893 ^ n2633 ;
  assign n3895 = n3894 ^ n683 ;
  assign n3901 = n3900 ^ n3895 ;
  assign n3903 = n3902 ^ n3901 ;
  assign n3904 = n3890 & n3903 ;
  assign n3874 = n3873 ^ n3709 ;
  assign n3905 = n3904 ^ n3874 ;
  assign n3906 = n3703 ^ n3685 ;
  assign n3924 = n514 ^ n365 ;
  assign n3920 = n497 ^ n343 ;
  assign n3921 = n3920 ^ n375 ;
  assign n3922 = n3921 ^ n2272 ;
  assign n3923 = n3922 ^ n2385 ;
  assign n3925 = n3924 ^ n3923 ;
  assign n3926 = n3925 ^ n262 ;
  assign n3907 = n558 ^ n321 ;
  assign n3908 = n3907 ^ n2599 ;
  assign n3909 = n3908 ^ n899 ;
  assign n3917 = n97 & n332 ;
  assign n3914 = n543 ^ n219 ;
  assign n3915 = n3914 ^ n2468 ;
  assign n3910 = n247 ^ n204 ;
  assign n3911 = n3910 ^ n404 ;
  assign n3912 = n3911 ^ n2431 ;
  assign n3913 = n3912 ^ n2551 ;
  assign n3916 = n3915 ^ n3913 ;
  assign n3918 = n3917 ^ n3916 ;
  assign n3919 = n3909 & ~n3918 ;
  assign n3927 = n3926 ^ n3919 ;
  assign n3957 = n671 ^ n451 ;
  assign n3958 = n3957 ^ n226 ;
  assign n3956 = n427 ^ n354 ;
  assign n3959 = n3958 ^ n3956 ;
  assign n3953 = n596 ^ n247 ;
  assign n3951 = n557 ^ n322 ;
  assign n3952 = n3951 ^ n161 ;
  assign n3954 = n3953 ^ n3952 ;
  assign n3950 = n2463 ^ n636 ;
  assign n3955 = n3954 ^ n3950 ;
  assign n3960 = n3959 ^ n3955 ;
  assign n3946 = ~n231 & ~n505 ;
  assign n3947 = n3946 ^ n865 ;
  assign n3943 = n392 ^ n103 ;
  assign n3944 = n3943 ^ n2634 ;
  assign n3945 = n3944 ^ n1043 ;
  assign n3948 = n3947 ^ n3945 ;
  assign n3949 = n3948 ^ n2480 ;
  assign n3961 = n3960 ^ n3949 ;
  assign n3935 = n850 ^ n386 ;
  assign n3938 = n3937 ^ n3935 ;
  assign n3939 = n3938 ^ n2538 ;
  assign n3940 = n3939 ^ n1278 ;
  assign n3930 = n289 ^ n211 ;
  assign n3931 = n3930 ^ n280 ;
  assign n3932 = n348 ^ n98 ;
  assign n3933 = n3932 ^ n3930 ;
  assign n3934 = ~n3931 & ~n3933 ;
  assign n3941 = n3940 ^ n3934 ;
  assign n3928 = n892 ^ n415 ;
  assign n3929 = n3928 ^ n110 ;
  assign n3942 = n3941 ^ n3929 ;
  assign n3962 = n3961 ^ n3942 ;
  assign n3963 = ~n3683 & n3927 ;
  assign n3964 = n3962 & ~n3963 ;
  assign n3984 = n3962 ^ n3473 ;
  assign n3985 = n3984 ^ n3963 ;
  assign n3993 = n3985 ^ n3473 ;
  assign n3989 = n3984 ^ n3906 ;
  assign n3991 = n3989 ^ n3473 ;
  assign n3994 = n3993 ^ n3991 ;
  assign n3995 = n3994 ^ n3473 ;
  assign n3965 = n3906 ^ n3473 ;
  assign n3966 = n3965 ^ n3962 ;
  assign n3967 = n3963 ^ n3962 ;
  assign n3969 = n3967 ^ n3963 ;
  assign n3970 = ~n3966 & n3969 ;
  assign n3972 = n3970 ^ n3963 ;
  assign n3973 = n3703 & ~n3972 ;
  assign n3980 = n3973 ^ n3970 ;
  assign n3974 = n3973 ^ n3967 ;
  assign n3979 = n3906 & ~n3974 ;
  assign n3981 = n3980 ^ n3979 ;
  assign n3982 = n3981 ^ n3966 ;
  assign n3983 = n3982 ^ n3963 ;
  assign n3996 = n3995 ^ n3983 ;
  assign n3997 = n3996 ^ n3985 ;
  assign n4000 = n3967 ^ n3683 ;
  assign n4001 = n4000 ^ n3964 ;
  assign n4002 = n4001 ^ n3683 ;
  assign n4003 = n3703 & ~n4002 ;
  assign n4004 = n4003 ^ n3683 ;
  assign n4005 = ~n3906 & ~n4004 ;
  assign n4006 = n4005 ^ n3683 ;
  assign n4007 = ~n3473 & ~n4006 ;
  assign n4008 = n4007 ^ n3473 ;
  assign n4009 = ~n3997 & n4008 ;
  assign n4010 = ~n3927 & n4009 ;
  assign n4011 = n3683 & n4010 ;
  assign n4014 = n4011 ^ n4009 ;
  assign n4015 = n4014 ^ n4008 ;
  assign n4012 = n3685 & n3703 ;
  assign n4013 = n4011 & n4012 ;
  assign n4016 = n4015 ^ n4013 ;
  assign n4017 = n3964 & ~n4016 ;
  assign n4018 = n3927 & n4017 ;
  assign n4019 = n3906 & n4018 ;
  assign n4020 = n4019 ^ n4017 ;
  assign n4021 = n4020 ^ n4016 ;
  assign n4022 = n4021 ^ n3904 ;
  assign n4023 = n3905 & n4022 ;
  assign n4024 = n4023 ^ n3905 ;
  assign n4193 = n4192 ^ n4024 ;
  assign n4355 = n476 ^ n228 ;
  assign n4208 = n204 ^ n182 ;
  assign n4209 = n4208 ^ n316 ;
  assign n4352 = n4209 ^ n2679 ;
  assign n4353 = n4352 ^ n3899 ;
  assign n4354 = n2332 & ~n4353 ;
  assign n4356 = n4355 ^ n4354 ;
  assign n4348 = n392 ^ n223 ;
  assign n4347 = n512 ^ n449 ;
  assign n4349 = n4348 ^ n4347 ;
  assign n4343 = ~n98 & n2642 ;
  assign n4342 = n3920 ^ n295 ;
  assign n4344 = n4343 ^ n4342 ;
  assign n4339 = n850 ^ n649 ;
  assign n4337 = n508 ^ n321 ;
  assign n4338 = n4337 ^ n350 ;
  assign n4340 = n4339 ^ n4338 ;
  assign n4341 = n4340 ^ n2653 ;
  assign n4345 = n4344 ^ n4341 ;
  assign n4346 = n4345 ^ n2349 ;
  assign n4350 = n4349 ^ n4346 ;
  assign n4351 = n4350 ^ n3888 ;
  assign n4357 = n4356 ^ n4351 ;
  assign n4331 = n4179 ^ n4151 ;
  assign n4332 = ~n4156 & ~n4331 ;
  assign n4333 = n4332 ^ n4151 ;
  assign n4324 = n4148 ^ n4143 ;
  assign n4325 = ~n4144 & n4324 ;
  assign n4326 = n4325 ^ n4148 ;
  assign n4319 = n1310 & ~n3184 ;
  assign n4320 = n2719 ^ n829 ;
  assign n4321 = n4319 & n4320 ;
  assign n4309 = n4142 ^ n2706 ;
  assign n4312 = ~n4132 & ~n4309 ;
  assign n4313 = n4312 ^ n2706 ;
  assign n4314 = ~n696 & n4313 ;
  assign n4315 = n4314 ^ n2705 ;
  assign n4316 = ~n696 & ~n4315 ;
  assign n4294 = n753 ^ n738 ;
  assign n4303 = n739 & n2704 ;
  assign n4304 = n4303 ^ n2703 ;
  assign n4305 = n4294 & n4304 ;
  assign n4295 = n739 & ~n3066 ;
  assign n4296 = n4295 ^ n2702 ;
  assign n4297 = n4296 ^ n2703 ;
  assign n4306 = n4305 ^ n4297 ;
  assign n4307 = ~n754 & ~n4306 ;
  assign n4308 = n4307 ^ n4296 ;
  assign n4317 = n4316 ^ n4308 ;
  assign n4286 = n753 & n1310 ;
  assign n4287 = ~n3183 & n4286 ;
  assign n4318 = n4317 ^ n4287 ;
  assign n4322 = n4321 ^ n4318 ;
  assign n4283 = ~n2701 & n2906 ;
  assign n4282 = ~n2700 & n2901 ;
  assign n4284 = n4283 ^ n4282 ;
  assign n4285 = n4284 ^ n753 ;
  assign n4288 = n4287 ^ n4284 ;
  assign n4289 = n1310 & n3185 ;
  assign n4290 = n4289 ^ n4284 ;
  assign n4291 = ~n4288 & ~n4290 ;
  assign n4292 = n4291 ^ n4284 ;
  assign n4293 = ~n4285 & n4292 ;
  assign n4323 = n4322 ^ n4293 ;
  assign n4327 = n4326 ^ n4323 ;
  assign n4266 = ~n2721 & n2871 ;
  assign n4265 = n2737 & ~n2865 ;
  assign n4267 = n4266 ^ n4265 ;
  assign n4268 = n4267 ^ n1017 ;
  assign n4270 = n1773 & ~n2816 ;
  assign n4271 = n4268 & n4270 ;
  assign n4262 = n1773 & ~n2813 ;
  assign n4263 = n2820 ^ n1021 ;
  assign n4264 = n4262 & n4263 ;
  assign n4269 = n4268 ^ n4264 ;
  assign n4272 = n4271 ^ n4269 ;
  assign n4273 = ~n1017 & ~n4272 ;
  assign n4274 = n4267 ^ n1773 ;
  assign n4275 = n4274 ^ n4267 ;
  assign n4276 = n4267 ^ n2828 ;
  assign n4277 = n4276 ^ n4267 ;
  assign n4278 = n4275 & n4277 ;
  assign n4279 = n4278 ^ n4267 ;
  assign n4280 = n4273 & n4279 ;
  assign n4281 = n4280 ^ n4272 ;
  assign n4328 = n4327 ^ n4281 ;
  assign n4259 = n4076 ^ n4073 ;
  assign n4260 = ~n4150 & ~n4259 ;
  assign n4261 = n4260 ^ n4076 ;
  assign n4329 = n4328 ^ n4261 ;
  assign n4256 = n2754 ^ n2659 ;
  assign n4257 = n2803 & ~n4256 ;
  assign n4251 = ~n1581 & n2754 ;
  assign n4249 = n3710 ^ n2662 ;
  assign n4250 = n4249 ^ n3715 ;
  assign n4252 = n4251 ^ n4250 ;
  assign n4253 = ~n2796 & ~n4252 ;
  assign n4248 = n2801 ^ n2662 ;
  assign n4254 = n4253 ^ n4248 ;
  assign n4241 = n2689 ^ n1483 ;
  assign n4245 = ~n2754 & ~n2796 ;
  assign n4246 = n4245 ^ n2797 ;
  assign n4247 = ~n4241 & n4246 ;
  assign n4255 = n4254 ^ n4247 ;
  assign n4258 = n4257 ^ n4255 ;
  assign n4330 = n4329 ^ n4258 ;
  assign n4334 = n4333 ^ n4330 ;
  assign n4235 = x2 & n3729 ;
  assign n4236 = n4235 ^ n4041 ;
  assign n4237 = ~x1 & ~n4236 ;
  assign n4221 = n903 ^ n189 ;
  assign n4222 = ~n62 & n4221 ;
  assign n4217 = n2269 ^ n309 ;
  assign n4218 = n4217 ^ n129 ;
  assign n4219 = n4218 ^ n449 ;
  assign n4220 = n4219 ^ n712 ;
  assign n4223 = n4222 ^ n4220 ;
  assign n4224 = n900 & ~n4223 ;
  assign n4215 = n545 ^ n355 ;
  assign n4211 = n211 ^ n78 ;
  assign n4212 = n4211 ^ n201 ;
  assign n4213 = n112 & n4212 ;
  assign n4210 = n4209 ^ n1428 ;
  assign n4214 = n4213 ^ n4210 ;
  assign n4216 = n4215 ^ n4214 ;
  assign n4225 = n4224 ^ n4216 ;
  assign n4226 = n2462 & ~n4225 ;
  assign n4205 = n4041 & ~n4043 ;
  assign n4204 = ~n4041 & ~n4042 ;
  assign n4206 = n4205 ^ n4204 ;
  assign n4207 = n27 & ~n4206 ;
  assign n4227 = n4226 ^ n4207 ;
  assign n4229 = n4227 ^ n4041 ;
  assign n4238 = n4237 ^ n4229 ;
  assign n4239 = ~x0 & n4238 ;
  assign n4228 = ~n4574 ^ n4227 ;
  assign n4240 = n4239 ^ n4228 ;
  assign n4335 = n4334 ^ n4240 ;
  assign n4201 = n4059 ^ n4027 ;
  assign n4202 = n4181 & n4201 ;
  assign n4203 = n4202 ^ n4059 ;
  assign n4336 = n4335 ^ n4203 ;
  assign n4358 = n4357 ^ n4336 ;
  assign n4199 = n4182 & n4191 ;
  assign n4200 = n4199 ^ n4192 ;
  assign n4359 = n4358 ^ n4200 ;
  assign n4197 = n3874 & n4024 ;
  assign n4198 = n4197 ^ n4024 ;
  assign n4360 = n4359 ^ n4198 ;
  assign n4194 = x23 ^ x22 ;
  assign n4195 = n4194 ^ n4024 ;
  assign n4196 = ~n4193 & ~n4195 ;
  assign n4361 = n4360 ^ n4196 ;
  assign n4522 = ~n4192 & n4358 ;
  assign n4362 = n4023 ^ n4021 ;
  assign n4519 = ~n4199 & ~n4362 ;
  assign n4528 = n4522 ^ n4519 ;
  assign n4529 = n4197 & ~n4528 ;
  assign n4363 = n4192 & ~n4198 ;
  assign n4364 = n4362 & n4363 ;
  assign n4527 = ~n4358 & n4364 ;
  assign n4530 = n4529 ^ n4527 ;
  assign n4523 = n4522 ^ n4200 ;
  assign n4524 = n4198 & ~n4523 ;
  assign n4518 = n4200 & ~n4358 ;
  assign n4520 = ~n4197 & n4519 ;
  assign n4521 = n4518 & n4520 ;
  assign n4525 = n4524 ^ n4521 ;
  assign n4531 = n4530 ^ n4525 ;
  assign n4532 = ~n4194 & ~n4531 ;
  assign n4514 = n574 ^ n194 ;
  assign n4515 = ~n62 & n4514 ;
  assign n4487 = n2662 & n2806 ;
  assign n4486 = ~n2689 & ~n2793 ;
  assign n4488 = n4487 ^ n4486 ;
  assign n4480 = n4241 ^ n2689 ;
  assign n4481 = n1581 & n2662 ;
  assign n4482 = n4481 ^ n2689 ;
  assign n4483 = ~n4480 & ~n4482 ;
  assign n4484 = n4483 ^ n2689 ;
  assign n4485 = ~n2781 & ~n4484 ;
  assign n4489 = n4488 ^ n4485 ;
  assign n4490 = n4489 ^ n1581 ;
  assign n4478 = n4044 ^ n3714 ;
  assign n4479 = n3229 & n4478 ;
  assign n4491 = n4490 ^ n4479 ;
  assign n4474 = n2790 ^ n2789 ;
  assign n4475 = n4044 ^ n3712 ;
  assign n4476 = n4475 ^ n3730 ;
  assign n4477 = ~n4474 & n4476 ;
  assign n4492 = n4491 ^ n4477 ;
  assign n4497 = ~n3715 & ~n4489 ;
  assign n4498 = n4497 ^ n2789 ;
  assign n4499 = n1581 & ~n4498 ;
  assign n4500 = n4499 ^ n2789 ;
  assign n4501 = n3730 ^ n3729 ;
  assign n4504 = n3729 ^ n1483 ;
  assign n4505 = n4504 ^ n3729 ;
  assign n4506 = ~n4501 & n4505 ;
  assign n4507 = n4506 ^ n3729 ;
  assign n4508 = ~n4500 & n4507 ;
  assign n4509 = ~n4492 & ~n4508 ;
  assign n4469 = n4226 ^ n1460 ;
  assign n4464 = n4206 & n4226 ;
  assign n4465 = n4464 ^ n4206 ;
  assign n4466 = n4465 ^ n4204 ;
  assign n4467 = n27 & ~n4466 ;
  assign n4468 = n4467 ^ n2672 ;
  assign n4470 = n4469 ^ n4468 ;
  assign n4461 = x2 & ~n4041 ;
  assign n4456 = n4226 ^ x22 ;
  assign n4462 = n4461 ^ n4456 ;
  assign n4463 = ~x1 & n4462 ;
  assign n4471 = n4470 ^ n4463 ;
  assign n4472 = ~x0 & ~n4471 ;
  assign n4473 = n4472 ^ n4468 ;
  assign n4510 = n4509 ^ n4473 ;
  assign n4449 = n4326 ^ n4317 ;
  assign n4450 = n4323 & ~n4449 ;
  assign n4451 = n4450 ^ n4317 ;
  assign n4443 = n4314 ^ n4308 ;
  assign n4444 = n4308 ^ n2705 ;
  assign n4445 = ~n4443 & n4444 ;
  assign n4446 = n4445 ^ n2992 ;
  assign n4447 = ~n696 & ~n4446 ;
  assign n4439 = n2703 & n3149 ;
  assign n4438 = ~n2702 & n3142 ;
  assign n4440 = n4439 ^ n4438 ;
  assign n4433 = n2701 ^ n739 ;
  assign n4434 = n4433 ^ n2701 ;
  assign n4435 = ~n3511 & n4434 ;
  assign n4436 = n4435 ^ n2701 ;
  assign n4437 = n754 & ~n4436 ;
  assign n4441 = n4440 ^ n4437 ;
  assign n4429 = n2721 ^ n829 ;
  assign n4430 = n1310 & ~n3186 ;
  assign n4431 = n4429 & n4430 ;
  assign n4417 = ~n2700 & n2906 ;
  assign n4416 = ~n2719 & n2901 ;
  assign n4418 = n4417 ^ n4416 ;
  assign n4419 = n4418 ^ n753 ;
  assign n4424 = n3206 ^ n3190 ;
  assign n4425 = ~n4419 & ~n4424 ;
  assign n4426 = n4425 ^ n3190 ;
  assign n4427 = n1310 & ~n4426 ;
  assign n4428 = n4427 ^ n4419 ;
  assign n4432 = n4431 ^ n4428 ;
  assign n4442 = n4441 ^ n4432 ;
  assign n4448 = n4447 ^ n4442 ;
  assign n4452 = n4451 ^ n4448 ;
  assign n4394 = n1021 & n2820 ;
  assign n4408 = ~n2737 & n2871 ;
  assign n4405 = n1017 & n2820 ;
  assign n4406 = n1021 & n2862 ;
  assign n4407 = ~n4405 & n4406 ;
  assign n4409 = n4408 ^ n4407 ;
  assign n4410 = n4409 ^ n2862 ;
  assign n4397 = n2659 ^ n1017 ;
  assign n4400 = n4397 ^ n2815 ;
  assign n4401 = n4400 ^ n4397 ;
  assign n4402 = ~n1022 & n4401 ;
  assign n4403 = n4402 ^ n4397 ;
  assign n4404 = n1773 & ~n4403 ;
  assign n4411 = n4410 ^ n4404 ;
  assign n4395 = n2820 ^ n1017 ;
  assign n4396 = ~n2865 & ~n4395 ;
  assign n4412 = n4411 ^ n4396 ;
  assign n4413 = n4412 ^ n4411 ;
  assign n4414 = n4394 & n4413 ;
  assign n4415 = n4414 ^ n4412 ;
  assign n4453 = n4452 ^ n4415 ;
  assign n4391 = n4281 ^ n4261 ;
  assign n4392 = n4328 & ~n4391 ;
  assign n4393 = n4392 ^ n4281 ;
  assign n4454 = n4453 ^ n4393 ;
  assign n4388 = n4333 ^ n4258 ;
  assign n4389 = n4330 & ~n4388 ;
  assign n4390 = n4389 ^ n4333 ;
  assign n4455 = n4454 ^ n4390 ;
  assign n4511 = n4510 ^ n4455 ;
  assign n4385 = n4240 ^ n4203 ;
  assign n4386 = ~n4335 & n4385 ;
  assign n4387 = n4386 ^ n4240 ;
  assign n4512 = n4511 ^ n4387 ;
  assign n4380 = n465 ^ n406 ;
  assign n4376 = n247 ^ n175 ;
  assign n4377 = n4376 ^ n864 ;
  assign n4378 = n4377 ^ n416 ;
  assign n4379 = n4378 ^ n1112 ;
  assign n4381 = n4380 ^ n4379 ;
  assign n4373 = n592 ^ n212 ;
  assign n4374 = n4373 ^ n295 ;
  assign n4371 = n557 ^ n166 ;
  assign n4372 = n4371 ^ n226 ;
  assign n4375 = n4374 ^ n4372 ;
  assign n4382 = n4381 ^ n4375 ;
  assign n4383 = n4382 ^ n916 ;
  assign n4384 = n4383 ^ n3926 ;
  assign n4513 = n4512 ^ n4384 ;
  assign n4516 = n4515 ^ n4513 ;
  assign n4366 = n4363 ^ n4192 ;
  assign n4365 = n4364 ^ n4199 ;
  assign n4367 = n4366 ^ n4365 ;
  assign n4368 = n4367 ^ n4336 ;
  assign n4369 = ~n4358 & n4368 ;
  assign n4370 = n4369 ^ n4357 ;
  assign n4517 = n4516 ^ n4370 ;
  assign n4526 = n4525 ^ n4517 ;
  assign n4533 = n4532 ^ n4526 ;
  assign n4700 = ~n4517 & n4530 ;
  assign n4701 = ~n4194 & ~n4700 ;
  assign n4534 = n4512 ^ n4370 ;
  assign n4535 = n4516 & n4534 ;
  assign n4536 = n4535 ^ n4512 ;
  assign n4689 = n4415 ^ n4393 ;
  assign n4690 = ~n4453 & n4689 ;
  assign n4691 = n4690 ^ n4415 ;
  assign n4673 = n2737 ^ n829 ;
  assign n4674 = n1310 & ~n2836 ;
  assign n4675 = n4673 & n4674 ;
  assign n4668 = ~n2719 & n2906 ;
  assign n4667 = ~n2721 & n2901 ;
  assign n4669 = n4668 ^ n4667 ;
  assign n4670 = n4669 ^ n753 ;
  assign n4676 = n4675 ^ n4670 ;
  assign n4666 = n2813 ^ n2722 ;
  assign n4671 = n1310 & n4670 ;
  assign n4672 = n4666 & n4671 ;
  assign n4677 = n4676 ^ n4672 ;
  assign n4678 = ~n753 & ~n4677 ;
  assign n4679 = n4669 ^ n1310 ;
  assign n4680 = n4679 ^ n4669 ;
  assign n4681 = n4669 ^ n2812 ;
  assign n4682 = n4681 ^ n4669 ;
  assign n4683 = n4680 & ~n4682 ;
  assign n4684 = n4683 ^ n4669 ;
  assign n4685 = n4678 & n4684 ;
  assign n4686 = n4685 ^ n4677 ;
  assign n4660 = n4441 ^ n2704 ;
  assign n4661 = n4446 & ~n4660 ;
  assign n4662 = n4661 ^ n2704 ;
  assign n4663 = n4662 ^ n2703 ;
  assign n4664 = ~n696 & ~n4663 ;
  assign n4656 = ~n2702 & n3149 ;
  assign n4655 = ~n2701 & n3142 ;
  assign n4657 = n4656 ^ n4655 ;
  assign n4650 = n2700 ^ n739 ;
  assign n4651 = n4650 ^ n2700 ;
  assign n4652 = ~n2855 & n4651 ;
  assign n4653 = n4652 ^ n2700 ;
  assign n4654 = n754 & ~n4653 ;
  assign n4658 = n4657 ^ n4654 ;
  assign n4645 = n4451 ^ n4432 ;
  assign n4646 = ~n4448 & ~n4645 ;
  assign n4647 = n4646 ^ n4451 ;
  assign n4659 = n4658 ^ n4647 ;
  assign n4665 = n4664 ^ n4659 ;
  assign n4687 = n4686 ^ n4665 ;
  assign n4616 = ~n1017 & ~n2863 ;
  assign n4631 = n4405 ^ n4397 ;
  assign n4632 = n4397 ^ n1581 ;
  assign n4633 = n4632 ^ n4397 ;
  assign n4634 = ~n4631 & ~n4633 ;
  assign n4635 = n4634 ^ n4397 ;
  assign n4636 = ~n1773 & n4635 ;
  assign n4625 = n2820 ^ n1581 ;
  assign n4626 = n4625 ^ n2820 ;
  assign n4627 = ~n3694 & ~n4626 ;
  assign n4628 = n4627 ^ n2820 ;
  assign n4629 = n2870 & n4628 ;
  assign n4638 = n4636 ^ n4629 ;
  assign n4639 = n1021 & n4638 ;
  assign n4617 = n2662 ^ n1017 ;
  assign n4620 = n4617 ^ n3688 ;
  assign n4621 = n4620 ^ n4617 ;
  assign n4622 = ~n1022 & ~n4621 ;
  assign n4623 = n4622 ^ n4617 ;
  assign n4624 = n1773 & ~n4623 ;
  assign n4630 = n4629 ^ n4624 ;
  assign n4640 = n4639 ^ n4630 ;
  assign n4641 = n4640 ^ n4624 ;
  assign n4642 = n2659 & ~n4641 ;
  assign n4643 = n4616 & n4642 ;
  assign n4644 = n4643 ^ n4640 ;
  assign n4688 = n4687 ^ n4644 ;
  assign n4692 = n4691 ^ n4688 ;
  assign n4576 = n2789 ^ n1581 ;
  assign n4586 = ~n2689 & n2806 ;
  assign n4585 = ~n2793 & n3729 ;
  assign n4587 = n4586 ^ n4585 ;
  assign n4579 = n2805 ^ n2781 ;
  assign n4582 = ~n4048 & ~n4505 ;
  assign n4583 = n4582 ^ n3729 ;
  assign n4584 = ~n4579 & n4583 ;
  assign n4588 = n4587 ^ n4584 ;
  assign n4589 = n1581 & n4588 ;
  assign n4577 = ~n4041 & ~n4474 ;
  assign n4578 = ~n4044 & n4577 ;
  assign n4590 = n4589 ^ n4578 ;
  assign n4591 = n4588 ^ n2789 ;
  assign n4592 = n4591 ^ n4588 ;
  assign n4593 = n4588 ^ n4044 ;
  assign n4594 = n4593 ^ n4588 ;
  assign n4595 = ~n4592 & ~n4594 ;
  assign n4596 = n4595 ^ n4588 ;
  assign n4597 = n1581 & ~n4596 ;
  assign n4598 = n4597 ^ n4588 ;
  assign n4603 = n1483 & ~n4044 ;
  assign n4604 = n4603 ^ n4041 ;
  assign n4605 = ~n4598 & n4604 ;
  assign n4606 = ~n4590 & ~n4605 ;
  assign n4607 = n4576 & n4606 ;
  assign n4608 = n4206 ^ n4043 ;
  assign n4609 = n4608 ^ n4588 ;
  assign n4610 = n4588 ^ n1581 ;
  assign n4611 = n4610 ^ n4588 ;
  assign n4612 = n4609 & n4611 ;
  assign n4613 = n4612 ^ n4588 ;
  assign n4614 = n4607 & ~n4613 ;
  assign n4615 = n4614 ^ n4606 ;
  assign n4693 = n4692 ^ n4615 ;
  assign n4570 = n2768 & ~n4205 ;
  assign n4571 = n4570 ^ n3502 ;
  assign n4572 = ~n4226 & ~n4571 ;
  assign n4575 = n4574 ^ n4572 ;
  assign n4694 = n4693 ^ n4575 ;
  assign n4563 = n3959 ^ n644 ;
  assign n4564 = ~n877 & n4563 ;
  assign n4558 = n389 ^ n146 ;
  assign n4557 = n4348 ^ n344 ;
  assign n4559 = n4558 ^ n4557 ;
  assign n4554 = n508 ^ n404 ;
  assign n4555 = n4554 ^ n402 ;
  assign n4556 = n4555 ^ n1123 ;
  assign n4560 = n4559 ^ n4556 ;
  assign n4561 = n4560 ^ n481 ;
  assign n4562 = n4561 ^ n1421 ;
  assign n4565 = n4564 ^ n4562 ;
  assign n4695 = n4694 ^ n4565 ;
  assign n4550 = n4509 ^ n4454 ;
  assign n4551 = n4454 ^ n4387 ;
  assign n4547 = n4473 ^ n4390 ;
  assign n4552 = n4551 ^ n4547 ;
  assign n4553 = ~n4550 & n4552 ;
  assign n4696 = n4695 ^ n4553 ;
  assign n4548 = n4473 ^ n4387 ;
  assign n4549 = ~n4547 & ~n4548 ;
  assign n4697 = n4696 ^ n4549 ;
  assign n4538 = n4194 & ~n4536 ;
  assign n4698 = n4697 ^ n4538 ;
  assign n4537 = n4536 ^ n4530 ;
  assign n4539 = n4538 ^ n4537 ;
  assign n4540 = n4539 ^ n4530 ;
  assign n4541 = n4530 ^ n4526 ;
  assign n4542 = n4540 & ~n4541 ;
  assign n4543 = n4542 ^ n4530 ;
  assign n4544 = n4538 ^ n4536 ;
  assign n4545 = n4544 ^ n4517 ;
  assign n4546 = n4543 & ~n4545 ;
  assign n4699 = n4698 ^ n4546 ;
  assign n4702 = n4699 ^ n4697 ;
  assign n4703 = n4536 & ~n4702 ;
  assign n4704 = n4701 & n4703 ;
  assign n4705 = n4704 ^ n4699 ;
  assign n4833 = ~n4390 & ~n4454 ;
  assign n4834 = n4551 ^ n4390 ;
  assign n4835 = ~n4473 & ~n4509 ;
  assign n4836 = n4835 ^ n4551 ;
  assign n4837 = n4836 ^ n4510 ;
  assign n4838 = n4837 ^ n4551 ;
  assign n4839 = ~n4834 & n4838 ;
  assign n4840 = n4839 ^ n4551 ;
  assign n4841 = n4455 & n4840 ;
  assign n4842 = n4841 ^ n4454 ;
  assign n4843 = n4694 ^ n4387 ;
  assign n4844 = n4843 ^ n4694 ;
  assign n4845 = n4835 ^ n4694 ;
  assign n4846 = n4845 ^ n4694 ;
  assign n4847 = ~n4844 & n4846 ;
  assign n4848 = n4847 ^ n4694 ;
  assign n4849 = ~n4842 & ~n4848 ;
  assign n4854 = n4510 & ~n4548 ;
  assign n4855 = n4854 ^ n4509 ;
  assign n4856 = ~n4849 & ~n4855 ;
  assign n4857 = ~n4694 & n4856 ;
  assign n4860 = n4857 ^ n4856 ;
  assign n4861 = n4833 & n4860 ;
  assign n4858 = n4857 ^ n4849 ;
  assign n4862 = n4861 ^ n4858 ;
  assign n4753 = n4691 ^ n4644 ;
  assign n4754 = ~n4688 & ~n4753 ;
  assign n4755 = n4754 ^ n4691 ;
  assign n4820 = n1021 & ~n2862 ;
  assign n4821 = ~n2754 & n4820 ;
  assign n4819 = n2871 & n4256 ;
  assign n4822 = n4821 ^ n4819 ;
  assign n4823 = n4822 ^ n4617 ;
  assign n4816 = ~n1017 & ~n2754 ;
  assign n4817 = n4816 ^ n2662 ;
  assign n4818 = n2865 & n4817 ;
  assign n4824 = n4823 ^ n4818 ;
  assign n4812 = n1773 & ~n2689 ;
  assign n4825 = n4824 ^ n4812 ;
  assign n4795 = n4658 ^ n2703 ;
  assign n4796 = n4658 ^ n696 ;
  assign n4797 = n4796 ^ n4658 ;
  assign n4800 = n4662 & ~n4797 ;
  assign n4801 = n4800 ^ n4658 ;
  assign n4802 = ~n4795 & n4801 ;
  assign n4803 = n4802 ^ n2703 ;
  assign n4804 = n4803 ^ n2702 ;
  assign n4805 = ~n696 & ~n4804 ;
  assign n4781 = ~n2721 & n2906 ;
  assign n4780 = n2737 & n2901 ;
  assign n4782 = n4781 ^ n4780 ;
  assign n4791 = n4782 ^ n753 ;
  assign n4788 = n2820 ^ n829 ;
  assign n4789 = n1310 & ~n2813 ;
  assign n4790 = n4788 & n4789 ;
  assign n4792 = n4791 ^ n4790 ;
  assign n4783 = ~n2816 & ~n4782 ;
  assign n4784 = n4783 ^ n2828 ;
  assign n4785 = ~n753 & n4784 ;
  assign n4786 = n4785 ^ n2828 ;
  assign n4787 = n1310 & n4786 ;
  assign n4793 = n4792 ^ n4787 ;
  assign n4762 = ~n2700 & n3142 ;
  assign n4760 = ~n2701 & n3149 ;
  assign n4758 = n754 & ~n3184 ;
  assign n4756 = n754 & n3185 ;
  assign n4757 = n4756 ^ n696 ;
  assign n4759 = n4758 ^ n4757 ;
  assign n4761 = n4760 ^ n4759 ;
  assign n4763 = n4762 ^ n4761 ;
  assign n4764 = n2719 ^ n738 ;
  assign n4765 = n4764 ^ n4756 ;
  assign n4766 = n4758 & n4765 ;
  assign n4770 = n4766 ^ n4756 ;
  assign n4772 = ~n696 & n4770 ;
  assign n4773 = n4772 ^ n4756 ;
  assign n4774 = n4763 & ~n4773 ;
  assign n4767 = n4766 ^ n4764 ;
  assign n4775 = n4774 ^ n4767 ;
  assign n4776 = n4775 ^ n4764 ;
  assign n4777 = n4776 ^ ~n4574 ;
  assign n4794 = n4793 ^ n4777 ;
  assign n4806 = n4805 ^ n4794 ;
  assign n4808 = n4806 ^ n4686 ;
  assign n4807 = n4806 ^ n4647 ;
  assign n4809 = n4808 ^ n4807 ;
  assign n4810 = n4665 & ~n4809 ;
  assign n4811 = n4810 ^ n4808 ;
  assign n4826 = n4825 ^ n4811 ;
  assign n4828 = ~n4755 & n4826 ;
  assign n4723 = n4615 ^ n4575 ;
  assign n4724 = n4693 & ~n4723 ;
  assign n4725 = n4724 ^ n4615 ;
  assign n4748 = ~n3189 & ~n4206 ;
  assign n4746 = ~n2789 & n4226 ;
  assign n4727 = n4041 ^ n2789 ;
  assign n4741 = n4727 ^ n1581 ;
  assign n4740 = n2806 & n3729 ;
  assign n4742 = n4741 ^ n4740 ;
  assign n4739 = n2795 & ~n4041 ;
  assign n4743 = n4742 ^ n4739 ;
  assign n4736 = n1581 & n3729 ;
  assign n4737 = n4736 ^ n4041 ;
  assign n4738 = n2792 & ~n4737 ;
  assign n4744 = n4743 ^ n4738 ;
  assign n4726 = n4206 ^ n4041 ;
  assign n4729 = ~n2789 & n4726 ;
  assign n4730 = n4729 ^ n4041 ;
  assign n4731 = ~n1483 & ~n4730 ;
  assign n4745 = n4744 ^ n4731 ;
  assign n4747 = n4746 ^ n4745 ;
  assign n4749 = n4748 ^ n4747 ;
  assign n4751 = n4725 & n4749 ;
  assign n4831 = n4828 ^ n4751 ;
  assign n4827 = n4826 ^ n4755 ;
  assign n4829 = n4828 ^ n4827 ;
  assign n4750 = n4749 ^ n4725 ;
  assign n4752 = n4751 ^ n4750 ;
  assign n4830 = n4829 ^ n4752 ;
  assign n4832 = n4831 ^ n4830 ;
  assign n4863 = n4862 ^ n4832 ;
  assign n4718 = n170 ^ n155 ;
  assign n4719 = n4718 ^ n535 ;
  assign n4716 = n2605 ^ n324 ;
  assign n4715 = n1117 ^ n896 ;
  assign n4717 = n4716 ^ n4715 ;
  assign n4720 = n4719 ^ n4717 ;
  assign n4721 = n1045 & n4720 ;
  assign n4714 = n2490 ^ n846 ;
  assign n4722 = n4721 ^ n4714 ;
  assign n4871 = n4863 ^ n4722 ;
  assign n4864 = n4722 & n4863 ;
  assign n4872 = n4871 ^ n4864 ;
  assign n4865 = n4565 ^ n4536 ;
  assign n4866 = ~n4697 & ~n4865 ;
  assign n4867 = n4866 ^ n4536 ;
  assign n4869 = n4867 ^ n4864 ;
  assign n4868 = n4864 & n4867 ;
  assign n4870 = n4869 ^ n4868 ;
  assign n4873 = n4872 ^ n4870 ;
  assign n4874 = n4873 ^ n4868 ;
  assign n4706 = n4697 ^ n4536 ;
  assign n4711 = n4700 & ~n4706 ;
  assign n4712 = ~n4194 & ~n4711 ;
  assign n4707 = n4517 & n4525 ;
  assign n4708 = n4706 & n4707 ;
  assign n4709 = n4194 & ~n4708 ;
  assign n4710 = n4709 ^ n4194 ;
  assign n4713 = n4712 ^ n4710 ;
  assign n4875 = n4874 ^ n4713 ;
  assign n5009 = n4870 & n4872 ;
  assign n5011 = n5009 ^ n4709 ;
  assign n5004 = n599 ^ n110 ;
  assign n5005 = ~n531 & n5004 ;
  assign n4999 = n1100 ^ n206 ;
  assign n4998 = n3891 ^ n2367 ;
  assign n5000 = n4999 ^ n4998 ;
  assign n4995 = n635 ^ n304 ;
  assign n4996 = n4995 ^ n402 ;
  assign n4997 = n4996 ^ n2389 ;
  assign n5001 = n5000 ^ n4997 ;
  assign n5002 = n5001 ^ n4223 ;
  assign n5003 = n5002 ^ n4356 ;
  assign n5006 = n5005 ^ n5003 ;
  assign n5007 = n2644 & ~n5006 ;
  assign n4966 = n2796 & ~n4226 ;
  assign n4967 = n4966 ^ n1581 ;
  assign n4968 = n4967 ^ n1483 ;
  assign n4973 = ~n4574 ^ n4466 ;
  assign n4974 = n4973 ^ n4466 ;
  assign n4975 = n4967 & ~n4974 ;
  assign n4976 = ~n4041 & n4975 ;
  assign n4977 = n4976 ^ n4041 ;
  assign n4969 = n4466 ^ n4041 ;
  assign n4978 = n4977 ^ n4969 ;
  assign n4979 = n2789 & n4978 ;
  assign n4980 = n4979 ^ n4466 ;
  assign n4981 = n4968 & ~n4980 ;
  assign n4982 = n4981 ^ n1483 ;
  assign n4983 = ~n1581 & ~n4982 ;
  assign n4984 = n4966 ^ n2803 ;
  assign n4985 = n4984 ^ n4966 ;
  assign n4988 = ~n4041 & n4985 ;
  assign n4989 = n4988 ^ n4966 ;
  assign n4990 = n4983 & n4989 ;
  assign n4991 = n4990 ^ n4982 ;
  assign n4957 = n1773 & n3729 ;
  assign n4949 = n3715 ^ n2689 ;
  assign n4950 = n4949 ^ n2689 ;
  assign n4953 = n1017 & ~n4950 ;
  assign n4954 = n4953 ^ n2689 ;
  assign n4955 = n2865 & ~n4954 ;
  assign n4951 = n2689 ^ n1017 ;
  assign n4956 = n4955 ^ n4951 ;
  assign n4958 = n4957 ^ n4956 ;
  assign n4947 = ~n3715 & n4062 ;
  assign n4945 = n3715 ^ n2662 ;
  assign n4946 = n2871 & ~n4945 ;
  assign n4948 = n4947 ^ n4946 ;
  assign n4959 = n4958 ^ n4948 ;
  assign n4939 = n4777 & n4793 ;
  assign n4936 = n4803 ^ n4793 ;
  assign n4932 = n4793 ^ n696 ;
  assign n4933 = n4932 ^ n4777 ;
  assign n4937 = n4933 ^ n2702 ;
  assign n4938 = n4936 & n4937 ;
  assign n4940 = n4939 ^ n4938 ;
  assign n4941 = ~n696 & n4940 ;
  assign n4942 = n4941 ^ n4939 ;
  assign n4943 = n4942 ^ n4793 ;
  assign n4926 = ~n696 & ~n2701 ;
  assign n4921 = n4574 & ~n4776 ;
  assign n4923 = n4921 ^ n4777 ;
  assign n4927 = n4926 ^ n4923 ;
  assign n4920 = ~n696 & ~n2702 ;
  assign n4922 = ~n2702 & n4921 ;
  assign n4924 = n4923 ^ n4922 ;
  assign n4925 = n4920 & ~n4924 ;
  assign n4928 = n4927 ^ n4925 ;
  assign n4909 = n2721 ^ n738 ;
  assign n4910 = n754 & ~n3186 ;
  assign n4911 = n4909 & n4910 ;
  assign n4898 = ~n738 & n2719 ;
  assign n4900 = ~n2612 & ~n4898 ;
  assign n4903 = ~n2700 & ~n3145 ;
  assign n4904 = n4900 & n4903 ;
  assign n4899 = n4898 ^ n696 ;
  assign n4901 = n4900 ^ n4899 ;
  assign n4891 = ~n696 & ~n2700 ;
  assign n4892 = n4891 ^ n2700 ;
  assign n4893 = n4892 ^ n2719 ;
  assign n4895 = ~n738 & n4893 ;
  assign n4896 = n4895 ^ n2719 ;
  assign n4897 = n799 & ~n4896 ;
  assign n4902 = n4901 ^ n4897 ;
  assign n4905 = n4904 ^ n4902 ;
  assign n4912 = n4911 ^ n4905 ;
  assign n4906 = n800 ^ n696 ;
  assign n4907 = n4906 ^ n3148 ;
  assign n4908 = ~n3190 & n4907 ;
  assign n4913 = n4912 ^ n4908 ;
  assign n4929 = n4928 ^ n4913 ;
  assign n4914 = n4913 ^ n696 ;
  assign n4915 = n754 & n3206 ;
  assign n4916 = n4915 ^ n696 ;
  assign n4917 = n4914 & ~n4916 ;
  assign n4918 = n4917 ^ n696 ;
  assign n4919 = n4905 & ~n4918 ;
  assign n4930 = n4929 ^ n4919 ;
  assign n4886 = n1537 & n2815 ;
  assign n4880 = ~n2820 & n2901 ;
  assign n4879 = n2737 & n2906 ;
  assign n4881 = n4880 ^ n4879 ;
  assign n4883 = n4881 ^ n2659 ;
  assign n4884 = ~n753 & ~n4883 ;
  assign n4885 = n4881 & n4884 ;
  assign n4887 = n4886 ^ n4885 ;
  assign n4888 = n4887 ^ n4883 ;
  assign n4889 = n1310 & ~n4888 ;
  assign n4882 = n4881 ^ n753 ;
  assign n4890 = n4889 ^ n4882 ;
  assign n4931 = n4930 ^ n4890 ;
  assign n4944 = n4943 ^ n4931 ;
  assign n4960 = n4959 ^ n4944 ;
  assign n4962 = n4960 ^ n4806 ;
  assign n4961 = n4960 ^ n4825 ;
  assign n4963 = n4962 ^ n4961 ;
  assign n4964 = ~n4811 & ~n4963 ;
  assign n4965 = n4964 ^ n4962 ;
  assign n4992 = n4991 ^ n4965 ;
  assign n4993 = n4992 ^ n4831 ;
  assign n4876 = n4862 ^ n4827 ;
  assign n4877 = n4827 ^ n4750 ;
  assign n4878 = ~n4876 & ~n4877 ;
  assign n4994 = n4993 ^ n4878 ;
  assign n5008 = n5007 ^ n4994 ;
  assign n5012 = n5011 ^ n5008 ;
  assign n5010 = n5009 ^ n5008 ;
  assign n5013 = n5012 ^ n5010 ;
  assign n5014 = n4871 ^ n4867 ;
  assign n5015 = ~n4712 & ~n5014 ;
  assign n5016 = ~n5013 & n5015 ;
  assign n5017 = n5016 ^ n5012 ;
  assign n5018 = n4867 ^ n4863 ;
  assign n5019 = n5018 ^ n4722 ;
  assign n5020 = n4711 & ~n5019 ;
  assign n5021 = n5008 ^ n4867 ;
  assign n5022 = n5021 ^ n5008 ;
  assign n5023 = n5008 ^ n4722 ;
  assign n5024 = n5023 ^ n5008 ;
  assign n5025 = ~n5022 & ~n5024 ;
  assign n5026 = n5025 ^ n5008 ;
  assign n5027 = n5020 & ~n5026 ;
  assign n5176 = n4194 & ~n5027 ;
  assign n5181 = n4874 & ~n5008 ;
  assign n5182 = n5181 ^ n4868 ;
  assign n5183 = n4708 & n5182 ;
  assign n5184 = n5176 & ~n5183 ;
  assign n5166 = n358 ^ n247 ;
  assign n5167 = n5166 ^ n675 ;
  assign n5168 = n5167 ^ n482 ;
  assign n5164 = n2679 ^ n140 ;
  assign n5165 = n5164 ^ n310 ;
  assign n5169 = n5168 ^ n5165 ;
  assign n5159 = n2367 ^ n477 ;
  assign n5160 = n5159 ^ n627 ;
  assign n5161 = n5160 ^ n2457 ;
  assign n5158 = n4348 ^ n4209 ;
  assign n5162 = n5161 ^ n5158 ;
  assign n5150 = n98 ^ n63 ;
  assign n5155 = ~n42 & n611 ;
  assign n5156 = n5155 ^ n194 ;
  assign n5157 = ~n5150 & n5156 ;
  assign n5163 = n5162 ^ n5157 ;
  assign n5170 = n5169 ^ n5163 ;
  assign n5171 = n5170 ^ n2485 ;
  assign n5172 = n3890 & n5171 ;
  assign n5130 = n4992 ^ n4751 ;
  assign n5131 = n4992 ^ n4752 ;
  assign n5132 = n5131 ^ n4826 ;
  assign n5133 = n5132 ^ n4755 ;
  assign n5134 = n5133 ^ n5131 ;
  assign n5135 = n4755 & n4992 ;
  assign n5136 = n5135 ^ n5131 ;
  assign n5137 = n5134 & ~n5136 ;
  assign n5138 = n5137 ^ n5131 ;
  assign n5139 = ~n4862 & ~n5138 ;
  assign n5140 = n5139 ^ n4828 ;
  assign n5141 = ~n5130 & ~n5140 ;
  assign n5142 = n4862 ^ n4749 ;
  assign n5143 = n4750 & n5142 ;
  assign n5144 = n5143 ^ n4749 ;
  assign n5145 = ~n5141 & n5144 ;
  assign n5147 = n5145 ^ n5141 ;
  assign n5129 = ~n4829 & n4992 ;
  assign n5146 = n5129 & n5145 ;
  assign n5148 = n5147 ^ n5146 ;
  assign n5123 = n1773 & ~n4041 ;
  assign n5117 = n3729 ^ n1017 ;
  assign n5118 = n5117 ^ n3729 ;
  assign n5119 = ~n4044 & n5118 ;
  assign n5120 = n5119 ^ n3729 ;
  assign n5121 = n2865 & n5120 ;
  assign n5122 = n5121 ^ n5117 ;
  assign n5124 = n5123 ^ n5122 ;
  assign n5113 = ~n4044 & n4062 ;
  assign n5111 = n4044 ^ n2689 ;
  assign n5112 = n2871 & n5111 ;
  assign n5114 = n5113 ^ n5112 ;
  assign n5125 = n5124 ^ n5114 ;
  assign n5085 = n1310 & ~n3688 ;
  assign n5092 = n2662 ^ n829 ;
  assign n5088 = ~n2820 & n2906 ;
  assign n5087 = ~n2659 & n2901 ;
  assign n5089 = n5088 ^ n5087 ;
  assign n5090 = n5089 ^ n753 ;
  assign n5086 = n1310 & n2662 ;
  assign n5091 = n5090 ^ n5086 ;
  assign n5093 = n5092 ^ n5091 ;
  assign n5094 = n5085 & n5093 ;
  assign n5095 = n5094 ^ n5091 ;
  assign n5078 = n2721 ^ n696 ;
  assign n5079 = n3144 ^ n3141 ;
  assign n5075 = ~n696 & ~n2721 ;
  assign n5076 = n2612 & n5075 ;
  assign n5072 = n3147 & n4898 ;
  assign n5070 = ~n696 & n2719 ;
  assign n5071 = ~n2615 & ~n5070 ;
  assign n5073 = n5072 ^ n5071 ;
  assign n5061 = n4924 ^ n4920 ;
  assign n5062 = n5061 ^ n4924 ;
  assign n5066 = ~n4923 & n5062 ;
  assign n5067 = n5066 ^ n4924 ;
  assign n5068 = ~n4926 & ~n5067 ;
  assign n5063 = n4922 ^ n4891 ;
  assign n5069 = n5068 ^ n5063 ;
  assign n5074 = n5073 ^ n5069 ;
  assign n5077 = n5076 ^ n5074 ;
  assign n5080 = n5077 ^ n5069 ;
  assign n5081 = n5079 & ~n5080 ;
  assign n5082 = ~n5078 & n5081 ;
  assign n5083 = n5082 ^ n5077 ;
  assign n5053 = n2737 ^ n738 ;
  assign n5056 = n5053 ^ n2836 ;
  assign n5057 = n5056 ^ n5053 ;
  assign n5058 = n739 & n5057 ;
  assign n5059 = n5058 ^ n5053 ;
  assign n5060 = n754 & n5059 ;
  assign n5084 = n5083 ^ n5060 ;
  assign n5105 = n5095 ^ n5084 ;
  assign n5106 = n5105 ^ n4928 ;
  assign n5107 = n5106 ^ n4890 ;
  assign n5108 = n5107 ^ n5105 ;
  assign n5109 = ~n4930 & ~n5108 ;
  assign n5110 = n5109 ^ n5106 ;
  assign n5126 = n5125 ^ n5110 ;
  assign n5050 = n4959 ^ n4943 ;
  assign n5051 = n4944 & ~n5050 ;
  assign n5052 = n5051 ^ n4959 ;
  assign n5127 = n5126 ^ n5052 ;
  assign n5046 = n4991 ^ n4960 ;
  assign n5047 = ~n4965 & n5046 ;
  assign n5048 = n5047 ^ n4960 ;
  assign n5033 = ~n1483 & ~n4226 ;
  assign n5034 = n5033 ^ n1581 ;
  assign n5035 = ~n4205 & ~n5034 ;
  assign n5036 = n5035 ^ n1581 ;
  assign n5037 = n3550 & ~n5036 ;
  assign n5038 = n2781 ^ n1581 ;
  assign n5041 = n1835 & ~n4226 ;
  assign n5042 = n5038 & n5041 ;
  assign n5043 = n5042 ^ n5038 ;
  assign n5044 = n5043 ^ n2781 ;
  assign n5045 = ~n5037 & n5044 ;
  assign n5049 = n5048 ^ n5045 ;
  assign n5128 = n5127 ^ n5049 ;
  assign n5149 = n5148 ^ n5128 ;
  assign n5173 = n5172 ^ n5149 ;
  assign n5028 = n5009 ^ n4994 ;
  assign n5029 = n5008 & ~n5028 ;
  assign n5030 = n5029 ^ n5009 ;
  assign n5174 = n5173 ^ n5030 ;
  assign n5175 = n5174 ^ n5027 ;
  assign n5185 = n5184 ^ n5175 ;
  assign n5186 = n5027 & ~n5174 ;
  assign n5187 = ~n4194 & ~n5186 ;
  assign n5287 = n5174 & n5183 ;
  assign n5290 = n5187 & ~n5287 ;
  assign n5282 = n5148 ^ n5127 ;
  assign n5283 = ~n5128 & ~n5282 ;
  assign n5274 = n4206 ^ n3729 ;
  assign n5275 = n2871 & ~n5274 ;
  assign n5273 = ~n4206 & n4820 ;
  assign n5276 = n5275 ^ n5273 ;
  assign n5268 = n4041 ^ n1017 ;
  assign n5277 = n5276 ^ n5268 ;
  assign n5270 = ~n1017 & ~n4206 ;
  assign n5271 = n5270 ^ n4041 ;
  assign n5272 = n2865 & ~n5271 ;
  assign n5278 = n5277 ^ n5272 ;
  assign n5266 = n1773 & ~n4226 ;
  assign n5279 = n5278 ^ n5266 ;
  assign n5240 = ~n2721 & n3149 ;
  assign n5239 = n754 & ~n2820 ;
  assign n5241 = n5240 ^ n5239 ;
  assign n5237 = n2737 & n3142 ;
  assign n5955 = n739 & n754 ;
  assign n5236 = ~n2813 & n5955 ;
  assign n5238 = n5237 ^ n5236 ;
  assign n5242 = n5241 ^ n5238 ;
  assign n5255 = n5242 ^ n1581 ;
  assign n5219 = ~n2700 & n4574 ;
  assign n5220 = ~n2701 & ~n2702 ;
  assign n5221 = ~n4776 & n5220 ;
  assign n5222 = n5219 & n5221 ;
  assign n5228 = n5070 ^ ~n4574 ;
  assign n5224 = ~n4777 & ~n4920 ;
  assign n5225 = ~n4891 & ~n4926 ;
  assign n5226 = n5224 & n5225 ;
  assign n5227 = ~n4574 & ~n5226 ;
  assign n5229 = n5228 ^ n5227 ;
  assign n5230 = ~n5222 & n5229 ;
  assign n5256 = n5255 ^ n5230 ;
  assign n5252 = n5095 ^ n5069 ;
  assign n5253 = n5084 & n5252 ;
  assign n5254 = n5253 ^ n5095 ;
  assign n5257 = n5256 ^ n5254 ;
  assign n5243 = n5230 ^ n4923 ;
  assign n5244 = n5243 ^ n5230 ;
  assign n5247 = n696 & n5244 ;
  assign n5248 = n5247 ^ n5230 ;
  assign n5249 = ~n5242 & ~n5248 ;
  assign n5258 = n5257 ^ n5249 ;
  assign n5223 = n5222 ^ n2719 ;
  assign n5250 = ~n5230 & n5249 ;
  assign n5251 = ~n5223 & n5250 ;
  assign n5259 = n5258 ^ n5251 ;
  assign n5213 = ~n753 & ~n2754 ;
  assign n5214 = n5213 ^ n2689 ;
  assign n5215 = n1310 & ~n5214 ;
  assign n5216 = n5215 ^ n753 ;
  assign n5208 = ~n2659 & n2906 ;
  assign n5217 = n5216 ^ n5208 ;
  assign n5206 = n2662 & n2901 ;
  assign n5205 = ~n2754 & n2897 ;
  assign n5207 = n5206 ^ n5205 ;
  assign n5218 = n5217 ^ n5207 ;
  assign n5260 = n5259 ^ n5218 ;
  assign n5262 = n5260 ^ n5105 ;
  assign n5261 = n5260 ^ n5125 ;
  assign n5263 = n5262 ^ n5261 ;
  assign n5264 = ~n5110 & ~n5263 ;
  assign n5265 = n5264 ^ n5261 ;
  assign n5280 = n5279 ^ n5265 ;
  assign n5202 = n5045 & n5048 ;
  assign n5203 = n5202 ^ n5049 ;
  assign n5200 = n5052 & ~n5126 ;
  assign n5201 = n5200 ^ n5049 ;
  assign n5204 = n5203 ^ n5201 ;
  assign n5281 = n5280 ^ n5204 ;
  assign n5284 = n5283 ^ n5281 ;
  assign n5197 = n188 & ~n3948 ;
  assign n5195 = ~n307 & n699 ;
  assign n5192 = n4996 ^ n176 ;
  assign n5191 = n856 ^ n385 ;
  assign n5193 = n5192 ^ n5191 ;
  assign n5194 = n5193 ^ n5163 ;
  assign n5196 = n5195 ^ n5194 ;
  assign n5198 = n5197 ^ n5196 ;
  assign n5199 = n2354 & n5198 ;
  assign n5285 = n5284 ^ n5199 ;
  assign n5188 = n5149 ^ n5030 ;
  assign n5189 = n5173 & n5188 ;
  assign n5190 = n5189 ^ n5149 ;
  assign n5286 = n5285 ^ n5190 ;
  assign n5288 = n5287 ^ n5286 ;
  assign n5291 = n5290 ^ n5288 ;
  assign n5426 = n527 ^ n358 ;
  assign n5425 = n2636 ^ n2465 ;
  assign n5427 = n5426 ^ n5425 ;
  assign n5423 = n709 ^ n388 ;
  assign n5422 = n1029 ^ n864 ;
  assign n5424 = n5423 ^ n5422 ;
  assign n5428 = n5427 ^ n5424 ;
  assign n5419 = n333 ^ n139 ;
  assign n5420 = ~n61 & n5419 ;
  assign n5415 = n432 ^ n109 ;
  assign n5416 = n5415 ^ n591 ;
  assign n5417 = n5416 ^ n457 ;
  assign n5418 = n5417 ^ n3902 ;
  assign n5421 = n5420 ^ n5418 ;
  assign n5429 = n5428 ^ n5421 ;
  assign n5430 = n3942 & n5429 ;
  assign n5409 = n5254 ^ n5218 ;
  assign n5410 = ~n5259 & n5409 ;
  assign n5411 = n5410 ^ n5218 ;
  assign n5401 = n1773 & n4466 ;
  assign n5403 = n2871 & ~n4041 ;
  assign n5402 = ~n2865 & ~n4226 ;
  assign n5404 = n5403 ^ n5402 ;
  assign n5405 = n5404 ^ n1017 ;
  assign n5406 = n5405 ^ n1021 ;
  assign n5407 = n5401 & ~n5406 ;
  assign n5408 = n5407 ^ n5405 ;
  assign n5412 = n5411 ^ n5408 ;
  assign n5387 = n2659 ^ n738 ;
  assign n5388 = n754 & n2815 ;
  assign n5389 = ~n5387 & n5388 ;
  assign n5374 = ~n2820 & n3142 ;
  assign n5373 = n2737 & n3149 ;
  assign n5375 = n5374 ^ n5373 ;
  assign n5376 = n5375 ^ n2659 ;
  assign n5377 = n5376 ^ n5375 ;
  assign n5380 = n5375 ^ n2815 ;
  assign n5381 = n5380 ^ n5375 ;
  assign n5382 = n754 & ~n5381 ;
  assign n5383 = ~n5377 & n5382 ;
  assign n5384 = n5383 ^ n5377 ;
  assign n5385 = n5384 ^ n5376 ;
  assign n5386 = ~n696 & n5385 ;
  assign n5390 = n5389 ^ n5386 ;
  assign n5391 = n5375 ^ n696 ;
  assign n5392 = ~n5390 & n5391 ;
  assign n5395 = n5392 ^ n5390 ;
  assign n5393 = n754 & n3753 ;
  assign n5394 = n5392 & n5393 ;
  assign n5396 = n5395 ^ n5394 ;
  assign n5367 = ~n4574 ^ n1581 ;
  assign n5368 = ~n4574 ^ n696 ;
  assign n5369 = n5368 ^ n5070 ;
  assign n5370 = n5367 & ~n5369 ;
  assign n5371 = n5370 ^ n1581 ;
  assign n5372 = n5371 ^ n5075 ;
  assign n5397 = n5396 ^ n5372 ;
  assign n5357 = n4891 & n5221 ;
  assign n5358 = ~n5227 & n5357 ;
  assign n5359 = n5358 ^ n5227 ;
  assign n5360 = n5359 ^ n5070 ;
  assign n5361 = n5228 & n5360 ;
  assign n5355 = n1581 ^ n696 ;
  assign n5356 = n5355 ^ ~n4574 ;
  assign n5362 = n5361 ^ n5356 ;
  assign n5363 = n5359 ^ n5242 ;
  assign n5364 = n5363 ^ n696 ;
  assign n5365 = ~n5362 & ~n5364 ;
  assign n5366 = n5365 ^ n5359 ;
  assign n5398 = n5397 ^ n5366 ;
  assign n5338 = n2905 & n4476 ;
  assign n5329 = n2662 & n2906 ;
  assign n5328 = ~n2689 & n2901 ;
  assign n5330 = n5329 ^ n5328 ;
  assign n5331 = n5330 ^ n753 ;
  assign n5334 = ~n829 & ~n4501 ;
  assign n5335 = n5334 ^ n3729 ;
  assign n5336 = n1310 & n5335 ;
  assign n5337 = n5331 & ~n5336 ;
  assign n5339 = n5338 ^ n5337 ;
  assign n5341 = n5330 ^ n1310 ;
  assign n5340 = n1310 & n4475 ;
  assign n5342 = n5341 ^ n5340 ;
  assign n5343 = n5342 ^ n3729 ;
  assign n5344 = n5343 ^ n5342 ;
  assign n5346 = n5342 ^ n5341 ;
  assign n5349 = ~n829 & n5346 ;
  assign n5350 = n5344 & n5349 ;
  assign n5351 = n5350 ^ n5344 ;
  assign n5352 = n5351 ^ n5343 ;
  assign n5353 = ~n753 & n5352 ;
  assign n5354 = ~n5339 & ~n5353 ;
  assign n5399 = n5398 ^ n5354 ;
  assign n5325 = n5279 ^ n5260 ;
  assign n5326 = n5265 & ~n5325 ;
  assign n5327 = n5326 ^ n5260 ;
  assign n5400 = n5399 ^ n5327 ;
  assign n5413 = n5412 ^ n5400 ;
  assign n5301 = ~n5202 & n5280 ;
  assign n5302 = n5200 ^ n5127 ;
  assign n5303 = n5302 ^ n5280 ;
  assign n5304 = n5148 ^ n5048 ;
  assign n5305 = n5049 ^ n5048 ;
  assign n5306 = n5305 ^ n5048 ;
  assign n5307 = n5304 & n5306 ;
  assign n5308 = n5307 ^ n5048 ;
  assign n5309 = ~n5303 & n5308 ;
  assign n5310 = n5280 ^ n5203 ;
  assign n5311 = n5310 ^ n5126 ;
  assign n5312 = n5311 ^ n5052 ;
  assign n5313 = n5312 ^ n5310 ;
  assign n5315 = ~n5052 & n5280 ;
  assign n5316 = n5315 ^ n5310 ;
  assign n5317 = n5313 & ~n5316 ;
  assign n5318 = n5317 ^ n5310 ;
  assign n5319 = ~n5148 & ~n5318 ;
  assign n5320 = n5319 ^ n5200 ;
  assign n5321 = ~n5309 & n5320 ;
  assign n5322 = n5321 ^ n5309 ;
  assign n5323 = n5301 & ~n5322 ;
  assign n5324 = n5323 ^ n5321 ;
  assign n5414 = n5413 ^ n5324 ;
  assign n5431 = n5430 ^ n5414 ;
  assign n5298 = n5284 ^ n5190 ;
  assign n5299 = ~n5285 & ~n5298 ;
  assign n5300 = n5299 ^ n5284 ;
  assign n5432 = n5431 ^ n5300 ;
  assign n5295 = ~n5286 & n5287 ;
  assign n5296 = n4194 & ~n5295 ;
  assign n5292 = n5186 & n5286 ;
  assign n5293 = ~n4194 & ~n5292 ;
  assign n5294 = n5293 ^ n4194 ;
  assign n5297 = n5296 ^ n5294 ;
  assign n5433 = n5432 ^ n5297 ;
  assign n5537 = ~n5414 & ~n5430 ;
  assign n5528 = n5327 & n5399 ;
  assign n5525 = n5400 ^ n5324 ;
  assign n5526 = n5413 & n5525 ;
  assign n5523 = n5408 & n5411 ;
  assign n5517 = n2737 ^ n2721 ;
  assign n5518 = ~n696 & n5517 ;
  assign n5506 = n5075 ^ n3694 ;
  assign n5504 = n2820 ^ n2721 ;
  assign n5505 = ~n696 & n5504 ;
  assign n5507 = n5506 ^ n5505 ;
  assign n5508 = n753 & n5507 ;
  assign n5509 = n5508 ^ n2659 ;
  assign n5510 = ~n738 & ~n5509 ;
  assign n5512 = ~n2659 & n3141 ;
  assign n5511 = ~n2820 & n5847 ;
  assign n5513 = n5512 ^ n5511 ;
  assign n5514 = n5513 ^ n754 ;
  assign n5515 = ~n5510 & ~n5514 ;
  assign n5501 = n739 & ~n3688 ;
  assign n5502 = n5501 ^ n2662 ;
  assign n5503 = n754 & ~n5502 ;
  assign n5516 = n5515 ^ n5503 ;
  assign n5519 = n5518 ^ n5516 ;
  assign n5468 = ~n2689 & n2906 ;
  assign n5467 = n2901 & n3729 ;
  assign n5469 = n5468 ^ n5467 ;
  assign n5470 = n5469 ^ n1310 ;
  assign n5471 = n5470 ^ n5469 ;
  assign n5472 = n5469 ^ n4608 ;
  assign n5473 = n5472 ^ n5469 ;
  assign n5474 = n5471 & ~n5473 ;
  assign n5475 = n5474 ^ n5469 ;
  assign n5476 = ~n753 & n5475 ;
  assign n5480 = n5469 ^ n753 ;
  assign n5477 = n4041 ^ n829 ;
  assign n5478 = n1310 & ~n4044 ;
  assign n5479 = ~n5477 & n5478 ;
  assign n5481 = n5480 ^ n5479 ;
  assign n5486 = n5481 ^ n1310 ;
  assign n5487 = n5486 ^ n5481 ;
  assign n5488 = n4206 ^ n4042 ;
  assign n5491 = n5487 & n5488 ;
  assign n5492 = n5480 & n5491 ;
  assign n5493 = n5492 ^ n5480 ;
  assign n5484 = n5481 ^ n5480 ;
  assign n5494 = n5493 ^ n5484 ;
  assign n5495 = ~n5476 & ~n5494 ;
  assign n5463 = n5396 ^ n5371 ;
  assign n5464 = n5396 ^ n5075 ;
  assign n5465 = ~n5463 & n5464 ;
  assign n5466 = n5465 ^ n5075 ;
  assign n5496 = n5495 ^ n5466 ;
  assign n5520 = n5519 ^ n5496 ;
  assign n5448 = n1021 & ~n4226 ;
  assign n5449 = n5448 ^ n1017 ;
  assign n5450 = ~n4205 & ~n5449 ;
  assign n5451 = n5450 ^ n1017 ;
  assign n5452 = ~n2862 & ~n5451 ;
  assign n5453 = n2863 ^ n1017 ;
  assign n5457 = ~n1022 & ~n4226 ;
  assign n5458 = n5453 & n5457 ;
  assign n5459 = n5458 ^ n5453 ;
  assign n5460 = n5459 ^ n2863 ;
  assign n5461 = ~n5452 & n5460 ;
  assign n5443 = n5366 ^ n5354 ;
  assign n5444 = ~n5398 & ~n5443 ;
  assign n5445 = n5444 ^ n5366 ;
  assign n5462 = n5461 ^ n5445 ;
  assign n5521 = n5520 ^ n5462 ;
  assign n5522 = n5521 ^ n5412 ;
  assign n5524 = n5523 ^ n5522 ;
  assign n5527 = n5526 ^ n5524 ;
  assign n5529 = n5528 ^ n5527 ;
  assign n5437 = n322 ^ n171 ;
  assign n5435 = n2381 ^ n109 ;
  assign n5436 = n5435 ^ n268 ;
  assign n5438 = n5437 ^ n5436 ;
  assign n5439 = n5438 ^ n4344 ;
  assign n5434 = n5165 ^ n858 ;
  assign n5440 = n5439 ^ n5434 ;
  assign n5441 = n5440 ^ n3895 ;
  assign n5442 = n2462 & ~n5441 ;
  assign n5530 = n5529 ^ n5442 ;
  assign n5531 = n5530 ^ n5293 ;
  assign n5532 = n5531 ^ n5296 ;
  assign n5533 = n5532 ^ n5530 ;
  assign n5534 = n5533 ^ n5300 ;
  assign n5535 = ~n5432 & ~n5534 ;
  assign n5536 = n5535 ^ n5531 ;
  assign n5538 = n5537 ^ n5536 ;
  assign n5539 = n5295 & ~n5432 ;
  assign n5540 = n5530 ^ n5430 ;
  assign n5541 = n5540 ^ n5530 ;
  assign n5542 = n5530 ^ n5300 ;
  assign n5543 = n5542 ^ n5530 ;
  assign n5544 = n5541 & ~n5543 ;
  assign n5545 = n5544 ^ n5530 ;
  assign n5546 = n5539 & ~n5545 ;
  assign n5658 = ~n4194 & ~n5546 ;
  assign n5659 = n5292 & n5432 ;
  assign n5660 = ~n5541 & n5543 ;
  assign n5661 = n5660 ^ n5530 ;
  assign n5662 = n5659 & ~n5661 ;
  assign n5663 = n5658 & ~n5662 ;
  assign n5648 = n3936 ^ n511 ;
  assign n5649 = n5648 ^ n180 ;
  assign n5647 = n2499 ^ n254 ;
  assign n5650 = n5649 ^ n5647 ;
  assign n5651 = n5650 ^ n4353 ;
  assign n5652 = ~n504 & ~n5651 ;
  assign n5653 = n3960 ^ n1226 ;
  assign n5654 = n5652 & n5653 ;
  assign n5611 = ~n2662 & n3146 ;
  assign n5628 = n2662 ^ n2659 ;
  assign n5629 = n5628 ^ n751 ;
  assign n5630 = n5629 ^ n696 ;
  assign n5631 = n5630 ^ n5628 ;
  assign n5632 = n696 & ~n2662 ;
  assign n5633 = n5632 ^ n5628 ;
  assign n5634 = n5631 & n5633 ;
  assign n5635 = n5634 ^ n5628 ;
  assign n5636 = ~n754 & n5635 ;
  assign n5637 = n5636 ^ n754 ;
  assign n5638 = n738 & ~n5637 ;
  assign n5626 = n2659 & n3147 ;
  assign n5620 = n2662 ^ n696 ;
  assign n5612 = n2689 ^ n696 ;
  assign n5615 = n5612 ^ n2754 ;
  assign n5616 = n5615 ^ n5612 ;
  assign n5617 = n739 & ~n5616 ;
  assign n5618 = n5617 ^ n5612 ;
  assign n5619 = n754 & n5618 ;
  assign n5621 = n5619 ^ n754 ;
  assign n5622 = n5621 ^ n799 ;
  assign n5623 = n5622 ^ n5619 ;
  assign n5624 = n5620 & ~n5623 ;
  assign n5625 = n5624 ^ n5621 ;
  assign n5627 = n5626 ^ n5625 ;
  assign n5639 = n5638 ^ n5627 ;
  assign n5640 = n5639 ^ n5619 ;
  assign n5641 = n5611 & n5640 ;
  assign n5642 = n5641 ^ n5639 ;
  assign n5607 = n5516 ^ n2737 ;
  assign n5608 = ~n5517 & n5607 ;
  assign n5609 = ~n696 & n5608 ;
  assign n5603 = n5505 ^ n1017 ;
  assign n5602 = n5516 ^ n696 ;
  assign n5604 = n5603 ^ n5602 ;
  assign n5610 = n5609 ^ n5604 ;
  assign n5643 = n5642 ^ n5610 ;
  assign n5599 = n5519 ^ n5466 ;
  assign n5600 = ~n5496 & ~n5599 ;
  assign n5601 = n5600 ^ n5519 ;
  assign n5644 = n5643 ^ n5601 ;
  assign n5586 = n2901 & ~n4041 ;
  assign n5585 = n2906 & n3729 ;
  assign n5587 = n5586 ^ n5585 ;
  assign n5591 = n5587 ^ n753 ;
  assign n5588 = n753 & n5587 ;
  assign n5592 = n5591 ^ n5588 ;
  assign n5595 = n1310 & ~n4464 ;
  assign n5596 = ~n5592 & n5595 ;
  assign n5582 = n4226 ^ n829 ;
  assign n5583 = n1310 & ~n4206 ;
  assign n5584 = n5582 & n5583 ;
  assign n5589 = n5588 ^ n5584 ;
  assign n5581 = n4286 & n4465 ;
  assign n5590 = n5589 ^ n5581 ;
  assign n5593 = n5592 ^ n5590 ;
  assign n5597 = n5596 ^ n5593 ;
  assign n5578 = n5520 ^ n5445 ;
  assign n5579 = ~n5462 & n5578 ;
  assign n5580 = n5579 ^ n5520 ;
  assign n5598 = n5597 ^ n5580 ;
  assign n5645 = n5644 ^ n5598 ;
  assign n5560 = n5521 ^ n5408 ;
  assign n5557 = ~n5327 & ~n5399 ;
  assign n5559 = n5557 ^ n5400 ;
  assign n5561 = n5560 ^ n5559 ;
  assign n5562 = n5561 ^ n5411 ;
  assign n5563 = ~n5408 & ~n5411 ;
  assign n5564 = n5563 ^ n5521 ;
  assign n5565 = ~n5562 & ~n5564 ;
  assign n5566 = n5565 ^ n5521 ;
  assign n5558 = ~n5523 & n5557 ;
  assign n5567 = n5566 ^ n5558 ;
  assign n5568 = n5324 & ~n5567 ;
  assign n5569 = n5521 ^ n5399 ;
  assign n5570 = n5569 ^ n5522 ;
  assign n5571 = n5521 ^ n5327 ;
  assign n5572 = n5571 ^ n5522 ;
  assign n5573 = ~n5570 & ~n5572 ;
  assign n5574 = n5573 ^ n5522 ;
  assign n5575 = ~n5564 & ~n5574 ;
  assign n5576 = n5575 ^ n5521 ;
  assign n5577 = ~n5568 & n5576 ;
  assign n5646 = n5645 ^ n5577 ;
  assign n5655 = n5654 ^ n5646 ;
  assign n5547 = n5529 ^ n5414 ;
  assign n5548 = n5547 ^ n5300 ;
  assign n5549 = n5548 ^ n5430 ;
  assign n5550 = n5549 ^ n5547 ;
  assign n5551 = n5442 ^ n5300 ;
  assign n5552 = n5551 ^ n5547 ;
  assign n5553 = n5550 & ~n5552 ;
  assign n5554 = n5553 ^ n5547 ;
  assign n5555 = ~n5530 & ~n5554 ;
  assign n5556 = n5555 ^ n5529 ;
  assign n5656 = n5655 ^ n5556 ;
  assign n5657 = n5656 ^ n5546 ;
  assign n5664 = n5663 ^ n5657 ;
  assign n5665 = ~n5656 & n5662 ;
  assign n5666 = ~n4194 & ~n5665 ;
  assign n5722 = n5546 & n5656 ;
  assign n5725 = n5666 & ~n5722 ;
  assign n5716 = n1117 ^ n1042 ;
  assign n5713 = n421 ^ n316 ;
  assign n5714 = n5713 ^ n328 ;
  assign n5715 = n5714 ^ n705 ;
  assign n5717 = n5716 ^ n5715 ;
  assign n5712 = n4034 ^ n1110 ;
  assign n5718 = n5717 ^ n5712 ;
  assign n5719 = n616 & n5718 ;
  assign n5709 = n5598 ^ n5577 ;
  assign n5710 = n5645 & n5709 ;
  assign n5704 = n1310 & n1537 ;
  assign n5705 = n4466 & n5704 ;
  assign n5701 = n2906 & ~n4041 ;
  assign n5700 = n2901 & ~n4226 ;
  assign n5702 = n5701 ^ n5700 ;
  assign n5703 = n5702 ^ n753 ;
  assign n5706 = n5705 ^ n5703 ;
  assign n5690 = ~n3715 & n5689 ;
  assign n5687 = n3149 & ~n4945 ;
  assign n5688 = n5687 ^ n5612 ;
  assign n5691 = n5690 ^ n5688 ;
  assign n5684 = ~n696 & ~n4950 ;
  assign n5685 = n5684 ^ n2689 ;
  assign n5686 = ~n3142 & ~n5685 ;
  assign n5692 = n5691 ^ n5686 ;
  assign n5682 = n754 & n3729 ;
  assign n5693 = n5692 ^ n5682 ;
  assign n5674 = n2721 ^ n1017 ;
  assign n5675 = ~n5504 & n5674 ;
  assign n5676 = n5675 ^ n1017 ;
  assign n5677 = ~n2659 & ~n5676 ;
  assign n5678 = n5676 ^ n2659 ;
  assign n5679 = n5678 ^ n5677 ;
  assign n5680 = ~n696 & n5679 ;
  assign n5681 = ~n5677 & n5680 ;
  assign n5694 = n5693 ^ n5681 ;
  assign n5696 = n5694 ^ n5603 ;
  assign n5695 = n5694 ^ n5642 ;
  assign n5697 = n5696 ^ n5695 ;
  assign n5698 = ~n5610 & n5697 ;
  assign n5699 = n5698 ^ n5696 ;
  assign n5707 = n5706 ^ n5699 ;
  assign n5672 = n5601 & n5643 ;
  assign n5670 = n5580 & n5597 ;
  assign n5671 = n5670 ^ n5598 ;
  assign n5673 = n5672 ^ n5671 ;
  assign n5708 = n5707 ^ n5673 ;
  assign n5711 = n5710 ^ n5708 ;
  assign n5720 = n5719 ^ n5711 ;
  assign n5667 = n5646 ^ n5556 ;
  assign n5668 = ~n5655 & n5667 ;
  assign n5669 = n5668 ^ n5646 ;
  assign n5721 = n5720 ^ n5669 ;
  assign n5723 = n5722 ^ n5721 ;
  assign n5726 = n5725 ^ n5723 ;
  assign n5727 = n5665 & ~n5721 ;
  assign n5728 = ~n4194 & ~n5727 ;
  assign n5808 = n5721 & n5722 ;
  assign n5795 = n2561 ^ n290 ;
  assign n5796 = n5795 ^ n159 ;
  assign n5797 = n5796 ^ n1123 ;
  assign n5798 = n5797 ^ n4381 ;
  assign n5799 = n5798 ^ n2312 ;
  assign n5800 = ~n2543 & n5799 ;
  assign n5803 = ~n251 & n1092 ;
  assign n5801 = n389 ^ n238 ;
  assign n5802 = n5801 ^ n384 ;
  assign n5804 = n5803 ^ n5802 ;
  assign n5805 = n5800 & ~n5804 ;
  assign n5790 = n5706 ^ n5694 ;
  assign n5791 = n5699 & ~n5790 ;
  assign n5792 = n5791 ^ n5694 ;
  assign n5788 = ~n5680 & ~n5693 ;
  assign n5785 = n5677 & n5693 ;
  assign n5786 = n5785 ^ n2662 ;
  assign n5787 = ~n696 & n5786 ;
  assign n5789 = n5788 ^ n5787 ;
  assign n5793 = n5792 ^ n5789 ;
  assign n5765 = n5672 ^ n5644 ;
  assign n5766 = n5707 ^ n5670 ;
  assign n5767 = n5765 & n5766 ;
  assign n5768 = ~n5577 & n5767 ;
  assign n5769 = n5707 ^ n5672 ;
  assign n5770 = n5769 ^ n5707 ;
  assign n5771 = n5707 ^ n5671 ;
  assign n5772 = n5771 ^ n5707 ;
  assign n5773 = ~n5770 & ~n5772 ;
  assign n5774 = n5773 ^ n5707 ;
  assign n5775 = n5768 & ~n5774 ;
  assign n5776 = n5775 ^ n5767 ;
  assign n5777 = n5580 ^ n5577 ;
  assign n5778 = n5598 & n5777 ;
  assign n5779 = n5778 ^ n5580 ;
  assign n5780 = ~n5776 & n5779 ;
  assign n5782 = n5780 ^ n5776 ;
  assign n5764 = ~n5672 & ~n5707 ;
  assign n5781 = n5764 & n5780 ;
  assign n5783 = n5782 ^ n5781 ;
  assign n5751 = ~n2689 & n3149 ;
  assign n5750 = n3142 & n3729 ;
  assign n5752 = n5751 ^ n5750 ;
  assign n5756 = n5752 ^ n696 ;
  assign n5753 = n696 & n5752 ;
  assign n5757 = n5756 ^ n5753 ;
  assign n5760 = n754 & n5488 ;
  assign n5761 = ~n5757 & n5760 ;
  assign n5747 = n4041 ^ n738 ;
  assign n5748 = n754 & ~n4044 ;
  assign n5749 = n5747 & n5748 ;
  assign n5754 = n5753 ^ n5749 ;
  assign n5746 = ~n4608 & n4907 ;
  assign n5755 = n5754 ^ n5746 ;
  assign n5758 = n5757 ^ n5755 ;
  assign n5762 = n5761 ^ n5758 ;
  assign n5734 = ~n829 & ~n4226 ;
  assign n5735 = n5734 ^ n753 ;
  assign n5736 = ~n4205 & ~n5735 ;
  assign n5737 = n5736 ^ n753 ;
  assign n5738 = ~n2899 & ~n5737 ;
  assign n5743 = n2904 & ~n4226 ;
  assign n5744 = n5743 ^ n753 ;
  assign n5745 = ~n5738 & n5744 ;
  assign n5763 = n5762 ^ n5745 ;
  assign n5784 = n5783 ^ n5763 ;
  assign n5794 = n5793 ^ n5784 ;
  assign n5806 = n5805 ^ n5794 ;
  assign n5729 = n5711 ^ n5669 ;
  assign n5730 = ~n5720 & n5729 ;
  assign n5731 = n5730 ^ n5711 ;
  assign n5807 = n5806 ^ n5731 ;
  assign n5809 = n5808 ^ n5807 ;
  assign n5810 = n5809 ^ n5807 ;
  assign n5811 = n5728 & ~n5810 ;
  assign n5812 = n5811 ^ n5809 ;
  assign n5813 = n5727 & ~n5807 ;
  assign n5814 = ~n4194 & ~n5813 ;
  assign n5902 = n5807 & n5808 ;
  assign n5905 = n5814 & ~n5902 ;
  assign n5895 = ~n297 & n1105 ;
  assign n5891 = n2415 ^ n376 ;
  assign n5890 = n649 ^ n324 ;
  assign n5892 = n5891 ^ n5890 ;
  assign n5889 = n3947 ^ n1211 ;
  assign n5893 = n5892 ^ n5889 ;
  assign n5886 = n627 ^ n204 ;
  assign n5887 = n5886 ^ n2676 ;
  assign n5884 = n415 ^ n356 ;
  assign n5885 = n5884 ^ n443 ;
  assign n5888 = n5887 ^ n5885 ;
  assign n5894 = n5893 ^ n5888 ;
  assign n5896 = n5895 ^ n5894 ;
  assign n5897 = n438 & ~n5896 ;
  assign n5898 = n3925 & n5897 ;
  assign n5899 = ~n4356 & n5898 ;
  assign n5834 = n4226 ^ n738 ;
  assign n5835 = ~n4206 & n5834 ;
  assign n5853 = n5835 ^ n4465 ;
  assign n5854 = n4907 & n5853 ;
  assign n5231 = n3148 ^ n3141 ;
  assign n5232 = n5231 ^ n3149 ;
  assign n5832 = ~n4041 & ~n5232 ;
  assign n5830 = ~n696 & ~n3729 ;
  assign n5831 = ~n2616 & ~n5830 ;
  assign n5833 = n5832 ^ n5831 ;
  assign n5836 = n5835 ^ n4464 ;
  assign n5837 = ~n5833 & n5836 ;
  assign n5838 = n4041 ^ n696 ;
  assign n5850 = n2612 & n5838 ;
  assign n5848 = ~n3729 & n5847 ;
  assign n5842 = n696 & ~n3729 ;
  assign n5843 = n5842 ^ n5838 ;
  assign n5844 = ~n738 & ~n5843 ;
  assign n5845 = n5844 ^ n5838 ;
  assign n5846 = n799 & n5845 ;
  assign n5849 = n5848 ^ n5846 ;
  assign n5851 = n5850 ^ n5849 ;
  assign n5852 = ~n5837 & ~n5851 ;
  assign n5855 = n5854 ^ n5852 ;
  assign n5856 = n5855 ^ n753 ;
  assign n5825 = ~n2662 & n2687 ;
  assign n5826 = n5825 ^ n2662 ;
  assign n5827 = n5826 ^ n2689 ;
  assign n5828 = ~n696 & ~n5825 ;
  assign n5829 = ~n5827 & n5828 ;
  assign n5857 = n5856 ^ n5829 ;
  assign n5821 = ~n696 & n2662 ;
  assign n5822 = ~n5785 & ~n5788 ;
  assign n5823 = n5821 & n5822 ;
  assign n5824 = n5823 ^ n5788 ;
  assign n5858 = n5857 ^ n5824 ;
  assign n5818 = n5789 & ~n5792 ;
  assign n5878 = n5858 ^ n5818 ;
  assign n5859 = ~n5818 & n5858 ;
  assign n5879 = n5878 ^ n5859 ;
  assign n5869 = ~n5793 & ~n5858 ;
  assign n5880 = n5879 ^ n5869 ;
  assign n5868 = n5793 ^ n5783 ;
  assign n5861 = ~n5745 & n5762 ;
  assign n5872 = n5869 ^ n5861 ;
  assign n5873 = n5872 ^ n5763 ;
  assign n5874 = n5869 & n5873 ;
  assign n5875 = n5874 ^ n5763 ;
  assign n5876 = n5868 & ~n5875 ;
  assign n5877 = n5876 ^ n5872 ;
  assign n5881 = n5880 ^ n5877 ;
  assign n5882 = n5881 ^ n5859 ;
  assign n5819 = n5818 ^ n5793 ;
  assign n5820 = n5783 & ~n5819 ;
  assign n5860 = n5859 ^ n5818 ;
  assign n5862 = n5861 ^ n5763 ;
  assign n5865 = ~n5860 & ~n5862 ;
  assign n5866 = n5865 ^ n5818 ;
  assign n5867 = n5820 & ~n5866 ;
  assign n5883 = n5882 ^ n5867 ;
  assign n5900 = n5899 ^ n5883 ;
  assign n5815 = n5794 ^ n5731 ;
  assign n5816 = ~n5806 & n5815 ;
  assign n5817 = n5816 ^ n5794 ;
  assign n5901 = n5900 ^ n5817 ;
  assign n5903 = n5902 ^ n5901 ;
  assign n5906 = n5905 ^ n5903 ;
  assign n5907 = n5813 & ~n5901 ;
  assign n5908 = ~n4194 & ~n5907 ;
  assign n5970 = n5901 & n5902 ;
  assign n5973 = n5908 & ~n5970 ;
  assign n5959 = ~n753 & ~n5825 ;
  assign n5960 = ~n5827 & n5959 ;
  assign n5961 = n5960 ^ n5827 ;
  assign n5962 = n5961 ^ n3729 ;
  assign n5963 = ~n696 & ~n5962 ;
  assign n5956 = n4466 & n5955 ;
  assign n5947 = ~n696 & n4041 ;
  assign n5948 = n5947 ^ n696 ;
  assign n5949 = n5948 ^ n4226 ;
  assign n5950 = n738 & n5949 ;
  assign n5951 = n5950 ^ n4226 ;
  assign n5952 = ~n800 & n5951 ;
  assign n5953 = n5952 ^ n754 ;
  assign n5942 = n696 & ~n4041 ;
  assign n5943 = n5942 ^ n4226 ;
  assign n5944 = ~n738 & ~n5943 ;
  assign n5945 = n5944 ^ n4226 ;
  assign n5946 = n799 & n5945 ;
  assign n5954 = n5953 ^ n5946 ;
  assign n5957 = n5956 ^ n5954 ;
  assign n5938 = n5855 ^ n5824 ;
  assign n5939 = n5857 & n5938 ;
  assign n5940 = n5939 ^ n5855 ;
  assign n5958 = n5957 ^ n5940 ;
  assign n5964 = n5963 ^ n5958 ;
  assign n5922 = n5880 ^ n5861 ;
  assign n5923 = n5880 ^ n5859 ;
  assign n5924 = n5923 ^ n5880 ;
  assign n5925 = n5880 ^ n5783 ;
  assign n5926 = n5925 ^ n5880 ;
  assign n5927 = ~n5924 & n5926 ;
  assign n5928 = n5927 ^ n5880 ;
  assign n5929 = ~n5922 & ~n5928 ;
  assign n5930 = n5929 ^ n5861 ;
  assign n5931 = n5862 ^ n5858 ;
  assign n5932 = ~n5878 & ~n5931 ;
  assign n5933 = n5932 ^ n5858 ;
  assign n5934 = n5930 & n5933 ;
  assign n5935 = n5820 & n5862 ;
  assign n5936 = n5934 & n5935 ;
  assign n5937 = n5936 ^ n5934 ;
  assign n5965 = n5964 ^ n5937 ;
  assign n5916 = n243 ^ n226 ;
  assign n5917 = n5916 ^ n539 ;
  assign n5918 = n5917 ^ n2679 ;
  assign n5914 = n327 ^ n223 ;
  assign n5915 = n5914 ^ n2561 ;
  assign n5919 = n5918 ^ n5915 ;
  assign n5920 = n5919 ^ n1064 ;
  assign n5921 = n5920 ^ n1432 ;
  assign n5966 = n5965 ^ n5921 ;
  assign n5913 = ~n102 & n5419 ;
  assign n5967 = n5966 ^ n5913 ;
  assign n5912 = n470 & ~n2281 ;
  assign n5968 = n5967 ^ n5912 ;
  assign n5909 = n5883 ^ n5817 ;
  assign n5910 = ~n5900 & n5909 ;
  assign n5911 = n5910 ^ n5883 ;
  assign n5969 = n5968 ^ n5911 ;
  assign n5971 = n5970 ^ n5969 ;
  assign n5974 = n5973 ^ n5971 ;
  assign n5975 = n5969 & n5970 ;
  assign n5976 = n4194 & ~n5975 ;
  assign n6053 = n5907 & ~n5969 ;
  assign n6041 = n5916 ^ n435 ;
  assign n6042 = n6041 ^ n427 ;
  assign n6037 = n3876 ^ n291 ;
  assign n6038 = n6037 ^ n398 ;
  assign n6039 = n6038 ^ n1039 ;
  assign n6040 = n6039 ^ n268 ;
  assign n6043 = n6042 ^ n6040 ;
  assign n6044 = n6043 ^ n3914 ;
  assign n6045 = n6044 ^ n1195 ;
  assign n6046 = n6045 ^ n2565 ;
  assign n6047 = n1056 ^ n310 ;
  assign n6048 = n6047 ^ n1280 ;
  assign n6049 = n6046 & n6048 ;
  assign n6050 = ~n5804 & n6049 ;
  assign n5233 = ~n5689 ^ n696 ;
  assign n5234 = n5233 ^ n5232 ;
  assign n5981 = ~n4226 & ~n5234 ;
  assign n5982 = n754 & n4205 ;
  assign n5983 = n5981 & n5982 ;
  assign n5984 = n5983 ^ n5981 ;
  assign n5991 = n3729 & ~n5948 ;
  assign n6030 = ~n5984 & n5991 ;
  assign n5980 = ~n3729 & n4041 ;
  assign n5985 = n5984 ^ n5980 ;
  assign n5986 = n5985 ^ n696 ;
  assign n5987 = n5986 ^ n5984 ;
  assign n5988 = n5987 ^ n5957 ;
  assign n5989 = n5988 ^ n5980 ;
  assign n5990 = n5989 ^ n5988 ;
  assign n5992 = n5957 ^ n696 ;
  assign n5994 = n5992 ^ n5961 ;
  assign n5995 = n5962 & n5994 ;
  assign n5996 = ~n696 & n5995 ;
  assign n5997 = n5996 ^ n5992 ;
  assign n5998 = ~n5991 & n5997 ;
  assign n6001 = ~n5990 & ~n5998 ;
  assign n6002 = n6001 ^ n5988 ;
  assign n6003 = ~n5985 & n6002 ;
  assign n6026 = n5986 & ~n6003 ;
  assign n6027 = n5980 ^ n5957 ;
  assign n6028 = n6026 & ~n6027 ;
  assign n6007 = ~n3729 & ~n5984 ;
  assign n6012 = ~n5957 & ~n5961 ;
  assign n6013 = n6012 ^ n5947 ;
  assign n6014 = n6007 & n6013 ;
  assign n6004 = n5998 ^ n5997 ;
  assign n6015 = n6014 ^ n6004 ;
  assign n6020 = ~n5980 & n5984 ;
  assign n6021 = n5997 & n6020 ;
  assign n6022 = n6021 ^ n5997 ;
  assign n6016 = n5948 ^ n5830 ;
  assign n6017 = ~n5984 & ~n6016 ;
  assign n6018 = n6017 ^ n5984 ;
  assign n6019 = ~n5997 & n6018 ;
  assign n6023 = n6022 ^ n6019 ;
  assign n6024 = ~n6015 & n6023 ;
  assign n6005 = n6004 ^ n5988 ;
  assign n6006 = n6005 ^ n6003 ;
  assign n6025 = n6024 ^ n6006 ;
  assign n6029 = n6028 ^ n6025 ;
  assign n6031 = n6030 ^ n6029 ;
  assign n6032 = n5940 ^ n5937 ;
  assign n6033 = n5964 & n6032 ;
  assign n6034 = n6033 ^ n5937 ;
  assign n6035 = n6031 & n6034 ;
  assign n6036 = n6035 ^ n6024 ;
  assign n6051 = n6050 ^ n6036 ;
  assign n5977 = n5965 ^ n5911 ;
  assign n5978 = ~n5968 & n5977 ;
  assign n5979 = n5978 ^ n5965 ;
  assign n6052 = n6051 ^ n5979 ;
  assign n6054 = n6053 ^ n6052 ;
  assign n6055 = n6054 ^ n6052 ;
  assign n6056 = n5976 & ~n6055 ;
  assign n6057 = n6056 ^ n6054 ;
  assign n6058 = ~n6052 & n6053 ;
  assign n6059 = ~n4194 & ~n6058 ;
  assign n6125 = n5975 & n6052 ;
  assign n6128 = n6059 & ~n6125 ;
  assign n6071 = n4226 ^ n4041 ;
  assign n6073 = n4226 ^ n3729 ;
  assign n6076 = n6073 ^ n6071 ;
  assign n6081 = n6076 ^ n3729 ;
  assign n6072 = n6071 ^ n5848 ;
  assign n6074 = n6073 ^ n6072 ;
  assign n6082 = n6081 ^ n6074 ;
  assign n6083 = n6082 ^ n6071 ;
  assign n6085 = ~n6081 & ~n6083 ;
  assign n6075 = n6074 ^ n696 ;
  assign n6078 = n6074 ^ n6071 ;
  assign n6077 = n6076 ^ n696 ;
  assign n6079 = n6078 ^ n6077 ;
  assign n6080 = ~n6075 & ~n6079 ;
  assign n6086 = n6085 ^ n6080 ;
  assign n6087 = n6086 ^ n6078 ;
  assign n6088 = n6085 ^ n6076 ;
  assign n6089 = n6088 ^ n6078 ;
  assign n6090 = n6087 & ~n6089 ;
  assign n6091 = ~n6071 & n6090 ;
  assign n6092 = n6091 ^ n6085 ;
  assign n6093 = n6092 ^ n6083 ;
  assign n6106 = n6093 ^ n4226 ;
  assign n6107 = n6106 ^ n3729 ;
  assign n6114 = n696 & ~n5984 ;
  assign n6115 = n6107 & n6114 ;
  assign n6108 = n6107 ^ n6019 ;
  assign n6109 = n6108 ^ n6107 ;
  assign n6110 = n6022 ^ n6017 ;
  assign n6111 = n6034 & ~n6110 ;
  assign n6112 = ~n6109 & n6111 ;
  assign n6113 = n6112 ^ n6108 ;
  assign n6116 = n6115 ^ n6113 ;
  assign n6064 = n3924 ^ n226 ;
  assign n6063 = n286 ^ n280 ;
  assign n6065 = n6064 ^ n6063 ;
  assign n6066 = n6065 ^ n2636 ;
  assign n6067 = n6066 ^ n3885 ;
  assign n6068 = n6067 ^ n5892 ;
  assign n6069 = n6068 ^ n3909 ;
  assign n6070 = n6069 ^ n1116 ;
  assign n6117 = n6116 ^ n6070 ;
  assign n6118 = n6117 ^ n6116 ;
  assign n6119 = ~n2421 & ~n6118 ;
  assign n6121 = n98 & n2323 ;
  assign n6122 = n6119 & n6121 ;
  assign n6120 = n6119 ^ n6117 ;
  assign n6123 = n6122 ^ n6120 ;
  assign n6060 = n6036 ^ n5979 ;
  assign n6061 = ~n6051 & n6060 ;
  assign n6062 = n6061 ^ n6036 ;
  assign n6124 = n6123 ^ n6062 ;
  assign n6126 = n6125 ^ n6124 ;
  assign n6129 = n6128 ^ n6126 ;
  assign n6145 = n626 ^ n78 ;
  assign n6146 = ~n251 & n6145 ;
  assign n6140 = n868 ^ n492 ;
  assign n6141 = n6140 ^ n5886 ;
  assign n6137 = n338 ^ n161 ;
  assign n6138 = n6137 ^ n2600 ;
  assign n6139 = n6138 ^ n136 ;
  assign n6142 = n6141 ^ n6139 ;
  assign n6143 = n6142 ^ n687 ;
  assign n6144 = n6143 ^ n2644 ;
  assign n6147 = n6146 ^ n6144 ;
  assign n6134 = n6116 ^ n6062 ;
  assign n6135 = n6123 & n6134 ;
  assign n6136 = n6135 ^ n6116 ;
  assign n6148 = n6147 ^ n6136 ;
  assign n6132 = n6058 & n6124 ;
  assign n6149 = n6148 ^ n6132 ;
  assign n6130 = ~n6124 & n6125 ;
  assign n6131 = n4194 & ~n6130 ;
  assign n6133 = n6131 & ~n6132 ;
  assign n6150 = n6149 ^ n6133 ;
  assign n6165 = ~n6136 & ~n6147 ;
  assign n6158 = n4558 ^ n3882 ;
  assign n6157 = n1032 ^ n592 ;
  assign n6159 = n6158 ^ n6157 ;
  assign n6160 = n6159 ^ n1244 ;
  assign n6156 = n1054 ^ n423 ;
  assign n6161 = n6160 ^ n6156 ;
  assign n6162 = n6161 ^ n633 ;
  assign n6163 = n6162 ^ n1188 ;
  assign n6164 = n3941 & ~n6163 ;
  assign n6166 = n6165 ^ n6164 ;
  assign n6151 = n6148 ^ n4194 ;
  assign n6152 = n6132 ^ n6130 ;
  assign n6153 = n6148 & n6152 ;
  assign n6154 = n6153 ^ n6130 ;
  assign n6155 = n6151 & ~n6154 ;
  assign n6167 = n6166 ^ n6155 ;
  assign n6181 = n218 ^ n132 ;
  assign n6182 = n6181 ^ n533 ;
  assign n6183 = n6182 ^ n135 ;
  assign n6179 = n428 ^ n415 ;
  assign n6180 = n6179 ^ n2459 ;
  assign n6184 = n6183 ^ n6180 ;
  assign n6185 = n6184 ^ n4996 ;
  assign n6186 = ~n342 & n6185 ;
  assign n6187 = n1082 & n6186 ;
  assign n6188 = n6048 & n6187 ;
  assign n6175 = n6136 ^ n6132 ;
  assign n6176 = n6148 & n6175 ;
  assign n6177 = n6176 ^ n6136 ;
  assign n6178 = ~n6164 & n6177 ;
  assign n6189 = n6188 ^ n6178 ;
  assign n6171 = n6130 & n6165 ;
  assign n6172 = n6171 ^ n6164 ;
  assign n6173 = n6154 & ~n6172 ;
  assign n6174 = n4194 & ~n6173 ;
  assign n6190 = n6189 ^ n6174 ;
  assign n6197 = n372 ^ n61 ;
  assign n6196 = n516 ^ n166 ;
  assign n6198 = n6197 ^ n6196 ;
  assign n6194 = n4211 ^ n132 ;
  assign n6195 = n509 & n6194 ;
  assign n6199 = n6198 ^ n6195 ;
  assign n6200 = ~n4998 & n6199 ;
  assign n6201 = n6200 ^ n2674 ;
  assign n6202 = n1066 & n6201 ;
  assign n6203 = n5421 & n6202 ;
  assign n6204 = n6203 ^ n4194 ;
  assign n6191 = n6174 ^ n4194 ;
  assign n6192 = n6191 ^ n6178 ;
  assign n6193 = n6189 & n6192 ;
  assign n6205 = n6204 ^ n6193 ;
  assign n6214 = n6203 ^ n6188 ;
  assign n6215 = n6193 & ~n6214 ;
  assign n6206 = n116 ^ n101 ;
  assign n6207 = n653 ^ n357 ;
  assign n6208 = n6207 ^ n727 ;
  assign n6209 = n6208 ^ n3723 ;
  assign n6210 = ~n688 & ~n6209 ;
  assign n6211 = n6206 & n6210 ;
  assign n6212 = n6211 ^ n6209 ;
  assign n6213 = n6212 ^ n4194 ;
  assign n6216 = n6215 ^ n6213 ;
  assign n6224 = ~n6188 & ~n6203 ;
  assign n6225 = n6178 & n6212 ;
  assign n6226 = n6224 & n6225 ;
  assign n6223 = n1144 & ~n3719 ;
  assign n6227 = n6226 ^ n6223 ;
  assign n6217 = n6212 ^ n6203 ;
  assign n6218 = n6173 & n6217 ;
  assign n6219 = n6212 ^ n6178 ;
  assign n6220 = n6189 & ~n6219 ;
  assign n6221 = n6218 & n6220 ;
  assign n6222 = n4194 & ~n6221 ;
  assign n6228 = n6227 ^ n6222 ;
  assign n6229 = n6223 & ~n6226 ;
  assign n6230 = n6229 ^ n6227 ;
  assign n6231 = ~n6191 & n6230 ;
  assign n6232 = n6231 ^ n4194 ;
  assign n6233 = ~x21 & ~x22 ;
  assign n6234 = n6229 & ~n6233 ;
  assign n6235 = n6221 & n6234 ;
  assign n6238 = n6235 ^ n6233 ;
  assign n6239 = n6238 ^ n6235 ;
  assign n6240 = n944 & n6239 ;
  assign n6241 = n6240 ^ n6235 ;
  assign n6242 = ~n6232 & ~n6241 ;
  assign n6243 = n6242 ^ n6235 ;
  assign n6244 = n4194 & ~n6235 ;
  assign y0 = ~n4193 ;
  assign y1 = ~n4361 ;
  assign y2 = n4533 ;
  assign y3 = ~n4705 ;
  assign y4 = n4875 ;
  assign y5 = n5017 ;
  assign y6 = ~n5185 ;
  assign y7 = ~n5291 ;
  assign y8 = ~n5433 ;
  assign y9 = n5538 ;
  assign y10 = n5664 ;
  assign y11 = n5726 ;
  assign y12 = n5812 ;
  assign y13 = n5906 ;
  assign y14 = n5974 ;
  assign y15 = ~n6057 ;
  assign y16 = ~n6129 ;
  assign y17 = n6150 ;
  assign y18 = n6167 ;
  assign y19 = ~n6190 ;
  assign y20 = ~n6205 ;
  assign y21 = n6216 ;
  assign y22 = ~n6228 ;
  assign y23 = ~n6243 ;
  assign y24 = n6244 ;
endmodule
