module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n212 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n279 , n280 , n281 , n282 , n283 , n284 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n328 , n329 , n330 , n331 , n332 , n333 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n383 , n384 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n501 , n502 , n503 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n563 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2535 , n2536 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2556 , n2557 , n2558 , n2559 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3820 , n3821 , n3822 , n3823 , n3825 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4562 , n4563 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5138 , n5139 , n5140 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5367 , n5368 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6305 , n6306 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6929 , n6930 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7358 , n7359 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8078 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8800 , n8801 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9153 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10321 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11054 , n11055 , n11058 , n11059 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11078 , n11079 , n11080 , n11081 , n11083 , n11084 , n11085 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11501 , n11502 , n11503 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11605 , n11606 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12005 , n12006 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14159 , n14160 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15117 , n15118 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15159 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15610 , n15611 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 ;
  assign n130 = ~x126 & ~x127 ;
  assign n131 = ~x125 & n130 ;
  assign n132 = ~x124 & n131 ;
  assign n133 = ~x123 & n132 ;
  assign n134 = ~x122 & n133 ;
  assign n135 = ~x121 & n134 ;
  assign n136 = ~x120 & n135 ;
  assign n137 = ~x119 & n136 ;
  assign n138 = ~x118 & n137 ;
  assign n139 = ~x117 & n138 ;
  assign n140 = ~x116 & n139 ;
  assign n141 = ~x115 & n140 ;
  assign n142 = ~x114 & n141 ;
  assign n143 = ~x111 & ~x112 ;
  assign n144 = ~x113 & ~x114 ;
  assign n145 = n143 & n144 ;
  assign n146 = n141 & n145 ;
  assign n147 = ~x110 & n146 ;
  assign n148 = ~x109 & n147 ;
  assign n6318 = ~x108 & n148 ;
  assign n149 = ~x106 & ~x107 ;
  assign n6319 = n149 & n6318 ;
  assign n150 = ~x104 & ~x105 ;
  assign n151 = ~x108 & n150 ;
  assign n152 = n149 & n151 ;
  assign n153 = n148 & n152 ;
  assign n154 = ~x103 & n153 ;
  assign n155 = ~x102 & n154 ;
  assign n156 = ~x101 & n155 ;
  assign n157 = ~x100 & n156 ;
  assign n158 = ~x99 & n157 ;
  assign n159 = ~x98 & n158 ;
  assign n160 = ~x97 & n159 ;
  assign n161 = ~x96 & n160 ;
  assign n162 = ~x95 & n161 ;
  assign n163 = ~x94 & n162 ;
  assign n164 = ~x93 & n163 ;
  assign n165 = ~x92 & n164 ;
  assign n168 = ~x91 & n165 ;
  assign n169 = ~x90 & n168 ;
  assign n170 = ~x89 & n169 ;
  assign n171 = ~x88 & n170 ;
  assign n172 = ~x87 & n171 ;
  assign n173 = ~x85 & ~x86 ;
  assign n174 = n172 & n173 ;
  assign n175 = ~x84 & ~x87 ;
  assign n176 = n173 & n175 ;
  assign n177 = n171 & n176 ;
  assign n178 = ~x83 & n177 ;
  assign n179 = ~x82 & n178 ;
  assign n180 = ~x81 & n179 ;
  assign n181 = ~x80 & n180 ;
  assign n182 = ~x79 & n181 ;
  assign n183 = ~x78 & n182 ;
  assign n184 = ~x77 & n183 ;
  assign n185 = ~x76 & n184 ;
  assign n186 = ~x75 & n185 ;
  assign n187 = ~x74 & n186 ;
  assign n188 = ~x73 & n187 ;
  assign n189 = ~x72 & n188 ;
  assign n240 = x65 ^ x61 ;
  assign n239 = x61 & ~x65 ;
  assign n241 = n240 ^ n239 ;
  assign n190 = ~x71 & n189 ;
  assign n191 = ~x70 & n190 ;
  assign n192 = ~x69 & n191 ;
  assign n193 = ~x68 & n192 ;
  assign n194 = ~x67 & n193 ;
  assign n217 = ~x66 & n194 ;
  assign n218 = ~x63 & x65 ;
  assign n219 = n217 & n218 ;
  assign n220 = n219 ^ n217 ;
  assign n237 = x64 & n220 ;
  assign n238 = n237 ^ x62 ;
  assign n245 = n241 ^ n238 ;
  assign n242 = n237 & n241 ;
  assign n243 = n238 & n242 ;
  assign n244 = n243 ^ n238 ;
  assign n246 = n245 ^ n244 ;
  assign n247 = x65 ^ x60 ;
  assign n196 = x65 ^ x64 ;
  assign n197 = ~x66 & ~n196 ;
  assign n198 = x65 & n197 ;
  assign n199 = x62 & n198 ;
  assign n200 = n199 ^ n197 ;
  assign n201 = n200 ^ x66 ;
  assign n248 = x63 & n201 ;
  assign n249 = n248 ^ x66 ;
  assign n212 = n240 ^ x62 ;
  assign n215 = x64 & ~n212 ;
  assign n216 = n215 ^ x62 ;
  assign n223 = n215 ^ x64 ;
  assign n224 = ~n220 & n223 ;
  assign n221 = n220 ^ n196 ;
  assign n225 = n224 ^ n221 ;
  assign n226 = n225 ^ n220 ;
  assign n227 = ~n216 & n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n228 ^ x65 ;
  assign n230 = n229 ^ n196 ;
  assign n250 = n230 ^ x63 ;
  assign n251 = n250 ^ n194 ;
  assign n252 = ~n249 & n251 ;
  assign n253 = n252 ^ x63 ;
  assign n254 = n194 & n253 ;
  assign n255 = n254 ^ x61 ;
  assign n256 = n255 ^ x60 ;
  assign n257 = ~n247 & n256 ;
  assign n258 = n257 ^ x60 ;
  assign n259 = x64 & ~n258 ;
  assign n260 = ~n246 & ~n259 ;
  assign n261 = n260 ^ x66 ;
  assign n267 = ~x62 & n237 ;
  assign n268 = n267 ^ n244 ;
  assign n263 = n239 ^ x65 ;
  assign n264 = x64 & ~n263 ;
  assign n265 = n264 ^ x65 ;
  assign n266 = n254 & n265 ;
  assign n269 = n268 ^ n266 ;
  assign n270 = n269 ^ n260 ;
  assign n271 = ~n261 & ~n270 ;
  assign n272 = n271 ^ x66 ;
  assign n195 = x63 & n194 ;
  assign n233 = n201 & ~n230 ;
  assign n234 = n233 ^ x66 ;
  assign n235 = n195 & ~n234 ;
  assign n236 = n235 ^ x63 ;
  assign n374 = n194 & n236 ;
  assign n375 = ~n272 & n374 ;
  assign n273 = n272 ^ x67 ;
  assign n274 = n193 & n273 ;
  assign n275 = n236 & n274 ;
  assign n276 = n275 ^ n236 ;
  assign n277 = n192 & n276 ;
  assign n316 = x68 ^ x67 ;
  assign n279 = ~x67 & ~n235 ;
  assign n280 = n279 ^ x63 ;
  assign n281 = n273 ^ n193 ;
  assign n282 = n280 & ~n281 ;
  assign n283 = n282 ^ x67 ;
  assign n284 = n193 & ~n283 ;
  assign n311 = ~n261 & n284 ;
  assign n312 = n311 ^ n269 ;
  assign n293 = x65 & n284 ;
  assign n289 = ~x60 & n284 ;
  assign n290 = n289 ^ n254 ;
  assign n291 = x64 & n290 ;
  assign n292 = n291 ^ x61 ;
  assign n294 = n293 ^ n292 ;
  assign n295 = n294 ^ x66 ;
  assign n297 = x65 ^ x59 ;
  assign n298 = x64 ^ x60 ;
  assign n299 = n298 ^ x65 ;
  assign n300 = n299 ^ n284 ;
  assign n301 = ~n297 & n300 ;
  assign n296 = x60 & x65 ;
  assign n302 = n301 ^ n296 ;
  assign n305 = x64 & n302 ;
  assign n306 = n305 ^ n296 ;
  assign n307 = n306 ^ x65 ;
  assign n308 = n307 ^ n294 ;
  assign n309 = ~n295 & n308 ;
  assign n310 = n309 ^ x66 ;
  assign n313 = n312 ^ n310 ;
  assign n314 = n312 ^ x67 ;
  assign n315 = n313 & ~n314 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = n277 & n317 ;
  assign n319 = n318 ^ n276 ;
  assign n320 = x69 & ~n276 ;
  assign n321 = n191 & ~n320 ;
  assign n322 = n320 ^ x69 ;
  assign n323 = n322 ^ n319 ;
  assign n324 = n310 ^ x67 ;
  assign n325 = n276 ^ x68 ;
  assign n328 = n317 & ~n325 ;
  assign n329 = n328 ^ x68 ;
  assign n330 = n192 & ~n329 ;
  assign n331 = n324 & n330 ;
  assign n332 = n331 ^ n312 ;
  assign n333 = n332 ^ x68 ;
  assign n360 = n307 ^ x66 ;
  assign n361 = n330 & n360 ;
  assign n362 = n361 ^ n294 ;
  assign n342 = x65 & n330 ;
  assign n338 = ~x59 & n330 ;
  assign n339 = n338 ^ n284 ;
  assign n340 = x64 & n339 ;
  assign n341 = n340 ^ x60 ;
  assign n343 = n342 ^ n341 ;
  assign n344 = n343 ^ x66 ;
  assign n352 = x59 & x65 ;
  assign n349 = x65 ^ x58 ;
  assign n345 = x64 ^ x59 ;
  assign n346 = n345 ^ x65 ;
  assign n350 = n346 ^ n330 ;
  assign n351 = ~n349 & n350 ;
  assign n353 = n352 ^ n351 ;
  assign n354 = x64 & n353 ;
  assign n355 = n354 ^ n352 ;
  assign n356 = n355 ^ x65 ;
  assign n357 = n356 ^ n343 ;
  assign n358 = ~n344 & n357 ;
  assign n359 = n358 ^ x66 ;
  assign n363 = n362 ^ n359 ;
  assign n364 = n362 ^ x67 ;
  assign n365 = n363 & ~n364 ;
  assign n366 = n365 ^ n316 ;
  assign n369 = ~n333 & n366 ;
  assign n370 = n369 ^ x68 ;
  assign n371 = ~n323 & n370 ;
  assign n372 = n321 & ~n371 ;
  assign n373 = n319 & ~n372 ;
  assign n376 = n375 ^ n373 ;
  assign n377 = ~n189 & n376 ;
  assign n384 = n376 ^ x70 ;
  assign n422 = n366 & n372 ;
  assign n423 = n422 ^ n332 ;
  assign n415 = n359 ^ x67 ;
  assign n416 = n372 & n415 ;
  assign n417 = n416 ^ n362 ;
  assign n408 = n356 ^ x66 ;
  assign n409 = n372 & n408 ;
  assign n410 = n409 ^ n343 ;
  assign n390 = x64 & n330 ;
  assign n386 = ~x58 & x64 ;
  assign n387 = n386 ^ x65 ;
  assign n388 = n372 & n387 ;
  assign n389 = n388 ^ x59 ;
  assign n391 = n390 ^ n389 ;
  assign n392 = n391 ^ x66 ;
  assign n394 = x65 ^ x57 ;
  assign n395 = x64 ^ x58 ;
  assign n396 = n395 ^ x65 ;
  assign n397 = n396 ^ n372 ;
  assign n398 = ~n394 & n397 ;
  assign n393 = x58 & x65 ;
  assign n399 = n398 ^ n393 ;
  assign n402 = x64 & n399 ;
  assign n403 = n402 ^ n393 ;
  assign n404 = n403 ^ x65 ;
  assign n405 = n404 ^ n391 ;
  assign n406 = ~n392 & n405 ;
  assign n407 = n406 ^ x66 ;
  assign n411 = n410 ^ n407 ;
  assign n412 = n410 ^ x67 ;
  assign n413 = n411 & ~n412 ;
  assign n414 = n413 ^ x67 ;
  assign n418 = n417 ^ n414 ;
  assign n419 = n417 ^ x68 ;
  assign n420 = n418 & ~n419 ;
  assign n421 = n420 ^ x68 ;
  assign n424 = n423 ^ n421 ;
  assign n425 = n423 ^ x69 ;
  assign n426 = n424 & ~n425 ;
  assign n427 = n426 ^ x69 ;
  assign n428 = n427 ^ x70 ;
  assign n429 = ~n384 & n428 ;
  assign n430 = n429 ^ x70 ;
  assign n431 = n190 & ~n430 ;
  assign n378 = n376 ^ x71 ;
  assign n480 = x70 & n427 ;
  assign n471 = n421 ^ x69 ;
  assign n472 = n431 & n471 ;
  assign n473 = n472 ^ n423 ;
  assign n464 = n414 ^ x68 ;
  assign n465 = n431 & n464 ;
  assign n466 = n465 ^ n417 ;
  assign n457 = n407 ^ x67 ;
  assign n458 = n431 & n457 ;
  assign n459 = n458 ^ n410 ;
  assign n450 = n404 ^ x66 ;
  assign n451 = n431 & n450 ;
  assign n452 = n451 ^ n391 ;
  assign n442 = x64 & n372 ;
  assign n441 = x65 & n431 ;
  assign n443 = n442 ^ n441 ;
  assign n444 = n443 ^ x58 ;
  assign n439 = x64 & n431 ;
  assign n440 = ~x57 & n439 ;
  assign n445 = n444 ^ n440 ;
  assign n434 = x57 & x65 ;
  assign n383 = x65 ^ x56 ;
  assign n379 = x64 ^ x57 ;
  assign n380 = n379 ^ x65 ;
  assign n432 = n431 ^ n380 ;
  assign n433 = ~n383 & n432 ;
  assign n435 = n434 ^ n433 ;
  assign n436 = x64 & n435 ;
  assign n437 = n436 ^ n434 ;
  assign n438 = n437 ^ x65 ;
  assign n446 = n445 ^ n438 ;
  assign n447 = n445 ^ x66 ;
  assign n448 = n446 & ~n447 ;
  assign n449 = n448 ^ x66 ;
  assign n453 = n452 ^ n449 ;
  assign n454 = n452 ^ x67 ;
  assign n455 = n453 & ~n454 ;
  assign n456 = n455 ^ x67 ;
  assign n460 = n459 ^ n456 ;
  assign n461 = n459 ^ x68 ;
  assign n462 = n460 & ~n461 ;
  assign n463 = n462 ^ x68 ;
  assign n467 = n466 ^ n463 ;
  assign n468 = n466 ^ x69 ;
  assign n469 = n467 & ~n468 ;
  assign n470 = n469 ^ x69 ;
  assign n474 = n473 ^ n470 ;
  assign n475 = n473 ^ x70 ;
  assign n476 = n474 & ~n475 ;
  assign n477 = n476 ^ x70 ;
  assign n481 = n480 ^ n477 ;
  assign n482 = n376 & ~n481 ;
  assign n483 = n482 ^ n477 ;
  assign n484 = n378 & ~n483 ;
  assign n485 = n484 ^ n477 ;
  assign n486 = n189 & ~n485 ;
  assign n487 = n376 & ~n486 ;
  assign n488 = ~n431 & n487 ;
  assign n489 = n488 ^ n375 ;
  assign n490 = n489 ^ x72 ;
  assign n491 = n188 & ~n490 ;
  assign n544 = n470 ^ x70 ;
  assign n545 = n486 & n544 ;
  assign n546 = n545 ^ n473 ;
  assign n537 = n463 ^ x69 ;
  assign n538 = n486 & n537 ;
  assign n539 = n538 ^ n466 ;
  assign n530 = n456 ^ x68 ;
  assign n531 = n486 & n530 ;
  assign n532 = n531 ^ n459 ;
  assign n523 = n449 ^ x67 ;
  assign n524 = n486 & n523 ;
  assign n525 = n524 ^ n452 ;
  assign n516 = n438 ^ x66 ;
  assign n517 = n486 & n516 ;
  assign n518 = n517 ^ n445 ;
  assign n510 = n439 ^ x57 ;
  assign n507 = ~x56 & x64 ;
  assign n508 = n507 ^ x65 ;
  assign n509 = n486 & n508 ;
  assign n511 = n510 ^ n509 ;
  assign n493 = x65 ^ x55 ;
  assign n494 = x64 ^ x56 ;
  assign n495 = n494 ^ x65 ;
  assign n496 = n495 ^ n486 ;
  assign n497 = ~n493 & n496 ;
  assign n492 = x56 & x65 ;
  assign n498 = n497 ^ n492 ;
  assign n501 = x64 & n498 ;
  assign n502 = n501 ^ n492 ;
  assign n503 = n502 ^ x65 ;
  assign n512 = n511 ^ n503 ;
  assign n513 = n511 ^ x66 ;
  assign n514 = n512 & ~n513 ;
  assign n515 = n514 ^ x66 ;
  assign n519 = n518 ^ n515 ;
  assign n520 = n518 ^ x67 ;
  assign n521 = n519 & ~n520 ;
  assign n522 = n521 ^ x67 ;
  assign n526 = n525 ^ n522 ;
  assign n527 = n525 ^ x68 ;
  assign n528 = n526 & ~n527 ;
  assign n529 = n528 ^ x68 ;
  assign n533 = n532 ^ n529 ;
  assign n534 = n532 ^ x69 ;
  assign n535 = n533 & ~n534 ;
  assign n536 = n535 ^ x69 ;
  assign n540 = n539 ^ n536 ;
  assign n541 = n539 ^ x70 ;
  assign n542 = n540 & ~n541 ;
  assign n543 = n542 ^ x70 ;
  assign n547 = n546 ^ n543 ;
  assign n548 = n546 ^ x71 ;
  assign n549 = n547 & ~n548 ;
  assign n550 = n549 ^ x71 ;
  assign n551 = n491 & ~n550 ;
  assign n552 = n377 & ~n551 ;
  assign n554 = n189 & n489 ;
  assign n555 = n554 ^ n551 ;
  assign n615 = n543 ^ x71 ;
  assign n616 = n555 & n615 ;
  assign n617 = n616 ^ n546 ;
  assign n553 = n536 ^ x70 ;
  assign n556 = n553 & n555 ;
  assign n557 = n556 ^ n539 ;
  assign n558 = n557 ^ x71 ;
  assign n559 = n529 ^ x69 ;
  assign n560 = n555 & n559 ;
  assign n561 = n560 ^ n532 ;
  assign n706 = n561 ^ x71 ;
  assign n707 = n706 ^ x70 ;
  assign n602 = n522 ^ x68 ;
  assign n603 = n555 & n602 ;
  assign n604 = n603 ^ n525 ;
  assign n595 = n515 ^ x67 ;
  assign n596 = n555 & n595 ;
  assign n597 = n596 ^ n518 ;
  assign n588 = n503 ^ x66 ;
  assign n589 = n555 & n588 ;
  assign n590 = n589 ^ n511 ;
  assign n568 = x65 & n555 ;
  assign n567 = x64 & n486 ;
  assign n569 = n568 ^ n567 ;
  assign n570 = n569 ^ x56 ;
  assign n565 = x64 & n555 ;
  assign n566 = ~x55 & n565 ;
  assign n571 = n570 ^ n566 ;
  assign n572 = n571 ^ x66 ;
  assign n580 = x55 & x65 ;
  assign n577 = x65 ^ x54 ;
  assign n573 = x64 ^ x55 ;
  assign n574 = n573 ^ x65 ;
  assign n578 = n574 ^ n555 ;
  assign n579 = ~n577 & n578 ;
  assign n581 = n580 ^ n579 ;
  assign n582 = x64 & n581 ;
  assign n583 = n582 ^ n580 ;
  assign n584 = n583 ^ x65 ;
  assign n585 = n584 ^ n571 ;
  assign n586 = ~n572 & n585 ;
  assign n587 = n586 ^ x66 ;
  assign n591 = n590 ^ n587 ;
  assign n592 = n590 ^ x67 ;
  assign n593 = n591 & ~n592 ;
  assign n594 = n593 ^ x67 ;
  assign n598 = n597 ^ n594 ;
  assign n599 = n597 ^ x68 ;
  assign n600 = n598 & ~n599 ;
  assign n601 = n600 ^ x68 ;
  assign n605 = n604 ^ n601 ;
  assign n606 = n604 ^ x69 ;
  assign n607 = n605 & ~n606 ;
  assign n608 = n607 ^ x69 ;
  assign n708 = n707 ^ n608 ;
  assign n709 = n708 ^ n706 ;
  assign n711 = x71 ^ x70 ;
  assign n712 = n711 ^ n706 ;
  assign n611 = n709 & ~n712 ;
  assign n563 = n557 ^ x70 ;
  assign n612 = n611 ^ n563 ;
  assign n613 = ~n558 & n612 ;
  assign n614 = n613 ^ x71 ;
  assign n618 = n617 ^ n614 ;
  assign n619 = x73 ^ x72 ;
  assign n620 = n619 ^ n552 ;
  assign n621 = n620 ^ n617 ;
  assign n622 = n618 & ~n621 ;
  assign n628 = n621 ^ x73 ;
  assign n629 = n628 ^ n618 ;
  assign n630 = n629 ^ n614 ;
  assign n631 = ~n619 & n630 ;
  assign n632 = n620 & n631 ;
  assign n633 = n632 ^ n630 ;
  assign n634 = n633 ^ n619 ;
  assign n635 = n622 & ~n634 ;
  assign n636 = n635 ^ n632 ;
  assign n637 = n636 ^ n631 ;
  assign n638 = n637 ^ n620 ;
  assign n639 = n187 & ~n638 ;
  assign n640 = n552 & ~n639 ;
  assign n641 = n640 ^ n375 ;
  assign n642 = n641 ^ x74 ;
  assign n647 = n641 ^ x73 ;
  assign n643 = n614 ^ x72 ;
  assign n644 = n639 & n643 ;
  assign n645 = n644 ^ n617 ;
  assign n646 = n645 ^ n641 ;
  assign n648 = n647 ^ n646 ;
  assign n713 = ~n709 & ~n712 ;
  assign n714 = n713 ^ n706 ;
  assign n715 = n639 & ~n714 ;
  assign n716 = n715 ^ n557 ;
  assign n700 = n639 & n709 ;
  assign n701 = n700 ^ n561 ;
  assign n692 = n601 ^ x69 ;
  assign n693 = n639 & n692 ;
  assign n694 = n693 ^ n604 ;
  assign n685 = n594 ^ x68 ;
  assign n686 = n639 & n685 ;
  assign n687 = n686 ^ n597 ;
  assign n678 = n587 ^ x67 ;
  assign n679 = n639 & n678 ;
  assign n680 = n679 ^ n590 ;
  assign n671 = n584 ^ x66 ;
  assign n672 = n639 & n671 ;
  assign n673 = n672 ^ n571 ;
  assign n656 = x54 & x65 ;
  assign n653 = x65 ^ x53 ;
  assign n649 = x64 ^ x54 ;
  assign n650 = n649 ^ x65 ;
  assign n654 = n650 ^ n639 ;
  assign n655 = ~n653 & n654 ;
  assign n657 = n656 ^ n655 ;
  assign n658 = x64 & n657 ;
  assign n659 = n658 ^ n656 ;
  assign n660 = n659 ^ x65 ;
  assign n661 = n660 ^ x66 ;
  assign n666 = n565 ^ x55 ;
  assign n663 = ~x54 & x64 ;
  assign n664 = n663 ^ x65 ;
  assign n665 = n639 & n664 ;
  assign n667 = n666 ^ n665 ;
  assign n668 = n667 ^ n660 ;
  assign n669 = n661 & n668 ;
  assign n670 = n669 ^ x66 ;
  assign n674 = n673 ^ n670 ;
  assign n675 = n673 ^ x67 ;
  assign n676 = n674 & ~n675 ;
  assign n677 = n676 ^ x67 ;
  assign n681 = n680 ^ n677 ;
  assign n682 = n680 ^ x68 ;
  assign n683 = n681 & ~n682 ;
  assign n684 = n683 ^ x68 ;
  assign n688 = n687 ^ n684 ;
  assign n689 = n687 ^ x69 ;
  assign n690 = n688 & ~n689 ;
  assign n691 = n690 ^ x69 ;
  assign n695 = n694 ^ n691 ;
  assign n696 = n694 ^ x70 ;
  assign n697 = n695 & ~n696 ;
  assign n698 = n697 ^ x70 ;
  assign n702 = n701 ^ n698 ;
  assign n703 = n701 ^ x71 ;
  assign n704 = n702 & ~n703 ;
  assign n705 = n704 ^ x71 ;
  assign n717 = n716 ^ n705 ;
  assign n718 = n716 ^ x72 ;
  assign n719 = n717 & ~n718 ;
  assign n720 = n719 ^ x72 ;
  assign n799 = n720 ^ x73 ;
  assign n723 = ~n648 & n799 ;
  assign n724 = n723 ^ n647 ;
  assign n725 = ~n642 & n724 ;
  assign n726 = n725 ^ x74 ;
  assign n727 = n186 & ~n726 ;
  assign n728 = n727 ^ n375 ;
  assign n729 = n641 & ~n728 ;
  assign n730 = n185 & n729 ;
  assign n731 = x75 & n730 ;
  assign n800 = n727 & n799 ;
  assign n801 = n800 ^ n645 ;
  assign n792 = n705 ^ x72 ;
  assign n793 = n727 & n792 ;
  assign n794 = n793 ^ n716 ;
  assign n785 = n698 ^ x71 ;
  assign n786 = n727 & n785 ;
  assign n787 = n786 ^ n701 ;
  assign n778 = n691 ^ x70 ;
  assign n779 = n727 & n778 ;
  assign n780 = n779 ^ n694 ;
  assign n771 = n684 ^ x69 ;
  assign n772 = n727 & n771 ;
  assign n773 = n772 ^ n687 ;
  assign n764 = n677 ^ x68 ;
  assign n765 = n727 & n764 ;
  assign n766 = n765 ^ n680 ;
  assign n757 = n670 ^ x67 ;
  assign n758 = n727 & n757 ;
  assign n759 = n758 ^ n673 ;
  assign n751 = n661 & n727 ;
  assign n752 = n751 ^ n667 ;
  assign n732 = ~x52 & x64 ;
  assign n736 = n732 ^ x53 ;
  assign n735 = x64 & n727 ;
  assign n737 = n736 ^ n735 ;
  assign n738 = x65 & ~n737 ;
  assign n733 = n727 ^ x53 ;
  assign n734 = n732 & ~n733 ;
  assign n739 = n738 ^ n734 ;
  assign n740 = n739 ^ x66 ;
  assign n746 = x64 & n639 ;
  assign n742 = ~x53 & x64 ;
  assign n743 = n742 ^ x65 ;
  assign n744 = n727 & n743 ;
  assign n745 = n744 ^ x54 ;
  assign n747 = n746 ^ n745 ;
  assign n748 = n747 ^ n739 ;
  assign n749 = n740 & n748 ;
  assign n750 = n749 ^ x66 ;
  assign n753 = n752 ^ n750 ;
  assign n754 = n752 ^ x67 ;
  assign n755 = n753 & ~n754 ;
  assign n756 = n755 ^ x67 ;
  assign n760 = n759 ^ n756 ;
  assign n761 = n759 ^ x68 ;
  assign n762 = n760 & ~n761 ;
  assign n763 = n762 ^ x68 ;
  assign n767 = n766 ^ n763 ;
  assign n768 = n766 ^ x69 ;
  assign n769 = n767 & ~n768 ;
  assign n770 = n769 ^ x69 ;
  assign n774 = n773 ^ n770 ;
  assign n775 = n773 ^ x70 ;
  assign n776 = n774 & ~n775 ;
  assign n777 = n776 ^ x70 ;
  assign n781 = n780 ^ n777 ;
  assign n782 = n780 ^ x71 ;
  assign n783 = n781 & ~n782 ;
  assign n784 = n783 ^ x71 ;
  assign n788 = n787 ^ n784 ;
  assign n789 = n787 ^ x72 ;
  assign n790 = n788 & ~n789 ;
  assign n791 = n790 ^ x72 ;
  assign n795 = n794 ^ n791 ;
  assign n796 = n794 ^ x73 ;
  assign n797 = n795 & ~n796 ;
  assign n798 = n797 ^ x73 ;
  assign n802 = n801 ^ n798 ;
  assign n803 = n801 ^ x74 ;
  assign n804 = n802 & ~n803 ;
  assign n805 = n804 ^ x74 ;
  assign n806 = n731 & n805 ;
  assign n807 = n806 ^ n730 ;
  assign n808 = n807 ^ n729 ;
  assign n812 = n729 ^ x75 ;
  assign n813 = n805 ^ x75 ;
  assign n814 = ~n812 & n813 ;
  assign n815 = n814 ^ x75 ;
  assign n816 = n185 & ~n815 ;
  assign n884 = n798 ^ x74 ;
  assign n885 = n816 & n884 ;
  assign n886 = n885 ^ n801 ;
  assign n877 = n791 ^ x73 ;
  assign n878 = n816 & n877 ;
  assign n879 = n878 ^ n794 ;
  assign n870 = n784 ^ x72 ;
  assign n871 = n816 & n870 ;
  assign n872 = n871 ^ n787 ;
  assign n863 = n777 ^ x71 ;
  assign n864 = n816 & n863 ;
  assign n865 = n864 ^ n780 ;
  assign n856 = n770 ^ x70 ;
  assign n857 = n816 & n856 ;
  assign n858 = n857 ^ n773 ;
  assign n849 = n763 ^ x69 ;
  assign n850 = n816 & n849 ;
  assign n851 = n850 ^ n766 ;
  assign n842 = n756 ^ x68 ;
  assign n843 = n816 & n842 ;
  assign n844 = n843 ^ n759 ;
  assign n835 = n750 ^ x67 ;
  assign n836 = n816 & n835 ;
  assign n837 = n836 ^ n752 ;
  assign n829 = n740 & n816 ;
  assign n830 = n829 ^ n747 ;
  assign n809 = ~x51 & x64 ;
  assign n810 = n809 ^ x65 ;
  assign n817 = x64 & n816 ;
  assign n811 = n809 ^ x52 ;
  assign n818 = n817 ^ n811 ;
  assign n819 = n810 & n818 ;
  assign n820 = n819 ^ x65 ;
  assign n821 = n820 ^ x66 ;
  assign n823 = n732 ^ x65 ;
  assign n824 = n816 & n823 ;
  assign n822 = n735 ^ x53 ;
  assign n825 = n824 ^ n822 ;
  assign n826 = n825 ^ n820 ;
  assign n827 = n821 & n826 ;
  assign n828 = n827 ^ x66 ;
  assign n831 = n830 ^ n828 ;
  assign n832 = n830 ^ x67 ;
  assign n833 = n831 & ~n832 ;
  assign n834 = n833 ^ x67 ;
  assign n838 = n837 ^ n834 ;
  assign n839 = n837 ^ x68 ;
  assign n840 = n838 & ~n839 ;
  assign n841 = n840 ^ x68 ;
  assign n845 = n844 ^ n841 ;
  assign n846 = n844 ^ x69 ;
  assign n847 = n845 & ~n846 ;
  assign n848 = n847 ^ x69 ;
  assign n852 = n851 ^ n848 ;
  assign n853 = n851 ^ x70 ;
  assign n854 = n852 & ~n853 ;
  assign n855 = n854 ^ x70 ;
  assign n859 = n858 ^ n855 ;
  assign n860 = n858 ^ x71 ;
  assign n861 = n859 & ~n860 ;
  assign n862 = n861 ^ x71 ;
  assign n866 = n865 ^ n862 ;
  assign n867 = n865 ^ x72 ;
  assign n868 = n866 & ~n867 ;
  assign n869 = n868 ^ x72 ;
  assign n873 = n872 ^ n869 ;
  assign n874 = n872 ^ x73 ;
  assign n875 = n873 & ~n874 ;
  assign n876 = n875 ^ x73 ;
  assign n880 = n879 ^ n876 ;
  assign n881 = n879 ^ x74 ;
  assign n882 = n880 & ~n881 ;
  assign n883 = n882 ^ x74 ;
  assign n887 = n886 ^ n883 ;
  assign n888 = x76 ^ x75 ;
  assign n889 = n888 ^ n808 ;
  assign n890 = n889 ^ n886 ;
  assign n891 = n887 & ~n890 ;
  assign n897 = n890 ^ x76 ;
  assign n898 = n897 ^ n887 ;
  assign n899 = n898 ^ n883 ;
  assign n900 = ~n888 & n899 ;
  assign n901 = n889 & n900 ;
  assign n902 = n901 ^ n899 ;
  assign n903 = n902 ^ n888 ;
  assign n904 = n891 & ~n903 ;
  assign n905 = n904 ^ n901 ;
  assign n906 = n905 ^ n900 ;
  assign n907 = n906 ^ n889 ;
  assign n908 = n184 & ~n907 ;
  assign n909 = n808 & ~n908 ;
  assign n910 = ~n183 & n909 ;
  assign n911 = n909 ^ n375 ;
  assign n912 = n911 ^ x77 ;
  assign n917 = n911 ^ x76 ;
  assign n913 = n883 ^ x75 ;
  assign n914 = n908 & n913 ;
  assign n915 = n914 ^ n886 ;
  assign n916 = n915 ^ n911 ;
  assign n918 = n917 ^ n916 ;
  assign n991 = n876 ^ x74 ;
  assign n992 = n908 & n991 ;
  assign n993 = n992 ^ n879 ;
  assign n984 = n869 ^ x73 ;
  assign n985 = n908 & n984 ;
  assign n986 = n985 ^ n872 ;
  assign n977 = n862 ^ x72 ;
  assign n978 = n908 & n977 ;
  assign n979 = n978 ^ n865 ;
  assign n970 = n855 ^ x71 ;
  assign n971 = n908 & n970 ;
  assign n972 = n971 ^ n858 ;
  assign n963 = n848 ^ x70 ;
  assign n964 = n908 & n963 ;
  assign n965 = n964 ^ n851 ;
  assign n956 = n841 ^ x69 ;
  assign n957 = n908 & n956 ;
  assign n958 = n957 ^ n844 ;
  assign n949 = n834 ^ x68 ;
  assign n950 = n908 & n949 ;
  assign n951 = n950 ^ n837 ;
  assign n942 = n828 ^ x67 ;
  assign n943 = n908 & n942 ;
  assign n944 = n943 ^ n830 ;
  assign n936 = n821 & n908 ;
  assign n937 = n936 ^ n825 ;
  assign n920 = n810 & n908 ;
  assign n919 = n817 ^ x52 ;
  assign n921 = n920 ^ n919 ;
  assign n922 = n921 ^ x66 ;
  assign n926 = ~x64 & x65 ;
  assign n925 = x64 & n908 ;
  assign n927 = n926 ^ n925 ;
  assign n923 = x64 ^ x51 ;
  assign n924 = n923 ^ x65 ;
  assign n928 = n927 ^ n924 ;
  assign n929 = ~x50 & x64 ;
  assign n930 = n929 ^ x65 ;
  assign n931 = n928 & n930 ;
  assign n932 = n931 ^ x65 ;
  assign n933 = n932 ^ n921 ;
  assign n934 = ~n922 & n933 ;
  assign n935 = n934 ^ x66 ;
  assign n938 = n937 ^ n935 ;
  assign n939 = n937 ^ x67 ;
  assign n940 = n938 & ~n939 ;
  assign n941 = n940 ^ x67 ;
  assign n945 = n944 ^ n941 ;
  assign n946 = n944 ^ x68 ;
  assign n947 = n945 & ~n946 ;
  assign n948 = n947 ^ x68 ;
  assign n952 = n951 ^ n948 ;
  assign n953 = n951 ^ x69 ;
  assign n954 = n952 & ~n953 ;
  assign n955 = n954 ^ x69 ;
  assign n959 = n958 ^ n955 ;
  assign n960 = n958 ^ x70 ;
  assign n961 = n959 & ~n960 ;
  assign n962 = n961 ^ x70 ;
  assign n966 = n965 ^ n962 ;
  assign n967 = n965 ^ x71 ;
  assign n968 = n966 & ~n967 ;
  assign n969 = n968 ^ x71 ;
  assign n973 = n972 ^ n969 ;
  assign n974 = n972 ^ x72 ;
  assign n975 = n973 & ~n974 ;
  assign n976 = n975 ^ x72 ;
  assign n980 = n979 ^ n976 ;
  assign n981 = n979 ^ x73 ;
  assign n982 = n980 & ~n981 ;
  assign n983 = n982 ^ x73 ;
  assign n987 = n986 ^ n983 ;
  assign n988 = n986 ^ x74 ;
  assign n989 = n987 & ~n988 ;
  assign n990 = n989 ^ x74 ;
  assign n994 = n993 ^ n990 ;
  assign n995 = n993 ^ x75 ;
  assign n996 = n994 & ~n995 ;
  assign n997 = n996 ^ x75 ;
  assign n1096 = n997 ^ x76 ;
  assign n1000 = ~n918 & n1096 ;
  assign n1001 = n1000 ^ n917 ;
  assign n1002 = ~n912 & n1001 ;
  assign n1003 = n1002 ^ x77 ;
  assign n1004 = n183 & ~n1003 ;
  assign n1005 = n909 & ~n1004 ;
  assign n1006 = n1005 ^ n375 ;
  assign n1007 = n1006 ^ x78 ;
  assign n1008 = n182 & ~n1007 ;
  assign n1097 = n1004 & n1096 ;
  assign n1098 = n1097 ^ n915 ;
  assign n1089 = n990 ^ x75 ;
  assign n1090 = n1004 & n1089 ;
  assign n1091 = n1090 ^ n993 ;
  assign n1082 = n983 ^ x74 ;
  assign n1083 = n1004 & n1082 ;
  assign n1084 = n1083 ^ n986 ;
  assign n1075 = n976 ^ x73 ;
  assign n1076 = n1004 & n1075 ;
  assign n1077 = n1076 ^ n979 ;
  assign n1068 = n969 ^ x72 ;
  assign n1069 = n1004 & n1068 ;
  assign n1070 = n1069 ^ n972 ;
  assign n1061 = n962 ^ x71 ;
  assign n1062 = n1004 & n1061 ;
  assign n1063 = n1062 ^ n965 ;
  assign n1054 = n955 ^ x70 ;
  assign n1055 = n1004 & n1054 ;
  assign n1056 = n1055 ^ n958 ;
  assign n1047 = n948 ^ x69 ;
  assign n1048 = n1004 & n1047 ;
  assign n1049 = n1048 ^ n951 ;
  assign n1040 = n941 ^ x68 ;
  assign n1041 = n1004 & n1040 ;
  assign n1042 = n1041 ^ n944 ;
  assign n1033 = n935 ^ x67 ;
  assign n1034 = n1004 & n1033 ;
  assign n1035 = n1034 ^ n937 ;
  assign n1026 = n932 ^ x66 ;
  assign n1027 = n1004 & n1026 ;
  assign n1028 = n1027 ^ n921 ;
  assign n1020 = n925 ^ x51 ;
  assign n1019 = n930 & n1004 ;
  assign n1021 = n1020 ^ n1019 ;
  assign n1009 = ~x49 & x64 ;
  assign n1010 = n1009 ^ n1004 ;
  assign n1011 = n1010 ^ x50 ;
  assign n1015 = n1009 ^ x65 ;
  assign n1016 = ~n1011 & ~n1015 ;
  assign n1014 = ~n926 & n1004 ;
  assign n1017 = n1016 ^ n1014 ;
  assign n1018 = n1017 ^ x50 ;
  assign n1022 = n1021 ^ n1018 ;
  assign n1023 = n1021 ^ x66 ;
  assign n1024 = ~n1022 & ~n1023 ;
  assign n1025 = n1024 ^ x66 ;
  assign n1029 = n1028 ^ n1025 ;
  assign n1030 = n1028 ^ x67 ;
  assign n1031 = n1029 & ~n1030 ;
  assign n1032 = n1031 ^ x67 ;
  assign n1036 = n1035 ^ n1032 ;
  assign n1037 = n1035 ^ x68 ;
  assign n1038 = n1036 & ~n1037 ;
  assign n1039 = n1038 ^ x68 ;
  assign n1043 = n1042 ^ n1039 ;
  assign n1044 = n1042 ^ x69 ;
  assign n1045 = n1043 & ~n1044 ;
  assign n1046 = n1045 ^ x69 ;
  assign n1050 = n1049 ^ n1046 ;
  assign n1051 = n1049 ^ x70 ;
  assign n1052 = n1050 & ~n1051 ;
  assign n1053 = n1052 ^ x70 ;
  assign n1057 = n1056 ^ n1053 ;
  assign n1058 = n1056 ^ x71 ;
  assign n1059 = n1057 & ~n1058 ;
  assign n1060 = n1059 ^ x71 ;
  assign n1064 = n1063 ^ n1060 ;
  assign n1065 = n1063 ^ x72 ;
  assign n1066 = n1064 & ~n1065 ;
  assign n1067 = n1066 ^ x72 ;
  assign n1071 = n1070 ^ n1067 ;
  assign n1072 = n1070 ^ x73 ;
  assign n1073 = n1071 & ~n1072 ;
  assign n1074 = n1073 ^ x73 ;
  assign n1078 = n1077 ^ n1074 ;
  assign n1079 = n1077 ^ x74 ;
  assign n1080 = n1078 & ~n1079 ;
  assign n1081 = n1080 ^ x74 ;
  assign n1085 = n1084 ^ n1081 ;
  assign n1086 = n1084 ^ x75 ;
  assign n1087 = n1085 & ~n1086 ;
  assign n1088 = n1087 ^ x75 ;
  assign n1092 = n1091 ^ n1088 ;
  assign n1093 = n1091 ^ x76 ;
  assign n1094 = n1092 & ~n1093 ;
  assign n1095 = n1094 ^ x76 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1100 = n1098 ^ x77 ;
  assign n1101 = n1099 & ~n1100 ;
  assign n1102 = n1101 ^ x77 ;
  assign n1103 = n1008 & ~n1102 ;
  assign n1104 = n910 & ~n1103 ;
  assign n1105 = n1104 ^ n375 ;
  assign n1106 = n1105 ^ x79 ;
  assign n1110 = n183 & n1006 ;
  assign n1111 = n1110 ^ n1103 ;
  assign n1201 = n1095 ^ x77 ;
  assign n1202 = n1111 & n1201 ;
  assign n1203 = n1202 ^ n1098 ;
  assign n1194 = n1088 ^ x76 ;
  assign n1195 = n1111 & n1194 ;
  assign n1196 = n1195 ^ n1091 ;
  assign n1187 = n1081 ^ x75 ;
  assign n1188 = n1111 & n1187 ;
  assign n1189 = n1188 ^ n1084 ;
  assign n1180 = n1074 ^ x74 ;
  assign n1181 = n1111 & n1180 ;
  assign n1182 = n1181 ^ n1077 ;
  assign n1173 = n1067 ^ x73 ;
  assign n1174 = n1111 & n1173 ;
  assign n1175 = n1174 ^ n1070 ;
  assign n1166 = n1060 ^ x72 ;
  assign n1167 = n1111 & n1166 ;
  assign n1168 = n1167 ^ n1063 ;
  assign n1159 = n1053 ^ x71 ;
  assign n1160 = n1111 & n1159 ;
  assign n1161 = n1160 ^ n1056 ;
  assign n1152 = n1046 ^ x70 ;
  assign n1153 = n1111 & n1152 ;
  assign n1154 = n1153 ^ n1049 ;
  assign n1145 = n1039 ^ x69 ;
  assign n1146 = n1111 & n1145 ;
  assign n1147 = n1146 ^ n1042 ;
  assign n1138 = n1032 ^ x68 ;
  assign n1139 = n1111 & n1138 ;
  assign n1140 = n1139 ^ n1035 ;
  assign n1131 = n1025 ^ x67 ;
  assign n1132 = n1111 & n1131 ;
  assign n1133 = n1132 ^ n1028 ;
  assign n1124 = n1018 ^ x66 ;
  assign n1125 = n1111 & ~n1124 ;
  assign n1126 = n1125 ^ n1021 ;
  assign n1117 = x64 & n1004 ;
  assign n1116 = n1015 & n1111 ;
  assign n1118 = n1117 ^ n1116 ;
  assign n1119 = n1118 ^ x50 ;
  assign n1107 = ~x48 & x64 ;
  assign n1108 = n1107 ^ x65 ;
  assign n1112 = x64 & n1111 ;
  assign n1109 = n1107 ^ x49 ;
  assign n1113 = n1112 ^ n1109 ;
  assign n1114 = n1108 & n1113 ;
  assign n1115 = n1114 ^ x65 ;
  assign n1120 = n1119 ^ n1115 ;
  assign n1121 = n1119 ^ x66 ;
  assign n1122 = n1120 & ~n1121 ;
  assign n1123 = n1122 ^ x66 ;
  assign n1127 = n1126 ^ n1123 ;
  assign n1128 = n1126 ^ x67 ;
  assign n1129 = n1127 & ~n1128 ;
  assign n1130 = n1129 ^ x67 ;
  assign n1134 = n1133 ^ n1130 ;
  assign n1135 = n1133 ^ x68 ;
  assign n1136 = n1134 & ~n1135 ;
  assign n1137 = n1136 ^ x68 ;
  assign n1141 = n1140 ^ n1137 ;
  assign n1142 = n1140 ^ x69 ;
  assign n1143 = n1141 & ~n1142 ;
  assign n1144 = n1143 ^ x69 ;
  assign n1148 = n1147 ^ n1144 ;
  assign n1149 = n1147 ^ x70 ;
  assign n1150 = n1148 & ~n1149 ;
  assign n1151 = n1150 ^ x70 ;
  assign n1155 = n1154 ^ n1151 ;
  assign n1156 = n1154 ^ x71 ;
  assign n1157 = n1155 & ~n1156 ;
  assign n1158 = n1157 ^ x71 ;
  assign n1162 = n1161 ^ n1158 ;
  assign n1163 = n1161 ^ x72 ;
  assign n1164 = n1162 & ~n1163 ;
  assign n1165 = n1164 ^ x72 ;
  assign n1169 = n1168 ^ n1165 ;
  assign n1170 = n1168 ^ x73 ;
  assign n1171 = n1169 & ~n1170 ;
  assign n1172 = n1171 ^ x73 ;
  assign n1176 = n1175 ^ n1172 ;
  assign n1177 = n1175 ^ x74 ;
  assign n1178 = n1176 & ~n1177 ;
  assign n1179 = n1178 ^ x74 ;
  assign n1183 = n1182 ^ n1179 ;
  assign n1184 = n1182 ^ x75 ;
  assign n1185 = n1183 & ~n1184 ;
  assign n1186 = n1185 ^ x75 ;
  assign n1190 = n1189 ^ n1186 ;
  assign n1191 = n1189 ^ x76 ;
  assign n1192 = n1190 & ~n1191 ;
  assign n1193 = n1192 ^ x76 ;
  assign n1197 = n1196 ^ n1193 ;
  assign n1198 = n1196 ^ x77 ;
  assign n1199 = n1197 & ~n1198 ;
  assign n1200 = n1199 ^ x77 ;
  assign n1204 = n1203 ^ n1200 ;
  assign n1216 = n1200 ^ x78 ;
  assign n1208 = n1204 & n1216 ;
  assign n1205 = x79 ^ x78 ;
  assign n1209 = n1208 ^ n1205 ;
  assign n1210 = ~n1106 & n1209 ;
  assign n1211 = n1210 ^ x79 ;
  assign n1212 = n181 & ~n1211 ;
  assign n1213 = n1104 & ~n1212 ;
  assign n1214 = n1213 ^ n375 ;
  assign n1215 = n1214 ^ x80 ;
  assign n1220 = n1214 ^ x79 ;
  assign n1217 = n1212 & n1216 ;
  assign n1218 = n1217 ^ n1203 ;
  assign n1219 = n1218 ^ n1214 ;
  assign n1221 = n1220 ^ n1219 ;
  assign n1314 = n1193 ^ x77 ;
  assign n1315 = n1212 & n1314 ;
  assign n1316 = n1315 ^ n1196 ;
  assign n1307 = n1186 ^ x76 ;
  assign n1308 = n1212 & n1307 ;
  assign n1309 = n1308 ^ n1189 ;
  assign n1300 = n1179 ^ x75 ;
  assign n1301 = n1212 & n1300 ;
  assign n1302 = n1301 ^ n1182 ;
  assign n1293 = n1172 ^ x74 ;
  assign n1294 = n1212 & n1293 ;
  assign n1295 = n1294 ^ n1175 ;
  assign n1286 = n1165 ^ x73 ;
  assign n1287 = n1212 & n1286 ;
  assign n1288 = n1287 ^ n1168 ;
  assign n1279 = n1158 ^ x72 ;
  assign n1280 = n1212 & n1279 ;
  assign n1281 = n1280 ^ n1161 ;
  assign n1272 = n1151 ^ x71 ;
  assign n1273 = n1212 & n1272 ;
  assign n1274 = n1273 ^ n1154 ;
  assign n1265 = n1144 ^ x70 ;
  assign n1266 = n1212 & n1265 ;
  assign n1267 = n1266 ^ n1147 ;
  assign n1258 = n1137 ^ x69 ;
  assign n1259 = n1212 & n1258 ;
  assign n1260 = n1259 ^ n1140 ;
  assign n1251 = n1130 ^ x68 ;
  assign n1252 = n1212 & n1251 ;
  assign n1253 = n1252 ^ n1133 ;
  assign n1244 = n1123 ^ x67 ;
  assign n1245 = n1212 & n1244 ;
  assign n1246 = n1245 ^ n1126 ;
  assign n1222 = n1115 ^ x66 ;
  assign n1223 = n1212 & n1222 ;
  assign n1224 = n1223 ^ n1119 ;
  assign n1225 = n1224 ^ x67 ;
  assign n1226 = x64 & n1212 ;
  assign n1231 = n1226 ^ x48 ;
  assign n1232 = x65 & ~n1231 ;
  assign n1228 = x64 & x65 ;
  assign n1227 = n1226 ^ n1107 ;
  assign n1229 = n1228 ^ n1227 ;
  assign n1230 = ~x47 & n1229 ;
  assign n1233 = n1232 ^ n1230 ;
  assign n1234 = n1233 ^ x66 ;
  assign n1236 = n1112 ^ x49 ;
  assign n1235 = n1108 & n1212 ;
  assign n1237 = n1236 ^ n1235 ;
  assign n1238 = n1237 ^ n1233 ;
  assign n1239 = n1234 & n1238 ;
  assign n1240 = n1239 ^ x66 ;
  assign n1241 = n1240 ^ n1224 ;
  assign n1242 = ~n1225 & n1241 ;
  assign n1243 = n1242 ^ x67 ;
  assign n1247 = n1246 ^ n1243 ;
  assign n1248 = n1246 ^ x68 ;
  assign n1249 = n1247 & ~n1248 ;
  assign n1250 = n1249 ^ x68 ;
  assign n1254 = n1253 ^ n1250 ;
  assign n1255 = n1253 ^ x69 ;
  assign n1256 = n1254 & ~n1255 ;
  assign n1257 = n1256 ^ x69 ;
  assign n1261 = n1260 ^ n1257 ;
  assign n1262 = n1260 ^ x70 ;
  assign n1263 = n1261 & ~n1262 ;
  assign n1264 = n1263 ^ x70 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1269 = n1267 ^ x71 ;
  assign n1270 = n1268 & ~n1269 ;
  assign n1271 = n1270 ^ x71 ;
  assign n1275 = n1274 ^ n1271 ;
  assign n1276 = n1274 ^ x72 ;
  assign n1277 = n1275 & ~n1276 ;
  assign n1278 = n1277 ^ x72 ;
  assign n1282 = n1281 ^ n1278 ;
  assign n1283 = n1281 ^ x73 ;
  assign n1284 = n1282 & ~n1283 ;
  assign n1285 = n1284 ^ x73 ;
  assign n1289 = n1288 ^ n1285 ;
  assign n1290 = n1288 ^ x74 ;
  assign n1291 = n1289 & ~n1290 ;
  assign n1292 = n1291 ^ x74 ;
  assign n1296 = n1295 ^ n1292 ;
  assign n1297 = n1295 ^ x75 ;
  assign n1298 = n1296 & ~n1297 ;
  assign n1299 = n1298 ^ x75 ;
  assign n1303 = n1302 ^ n1299 ;
  assign n1304 = n1302 ^ x76 ;
  assign n1305 = n1303 & ~n1304 ;
  assign n1306 = n1305 ^ x76 ;
  assign n1310 = n1309 ^ n1306 ;
  assign n1311 = n1309 ^ x77 ;
  assign n1312 = n1310 & ~n1311 ;
  assign n1313 = n1312 ^ x77 ;
  assign n1317 = n1316 ^ n1313 ;
  assign n1318 = n1316 ^ x78 ;
  assign n1319 = n1317 & ~n1318 ;
  assign n1320 = n1319 ^ x78 ;
  assign n1321 = n1320 ^ n1214 ;
  assign n1322 = n1321 ^ n1220 ;
  assign n1323 = ~n1221 & n1322 ;
  assign n1324 = n1323 ^ n1220 ;
  assign n1325 = ~n1215 & n1324 ;
  assign n1326 = n1325 ^ x80 ;
  assign n1327 = n180 & ~n1326 ;
  assign n1328 = n1327 ^ n375 ;
  assign n1329 = n1214 & ~n1328 ;
  assign n1330 = n1329 ^ x81 ;
  assign n1331 = n179 & ~n1330 ;
  assign n1442 = n1320 ^ x79 ;
  assign n1443 = n1327 & n1442 ;
  assign n1444 = n1443 ^ n1218 ;
  assign n1435 = n1313 ^ x78 ;
  assign n1436 = n1327 & n1435 ;
  assign n1437 = n1436 ^ n1316 ;
  assign n1428 = n1306 ^ x77 ;
  assign n1429 = n1327 & n1428 ;
  assign n1430 = n1429 ^ n1309 ;
  assign n1421 = n1299 ^ x76 ;
  assign n1422 = n1327 & n1421 ;
  assign n1423 = n1422 ^ n1302 ;
  assign n1414 = n1292 ^ x75 ;
  assign n1415 = n1327 & n1414 ;
  assign n1416 = n1415 ^ n1295 ;
  assign n1407 = n1285 ^ x74 ;
  assign n1408 = n1327 & n1407 ;
  assign n1409 = n1408 ^ n1288 ;
  assign n1400 = n1278 ^ x73 ;
  assign n1401 = n1327 & n1400 ;
  assign n1402 = n1401 ^ n1281 ;
  assign n1393 = n1271 ^ x72 ;
  assign n1394 = n1327 & n1393 ;
  assign n1395 = n1394 ^ n1274 ;
  assign n1386 = n1264 ^ x71 ;
  assign n1387 = n1327 & n1386 ;
  assign n1388 = n1387 ^ n1267 ;
  assign n1379 = n1257 ^ x70 ;
  assign n1380 = n1327 & n1379 ;
  assign n1381 = n1380 ^ n1260 ;
  assign n1372 = n1250 ^ x69 ;
  assign n1373 = n1327 & n1372 ;
  assign n1374 = n1373 ^ n1253 ;
  assign n1365 = n1243 ^ x68 ;
  assign n1366 = n1327 & n1365 ;
  assign n1367 = n1366 ^ n1246 ;
  assign n1358 = n1240 ^ x67 ;
  assign n1359 = n1327 & n1358 ;
  assign n1360 = n1359 ^ n1224 ;
  assign n1352 = n1234 & n1327 ;
  assign n1353 = n1352 ^ n1237 ;
  assign n1340 = x65 ^ x46 ;
  assign n1344 = x64 & n1327 ;
  assign n1345 = ~n1340 & ~n1344 ;
  assign n1338 = ~x46 & x64 ;
  assign n1339 = n1338 ^ x65 ;
  assign n1342 = x65 ^ x47 ;
  assign n1343 = n1339 & ~n1342 ;
  assign n1346 = n1345 ^ n1343 ;
  assign n1347 = n1346 ^ x46 ;
  assign n1334 = ~x47 & x64 ;
  assign n1335 = n1334 ^ x65 ;
  assign n1336 = n1327 & n1335 ;
  assign n1337 = n1336 ^ n1231 ;
  assign n1348 = n1347 ^ n1337 ;
  assign n1349 = n1347 ^ x66 ;
  assign n1350 = ~n1348 & ~n1349 ;
  assign n1351 = n1350 ^ x66 ;
  assign n1354 = n1353 ^ n1351 ;
  assign n1355 = n1353 ^ x67 ;
  assign n1356 = n1354 & ~n1355 ;
  assign n1357 = n1356 ^ x67 ;
  assign n1361 = n1360 ^ n1357 ;
  assign n1362 = n1360 ^ x68 ;
  assign n1363 = n1361 & ~n1362 ;
  assign n1364 = n1363 ^ x68 ;
  assign n1368 = n1367 ^ n1364 ;
  assign n1369 = n1367 ^ x69 ;
  assign n1370 = n1368 & ~n1369 ;
  assign n1371 = n1370 ^ x69 ;
  assign n1375 = n1374 ^ n1371 ;
  assign n1376 = n1374 ^ x70 ;
  assign n1377 = n1375 & ~n1376 ;
  assign n1378 = n1377 ^ x70 ;
  assign n1382 = n1381 ^ n1378 ;
  assign n1383 = n1381 ^ x71 ;
  assign n1384 = n1382 & ~n1383 ;
  assign n1385 = n1384 ^ x71 ;
  assign n1389 = n1388 ^ n1385 ;
  assign n1390 = n1388 ^ x72 ;
  assign n1391 = n1389 & ~n1390 ;
  assign n1392 = n1391 ^ x72 ;
  assign n1396 = n1395 ^ n1392 ;
  assign n1397 = n1395 ^ x73 ;
  assign n1398 = n1396 & ~n1397 ;
  assign n1399 = n1398 ^ x73 ;
  assign n1403 = n1402 ^ n1399 ;
  assign n1404 = n1402 ^ x74 ;
  assign n1405 = n1403 & ~n1404 ;
  assign n1406 = n1405 ^ x74 ;
  assign n1410 = n1409 ^ n1406 ;
  assign n1411 = n1409 ^ x75 ;
  assign n1412 = n1410 & ~n1411 ;
  assign n1413 = n1412 ^ x75 ;
  assign n1417 = n1416 ^ n1413 ;
  assign n1418 = n1416 ^ x76 ;
  assign n1419 = n1417 & ~n1418 ;
  assign n1420 = n1419 ^ x76 ;
  assign n1424 = n1423 ^ n1420 ;
  assign n1425 = n1423 ^ x77 ;
  assign n1426 = n1424 & ~n1425 ;
  assign n1427 = n1426 ^ x77 ;
  assign n1431 = n1430 ^ n1427 ;
  assign n1432 = n1430 ^ x78 ;
  assign n1433 = n1431 & ~n1432 ;
  assign n1434 = n1433 ^ x78 ;
  assign n1438 = n1437 ^ n1434 ;
  assign n1439 = n1437 ^ x79 ;
  assign n1440 = n1438 & ~n1439 ;
  assign n1441 = n1440 ^ x79 ;
  assign n1445 = n1444 ^ n1441 ;
  assign n1446 = n1444 ^ x80 ;
  assign n1447 = n1445 & ~n1446 ;
  assign n1448 = n1447 ^ x80 ;
  assign n1449 = n1331 & ~n1448 ;
  assign n1450 = ~n180 & n1213 ;
  assign n1451 = ~n1449 & n1450 ;
  assign n1452 = n1451 ^ n375 ;
  assign n1453 = n1452 ^ x82 ;
  assign n1460 = n1452 ^ x81 ;
  assign n1454 = n1441 ^ x80 ;
  assign n1455 = n180 & n1329 ;
  assign n1456 = n1455 ^ n1449 ;
  assign n1457 = n1454 & n1456 ;
  assign n1458 = n1457 ^ n1444 ;
  assign n1459 = n1458 ^ n1452 ;
  assign n1461 = n1460 ^ n1459 ;
  assign n1568 = n1434 ^ x79 ;
  assign n1569 = n1456 & n1568 ;
  assign n1570 = n1569 ^ n1437 ;
  assign n1561 = n1427 ^ x78 ;
  assign n1562 = n1456 & n1561 ;
  assign n1563 = n1562 ^ n1430 ;
  assign n1554 = n1420 ^ x77 ;
  assign n1555 = n1456 & n1554 ;
  assign n1556 = n1555 ^ n1423 ;
  assign n1547 = n1413 ^ x76 ;
  assign n1548 = n1456 & n1547 ;
  assign n1549 = n1548 ^ n1416 ;
  assign n1540 = n1406 ^ x75 ;
  assign n1541 = n1456 & n1540 ;
  assign n1542 = n1541 ^ n1409 ;
  assign n1533 = n1399 ^ x74 ;
  assign n1534 = n1456 & n1533 ;
  assign n1535 = n1534 ^ n1402 ;
  assign n1526 = n1392 ^ x73 ;
  assign n1527 = n1456 & n1526 ;
  assign n1528 = n1527 ^ n1395 ;
  assign n1519 = n1385 ^ x72 ;
  assign n1520 = n1456 & n1519 ;
  assign n1521 = n1520 ^ n1388 ;
  assign n1512 = n1378 ^ x71 ;
  assign n1513 = n1456 & n1512 ;
  assign n1514 = n1513 ^ n1381 ;
  assign n1505 = n1371 ^ x70 ;
  assign n1506 = n1456 & n1505 ;
  assign n1507 = n1506 ^ n1374 ;
  assign n1498 = n1364 ^ x69 ;
  assign n1499 = n1456 & n1498 ;
  assign n1500 = n1499 ^ n1367 ;
  assign n1462 = n1357 ^ x68 ;
  assign n1463 = n1456 & n1462 ;
  assign n1464 = n1463 ^ n1360 ;
  assign n1465 = n1464 ^ x69 ;
  assign n1470 = n1464 ^ x68 ;
  assign n1466 = n1351 ^ x67 ;
  assign n1467 = n1456 & n1466 ;
  assign n1468 = n1467 ^ n1353 ;
  assign n1469 = n1468 ^ n1464 ;
  assign n1471 = n1470 ^ n1469 ;
  assign n1477 = ~x45 & x64 ;
  assign n1478 = n1477 ^ x65 ;
  assign n1479 = x64 & n1456 ;
  assign n1480 = n1479 ^ x46 ;
  assign n1481 = n1480 ^ n1477 ;
  assign n1482 = n1478 & n1481 ;
  assign n1483 = n1482 ^ x65 ;
  assign n1475 = n1339 & n1456 ;
  assign n1474 = n1344 ^ x47 ;
  assign n1476 = n1475 ^ n1474 ;
  assign n1484 = n1483 ^ n1476 ;
  assign n1485 = n1483 ^ x66 ;
  assign n1486 = n1484 & n1485 ;
  assign n1487 = n1486 ^ x66 ;
  assign n1472 = ~n1349 & n1456 ;
  assign n1473 = n1472 ^ n1337 ;
  assign n1488 = n1487 ^ n1473 ;
  assign n1489 = n1487 ^ x67 ;
  assign n1490 = n1488 & n1489 ;
  assign n1491 = n1490 ^ x67 ;
  assign n1492 = n1491 ^ n1464 ;
  assign n1493 = n1492 ^ n1470 ;
  assign n1494 = ~n1471 & n1493 ;
  assign n1495 = n1494 ^ n1470 ;
  assign n1496 = ~n1465 & n1495 ;
  assign n1497 = n1496 ^ x69 ;
  assign n1501 = n1500 ^ n1497 ;
  assign n1502 = n1500 ^ x70 ;
  assign n1503 = n1501 & ~n1502 ;
  assign n1504 = n1503 ^ x70 ;
  assign n1508 = n1507 ^ n1504 ;
  assign n1509 = n1507 ^ x71 ;
  assign n1510 = n1508 & ~n1509 ;
  assign n1511 = n1510 ^ x71 ;
  assign n1515 = n1514 ^ n1511 ;
  assign n1516 = n1514 ^ x72 ;
  assign n1517 = n1515 & ~n1516 ;
  assign n1518 = n1517 ^ x72 ;
  assign n1522 = n1521 ^ n1518 ;
  assign n1523 = n1521 ^ x73 ;
  assign n1524 = n1522 & ~n1523 ;
  assign n1525 = n1524 ^ x73 ;
  assign n1529 = n1528 ^ n1525 ;
  assign n1530 = n1528 ^ x74 ;
  assign n1531 = n1529 & ~n1530 ;
  assign n1532 = n1531 ^ x74 ;
  assign n1536 = n1535 ^ n1532 ;
  assign n1537 = n1535 ^ x75 ;
  assign n1538 = n1536 & ~n1537 ;
  assign n1539 = n1538 ^ x75 ;
  assign n1543 = n1542 ^ n1539 ;
  assign n1544 = n1542 ^ x76 ;
  assign n1545 = n1543 & ~n1544 ;
  assign n1546 = n1545 ^ x76 ;
  assign n1550 = n1549 ^ n1546 ;
  assign n1551 = n1549 ^ x77 ;
  assign n1552 = n1550 & ~n1551 ;
  assign n1553 = n1552 ^ x77 ;
  assign n1557 = n1556 ^ n1553 ;
  assign n1558 = n1556 ^ x78 ;
  assign n1559 = n1557 & ~n1558 ;
  assign n1560 = n1559 ^ x78 ;
  assign n1564 = n1563 ^ n1560 ;
  assign n1565 = n1563 ^ x79 ;
  assign n1566 = n1564 & ~n1565 ;
  assign n1567 = n1566 ^ x79 ;
  assign n1571 = n1570 ^ n1567 ;
  assign n1572 = n1570 ^ x80 ;
  assign n1573 = n1571 & ~n1572 ;
  assign n1574 = n1573 ^ x80 ;
  assign n1575 = n1574 ^ n1452 ;
  assign n1576 = n1575 ^ n1460 ;
  assign n1577 = ~n1461 & n1576 ;
  assign n1578 = n1577 ^ n1460 ;
  assign n1579 = ~n1453 & n1578 ;
  assign n1580 = n1579 ^ x82 ;
  assign n1581 = n178 & ~n1580 ;
  assign n1582 = n1451 & ~n1581 ;
  assign n1583 = n1582 ^ n375 ;
  assign n1584 = n1583 ^ x83 ;
  assign n1589 = n1583 ^ x82 ;
  assign n1585 = n1574 ^ x81 ;
  assign n1586 = n1581 & n1585 ;
  assign n1587 = n1586 ^ n1458 ;
  assign n1588 = n1587 ^ n1583 ;
  assign n1590 = n1589 ^ n1588 ;
  assign n1713 = n1567 ^ x80 ;
  assign n1714 = n1581 & n1713 ;
  assign n1715 = n1714 ^ n1570 ;
  assign n1706 = n1560 ^ x79 ;
  assign n1707 = n1581 & n1706 ;
  assign n1708 = n1707 ^ n1563 ;
  assign n1699 = n1553 ^ x78 ;
  assign n1700 = n1581 & n1699 ;
  assign n1701 = n1700 ^ n1556 ;
  assign n1692 = n1546 ^ x77 ;
  assign n1693 = n1581 & n1692 ;
  assign n1694 = n1693 ^ n1549 ;
  assign n1685 = n1539 ^ x76 ;
  assign n1686 = n1581 & n1685 ;
  assign n1687 = n1686 ^ n1542 ;
  assign n1678 = n1532 ^ x75 ;
  assign n1679 = n1581 & n1678 ;
  assign n1680 = n1679 ^ n1535 ;
  assign n1671 = n1525 ^ x74 ;
  assign n1672 = n1581 & n1671 ;
  assign n1673 = n1672 ^ n1528 ;
  assign n1664 = n1518 ^ x73 ;
  assign n1665 = n1581 & n1664 ;
  assign n1666 = n1665 ^ n1521 ;
  assign n1657 = n1511 ^ x72 ;
  assign n1658 = n1581 & n1657 ;
  assign n1659 = n1658 ^ n1514 ;
  assign n1650 = n1504 ^ x71 ;
  assign n1651 = n1581 & n1650 ;
  assign n1652 = n1651 ^ n1507 ;
  assign n1643 = n1497 ^ x70 ;
  assign n1644 = n1581 & n1643 ;
  assign n1645 = n1644 ^ n1500 ;
  assign n1628 = n1468 ^ x69 ;
  assign n1629 = n1628 ^ n1491 ;
  assign n1630 = n1629 ^ x68 ;
  assign n1631 = n1630 ^ n1628 ;
  assign n1633 = n1491 ^ x69 ;
  assign n1634 = n1633 ^ n1628 ;
  assign n1635 = ~n1631 & ~n1634 ;
  assign n1636 = n1635 ^ n1628 ;
  assign n1637 = n1581 & ~n1636 ;
  assign n1638 = n1637 ^ n1464 ;
  assign n1621 = n1491 ^ x68 ;
  assign n1622 = n1581 & n1621 ;
  assign n1623 = n1622 ^ n1468 ;
  assign n1615 = n1489 & n1581 ;
  assign n1616 = n1615 ^ n1473 ;
  assign n1609 = n1485 & n1581 ;
  assign n1610 = n1609 ^ n1476 ;
  assign n1591 = n1478 & n1581 ;
  assign n1592 = n1591 ^ n1480 ;
  assign n1593 = n1592 ^ x66 ;
  assign n1595 = x65 ^ x44 ;
  assign n1596 = x64 ^ x45 ;
  assign n1597 = n1596 ^ x65 ;
  assign n1598 = n1597 ^ n1581 ;
  assign n1599 = ~n1595 & n1598 ;
  assign n1594 = x45 & x65 ;
  assign n1600 = n1599 ^ n1594 ;
  assign n1603 = x64 & n1600 ;
  assign n1604 = n1603 ^ n1594 ;
  assign n1605 = n1604 ^ x65 ;
  assign n1606 = n1605 ^ n1592 ;
  assign n1607 = ~n1593 & n1606 ;
  assign n1608 = n1607 ^ x66 ;
  assign n1611 = n1610 ^ n1608 ;
  assign n1612 = n1610 ^ x67 ;
  assign n1613 = n1611 & ~n1612 ;
  assign n1614 = n1613 ^ x67 ;
  assign n1617 = n1616 ^ n1614 ;
  assign n1618 = n1616 ^ x68 ;
  assign n1619 = n1617 & ~n1618 ;
  assign n1620 = n1619 ^ x68 ;
  assign n1624 = n1623 ^ n1620 ;
  assign n1625 = n1623 ^ x69 ;
  assign n1626 = n1624 & ~n1625 ;
  assign n1627 = n1626 ^ x69 ;
  assign n1639 = n1638 ^ n1627 ;
  assign n1640 = n1638 ^ x70 ;
  assign n1641 = n1639 & ~n1640 ;
  assign n1642 = n1641 ^ x70 ;
  assign n1646 = n1645 ^ n1642 ;
  assign n1647 = n1645 ^ x71 ;
  assign n1648 = n1646 & ~n1647 ;
  assign n1649 = n1648 ^ x71 ;
  assign n1653 = n1652 ^ n1649 ;
  assign n1654 = n1652 ^ x72 ;
  assign n1655 = n1653 & ~n1654 ;
  assign n1656 = n1655 ^ x72 ;
  assign n1660 = n1659 ^ n1656 ;
  assign n1661 = n1659 ^ x73 ;
  assign n1662 = n1660 & ~n1661 ;
  assign n1663 = n1662 ^ x73 ;
  assign n1667 = n1666 ^ n1663 ;
  assign n1668 = n1666 ^ x74 ;
  assign n1669 = n1667 & ~n1668 ;
  assign n1670 = n1669 ^ x74 ;
  assign n1674 = n1673 ^ n1670 ;
  assign n1675 = n1673 ^ x75 ;
  assign n1676 = n1674 & ~n1675 ;
  assign n1677 = n1676 ^ x75 ;
  assign n1681 = n1680 ^ n1677 ;
  assign n1682 = n1680 ^ x76 ;
  assign n1683 = n1681 & ~n1682 ;
  assign n1684 = n1683 ^ x76 ;
  assign n1688 = n1687 ^ n1684 ;
  assign n1689 = n1687 ^ x77 ;
  assign n1690 = n1688 & ~n1689 ;
  assign n1691 = n1690 ^ x77 ;
  assign n1695 = n1694 ^ n1691 ;
  assign n1696 = n1694 ^ x78 ;
  assign n1697 = n1695 & ~n1696 ;
  assign n1698 = n1697 ^ x78 ;
  assign n1702 = n1701 ^ n1698 ;
  assign n1703 = n1701 ^ x79 ;
  assign n1704 = n1702 & ~n1703 ;
  assign n1705 = n1704 ^ x79 ;
  assign n1709 = n1708 ^ n1705 ;
  assign n1710 = n1708 ^ x80 ;
  assign n1711 = n1709 & ~n1710 ;
  assign n1712 = n1711 ^ x80 ;
  assign n1716 = n1715 ^ n1712 ;
  assign n1717 = n1715 ^ x81 ;
  assign n1718 = n1716 & ~n1717 ;
  assign n1719 = n1718 ^ x81 ;
  assign n1720 = n1719 ^ n1583 ;
  assign n1721 = n1720 ^ n1589 ;
  assign n1722 = ~n1590 & n1721 ;
  assign n1723 = n1722 ^ n1589 ;
  assign n1724 = ~n1584 & n1723 ;
  assign n1725 = n1724 ^ x83 ;
  assign n1726 = n177 & ~n1725 ;
  assign n1727 = n1726 ^ n375 ;
  assign n1728 = n1583 & ~n1727 ;
  assign n1729 = n174 & n1728 ;
  assign n1730 = x84 & n1729 ;
  assign n1865 = n1719 ^ x82 ;
  assign n1866 = n1726 & n1865 ;
  assign n1867 = n1866 ^ n1587 ;
  assign n1858 = n1712 ^ x81 ;
  assign n1859 = n1726 & n1858 ;
  assign n1860 = n1859 ^ n1715 ;
  assign n1851 = n1705 ^ x80 ;
  assign n1852 = n1726 & n1851 ;
  assign n1853 = n1852 ^ n1708 ;
  assign n1844 = n1698 ^ x79 ;
  assign n1845 = n1726 & n1844 ;
  assign n1846 = n1845 ^ n1701 ;
  assign n1837 = n1691 ^ x78 ;
  assign n1838 = n1726 & n1837 ;
  assign n1839 = n1838 ^ n1694 ;
  assign n1830 = n1684 ^ x77 ;
  assign n1831 = n1726 & n1830 ;
  assign n1832 = n1831 ^ n1687 ;
  assign n1823 = n1677 ^ x76 ;
  assign n1824 = n1726 & n1823 ;
  assign n1825 = n1824 ^ n1680 ;
  assign n1816 = n1670 ^ x75 ;
  assign n1817 = n1726 & n1816 ;
  assign n1818 = n1817 ^ n1673 ;
  assign n1809 = n1663 ^ x74 ;
  assign n1810 = n1726 & n1809 ;
  assign n1811 = n1810 ^ n1666 ;
  assign n1802 = n1656 ^ x73 ;
  assign n1803 = n1726 & n1802 ;
  assign n1804 = n1803 ^ n1659 ;
  assign n1795 = n1649 ^ x72 ;
  assign n1796 = n1726 & n1795 ;
  assign n1797 = n1796 ^ n1652 ;
  assign n1788 = n1642 ^ x71 ;
  assign n1789 = n1726 & n1788 ;
  assign n1790 = n1789 ^ n1645 ;
  assign n1781 = n1627 ^ x70 ;
  assign n1782 = n1726 & n1781 ;
  assign n1783 = n1782 ^ n1638 ;
  assign n1774 = n1620 ^ x69 ;
  assign n1775 = n1726 & n1774 ;
  assign n1776 = n1775 ^ n1623 ;
  assign n1767 = n1614 ^ x68 ;
  assign n1768 = n1726 & n1767 ;
  assign n1769 = n1768 ^ n1616 ;
  assign n1760 = n1608 ^ x67 ;
  assign n1761 = n1726 & n1760 ;
  assign n1762 = n1761 ^ n1610 ;
  assign n1731 = n1605 ^ x66 ;
  assign n1732 = n1726 & n1731 ;
  assign n1733 = n1732 ^ n1592 ;
  assign n1734 = n1733 ^ x67 ;
  assign n1737 = ~x43 & x64 ;
  assign n1740 = n1726 ^ x44 ;
  assign n1741 = n1737 & ~n1740 ;
  assign n1735 = x64 & n1726 ;
  assign n1736 = n1735 ^ x44 ;
  assign n1738 = n1737 ^ n1736 ;
  assign n1739 = x65 & ~n1738 ;
  assign n1742 = n1741 ^ n1739 ;
  assign n1743 = n1742 ^ x66 ;
  assign n1752 = x65 & n1726 ;
  assign n1746 = n1581 ^ x44 ;
  assign n1747 = n1746 ^ n1581 ;
  assign n1748 = n1726 & ~n1747 ;
  assign n1749 = n1748 ^ n1581 ;
  assign n1750 = x64 & n1749 ;
  assign n1751 = n1750 ^ x45 ;
  assign n1753 = n1752 ^ n1751 ;
  assign n1754 = n1753 ^ n1742 ;
  assign n1755 = n1743 & n1754 ;
  assign n1756 = n1755 ^ x66 ;
  assign n1757 = n1756 ^ n1733 ;
  assign n1758 = ~n1734 & n1757 ;
  assign n1759 = n1758 ^ x67 ;
  assign n1763 = n1762 ^ n1759 ;
  assign n1764 = n1762 ^ x68 ;
  assign n1765 = n1763 & ~n1764 ;
  assign n1766 = n1765 ^ x68 ;
  assign n1770 = n1769 ^ n1766 ;
  assign n1771 = n1769 ^ x69 ;
  assign n1772 = n1770 & ~n1771 ;
  assign n1773 = n1772 ^ x69 ;
  assign n1777 = n1776 ^ n1773 ;
  assign n1778 = n1776 ^ x70 ;
  assign n1779 = n1777 & ~n1778 ;
  assign n1780 = n1779 ^ x70 ;
  assign n1784 = n1783 ^ n1780 ;
  assign n1785 = n1783 ^ x71 ;
  assign n1786 = n1784 & ~n1785 ;
  assign n1787 = n1786 ^ x71 ;
  assign n1791 = n1790 ^ n1787 ;
  assign n1792 = n1790 ^ x72 ;
  assign n1793 = n1791 & ~n1792 ;
  assign n1794 = n1793 ^ x72 ;
  assign n1798 = n1797 ^ n1794 ;
  assign n1799 = n1797 ^ x73 ;
  assign n1800 = n1798 & ~n1799 ;
  assign n1801 = n1800 ^ x73 ;
  assign n1805 = n1804 ^ n1801 ;
  assign n1806 = n1804 ^ x74 ;
  assign n1807 = n1805 & ~n1806 ;
  assign n1808 = n1807 ^ x74 ;
  assign n1812 = n1811 ^ n1808 ;
  assign n1813 = n1811 ^ x75 ;
  assign n1814 = n1812 & ~n1813 ;
  assign n1815 = n1814 ^ x75 ;
  assign n1819 = n1818 ^ n1815 ;
  assign n1820 = n1818 ^ x76 ;
  assign n1821 = n1819 & ~n1820 ;
  assign n1822 = n1821 ^ x76 ;
  assign n1826 = n1825 ^ n1822 ;
  assign n1827 = n1825 ^ x77 ;
  assign n1828 = n1826 & ~n1827 ;
  assign n1829 = n1828 ^ x77 ;
  assign n1833 = n1832 ^ n1829 ;
  assign n1834 = n1832 ^ x78 ;
  assign n1835 = n1833 & ~n1834 ;
  assign n1836 = n1835 ^ x78 ;
  assign n1840 = n1839 ^ n1836 ;
  assign n1841 = n1839 ^ x79 ;
  assign n1842 = n1840 & ~n1841 ;
  assign n1843 = n1842 ^ x79 ;
  assign n1847 = n1846 ^ n1843 ;
  assign n1848 = n1846 ^ x80 ;
  assign n1849 = n1847 & ~n1848 ;
  assign n1850 = n1849 ^ x80 ;
  assign n1854 = n1853 ^ n1850 ;
  assign n1855 = n1853 ^ x81 ;
  assign n1856 = n1854 & ~n1855 ;
  assign n1857 = n1856 ^ x81 ;
  assign n1861 = n1860 ^ n1857 ;
  assign n1862 = n1860 ^ x82 ;
  assign n1863 = n1861 & ~n1862 ;
  assign n1864 = n1863 ^ x82 ;
  assign n1868 = n1867 ^ n1864 ;
  assign n1869 = n1867 ^ x83 ;
  assign n1870 = n1868 & ~n1869 ;
  assign n1871 = n1870 ^ x83 ;
  assign n1872 = n1730 & n1871 ;
  assign n1873 = n1872 ^ n1729 ;
  assign n1874 = n1873 ^ n1728 ;
  assign n1875 = ~x86 & n172 ;
  assign n1876 = n1874 ^ x85 ;
  assign n1886 = n1874 ^ x84 ;
  assign n1877 = n1864 ^ x83 ;
  assign n1878 = n1728 ^ x84 ;
  assign n1879 = n1871 ^ x84 ;
  assign n1880 = ~n1878 & n1879 ;
  assign n1881 = n1880 ^ x84 ;
  assign n1882 = n174 & ~n1881 ;
  assign n1883 = n1877 & n1882 ;
  assign n1884 = n1883 ^ n1867 ;
  assign n1885 = n1884 ^ n1874 ;
  assign n1887 = n1886 ^ n1885 ;
  assign n2019 = n1857 ^ x82 ;
  assign n2020 = n1882 & n2019 ;
  assign n2021 = n2020 ^ n1860 ;
  assign n2012 = n1850 ^ x81 ;
  assign n2013 = n1882 & n2012 ;
  assign n2014 = n2013 ^ n1853 ;
  assign n2005 = n1843 ^ x80 ;
  assign n2006 = n1882 & n2005 ;
  assign n2007 = n2006 ^ n1846 ;
  assign n1998 = n1836 ^ x79 ;
  assign n1999 = n1882 & n1998 ;
  assign n2000 = n1999 ^ n1839 ;
  assign n1991 = n1829 ^ x78 ;
  assign n1992 = n1882 & n1991 ;
  assign n1993 = n1992 ^ n1832 ;
  assign n1984 = n1822 ^ x77 ;
  assign n1985 = n1882 & n1984 ;
  assign n1986 = n1985 ^ n1825 ;
  assign n1977 = n1815 ^ x76 ;
  assign n1978 = n1882 & n1977 ;
  assign n1979 = n1978 ^ n1818 ;
  assign n1888 = n1808 ^ x75 ;
  assign n1889 = n1882 & n1888 ;
  assign n1890 = n1889 ^ n1811 ;
  assign n1891 = n1890 ^ x76 ;
  assign n1892 = n1801 ^ x74 ;
  assign n1893 = n1882 & n1892 ;
  assign n1894 = n1893 ^ n1804 ;
  assign n1895 = n1894 ^ x75 ;
  assign n1964 = n1794 ^ x73 ;
  assign n1965 = n1882 & n1964 ;
  assign n1966 = n1965 ^ n1797 ;
  assign n1957 = n1787 ^ x72 ;
  assign n1958 = n1882 & n1957 ;
  assign n1959 = n1958 ^ n1790 ;
  assign n1950 = n1780 ^ x71 ;
  assign n1951 = n1882 & n1950 ;
  assign n1952 = n1951 ^ n1783 ;
  assign n1943 = n1773 ^ x70 ;
  assign n1944 = n1882 & n1943 ;
  assign n1945 = n1944 ^ n1776 ;
  assign n1936 = n1766 ^ x69 ;
  assign n1937 = n1882 & n1936 ;
  assign n1938 = n1937 ^ n1769 ;
  assign n1929 = n1759 ^ x68 ;
  assign n1930 = n1882 & n1929 ;
  assign n1931 = n1930 ^ n1762 ;
  assign n1922 = n1756 ^ x67 ;
  assign n1923 = n1882 & n1922 ;
  assign n1924 = n1923 ^ n1733 ;
  assign n1916 = n1743 & n1882 ;
  assign n1917 = n1916 ^ n1753 ;
  assign n1896 = n1737 ^ x65 ;
  assign n1897 = n1882 & n1896 ;
  assign n1898 = n1897 ^ n1736 ;
  assign n1899 = n1898 ^ x66 ;
  assign n1900 = ~x42 & x64 ;
  assign n1901 = n1900 ^ x43 ;
  assign n1908 = x65 & n1901 ;
  assign n1905 = n1900 ^ x65 ;
  assign n1906 = n1901 ^ n1882 ;
  assign n1907 = n1905 & n1906 ;
  assign n1909 = n1908 ^ n1907 ;
  assign n1910 = x64 & n1909 ;
  assign n1911 = n1910 ^ n1908 ;
  assign n1912 = n1911 ^ x65 ;
  assign n1913 = n1912 ^ n1898 ;
  assign n1914 = ~n1899 & n1913 ;
  assign n1915 = n1914 ^ x66 ;
  assign n1918 = n1917 ^ n1915 ;
  assign n1919 = n1917 ^ x67 ;
  assign n1920 = n1918 & ~n1919 ;
  assign n1921 = n1920 ^ x67 ;
  assign n1925 = n1924 ^ n1921 ;
  assign n1926 = n1924 ^ x68 ;
  assign n1927 = n1925 & ~n1926 ;
  assign n1928 = n1927 ^ x68 ;
  assign n1932 = n1931 ^ n1928 ;
  assign n1933 = n1931 ^ x69 ;
  assign n1934 = n1932 & ~n1933 ;
  assign n1935 = n1934 ^ x69 ;
  assign n1939 = n1938 ^ n1935 ;
  assign n1940 = n1938 ^ x70 ;
  assign n1941 = n1939 & ~n1940 ;
  assign n1942 = n1941 ^ x70 ;
  assign n1946 = n1945 ^ n1942 ;
  assign n1947 = n1945 ^ x71 ;
  assign n1948 = n1946 & ~n1947 ;
  assign n1949 = n1948 ^ x71 ;
  assign n1953 = n1952 ^ n1949 ;
  assign n1954 = n1952 ^ x72 ;
  assign n1955 = n1953 & ~n1954 ;
  assign n1956 = n1955 ^ x72 ;
  assign n1960 = n1959 ^ n1956 ;
  assign n1961 = n1959 ^ x73 ;
  assign n1962 = n1960 & ~n1961 ;
  assign n1963 = n1962 ^ x73 ;
  assign n1967 = n1966 ^ n1963 ;
  assign n1968 = n1966 ^ x74 ;
  assign n1969 = n1967 & ~n1968 ;
  assign n1970 = n1969 ^ x74 ;
  assign n1971 = n1970 ^ n1894 ;
  assign n1972 = ~n1895 & n1971 ;
  assign n1973 = n1972 ^ x75 ;
  assign n1974 = n1973 ^ n1890 ;
  assign n1975 = ~n1891 & n1974 ;
  assign n1976 = n1975 ^ x76 ;
  assign n1980 = n1979 ^ n1976 ;
  assign n1981 = n1979 ^ x77 ;
  assign n1982 = n1980 & ~n1981 ;
  assign n1983 = n1982 ^ x77 ;
  assign n1987 = n1986 ^ n1983 ;
  assign n1988 = n1986 ^ x78 ;
  assign n1989 = n1987 & ~n1988 ;
  assign n1990 = n1989 ^ x78 ;
  assign n1994 = n1993 ^ n1990 ;
  assign n1995 = n1993 ^ x79 ;
  assign n1996 = n1994 & ~n1995 ;
  assign n1997 = n1996 ^ x79 ;
  assign n2001 = n2000 ^ n1997 ;
  assign n2002 = n2000 ^ x80 ;
  assign n2003 = n2001 & ~n2002 ;
  assign n2004 = n2003 ^ x80 ;
  assign n2008 = n2007 ^ n2004 ;
  assign n2009 = n2007 ^ x81 ;
  assign n2010 = n2008 & ~n2009 ;
  assign n2011 = n2010 ^ x81 ;
  assign n2015 = n2014 ^ n2011 ;
  assign n2016 = n2014 ^ x82 ;
  assign n2017 = n2015 & ~n2016 ;
  assign n2018 = n2017 ^ x82 ;
  assign n2022 = n2021 ^ n2018 ;
  assign n2023 = n2021 ^ x83 ;
  assign n2024 = n2022 & ~n2023 ;
  assign n2025 = n2024 ^ x83 ;
  assign n2026 = n2025 ^ n1874 ;
  assign n2027 = n2026 ^ n1886 ;
  assign n2028 = ~n1887 & n2027 ;
  assign n2029 = n2028 ^ n1886 ;
  assign n2030 = ~n1876 & n2029 ;
  assign n2031 = n2030 ^ x85 ;
  assign n2032 = n1875 & ~n2031 ;
  assign n2033 = n1874 & ~n2032 ;
  assign n2034 = n2033 ^ n375 ;
  assign n2193 = n1875 & n2034 ;
  assign n2035 = n2025 ^ x84 ;
  assign n2036 = n2032 & n2035 ;
  assign n2037 = n2036 ^ n1884 ;
  assign n2038 = x85 & ~n2037 ;
  assign n2039 = n2034 ^ x86 ;
  assign n2040 = n172 & ~n2039 ;
  assign n2041 = ~n2038 & n2040 ;
  assign n2042 = n2018 ^ x83 ;
  assign n2043 = n2032 & n2042 ;
  assign n2044 = n2043 ^ n2021 ;
  assign n2045 = ~x84 & n2044 ;
  assign n2046 = n2037 ^ x85 ;
  assign n2047 = n2046 ^ n2038 ;
  assign n2048 = ~n2045 & ~n2047 ;
  assign n2049 = n2044 ^ x84 ;
  assign n2050 = n2049 ^ n2045 ;
  assign n2183 = n2011 ^ x82 ;
  assign n2184 = n2032 & n2183 ;
  assign n2185 = n2184 ^ n2014 ;
  assign n2176 = n2004 ^ x81 ;
  assign n2177 = n2032 & n2176 ;
  assign n2178 = n2177 ^ n2007 ;
  assign n2051 = n1997 ^ x80 ;
  assign n2052 = n2032 & n2051 ;
  assign n2053 = n2052 ^ n2000 ;
  assign n2054 = n2053 ^ x81 ;
  assign n2055 = n1990 ^ x79 ;
  assign n2056 = n2032 & n2055 ;
  assign n2057 = n2056 ^ n1993 ;
  assign n2058 = n2057 ^ x80 ;
  assign n2163 = n1983 ^ x78 ;
  assign n2164 = n2032 & n2163 ;
  assign n2165 = n2164 ^ n1986 ;
  assign n2156 = n1976 ^ x77 ;
  assign n2157 = n2032 & n2156 ;
  assign n2158 = n2157 ^ n1979 ;
  assign n2149 = n1973 ^ x76 ;
  assign n2150 = n2032 & n2149 ;
  assign n2151 = n2150 ^ n1890 ;
  assign n2142 = n1970 ^ x75 ;
  assign n2143 = n2032 & n2142 ;
  assign n2144 = n2143 ^ n1894 ;
  assign n2135 = n1963 ^ x74 ;
  assign n2136 = n2032 & n2135 ;
  assign n2137 = n2136 ^ n1966 ;
  assign n2128 = n1956 ^ x73 ;
  assign n2129 = n2032 & n2128 ;
  assign n2130 = n2129 ^ n1959 ;
  assign n2121 = n1949 ^ x72 ;
  assign n2122 = n2032 & n2121 ;
  assign n2123 = n2122 ^ n1952 ;
  assign n2114 = n1942 ^ x71 ;
  assign n2115 = n2032 & n2114 ;
  assign n2116 = n2115 ^ n1945 ;
  assign n2107 = n1935 ^ x70 ;
  assign n2108 = n2032 & n2107 ;
  assign n2109 = n2108 ^ n1938 ;
  assign n2100 = n1928 ^ x69 ;
  assign n2101 = n2032 & n2100 ;
  assign n2102 = n2101 ^ n1931 ;
  assign n2093 = n1921 ^ x68 ;
  assign n2094 = n2032 & n2093 ;
  assign n2095 = n2094 ^ n1924 ;
  assign n2086 = n1915 ^ x67 ;
  assign n2087 = n2032 & n2086 ;
  assign n2088 = n2087 ^ n1917 ;
  assign n2079 = n1912 ^ x66 ;
  assign n2080 = n2032 & n2079 ;
  assign n2081 = n2080 ^ n1898 ;
  assign n2072 = x64 & n1882 ;
  assign n2071 = n1905 & n2032 ;
  assign n2073 = n2072 ^ n2071 ;
  assign n2074 = n2073 ^ x43 ;
  assign n2066 = x42 & x65 ;
  assign n2063 = x65 ^ x41 ;
  assign n2059 = x64 ^ x42 ;
  assign n2060 = n2059 ^ x65 ;
  assign n2064 = n2060 ^ n2032 ;
  assign n2065 = ~n2063 & n2064 ;
  assign n2067 = n2066 ^ n2065 ;
  assign n2068 = x64 & n2067 ;
  assign n2069 = n2068 ^ n2066 ;
  assign n2070 = n2069 ^ x65 ;
  assign n2075 = n2074 ^ n2070 ;
  assign n2076 = n2074 ^ x66 ;
  assign n2077 = n2075 & ~n2076 ;
  assign n2078 = n2077 ^ x66 ;
  assign n2082 = n2081 ^ n2078 ;
  assign n2083 = n2081 ^ x67 ;
  assign n2084 = n2082 & ~n2083 ;
  assign n2085 = n2084 ^ x67 ;
  assign n2089 = n2088 ^ n2085 ;
  assign n2090 = n2088 ^ x68 ;
  assign n2091 = n2089 & ~n2090 ;
  assign n2092 = n2091 ^ x68 ;
  assign n2096 = n2095 ^ n2092 ;
  assign n2097 = n2095 ^ x69 ;
  assign n2098 = n2096 & ~n2097 ;
  assign n2099 = n2098 ^ x69 ;
  assign n2103 = n2102 ^ n2099 ;
  assign n2104 = n2102 ^ x70 ;
  assign n2105 = n2103 & ~n2104 ;
  assign n2106 = n2105 ^ x70 ;
  assign n2110 = n2109 ^ n2106 ;
  assign n2111 = n2109 ^ x71 ;
  assign n2112 = n2110 & ~n2111 ;
  assign n2113 = n2112 ^ x71 ;
  assign n2117 = n2116 ^ n2113 ;
  assign n2118 = n2116 ^ x72 ;
  assign n2119 = n2117 & ~n2118 ;
  assign n2120 = n2119 ^ x72 ;
  assign n2124 = n2123 ^ n2120 ;
  assign n2125 = n2123 ^ x73 ;
  assign n2126 = n2124 & ~n2125 ;
  assign n2127 = n2126 ^ x73 ;
  assign n2131 = n2130 ^ n2127 ;
  assign n2132 = n2130 ^ x74 ;
  assign n2133 = n2131 & ~n2132 ;
  assign n2134 = n2133 ^ x74 ;
  assign n2138 = n2137 ^ n2134 ;
  assign n2139 = n2137 ^ x75 ;
  assign n2140 = n2138 & ~n2139 ;
  assign n2141 = n2140 ^ x75 ;
  assign n2145 = n2144 ^ n2141 ;
  assign n2146 = n2144 ^ x76 ;
  assign n2147 = n2145 & ~n2146 ;
  assign n2148 = n2147 ^ x76 ;
  assign n2152 = n2151 ^ n2148 ;
  assign n2153 = n2151 ^ x77 ;
  assign n2154 = n2152 & ~n2153 ;
  assign n2155 = n2154 ^ x77 ;
  assign n2159 = n2158 ^ n2155 ;
  assign n2160 = n2158 ^ x78 ;
  assign n2161 = n2159 & ~n2160 ;
  assign n2162 = n2161 ^ x78 ;
  assign n2166 = n2165 ^ n2162 ;
  assign n2167 = n2165 ^ x79 ;
  assign n2168 = n2166 & ~n2167 ;
  assign n2169 = n2168 ^ x79 ;
  assign n2170 = n2169 ^ n2057 ;
  assign n2171 = ~n2058 & n2170 ;
  assign n2172 = n2171 ^ x80 ;
  assign n2173 = n2172 ^ n2053 ;
  assign n2174 = ~n2054 & n2173 ;
  assign n2175 = n2174 ^ x81 ;
  assign n2179 = n2178 ^ n2175 ;
  assign n2180 = n2178 ^ x82 ;
  assign n2181 = n2179 & ~n2180 ;
  assign n2182 = n2181 ^ x82 ;
  assign n2186 = n2185 ^ n2182 ;
  assign n2187 = n2185 ^ x83 ;
  assign n2188 = n2186 & ~n2187 ;
  assign n2189 = n2188 ^ x83 ;
  assign n2190 = ~n2050 & ~n2189 ;
  assign n2191 = n2048 & ~n2190 ;
  assign n2192 = n2041 & ~n2191 ;
  assign n2194 = n2193 ^ n2192 ;
  assign n2195 = n2194 ^ n375 ;
  assign n2196 = n2034 & ~n2195 ;
  assign n2543 = ~n172 & n2196 ;
  assign n2361 = ~n2045 & ~n2190 ;
  assign n2362 = n2361 ^ x85 ;
  assign n2363 = n2194 & n2362 ;
  assign n2364 = n2363 ^ n2037 ;
  assign n2348 = n2189 ^ x84 ;
  assign n2349 = n2194 & n2348 ;
  assign n2350 = n2349 ^ n2044 ;
  assign n2341 = n2182 ^ x83 ;
  assign n2342 = n2194 & n2341 ;
  assign n2343 = n2342 ^ n2185 ;
  assign n2334 = n2175 ^ x82 ;
  assign n2335 = n2194 & n2334 ;
  assign n2336 = n2335 ^ n2178 ;
  assign n2327 = n2172 ^ x81 ;
  assign n2328 = n2194 & n2327 ;
  assign n2329 = n2328 ^ n2053 ;
  assign n2320 = n2169 ^ x80 ;
  assign n2321 = n2194 & n2320 ;
  assign n2322 = n2321 ^ n2057 ;
  assign n2313 = n2162 ^ x79 ;
  assign n2314 = n2194 & n2313 ;
  assign n2315 = n2314 ^ n2165 ;
  assign n2306 = n2155 ^ x78 ;
  assign n2307 = n2194 & n2306 ;
  assign n2308 = n2307 ^ n2158 ;
  assign n2299 = n2148 ^ x77 ;
  assign n2300 = n2194 & n2299 ;
  assign n2301 = n2300 ^ n2151 ;
  assign n2292 = n2141 ^ x76 ;
  assign n2293 = n2194 & n2292 ;
  assign n2294 = n2293 ^ n2144 ;
  assign n2285 = n2134 ^ x75 ;
  assign n2286 = n2194 & n2285 ;
  assign n2287 = n2286 ^ n2137 ;
  assign n2278 = n2127 ^ x74 ;
  assign n2279 = n2194 & n2278 ;
  assign n2280 = n2279 ^ n2130 ;
  assign n2271 = n2120 ^ x73 ;
  assign n2272 = n2194 & n2271 ;
  assign n2273 = n2272 ^ n2123 ;
  assign n2264 = n2113 ^ x72 ;
  assign n2265 = n2194 & n2264 ;
  assign n2266 = n2265 ^ n2116 ;
  assign n2257 = n2106 ^ x71 ;
  assign n2258 = n2194 & n2257 ;
  assign n2259 = n2258 ^ n2109 ;
  assign n2250 = n2099 ^ x70 ;
  assign n2251 = n2194 & n2250 ;
  assign n2252 = n2251 ^ n2102 ;
  assign n2243 = n2092 ^ x69 ;
  assign n2244 = n2194 & n2243 ;
  assign n2245 = n2244 ^ n2095 ;
  assign n2200 = n2085 ^ x68 ;
  assign n2201 = n2194 & n2200 ;
  assign n2202 = n2201 ^ n2088 ;
  assign n2203 = n2202 ^ x69 ;
  assign n2204 = n2078 ^ x67 ;
  assign n2205 = n2194 & n2204 ;
  assign n2206 = n2205 ^ n2081 ;
  assign n2207 = n2206 ^ x68 ;
  assign n2230 = n2070 ^ x66 ;
  assign n2231 = n2194 & n2230 ;
  assign n2232 = n2231 ^ n2074 ;
  assign n2223 = x64 & n2032 ;
  assign n2221 = x65 ^ x42 ;
  assign n2215 = n2194 ^ x41 ;
  assign n2210 = x64 & n2194 ;
  assign n2219 = n2210 ^ x65 ;
  assign n2220 = n2215 & n2219 ;
  assign n2222 = n2221 ^ n2220 ;
  assign n2224 = n2223 ^ n2222 ;
  assign n2214 = ~x41 & x65 ;
  assign n2225 = n2224 ^ n2214 ;
  assign n2208 = ~x40 & x64 ;
  assign n2209 = n2208 ^ x65 ;
  assign n2211 = n2210 ^ n2063 ;
  assign n2212 = n2209 & ~n2211 ;
  assign n2213 = n2212 ^ x65 ;
  assign n2226 = n2225 ^ n2213 ;
  assign n2227 = n2225 ^ x66 ;
  assign n2228 = n2226 & ~n2227 ;
  assign n2229 = n2228 ^ x66 ;
  assign n2233 = n2232 ^ n2229 ;
  assign n2234 = n2232 ^ x67 ;
  assign n2235 = n2233 & ~n2234 ;
  assign n2236 = n2235 ^ x67 ;
  assign n2237 = n2236 ^ n2206 ;
  assign n2238 = ~n2207 & n2237 ;
  assign n2239 = n2238 ^ x68 ;
  assign n2240 = n2239 ^ n2202 ;
  assign n2241 = ~n2203 & n2240 ;
  assign n2242 = n2241 ^ x69 ;
  assign n2246 = n2245 ^ n2242 ;
  assign n2247 = n2245 ^ x70 ;
  assign n2248 = n2246 & ~n2247 ;
  assign n2249 = n2248 ^ x70 ;
  assign n2253 = n2252 ^ n2249 ;
  assign n2254 = n2252 ^ x71 ;
  assign n2255 = n2253 & ~n2254 ;
  assign n2256 = n2255 ^ x71 ;
  assign n2260 = n2259 ^ n2256 ;
  assign n2261 = n2259 ^ x72 ;
  assign n2262 = n2260 & ~n2261 ;
  assign n2263 = n2262 ^ x72 ;
  assign n2267 = n2266 ^ n2263 ;
  assign n2268 = n2266 ^ x73 ;
  assign n2269 = n2267 & ~n2268 ;
  assign n2270 = n2269 ^ x73 ;
  assign n2274 = n2273 ^ n2270 ;
  assign n2275 = n2273 ^ x74 ;
  assign n2276 = n2274 & ~n2275 ;
  assign n2277 = n2276 ^ x74 ;
  assign n2281 = n2280 ^ n2277 ;
  assign n2282 = n2280 ^ x75 ;
  assign n2283 = n2281 & ~n2282 ;
  assign n2284 = n2283 ^ x75 ;
  assign n2288 = n2287 ^ n2284 ;
  assign n2289 = n2287 ^ x76 ;
  assign n2290 = n2288 & ~n2289 ;
  assign n2291 = n2290 ^ x76 ;
  assign n2295 = n2294 ^ n2291 ;
  assign n2296 = n2294 ^ x77 ;
  assign n2297 = n2295 & ~n2296 ;
  assign n2298 = n2297 ^ x77 ;
  assign n2302 = n2301 ^ n2298 ;
  assign n2303 = n2301 ^ x78 ;
  assign n2304 = n2302 & ~n2303 ;
  assign n2305 = n2304 ^ x78 ;
  assign n2309 = n2308 ^ n2305 ;
  assign n2310 = n2308 ^ x79 ;
  assign n2311 = n2309 & ~n2310 ;
  assign n2312 = n2311 ^ x79 ;
  assign n2316 = n2315 ^ n2312 ;
  assign n2317 = n2315 ^ x80 ;
  assign n2318 = n2316 & ~n2317 ;
  assign n2319 = n2318 ^ x80 ;
  assign n2323 = n2322 ^ n2319 ;
  assign n2324 = n2322 ^ x81 ;
  assign n2325 = n2323 & ~n2324 ;
  assign n2326 = n2325 ^ x81 ;
  assign n2330 = n2329 ^ n2326 ;
  assign n2331 = n2329 ^ x82 ;
  assign n2332 = n2330 & ~n2331 ;
  assign n2333 = n2332 ^ x82 ;
  assign n2337 = n2336 ^ n2333 ;
  assign n2338 = n2336 ^ x83 ;
  assign n2339 = n2337 & ~n2338 ;
  assign n2340 = n2339 ^ x83 ;
  assign n2344 = n2343 ^ n2340 ;
  assign n2345 = n2343 ^ x84 ;
  assign n2346 = n2344 & ~n2345 ;
  assign n2347 = n2346 ^ x84 ;
  assign n2351 = n2350 ^ n2347 ;
  assign n2352 = n2350 ^ x85 ;
  assign n2353 = n2351 & ~n2352 ;
  assign n2354 = n2353 ^ x85 ;
  assign n2365 = n2364 ^ n2354 ;
  assign n2366 = n2364 ^ x86 ;
  assign n2367 = n2365 & ~n2366 ;
  assign n2368 = n2367 ^ x86 ;
  assign n2544 = n171 & ~n2368 ;
  assign n2545 = n2543 & ~n2544 ;
  assign n2197 = x88 & n170 ;
  assign n2198 = ~n2196 & n2197 ;
  assign n2199 = n2198 ^ n170 ;
  assign n2355 = n2354 ^ x86 ;
  assign n2356 = n2196 ^ x87 ;
  assign n2369 = n2368 ^ x87 ;
  assign n2370 = ~n2356 & n2369 ;
  assign n2371 = n2370 ^ x87 ;
  assign n2372 = n171 & ~n2371 ;
  assign n2373 = n2355 & n2372 ;
  assign n2374 = n2373 ^ n2364 ;
  assign n2375 = n2374 ^ x87 ;
  assign n2528 = n2347 ^ x85 ;
  assign n2529 = n2372 & n2528 ;
  assign n2530 = n2529 ^ n2350 ;
  assign n2521 = n2340 ^ x84 ;
  assign n2522 = n2372 & n2521 ;
  assign n2523 = n2522 ^ n2343 ;
  assign n2514 = n2333 ^ x83 ;
  assign n2515 = n2372 & n2514 ;
  assign n2516 = n2515 ^ n2336 ;
  assign n2507 = n2326 ^ x82 ;
  assign n2508 = n2372 & n2507 ;
  assign n2509 = n2508 ^ n2329 ;
  assign n2500 = n2319 ^ x81 ;
  assign n2501 = n2372 & n2500 ;
  assign n2502 = n2501 ^ n2322 ;
  assign n2493 = n2312 ^ x80 ;
  assign n2494 = n2372 & n2493 ;
  assign n2495 = n2494 ^ n2315 ;
  assign n2486 = n2305 ^ x79 ;
  assign n2487 = n2372 & n2486 ;
  assign n2488 = n2487 ^ n2308 ;
  assign n2479 = n2298 ^ x78 ;
  assign n2480 = n2372 & n2479 ;
  assign n2481 = n2480 ^ n2301 ;
  assign n2472 = n2291 ^ x77 ;
  assign n2473 = n2372 & n2472 ;
  assign n2474 = n2473 ^ n2294 ;
  assign n2465 = n2284 ^ x76 ;
  assign n2466 = n2372 & n2465 ;
  assign n2467 = n2466 ^ n2287 ;
  assign n2458 = n2277 ^ x75 ;
  assign n2459 = n2372 & n2458 ;
  assign n2460 = n2459 ^ n2280 ;
  assign n2451 = n2270 ^ x74 ;
  assign n2452 = n2372 & n2451 ;
  assign n2453 = n2452 ^ n2273 ;
  assign n2376 = n2263 ^ x73 ;
  assign n2377 = n2372 & n2376 ;
  assign n2378 = n2377 ^ n2266 ;
  assign n2379 = n2378 ^ x74 ;
  assign n2380 = n2256 ^ x72 ;
  assign n2381 = n2372 & n2380 ;
  assign n2382 = n2381 ^ n2259 ;
  assign n2383 = n2382 ^ x73 ;
  assign n2438 = n2249 ^ x71 ;
  assign n2439 = n2372 & n2438 ;
  assign n2440 = n2439 ^ n2252 ;
  assign n2431 = n2242 ^ x70 ;
  assign n2432 = n2372 & n2431 ;
  assign n2433 = n2432 ^ n2245 ;
  assign n2424 = n2239 ^ x69 ;
  assign n2425 = n2372 & n2424 ;
  assign n2426 = n2425 ^ n2202 ;
  assign n2417 = n2236 ^ x68 ;
  assign n2418 = n2372 & n2417 ;
  assign n2419 = n2418 ^ n2206 ;
  assign n2410 = n2229 ^ x67 ;
  assign n2411 = n2372 & n2410 ;
  assign n2412 = n2411 ^ n2232 ;
  assign n2403 = n2213 ^ x66 ;
  assign n2404 = n2372 & n2403 ;
  assign n2405 = n2404 ^ n2225 ;
  assign n2385 = n2209 & n2372 ;
  assign n2384 = n2210 ^ x41 ;
  assign n2386 = n2385 ^ n2384 ;
  assign n2387 = n2386 ^ x66 ;
  assign n2389 = x65 ^ x39 ;
  assign n2390 = x64 ^ x40 ;
  assign n2391 = n2390 ^ x65 ;
  assign n2392 = n2391 ^ n2372 ;
  assign n2393 = ~n2389 & n2392 ;
  assign n2388 = x40 & x65 ;
  assign n2394 = n2393 ^ n2388 ;
  assign n2397 = x64 & n2394 ;
  assign n2398 = n2397 ^ n2388 ;
  assign n2399 = n2398 ^ x65 ;
  assign n2400 = n2399 ^ n2386 ;
  assign n2401 = ~n2387 & n2400 ;
  assign n2402 = n2401 ^ x66 ;
  assign n2406 = n2405 ^ n2402 ;
  assign n2407 = n2405 ^ x67 ;
  assign n2408 = n2406 & ~n2407 ;
  assign n2409 = n2408 ^ x67 ;
  assign n2413 = n2412 ^ n2409 ;
  assign n2414 = n2412 ^ x68 ;
  assign n2415 = n2413 & ~n2414 ;
  assign n2416 = n2415 ^ x68 ;
  assign n2420 = n2419 ^ n2416 ;
  assign n2421 = n2419 ^ x69 ;
  assign n2422 = n2420 & ~n2421 ;
  assign n2423 = n2422 ^ x69 ;
  assign n2427 = n2426 ^ n2423 ;
  assign n2428 = n2426 ^ x70 ;
  assign n2429 = n2427 & ~n2428 ;
  assign n2430 = n2429 ^ x70 ;
  assign n2434 = n2433 ^ n2430 ;
  assign n2435 = n2433 ^ x71 ;
  assign n2436 = n2434 & ~n2435 ;
  assign n2437 = n2436 ^ x71 ;
  assign n2441 = n2440 ^ n2437 ;
  assign n2442 = n2440 ^ x72 ;
  assign n2443 = n2441 & ~n2442 ;
  assign n2444 = n2443 ^ x72 ;
  assign n2445 = n2444 ^ n2382 ;
  assign n2446 = ~n2383 & n2445 ;
  assign n2447 = n2446 ^ x73 ;
  assign n2448 = n2447 ^ n2378 ;
  assign n2449 = ~n2379 & n2448 ;
  assign n2450 = n2449 ^ x74 ;
  assign n2454 = n2453 ^ n2450 ;
  assign n2455 = n2453 ^ x75 ;
  assign n2456 = n2454 & ~n2455 ;
  assign n2457 = n2456 ^ x75 ;
  assign n2461 = n2460 ^ n2457 ;
  assign n2462 = n2460 ^ x76 ;
  assign n2463 = n2461 & ~n2462 ;
  assign n2464 = n2463 ^ x76 ;
  assign n2468 = n2467 ^ n2464 ;
  assign n2469 = n2467 ^ x77 ;
  assign n2470 = n2468 & ~n2469 ;
  assign n2471 = n2470 ^ x77 ;
  assign n2475 = n2474 ^ n2471 ;
  assign n2476 = n2474 ^ x78 ;
  assign n2477 = n2475 & ~n2476 ;
  assign n2478 = n2477 ^ x78 ;
  assign n2482 = n2481 ^ n2478 ;
  assign n2483 = n2481 ^ x79 ;
  assign n2484 = n2482 & ~n2483 ;
  assign n2485 = n2484 ^ x79 ;
  assign n2489 = n2488 ^ n2485 ;
  assign n2490 = n2488 ^ x80 ;
  assign n2491 = n2489 & ~n2490 ;
  assign n2492 = n2491 ^ x80 ;
  assign n2496 = n2495 ^ n2492 ;
  assign n2497 = n2495 ^ x81 ;
  assign n2498 = n2496 & ~n2497 ;
  assign n2499 = n2498 ^ x81 ;
  assign n2503 = n2502 ^ n2499 ;
  assign n2504 = n2502 ^ x82 ;
  assign n2505 = n2503 & ~n2504 ;
  assign n2506 = n2505 ^ x82 ;
  assign n2510 = n2509 ^ n2506 ;
  assign n2511 = n2509 ^ x83 ;
  assign n2512 = n2510 & ~n2511 ;
  assign n2513 = n2512 ^ x83 ;
  assign n2517 = n2516 ^ n2513 ;
  assign n2518 = n2516 ^ x84 ;
  assign n2519 = n2517 & ~n2518 ;
  assign n2520 = n2519 ^ x84 ;
  assign n2524 = n2523 ^ n2520 ;
  assign n2525 = n2523 ^ x85 ;
  assign n2526 = n2524 & ~n2525 ;
  assign n2527 = n2526 ^ x85 ;
  assign n2531 = n2530 ^ n2527 ;
  assign n2610 = n2527 ^ x86 ;
  assign n2535 = n2531 & n2610 ;
  assign n2532 = x87 ^ x86 ;
  assign n2536 = n2535 ^ n2532 ;
  assign n2539 = ~n2375 & n2536 ;
  assign n2540 = n2539 ^ x87 ;
  assign n2541 = n2199 & n2540 ;
  assign n2542 = n2198 ^ x88 ;
  assign n2546 = n2545 ^ n2542 ;
  assign n2547 = n2541 & ~n2546 ;
  assign n2548 = n2547 ^ n2199 ;
  assign n2602 = n2545 & ~n2548 ;
  assign n2603 = n2602 ^ n375 ;
  assign n2923 = n375 ^ n168 ;
  assign n2924 = n2603 & n2923 ;
  assign n2927 = n2924 ^ n2603 ;
  assign n2604 = n2603 ^ x89 ;
  assign n2608 = n2603 ^ x88 ;
  assign n2605 = n2536 & n2548 ;
  assign n2606 = n2605 ^ n2374 ;
  assign n2607 = n2606 ^ n2603 ;
  assign n2609 = n2608 ^ n2607 ;
  assign n2611 = n2548 & n2610 ;
  assign n2612 = n2611 ^ n2530 ;
  assign n2613 = n2612 ^ x87 ;
  assign n2719 = n2520 ^ x85 ;
  assign n2720 = n2548 & n2719 ;
  assign n2721 = n2720 ^ n2523 ;
  assign n2712 = n2513 ^ x84 ;
  assign n2713 = n2548 & n2712 ;
  assign n2714 = n2713 ^ n2516 ;
  assign n2705 = n2506 ^ x83 ;
  assign n2706 = n2548 & n2705 ;
  assign n2707 = n2706 ^ n2509 ;
  assign n2698 = n2499 ^ x82 ;
  assign n2699 = n2548 & n2698 ;
  assign n2700 = n2699 ^ n2502 ;
  assign n2691 = n2492 ^ x81 ;
  assign n2692 = n2548 & n2691 ;
  assign n2693 = n2692 ^ n2495 ;
  assign n2684 = n2485 ^ x80 ;
  assign n2685 = n2548 & n2684 ;
  assign n2686 = n2685 ^ n2488 ;
  assign n2677 = n2478 ^ x79 ;
  assign n2678 = n2548 & n2677 ;
  assign n2679 = n2678 ^ n2481 ;
  assign n2670 = n2471 ^ x78 ;
  assign n2671 = n2548 & n2670 ;
  assign n2672 = n2671 ^ n2474 ;
  assign n2663 = n2464 ^ x77 ;
  assign n2664 = n2548 & n2663 ;
  assign n2665 = n2664 ^ n2467 ;
  assign n2656 = n2457 ^ x76 ;
  assign n2657 = n2548 & n2656 ;
  assign n2658 = n2657 ^ n2460 ;
  assign n2649 = n2450 ^ x75 ;
  assign n2650 = n2548 & n2649 ;
  assign n2651 = n2650 ^ n2453 ;
  assign n2642 = n2447 ^ x74 ;
  assign n2643 = n2548 & n2642 ;
  assign n2644 = n2643 ^ n2378 ;
  assign n2635 = n2444 ^ x73 ;
  assign n2636 = n2548 & n2635 ;
  assign n2637 = n2636 ^ n2382 ;
  assign n2628 = n2437 ^ x72 ;
  assign n2629 = n2548 & n2628 ;
  assign n2630 = n2629 ^ n2440 ;
  assign n2621 = n2430 ^ x71 ;
  assign n2622 = n2548 & n2621 ;
  assign n2623 = n2622 ^ n2433 ;
  assign n2614 = n2423 ^ x70 ;
  assign n2615 = n2548 & n2614 ;
  assign n2616 = n2615 ^ n2426 ;
  assign n2594 = n2416 ^ x69 ;
  assign n2595 = n2548 & n2594 ;
  assign n2596 = n2595 ^ n2419 ;
  assign n2587 = n2409 ^ x68 ;
  assign n2588 = n2548 & n2587 ;
  assign n2589 = n2588 ^ n2412 ;
  assign n2580 = n2402 ^ x67 ;
  assign n2581 = n2548 & n2580 ;
  assign n2582 = n2581 ^ n2405 ;
  assign n2573 = n2399 ^ x66 ;
  assign n2574 = n2548 & n2573 ;
  assign n2575 = n2574 ^ n2386 ;
  assign n167 = x65 ^ x38 ;
  assign n2549 = x64 ^ x39 ;
  assign n2550 = n2549 ^ x65 ;
  assign n2551 = n2550 ^ n2548 ;
  assign n2552 = ~n167 & n2551 ;
  assign n166 = x39 & x65 ;
  assign n2553 = n2552 ^ n166 ;
  assign n2556 = x64 & n2553 ;
  assign n2557 = n2556 ^ n166 ;
  assign n2558 = n2557 ^ x65 ;
  assign n2559 = n2558 ^ x66 ;
  assign n2568 = x65 & n2548 ;
  assign n2562 = n2372 ^ x39 ;
  assign n2563 = n2562 ^ n2372 ;
  assign n2564 = n2548 & ~n2563 ;
  assign n2565 = n2564 ^ n2372 ;
  assign n2566 = x64 & n2565 ;
  assign n2567 = n2566 ^ x40 ;
  assign n2569 = n2568 ^ n2567 ;
  assign n2570 = n2569 ^ n2558 ;
  assign n2571 = n2559 & n2570 ;
  assign n2572 = n2571 ^ x66 ;
  assign n2576 = n2575 ^ n2572 ;
  assign n2577 = n2575 ^ x67 ;
  assign n2578 = n2576 & ~n2577 ;
  assign n2579 = n2578 ^ x67 ;
  assign n2583 = n2582 ^ n2579 ;
  assign n2584 = n2582 ^ x68 ;
  assign n2585 = n2583 & ~n2584 ;
  assign n2586 = n2585 ^ x68 ;
  assign n2590 = n2589 ^ n2586 ;
  assign n2591 = n2589 ^ x69 ;
  assign n2592 = n2590 & ~n2591 ;
  assign n2593 = n2592 ^ x69 ;
  assign n2597 = n2596 ^ n2593 ;
  assign n2598 = n2596 ^ x70 ;
  assign n2599 = n2597 & ~n2598 ;
  assign n2600 = n2599 ^ x70 ;
  assign n2617 = n2616 ^ n2600 ;
  assign n2618 = n2616 ^ x71 ;
  assign n2619 = n2617 & ~n2618 ;
  assign n2620 = n2619 ^ x71 ;
  assign n2624 = n2623 ^ n2620 ;
  assign n2625 = n2623 ^ x72 ;
  assign n2626 = n2624 & ~n2625 ;
  assign n2627 = n2626 ^ x72 ;
  assign n2631 = n2630 ^ n2627 ;
  assign n2632 = n2630 ^ x73 ;
  assign n2633 = n2631 & ~n2632 ;
  assign n2634 = n2633 ^ x73 ;
  assign n2638 = n2637 ^ n2634 ;
  assign n2639 = n2637 ^ x74 ;
  assign n2640 = n2638 & ~n2639 ;
  assign n2641 = n2640 ^ x74 ;
  assign n2645 = n2644 ^ n2641 ;
  assign n2646 = n2644 ^ x75 ;
  assign n2647 = n2645 & ~n2646 ;
  assign n2648 = n2647 ^ x75 ;
  assign n2652 = n2651 ^ n2648 ;
  assign n2653 = n2651 ^ x76 ;
  assign n2654 = n2652 & ~n2653 ;
  assign n2655 = n2654 ^ x76 ;
  assign n2659 = n2658 ^ n2655 ;
  assign n2660 = n2658 ^ x77 ;
  assign n2661 = n2659 & ~n2660 ;
  assign n2662 = n2661 ^ x77 ;
  assign n2666 = n2665 ^ n2662 ;
  assign n2667 = n2665 ^ x78 ;
  assign n2668 = n2666 & ~n2667 ;
  assign n2669 = n2668 ^ x78 ;
  assign n2673 = n2672 ^ n2669 ;
  assign n2674 = n2672 ^ x79 ;
  assign n2675 = n2673 & ~n2674 ;
  assign n2676 = n2675 ^ x79 ;
  assign n2680 = n2679 ^ n2676 ;
  assign n2681 = n2679 ^ x80 ;
  assign n2682 = n2680 & ~n2681 ;
  assign n2683 = n2682 ^ x80 ;
  assign n2687 = n2686 ^ n2683 ;
  assign n2688 = n2686 ^ x81 ;
  assign n2689 = n2687 & ~n2688 ;
  assign n2690 = n2689 ^ x81 ;
  assign n2694 = n2693 ^ n2690 ;
  assign n2695 = n2693 ^ x82 ;
  assign n2696 = n2694 & ~n2695 ;
  assign n2697 = n2696 ^ x82 ;
  assign n2701 = n2700 ^ n2697 ;
  assign n2702 = n2700 ^ x83 ;
  assign n2703 = n2701 & ~n2702 ;
  assign n2704 = n2703 ^ x83 ;
  assign n2708 = n2707 ^ n2704 ;
  assign n2709 = n2707 ^ x84 ;
  assign n2710 = n2708 & ~n2709 ;
  assign n2711 = n2710 ^ x84 ;
  assign n2715 = n2714 ^ n2711 ;
  assign n2716 = n2714 ^ x85 ;
  assign n2717 = n2715 & ~n2716 ;
  assign n2718 = n2717 ^ x85 ;
  assign n2722 = n2721 ^ n2718 ;
  assign n2723 = n2721 ^ x86 ;
  assign n2724 = n2722 & ~n2723 ;
  assign n2725 = n2724 ^ x86 ;
  assign n2726 = n2725 ^ n2612 ;
  assign n2727 = ~n2613 & n2726 ;
  assign n2728 = n2727 ^ x87 ;
  assign n2729 = n2728 ^ n2603 ;
  assign n2730 = n2729 ^ n2608 ;
  assign n2731 = ~n2609 & n2730 ;
  assign n2732 = n2731 ^ n2608 ;
  assign n2733 = ~n2604 & n2732 ;
  assign n2734 = n2733 ^ x89 ;
  assign n2735 = n169 & ~n2734 ;
  assign n2916 = n2728 ^ x88 ;
  assign n2917 = n2735 & n2916 ;
  assign n2918 = n2917 ^ n2606 ;
  assign n2909 = n2725 ^ x87 ;
  assign n2910 = n2735 & n2909 ;
  assign n2911 = n2910 ^ n2612 ;
  assign n2902 = n2718 ^ x86 ;
  assign n2903 = n2735 & n2902 ;
  assign n2904 = n2903 ^ n2721 ;
  assign n2895 = n2711 ^ x85 ;
  assign n2896 = n2735 & n2895 ;
  assign n2897 = n2896 ^ n2714 ;
  assign n2888 = n2704 ^ x84 ;
  assign n2889 = n2735 & n2888 ;
  assign n2890 = n2889 ^ n2707 ;
  assign n2881 = n2697 ^ x83 ;
  assign n2882 = n2735 & n2881 ;
  assign n2883 = n2882 ^ n2700 ;
  assign n2874 = n2690 ^ x82 ;
  assign n2875 = n2735 & n2874 ;
  assign n2876 = n2875 ^ n2693 ;
  assign n2867 = n2683 ^ x81 ;
  assign n2868 = n2735 & n2867 ;
  assign n2869 = n2868 ^ n2686 ;
  assign n2860 = n2676 ^ x80 ;
  assign n2861 = n2735 & n2860 ;
  assign n2862 = n2861 ^ n2679 ;
  assign n2853 = n2669 ^ x79 ;
  assign n2854 = n2735 & n2853 ;
  assign n2855 = n2854 ^ n2672 ;
  assign n2846 = n2662 ^ x78 ;
  assign n2847 = n2735 & n2846 ;
  assign n2848 = n2847 ^ n2665 ;
  assign n2839 = n2655 ^ x77 ;
  assign n2840 = n2735 & n2839 ;
  assign n2841 = n2840 ^ n2658 ;
  assign n2832 = n2648 ^ x76 ;
  assign n2833 = n2735 & n2832 ;
  assign n2834 = n2833 ^ n2651 ;
  assign n2825 = n2641 ^ x75 ;
  assign n2826 = n2735 & n2825 ;
  assign n2827 = n2826 ^ n2644 ;
  assign n2818 = n2634 ^ x74 ;
  assign n2819 = n2735 & n2818 ;
  assign n2820 = n2819 ^ n2637 ;
  assign n2811 = n2627 ^ x73 ;
  assign n2812 = n2735 & n2811 ;
  assign n2813 = n2812 ^ n2630 ;
  assign n2804 = n2620 ^ x72 ;
  assign n2805 = n2735 & n2804 ;
  assign n2806 = n2805 ^ n2623 ;
  assign n2601 = n2600 ^ x71 ;
  assign n2736 = n2601 & n2735 ;
  assign n2737 = n2736 ^ n2616 ;
  assign n2738 = n2737 ^ x72 ;
  assign n2743 = n2737 ^ x71 ;
  assign n2739 = n2593 ^ x70 ;
  assign n2740 = n2735 & n2739 ;
  assign n2741 = n2740 ^ n2596 ;
  assign n2742 = n2741 ^ n2737 ;
  assign n2744 = n2743 ^ n2742 ;
  assign n2791 = n2586 ^ x69 ;
  assign n2792 = n2735 & n2791 ;
  assign n2793 = n2792 ^ n2589 ;
  assign n2784 = n2579 ^ x68 ;
  assign n2785 = n2735 & n2784 ;
  assign n2786 = n2785 ^ n2582 ;
  assign n2777 = n2572 ^ x67 ;
  assign n2778 = n2735 & n2777 ;
  assign n2779 = n2778 ^ n2575 ;
  assign n2771 = n2559 & n2735 ;
  assign n2772 = n2771 ^ n2569 ;
  assign n2753 = x65 & n2735 ;
  assign n2745 = n2548 ^ x38 ;
  assign n2746 = n2745 ^ n2548 ;
  assign n2749 = n2735 & ~n2746 ;
  assign n2750 = n2749 ^ n2548 ;
  assign n2751 = x64 & n2750 ;
  assign n2752 = n2751 ^ x39 ;
  assign n2754 = n2753 ^ n2752 ;
  assign n2755 = n2754 ^ x66 ;
  assign n2763 = x38 & x65 ;
  assign n2760 = x65 ^ x37 ;
  assign n2756 = x64 ^ x38 ;
  assign n2757 = n2756 ^ x65 ;
  assign n2761 = n2757 ^ n2735 ;
  assign n2762 = ~n2760 & n2761 ;
  assign n2764 = n2763 ^ n2762 ;
  assign n2765 = x64 & n2764 ;
  assign n2766 = n2765 ^ n2763 ;
  assign n2767 = n2766 ^ x65 ;
  assign n2768 = n2767 ^ n2754 ;
  assign n2769 = ~n2755 & n2768 ;
  assign n2770 = n2769 ^ x66 ;
  assign n2773 = n2772 ^ n2770 ;
  assign n2774 = n2772 ^ x67 ;
  assign n2775 = n2773 & ~n2774 ;
  assign n2776 = n2775 ^ x67 ;
  assign n2780 = n2779 ^ n2776 ;
  assign n2781 = n2779 ^ x68 ;
  assign n2782 = n2780 & ~n2781 ;
  assign n2783 = n2782 ^ x68 ;
  assign n2787 = n2786 ^ n2783 ;
  assign n2788 = n2786 ^ x69 ;
  assign n2789 = n2787 & ~n2788 ;
  assign n2790 = n2789 ^ x69 ;
  assign n2794 = n2793 ^ n2790 ;
  assign n2795 = n2793 ^ x70 ;
  assign n2796 = n2794 & ~n2795 ;
  assign n2797 = n2796 ^ x70 ;
  assign n2798 = n2797 ^ n2737 ;
  assign n2799 = n2798 ^ n2743 ;
  assign n2800 = ~n2744 & n2799 ;
  assign n2801 = n2800 ^ n2743 ;
  assign n2802 = ~n2738 & n2801 ;
  assign n2803 = n2802 ^ x72 ;
  assign n2807 = n2806 ^ n2803 ;
  assign n2808 = n2806 ^ x73 ;
  assign n2809 = n2807 & ~n2808 ;
  assign n2810 = n2809 ^ x73 ;
  assign n2814 = n2813 ^ n2810 ;
  assign n2815 = n2813 ^ x74 ;
  assign n2816 = n2814 & ~n2815 ;
  assign n2817 = n2816 ^ x74 ;
  assign n2821 = n2820 ^ n2817 ;
  assign n2822 = n2820 ^ x75 ;
  assign n2823 = n2821 & ~n2822 ;
  assign n2824 = n2823 ^ x75 ;
  assign n2828 = n2827 ^ n2824 ;
  assign n2829 = n2827 ^ x76 ;
  assign n2830 = n2828 & ~n2829 ;
  assign n2831 = n2830 ^ x76 ;
  assign n2835 = n2834 ^ n2831 ;
  assign n2836 = n2834 ^ x77 ;
  assign n2837 = n2835 & ~n2836 ;
  assign n2838 = n2837 ^ x77 ;
  assign n2842 = n2841 ^ n2838 ;
  assign n2843 = n2841 ^ x78 ;
  assign n2844 = n2842 & ~n2843 ;
  assign n2845 = n2844 ^ x78 ;
  assign n2849 = n2848 ^ n2845 ;
  assign n2850 = n2848 ^ x79 ;
  assign n2851 = n2849 & ~n2850 ;
  assign n2852 = n2851 ^ x79 ;
  assign n2856 = n2855 ^ n2852 ;
  assign n2857 = n2855 ^ x80 ;
  assign n2858 = n2856 & ~n2857 ;
  assign n2859 = n2858 ^ x80 ;
  assign n2863 = n2862 ^ n2859 ;
  assign n2864 = n2862 ^ x81 ;
  assign n2865 = n2863 & ~n2864 ;
  assign n2866 = n2865 ^ x81 ;
  assign n2870 = n2869 ^ n2866 ;
  assign n2871 = n2869 ^ x82 ;
  assign n2872 = n2870 & ~n2871 ;
  assign n2873 = n2872 ^ x82 ;
  assign n2877 = n2876 ^ n2873 ;
  assign n2878 = n2876 ^ x83 ;
  assign n2879 = n2877 & ~n2878 ;
  assign n2880 = n2879 ^ x83 ;
  assign n2884 = n2883 ^ n2880 ;
  assign n2885 = n2883 ^ x84 ;
  assign n2886 = n2884 & ~n2885 ;
  assign n2887 = n2886 ^ x84 ;
  assign n2891 = n2890 ^ n2887 ;
  assign n2892 = n2890 ^ x85 ;
  assign n2893 = n2891 & ~n2892 ;
  assign n2894 = n2893 ^ x85 ;
  assign n2898 = n2897 ^ n2894 ;
  assign n2899 = n2897 ^ x86 ;
  assign n2900 = n2898 & ~n2899 ;
  assign n2901 = n2900 ^ x86 ;
  assign n2905 = n2904 ^ n2901 ;
  assign n2906 = n2904 ^ x87 ;
  assign n2907 = n2905 & ~n2906 ;
  assign n2908 = n2907 ^ x87 ;
  assign n2912 = n2911 ^ n2908 ;
  assign n2913 = n2911 ^ x88 ;
  assign n2914 = n2912 & ~n2913 ;
  assign n2915 = n2914 ^ x88 ;
  assign n2919 = n2918 ^ n2915 ;
  assign n2920 = n2918 ^ x89 ;
  assign n2921 = n2919 & ~n2920 ;
  assign n2922 = n2921 ^ x89 ;
  assign n2925 = x90 & n2924 ;
  assign n2926 = n2922 & n2925 ;
  assign n2928 = n2927 ^ n2926 ;
  assign n2929 = n2928 ^ x91 ;
  assign n3134 = n2928 ^ x90 ;
  assign n2930 = n2908 ^ x88 ;
  assign n2931 = n2922 ^ x90 ;
  assign n2935 = n2922 ^ n375 ;
  assign n2932 = n2734 ^ n375 ;
  assign n2936 = n2935 ^ n2932 ;
  assign n2937 = ~n2603 & ~n2936 ;
  assign n2938 = n2937 ^ n2932 ;
  assign n2939 = n2931 & ~n2938 ;
  assign n2940 = n2939 ^ x90 ;
  assign n2941 = n168 & ~n2940 ;
  assign n2942 = n2930 & n2941 ;
  assign n2943 = n2942 ^ n2911 ;
  assign n2944 = n2943 ^ x89 ;
  assign n3123 = n2901 ^ x87 ;
  assign n3124 = n2941 & n3123 ;
  assign n3125 = n3124 ^ n2904 ;
  assign n3116 = n2894 ^ x86 ;
  assign n3117 = n2941 & n3116 ;
  assign n3118 = n3117 ^ n2897 ;
  assign n3109 = n2887 ^ x85 ;
  assign n3110 = n2941 & n3109 ;
  assign n3111 = n3110 ^ n2890 ;
  assign n3102 = n2880 ^ x84 ;
  assign n3103 = n2941 & n3102 ;
  assign n3104 = n3103 ^ n2883 ;
  assign n3095 = n2873 ^ x83 ;
  assign n3096 = n2941 & n3095 ;
  assign n3097 = n3096 ^ n2876 ;
  assign n3088 = n2866 ^ x82 ;
  assign n3089 = n2941 & n3088 ;
  assign n3090 = n3089 ^ n2869 ;
  assign n3081 = n2859 ^ x81 ;
  assign n3082 = n2941 & n3081 ;
  assign n3083 = n3082 ^ n2862 ;
  assign n2945 = n2852 ^ x80 ;
  assign n2946 = n2941 & n2945 ;
  assign n2947 = n2946 ^ n2855 ;
  assign n2948 = n2947 ^ x81 ;
  assign n2949 = n2845 ^ x79 ;
  assign n2950 = n2941 & n2949 ;
  assign n2951 = n2950 ^ n2848 ;
  assign n2952 = n2951 ^ x80 ;
  assign n3068 = n2838 ^ x78 ;
  assign n3069 = n2941 & n3068 ;
  assign n3070 = n3069 ^ n2841 ;
  assign n3061 = n2831 ^ x77 ;
  assign n3062 = n2941 & n3061 ;
  assign n3063 = n3062 ^ n2834 ;
  assign n3054 = n2824 ^ x76 ;
  assign n3055 = n2941 & n3054 ;
  assign n3056 = n3055 ^ n2827 ;
  assign n3047 = n2817 ^ x75 ;
  assign n3048 = n2941 & n3047 ;
  assign n3049 = n3048 ^ n2820 ;
  assign n3040 = n2810 ^ x74 ;
  assign n3041 = n2941 & n3040 ;
  assign n3042 = n3041 ^ n2813 ;
  assign n3033 = n2803 ^ x73 ;
  assign n3034 = n2941 & n3033 ;
  assign n3035 = n3034 ^ n2806 ;
  assign n3018 = n2741 ^ x72 ;
  assign n3019 = n3018 ^ x71 ;
  assign n3020 = n3019 ^ n2797 ;
  assign n3021 = n3020 ^ n3018 ;
  assign n3023 = x72 ^ x71 ;
  assign n3024 = n3023 ^ n3018 ;
  assign n3025 = ~n3021 & ~n3024 ;
  assign n3026 = n3025 ^ n3018 ;
  assign n3027 = n2941 & ~n3026 ;
  assign n3028 = n3027 ^ n2737 ;
  assign n3011 = n2797 ^ x71 ;
  assign n3012 = n2941 & n3011 ;
  assign n3013 = n3012 ^ n2741 ;
  assign n3004 = n2790 ^ x70 ;
  assign n3005 = n2941 & n3004 ;
  assign n3006 = n3005 ^ n2793 ;
  assign n2997 = n2783 ^ x69 ;
  assign n2998 = n2941 & n2997 ;
  assign n2999 = n2998 ^ n2786 ;
  assign n2990 = n2776 ^ x68 ;
  assign n2991 = n2941 & n2990 ;
  assign n2992 = n2991 ^ n2779 ;
  assign n2983 = n2770 ^ x67 ;
  assign n2984 = n2941 & n2983 ;
  assign n2985 = n2984 ^ n2772 ;
  assign n2976 = n2767 ^ x66 ;
  assign n2977 = n2941 & n2976 ;
  assign n2978 = n2977 ^ n2754 ;
  assign n2958 = x64 & n2735 ;
  assign n2954 = ~x37 & x64 ;
  assign n2955 = n2954 ^ x65 ;
  assign n2956 = n2941 & n2955 ;
  assign n2957 = n2956 ^ x38 ;
  assign n2959 = n2958 ^ n2957 ;
  assign n2960 = n2959 ^ x66 ;
  assign n2968 = x37 & x65 ;
  assign n2965 = x65 ^ x36 ;
  assign n2961 = x64 ^ x37 ;
  assign n2962 = n2961 ^ x65 ;
  assign n2966 = n2962 ^ n2941 ;
  assign n2967 = ~n2965 & n2966 ;
  assign n2969 = n2968 ^ n2967 ;
  assign n2970 = x64 & n2969 ;
  assign n2971 = n2970 ^ n2968 ;
  assign n2972 = n2971 ^ x65 ;
  assign n2973 = n2972 ^ n2959 ;
  assign n2974 = ~n2960 & n2973 ;
  assign n2975 = n2974 ^ x66 ;
  assign n2979 = n2978 ^ n2975 ;
  assign n2980 = n2978 ^ x67 ;
  assign n2981 = n2979 & ~n2980 ;
  assign n2982 = n2981 ^ x67 ;
  assign n2986 = n2985 ^ n2982 ;
  assign n2987 = n2985 ^ x68 ;
  assign n2988 = n2986 & ~n2987 ;
  assign n2989 = n2988 ^ x68 ;
  assign n2993 = n2992 ^ n2989 ;
  assign n2994 = n2992 ^ x69 ;
  assign n2995 = n2993 & ~n2994 ;
  assign n2996 = n2995 ^ x69 ;
  assign n3000 = n2999 ^ n2996 ;
  assign n3001 = n2999 ^ x70 ;
  assign n3002 = n3000 & ~n3001 ;
  assign n3003 = n3002 ^ x70 ;
  assign n3007 = n3006 ^ n3003 ;
  assign n3008 = n3006 ^ x71 ;
  assign n3009 = n3007 & ~n3008 ;
  assign n3010 = n3009 ^ x71 ;
  assign n3014 = n3013 ^ n3010 ;
  assign n3015 = n3013 ^ x72 ;
  assign n3016 = n3014 & ~n3015 ;
  assign n3017 = n3016 ^ x72 ;
  assign n3029 = n3028 ^ n3017 ;
  assign n3030 = n3028 ^ x73 ;
  assign n3031 = n3029 & ~n3030 ;
  assign n3032 = n3031 ^ x73 ;
  assign n3036 = n3035 ^ n3032 ;
  assign n3037 = n3035 ^ x74 ;
  assign n3038 = n3036 & ~n3037 ;
  assign n3039 = n3038 ^ x74 ;
  assign n3043 = n3042 ^ n3039 ;
  assign n3044 = n3042 ^ x75 ;
  assign n3045 = n3043 & ~n3044 ;
  assign n3046 = n3045 ^ x75 ;
  assign n3050 = n3049 ^ n3046 ;
  assign n3051 = n3049 ^ x76 ;
  assign n3052 = n3050 & ~n3051 ;
  assign n3053 = n3052 ^ x76 ;
  assign n3057 = n3056 ^ n3053 ;
  assign n3058 = n3056 ^ x77 ;
  assign n3059 = n3057 & ~n3058 ;
  assign n3060 = n3059 ^ x77 ;
  assign n3064 = n3063 ^ n3060 ;
  assign n3065 = n3063 ^ x78 ;
  assign n3066 = n3064 & ~n3065 ;
  assign n3067 = n3066 ^ x78 ;
  assign n3071 = n3070 ^ n3067 ;
  assign n3072 = n3070 ^ x79 ;
  assign n3073 = n3071 & ~n3072 ;
  assign n3074 = n3073 ^ x79 ;
  assign n3075 = n3074 ^ n2951 ;
  assign n3076 = ~n2952 & n3075 ;
  assign n3077 = n3076 ^ x80 ;
  assign n3078 = n3077 ^ n2947 ;
  assign n3079 = ~n2948 & n3078 ;
  assign n3080 = n3079 ^ x81 ;
  assign n3084 = n3083 ^ n3080 ;
  assign n3085 = n3083 ^ x82 ;
  assign n3086 = n3084 & ~n3085 ;
  assign n3087 = n3086 ^ x82 ;
  assign n3091 = n3090 ^ n3087 ;
  assign n3092 = n3090 ^ x83 ;
  assign n3093 = n3091 & ~n3092 ;
  assign n3094 = n3093 ^ x83 ;
  assign n3098 = n3097 ^ n3094 ;
  assign n3099 = n3097 ^ x84 ;
  assign n3100 = n3098 & ~n3099 ;
  assign n3101 = n3100 ^ x84 ;
  assign n3105 = n3104 ^ n3101 ;
  assign n3106 = n3104 ^ x85 ;
  assign n3107 = n3105 & ~n3106 ;
  assign n3108 = n3107 ^ x85 ;
  assign n3112 = n3111 ^ n3108 ;
  assign n3113 = n3111 ^ x86 ;
  assign n3114 = n3112 & ~n3113 ;
  assign n3115 = n3114 ^ x86 ;
  assign n3119 = n3118 ^ n3115 ;
  assign n3120 = n3118 ^ x87 ;
  assign n3121 = n3119 & ~n3120 ;
  assign n3122 = n3121 ^ x87 ;
  assign n3126 = n3125 ^ n3122 ;
  assign n3127 = n3125 ^ x88 ;
  assign n3128 = n3126 & ~n3127 ;
  assign n3129 = n3128 ^ x88 ;
  assign n3130 = n3129 ^ n2943 ;
  assign n3131 = ~n2944 & n3130 ;
  assign n3132 = n3131 ^ x89 ;
  assign n3133 = n3132 ^ n2928 ;
  assign n3135 = n3134 ^ n3133 ;
  assign n3136 = n2915 ^ x89 ;
  assign n3137 = n2941 & n3136 ;
  assign n3138 = n3137 ^ n2918 ;
  assign n3139 = n3138 ^ n2928 ;
  assign n3140 = n3139 ^ n3134 ;
  assign n3141 = n3135 & ~n3140 ;
  assign n3142 = n3141 ^ n3134 ;
  assign n3143 = ~n2929 & n3142 ;
  assign n3144 = n3143 ^ x91 ;
  assign n3145 = n165 & ~n3144 ;
  assign n3152 = n2928 & ~n3145 ;
  assign n3153 = n3152 ^ n375 ;
  assign n3154 = n3153 ^ x92 ;
  assign n3146 = n3132 ^ x90 ;
  assign n3147 = n3145 & n3146 ;
  assign n3148 = n3147 ^ n3138 ;
  assign n3150 = n3148 ^ x91 ;
  assign n3149 = x91 & ~n3148 ;
  assign n3151 = n3150 ^ n3149 ;
  assign n3155 = n3154 ^ n3151 ;
  assign n3156 = n3129 ^ x89 ;
  assign n3157 = n3145 & n3156 ;
  assign n3158 = n3157 ^ n2943 ;
  assign n3159 = n3158 ^ x90 ;
  assign n3160 = n3122 ^ x88 ;
  assign n3161 = n3145 & n3160 ;
  assign n3162 = n3161 ^ n3125 ;
  assign n3163 = n3162 ^ x89 ;
  assign n3164 = n3115 ^ x87 ;
  assign n3165 = n3145 & n3164 ;
  assign n3166 = n3165 ^ n3118 ;
  assign n3167 = n3166 ^ x88 ;
  assign n3172 = n3166 ^ x87 ;
  assign n3168 = n3108 ^ x86 ;
  assign n3169 = n3145 & n3168 ;
  assign n3170 = n3169 ^ n3111 ;
  assign n3171 = n3170 ^ n3166 ;
  assign n3173 = n3172 ^ n3171 ;
  assign n3326 = n3101 ^ x85 ;
  assign n3327 = n3145 & n3326 ;
  assign n3328 = n3327 ^ n3104 ;
  assign n3319 = n3094 ^ x84 ;
  assign n3320 = n3145 & n3319 ;
  assign n3321 = n3320 ^ n3097 ;
  assign n3312 = n3087 ^ x83 ;
  assign n3313 = n3145 & n3312 ;
  assign n3314 = n3313 ^ n3090 ;
  assign n3305 = n3080 ^ x82 ;
  assign n3306 = n3145 & n3305 ;
  assign n3307 = n3306 ^ n3083 ;
  assign n3298 = n3077 ^ x81 ;
  assign n3299 = n3145 & n3298 ;
  assign n3300 = n3299 ^ n2947 ;
  assign n3291 = n3074 ^ x80 ;
  assign n3292 = n3145 & n3291 ;
  assign n3293 = n3292 ^ n2951 ;
  assign n3284 = n3067 ^ x79 ;
  assign n3285 = n3145 & n3284 ;
  assign n3286 = n3285 ^ n3070 ;
  assign n3277 = n3060 ^ x78 ;
  assign n3278 = n3145 & n3277 ;
  assign n3279 = n3278 ^ n3063 ;
  assign n3270 = n3053 ^ x77 ;
  assign n3271 = n3145 & n3270 ;
  assign n3272 = n3271 ^ n3056 ;
  assign n3263 = n3046 ^ x76 ;
  assign n3264 = n3145 & n3263 ;
  assign n3265 = n3264 ^ n3049 ;
  assign n3256 = n3039 ^ x75 ;
  assign n3257 = n3145 & n3256 ;
  assign n3258 = n3257 ^ n3042 ;
  assign n3249 = n3032 ^ x74 ;
  assign n3250 = n3145 & n3249 ;
  assign n3251 = n3250 ^ n3035 ;
  assign n3242 = n3017 ^ x73 ;
  assign n3243 = n3145 & n3242 ;
  assign n3244 = n3243 ^ n3028 ;
  assign n3235 = n3010 ^ x72 ;
  assign n3236 = n3145 & n3235 ;
  assign n3237 = n3236 ^ n3013 ;
  assign n3228 = n3003 ^ x71 ;
  assign n3229 = n3145 & n3228 ;
  assign n3230 = n3229 ^ n3006 ;
  assign n3221 = n2996 ^ x70 ;
  assign n3222 = n3145 & n3221 ;
  assign n3223 = n3222 ^ n2999 ;
  assign n3214 = n2989 ^ x69 ;
  assign n3215 = n3145 & n3214 ;
  assign n3216 = n3215 ^ n2992 ;
  assign n3174 = n2982 ^ x68 ;
  assign n3175 = n3145 & n3174 ;
  assign n3176 = n3175 ^ n2985 ;
  assign n3177 = n3176 ^ x69 ;
  assign n3182 = n3176 ^ x68 ;
  assign n3178 = n2975 ^ x67 ;
  assign n3179 = n3145 & n3178 ;
  assign n3180 = n3179 ^ n2978 ;
  assign n3181 = n3180 ^ n3176 ;
  assign n3183 = n3182 ^ n3181 ;
  assign n3201 = n2972 ^ x66 ;
  assign n3202 = n3145 & n3201 ;
  assign n3203 = n3202 ^ n2959 ;
  assign n3195 = x64 & n2941 ;
  assign n3191 = ~x36 & x64 ;
  assign n3192 = n3191 ^ x65 ;
  assign n3193 = n3145 & n3192 ;
  assign n3194 = n3193 ^ x37 ;
  assign n3196 = n3195 ^ n3194 ;
  assign n3184 = ~x35 & x64 ;
  assign n3185 = n3184 ^ x65 ;
  assign n3186 = x64 & n3145 ;
  assign n3187 = n3186 ^ n2965 ;
  assign n3188 = n3185 & ~n3187 ;
  assign n3189 = n3188 ^ x65 ;
  assign n3197 = n3196 ^ n3189 ;
  assign n3198 = n3196 ^ x66 ;
  assign n3199 = n3197 & ~n3198 ;
  assign n3200 = n3199 ^ x66 ;
  assign n3204 = n3203 ^ n3200 ;
  assign n3205 = n3203 ^ x67 ;
  assign n3206 = n3204 & ~n3205 ;
  assign n3207 = n3206 ^ x67 ;
  assign n3208 = n3207 ^ n3176 ;
  assign n3209 = n3208 ^ n3182 ;
  assign n3210 = ~n3183 & n3209 ;
  assign n3211 = n3210 ^ n3182 ;
  assign n3212 = ~n3177 & n3211 ;
  assign n3213 = n3212 ^ x69 ;
  assign n3217 = n3216 ^ n3213 ;
  assign n3218 = n3216 ^ x70 ;
  assign n3219 = n3217 & ~n3218 ;
  assign n3220 = n3219 ^ x70 ;
  assign n3224 = n3223 ^ n3220 ;
  assign n3225 = n3223 ^ x71 ;
  assign n3226 = n3224 & ~n3225 ;
  assign n3227 = n3226 ^ x71 ;
  assign n3231 = n3230 ^ n3227 ;
  assign n3232 = n3230 ^ x72 ;
  assign n3233 = n3231 & ~n3232 ;
  assign n3234 = n3233 ^ x72 ;
  assign n3238 = n3237 ^ n3234 ;
  assign n3239 = n3237 ^ x73 ;
  assign n3240 = n3238 & ~n3239 ;
  assign n3241 = n3240 ^ x73 ;
  assign n3245 = n3244 ^ n3241 ;
  assign n3246 = n3244 ^ x74 ;
  assign n3247 = n3245 & ~n3246 ;
  assign n3248 = n3247 ^ x74 ;
  assign n3252 = n3251 ^ n3248 ;
  assign n3253 = n3251 ^ x75 ;
  assign n3254 = n3252 & ~n3253 ;
  assign n3255 = n3254 ^ x75 ;
  assign n3259 = n3258 ^ n3255 ;
  assign n3260 = n3258 ^ x76 ;
  assign n3261 = n3259 & ~n3260 ;
  assign n3262 = n3261 ^ x76 ;
  assign n3266 = n3265 ^ n3262 ;
  assign n3267 = n3265 ^ x77 ;
  assign n3268 = n3266 & ~n3267 ;
  assign n3269 = n3268 ^ x77 ;
  assign n3273 = n3272 ^ n3269 ;
  assign n3274 = n3272 ^ x78 ;
  assign n3275 = n3273 & ~n3274 ;
  assign n3276 = n3275 ^ x78 ;
  assign n3280 = n3279 ^ n3276 ;
  assign n3281 = n3279 ^ x79 ;
  assign n3282 = n3280 & ~n3281 ;
  assign n3283 = n3282 ^ x79 ;
  assign n3287 = n3286 ^ n3283 ;
  assign n3288 = n3286 ^ x80 ;
  assign n3289 = n3287 & ~n3288 ;
  assign n3290 = n3289 ^ x80 ;
  assign n3294 = n3293 ^ n3290 ;
  assign n3295 = n3293 ^ x81 ;
  assign n3296 = n3294 & ~n3295 ;
  assign n3297 = n3296 ^ x81 ;
  assign n3301 = n3300 ^ n3297 ;
  assign n3302 = n3300 ^ x82 ;
  assign n3303 = n3301 & ~n3302 ;
  assign n3304 = n3303 ^ x82 ;
  assign n3308 = n3307 ^ n3304 ;
  assign n3309 = n3307 ^ x83 ;
  assign n3310 = n3308 & ~n3309 ;
  assign n3311 = n3310 ^ x83 ;
  assign n3315 = n3314 ^ n3311 ;
  assign n3316 = n3314 ^ x84 ;
  assign n3317 = n3315 & ~n3316 ;
  assign n3318 = n3317 ^ x84 ;
  assign n3322 = n3321 ^ n3318 ;
  assign n3323 = n3321 ^ x85 ;
  assign n3324 = n3322 & ~n3323 ;
  assign n3325 = n3324 ^ x85 ;
  assign n3329 = n3328 ^ n3325 ;
  assign n3330 = n3328 ^ x86 ;
  assign n3331 = n3329 & ~n3330 ;
  assign n3332 = n3331 ^ x86 ;
  assign n3333 = n3332 ^ n3166 ;
  assign n3334 = n3333 ^ n3172 ;
  assign n3335 = ~n3173 & n3334 ;
  assign n3336 = n3335 ^ n3172 ;
  assign n3337 = ~n3167 & n3336 ;
  assign n3338 = n3337 ^ x88 ;
  assign n3339 = n3338 ^ n3162 ;
  assign n3340 = ~n3163 & n3339 ;
  assign n3341 = n3340 ^ x89 ;
  assign n3342 = n3341 ^ n3158 ;
  assign n3343 = ~n3159 & n3342 ;
  assign n3344 = n3343 ^ x90 ;
  assign n3345 = ~n3155 & n3344 ;
  assign n3346 = n3149 ^ x92 ;
  assign n3347 = ~n3154 & n3346 ;
  assign n3348 = n3347 ^ x92 ;
  assign n3349 = n164 & ~n3348 ;
  assign n3350 = ~n3345 & n3349 ;
  assign n3352 = n3152 & ~n3350 ;
  assign n3353 = n3352 ^ n375 ;
  assign n3354 = ~n164 & n3353 ;
  assign n3569 = n3344 ^ x91 ;
  assign n3570 = n3350 & n3569 ;
  assign n3571 = n3570 ^ n3148 ;
  assign n3355 = n3341 ^ x90 ;
  assign n3356 = n3350 & n3355 ;
  assign n3357 = n3356 ^ n3158 ;
  assign n3358 = n3357 ^ x91 ;
  assign n3363 = n3357 ^ x90 ;
  assign n3359 = n3338 ^ x89 ;
  assign n3360 = n3350 & n3359 ;
  assign n3361 = n3360 ^ n3162 ;
  assign n3362 = n3361 ^ n3357 ;
  assign n3364 = n3363 ^ n3362 ;
  assign n3548 = n3170 ^ x88 ;
  assign n3549 = n3548 ^ x87 ;
  assign n3550 = n3549 ^ n3332 ;
  assign n3551 = n3550 ^ n3548 ;
  assign n3553 = x88 ^ x87 ;
  assign n3554 = n3553 ^ n3548 ;
  assign n3555 = ~n3551 & ~n3554 ;
  assign n3556 = n3555 ^ n3548 ;
  assign n3557 = n3350 & ~n3556 ;
  assign n3558 = n3557 ^ n3166 ;
  assign n3541 = n3332 ^ x87 ;
  assign n3542 = n3350 & n3541 ;
  assign n3543 = n3542 ^ n3170 ;
  assign n3534 = n3325 ^ x86 ;
  assign n3535 = n3350 & n3534 ;
  assign n3536 = n3535 ^ n3328 ;
  assign n3527 = n3318 ^ x85 ;
  assign n3528 = n3350 & n3527 ;
  assign n3529 = n3528 ^ n3321 ;
  assign n3520 = n3311 ^ x84 ;
  assign n3521 = n3350 & n3520 ;
  assign n3522 = n3521 ^ n3314 ;
  assign n3513 = n3304 ^ x83 ;
  assign n3514 = n3350 & n3513 ;
  assign n3515 = n3514 ^ n3307 ;
  assign n3506 = n3297 ^ x82 ;
  assign n3507 = n3350 & n3506 ;
  assign n3508 = n3507 ^ n3300 ;
  assign n3499 = n3290 ^ x81 ;
  assign n3500 = n3350 & n3499 ;
  assign n3501 = n3500 ^ n3293 ;
  assign n3492 = n3283 ^ x80 ;
  assign n3493 = n3350 & n3492 ;
  assign n3494 = n3493 ^ n3286 ;
  assign n3485 = n3276 ^ x79 ;
  assign n3486 = n3350 & n3485 ;
  assign n3487 = n3486 ^ n3279 ;
  assign n3478 = n3269 ^ x78 ;
  assign n3479 = n3350 & n3478 ;
  assign n3480 = n3479 ^ n3272 ;
  assign n3471 = n3262 ^ x77 ;
  assign n3472 = n3350 & n3471 ;
  assign n3473 = n3472 ^ n3265 ;
  assign n3365 = n3255 ^ x76 ;
  assign n3366 = n3350 & n3365 ;
  assign n3367 = n3366 ^ n3258 ;
  assign n3368 = n3367 ^ x77 ;
  assign n3373 = n3367 ^ x76 ;
  assign n3369 = n3248 ^ x75 ;
  assign n3370 = n3350 & n3369 ;
  assign n3371 = n3370 ^ n3251 ;
  assign n3372 = n3371 ^ n3367 ;
  assign n3374 = n3373 ^ n3372 ;
  assign n3458 = n3241 ^ x74 ;
  assign n3459 = n3350 & n3458 ;
  assign n3460 = n3459 ^ n3244 ;
  assign n3451 = n3234 ^ x73 ;
  assign n3452 = n3350 & n3451 ;
  assign n3453 = n3452 ^ n3237 ;
  assign n3444 = n3227 ^ x72 ;
  assign n3445 = n3350 & n3444 ;
  assign n3446 = n3445 ^ n3230 ;
  assign n3437 = n3220 ^ x71 ;
  assign n3438 = n3350 & n3437 ;
  assign n3439 = n3438 ^ n3223 ;
  assign n3430 = n3213 ^ x70 ;
  assign n3431 = n3350 & n3430 ;
  assign n3432 = n3431 ^ n3216 ;
  assign n3415 = n3180 ^ x69 ;
  assign n3416 = n3415 ^ x68 ;
  assign n3417 = n3416 ^ n3207 ;
  assign n3418 = n3417 ^ n3415 ;
  assign n3420 = x69 ^ x68 ;
  assign n3421 = n3420 ^ n3415 ;
  assign n3422 = ~n3418 & ~n3421 ;
  assign n3423 = n3422 ^ n3415 ;
  assign n3424 = n3350 & ~n3423 ;
  assign n3425 = n3424 ^ n3176 ;
  assign n3408 = n3207 ^ x68 ;
  assign n3409 = n3350 & n3408 ;
  assign n3410 = n3409 ^ n3180 ;
  assign n3401 = n3200 ^ x67 ;
  assign n3402 = n3350 & n3401 ;
  assign n3403 = n3402 ^ n3203 ;
  assign n3394 = n3189 ^ x66 ;
  assign n3395 = n3350 & n3394 ;
  assign n3396 = n3395 ^ n3196 ;
  assign n3388 = n3186 ^ x36 ;
  assign n3387 = n3185 & n3350 ;
  assign n3389 = n3388 ^ n3387 ;
  assign n3382 = x35 & x65 ;
  assign n3379 = x65 ^ x34 ;
  assign n3375 = x64 ^ x35 ;
  assign n3376 = n3375 ^ x65 ;
  assign n3380 = n3376 ^ n3350 ;
  assign n3381 = ~n3379 & n3380 ;
  assign n3383 = n3382 ^ n3381 ;
  assign n3384 = x64 & n3383 ;
  assign n3385 = n3384 ^ n3382 ;
  assign n3386 = n3385 ^ x65 ;
  assign n3390 = n3389 ^ n3386 ;
  assign n3391 = n3389 ^ x66 ;
  assign n3392 = n3390 & ~n3391 ;
  assign n3393 = n3392 ^ x66 ;
  assign n3397 = n3396 ^ n3393 ;
  assign n3398 = n3396 ^ x67 ;
  assign n3399 = n3397 & ~n3398 ;
  assign n3400 = n3399 ^ x67 ;
  assign n3404 = n3403 ^ n3400 ;
  assign n3405 = n3403 ^ x68 ;
  assign n3406 = n3404 & ~n3405 ;
  assign n3407 = n3406 ^ x68 ;
  assign n3411 = n3410 ^ n3407 ;
  assign n3412 = n3410 ^ x69 ;
  assign n3413 = n3411 & ~n3412 ;
  assign n3414 = n3413 ^ x69 ;
  assign n3426 = n3425 ^ n3414 ;
  assign n3427 = n3425 ^ x70 ;
  assign n3428 = n3426 & ~n3427 ;
  assign n3429 = n3428 ^ x70 ;
  assign n3433 = n3432 ^ n3429 ;
  assign n3434 = n3432 ^ x71 ;
  assign n3435 = n3433 & ~n3434 ;
  assign n3436 = n3435 ^ x71 ;
  assign n3440 = n3439 ^ n3436 ;
  assign n3441 = n3439 ^ x72 ;
  assign n3442 = n3440 & ~n3441 ;
  assign n3443 = n3442 ^ x72 ;
  assign n3447 = n3446 ^ n3443 ;
  assign n3448 = n3446 ^ x73 ;
  assign n3449 = n3447 & ~n3448 ;
  assign n3450 = n3449 ^ x73 ;
  assign n3454 = n3453 ^ n3450 ;
  assign n3455 = n3453 ^ x74 ;
  assign n3456 = n3454 & ~n3455 ;
  assign n3457 = n3456 ^ x74 ;
  assign n3461 = n3460 ^ n3457 ;
  assign n3462 = n3460 ^ x75 ;
  assign n3463 = n3461 & ~n3462 ;
  assign n3464 = n3463 ^ x75 ;
  assign n3465 = n3464 ^ n3367 ;
  assign n3466 = n3465 ^ n3373 ;
  assign n3467 = ~n3374 & n3466 ;
  assign n3468 = n3467 ^ n3373 ;
  assign n3469 = ~n3368 & n3468 ;
  assign n3470 = n3469 ^ x77 ;
  assign n3474 = n3473 ^ n3470 ;
  assign n3475 = n3473 ^ x78 ;
  assign n3476 = n3474 & ~n3475 ;
  assign n3477 = n3476 ^ x78 ;
  assign n3481 = n3480 ^ n3477 ;
  assign n3482 = n3480 ^ x79 ;
  assign n3483 = n3481 & ~n3482 ;
  assign n3484 = n3483 ^ x79 ;
  assign n3488 = n3487 ^ n3484 ;
  assign n3489 = n3487 ^ x80 ;
  assign n3490 = n3488 & ~n3489 ;
  assign n3491 = n3490 ^ x80 ;
  assign n3495 = n3494 ^ n3491 ;
  assign n3496 = n3494 ^ x81 ;
  assign n3497 = n3495 & ~n3496 ;
  assign n3498 = n3497 ^ x81 ;
  assign n3502 = n3501 ^ n3498 ;
  assign n3503 = n3501 ^ x82 ;
  assign n3504 = n3502 & ~n3503 ;
  assign n3505 = n3504 ^ x82 ;
  assign n3509 = n3508 ^ n3505 ;
  assign n3510 = n3508 ^ x83 ;
  assign n3511 = n3509 & ~n3510 ;
  assign n3512 = n3511 ^ x83 ;
  assign n3516 = n3515 ^ n3512 ;
  assign n3517 = n3515 ^ x84 ;
  assign n3518 = n3516 & ~n3517 ;
  assign n3519 = n3518 ^ x84 ;
  assign n3523 = n3522 ^ n3519 ;
  assign n3524 = n3522 ^ x85 ;
  assign n3525 = n3523 & ~n3524 ;
  assign n3526 = n3525 ^ x85 ;
  assign n3530 = n3529 ^ n3526 ;
  assign n3531 = n3529 ^ x86 ;
  assign n3532 = n3530 & ~n3531 ;
  assign n3533 = n3532 ^ x86 ;
  assign n3537 = n3536 ^ n3533 ;
  assign n3538 = n3536 ^ x87 ;
  assign n3539 = n3537 & ~n3538 ;
  assign n3540 = n3539 ^ x87 ;
  assign n3544 = n3543 ^ n3540 ;
  assign n3545 = n3543 ^ x88 ;
  assign n3546 = n3544 & ~n3545 ;
  assign n3547 = n3546 ^ x88 ;
  assign n3559 = n3558 ^ n3547 ;
  assign n3560 = n3558 ^ x89 ;
  assign n3561 = n3559 & ~n3560 ;
  assign n3562 = n3561 ^ x89 ;
  assign n3563 = n3562 ^ n3357 ;
  assign n3564 = n3563 ^ n3363 ;
  assign n3565 = ~n3364 & n3564 ;
  assign n3566 = n3565 ^ n3363 ;
  assign n3567 = ~n3358 & n3566 ;
  assign n3568 = n3567 ^ x91 ;
  assign n3572 = n3571 ^ n3568 ;
  assign n3573 = n3571 ^ x92 ;
  assign n3574 = n3572 & ~n3573 ;
  assign n3575 = n3574 ^ x92 ;
  assign n3576 = n163 & ~n3575 ;
  assign n3577 = n3354 & ~n3576 ;
  assign n3579 = n3353 ^ x93 ;
  assign n3580 = n3575 ^ x93 ;
  assign n3581 = ~n3579 & n3580 ;
  assign n3582 = n3581 ^ x93 ;
  assign n3583 = n163 & ~n3582 ;
  assign n3809 = n3568 ^ x92 ;
  assign n3810 = n3583 & n3809 ;
  assign n3811 = n3810 ^ n3571 ;
  assign n3791 = n3361 ^ x91 ;
  assign n3792 = n3791 ^ n3562 ;
  assign n3793 = n3792 ^ x90 ;
  assign n3794 = n3793 ^ n3791 ;
  assign n3796 = n3562 ^ x91 ;
  assign n3797 = n3796 ^ n3791 ;
  assign n3798 = ~n3794 & ~n3797 ;
  assign n3799 = n3798 ^ n3791 ;
  assign n3800 = n3583 & ~n3799 ;
  assign n3801 = n3800 ^ n3357 ;
  assign n3784 = n3562 ^ x90 ;
  assign n3785 = n3583 & n3784 ;
  assign n3786 = n3785 ^ n3361 ;
  assign n3777 = n3547 ^ x89 ;
  assign n3778 = n3583 & n3777 ;
  assign n3779 = n3778 ^ n3558 ;
  assign n3770 = n3540 ^ x88 ;
  assign n3771 = n3583 & n3770 ;
  assign n3772 = n3771 ^ n3543 ;
  assign n3763 = n3533 ^ x87 ;
  assign n3764 = n3583 & n3763 ;
  assign n3765 = n3764 ^ n3536 ;
  assign n3756 = n3526 ^ x86 ;
  assign n3757 = n3583 & n3756 ;
  assign n3758 = n3757 ^ n3529 ;
  assign n3749 = n3519 ^ x85 ;
  assign n3750 = n3583 & n3749 ;
  assign n3751 = n3750 ^ n3522 ;
  assign n3742 = n3512 ^ x84 ;
  assign n3743 = n3583 & n3742 ;
  assign n3744 = n3743 ^ n3515 ;
  assign n3578 = n3505 ^ x83 ;
  assign n3584 = n3578 & n3583 ;
  assign n3585 = n3584 ^ n3508 ;
  assign n3586 = n3585 ^ x84 ;
  assign n3591 = n3585 ^ x83 ;
  assign n3587 = n3498 ^ x82 ;
  assign n3588 = n3583 & n3587 ;
  assign n3589 = n3588 ^ n3501 ;
  assign n3590 = n3589 ^ n3585 ;
  assign n3592 = n3591 ^ n3590 ;
  assign n3729 = n3491 ^ x81 ;
  assign n3730 = n3583 & n3729 ;
  assign n3731 = n3730 ^ n3494 ;
  assign n3722 = n3484 ^ x80 ;
  assign n3723 = n3583 & n3722 ;
  assign n3724 = n3723 ^ n3487 ;
  assign n3715 = n3477 ^ x79 ;
  assign n3716 = n3583 & n3715 ;
  assign n3717 = n3716 ^ n3480 ;
  assign n3708 = n3470 ^ x78 ;
  assign n3709 = n3583 & n3708 ;
  assign n3710 = n3709 ^ n3473 ;
  assign n3693 = n3371 ^ x77 ;
  assign n3694 = n3693 ^ n3464 ;
  assign n3695 = n3694 ^ x76 ;
  assign n3696 = n3695 ^ n3693 ;
  assign n3698 = n3464 ^ x77 ;
  assign n3699 = n3698 ^ n3693 ;
  assign n3700 = ~n3696 & ~n3699 ;
  assign n3701 = n3700 ^ n3693 ;
  assign n3702 = n3583 & ~n3701 ;
  assign n3703 = n3702 ^ n3367 ;
  assign n3686 = n3464 ^ x76 ;
  assign n3687 = n3583 & n3686 ;
  assign n3688 = n3687 ^ n3371 ;
  assign n3679 = n3457 ^ x75 ;
  assign n3680 = n3583 & n3679 ;
  assign n3681 = n3680 ^ n3460 ;
  assign n3672 = n3450 ^ x74 ;
  assign n3673 = n3583 & n3672 ;
  assign n3674 = n3673 ^ n3453 ;
  assign n3665 = n3443 ^ x73 ;
  assign n3666 = n3583 & n3665 ;
  assign n3667 = n3666 ^ n3446 ;
  assign n3658 = n3436 ^ x72 ;
  assign n3659 = n3583 & n3658 ;
  assign n3660 = n3659 ^ n3439 ;
  assign n3651 = n3429 ^ x71 ;
  assign n3652 = n3583 & n3651 ;
  assign n3653 = n3652 ^ n3432 ;
  assign n3644 = n3414 ^ x70 ;
  assign n3645 = n3583 & n3644 ;
  assign n3646 = n3645 ^ n3425 ;
  assign n3637 = n3407 ^ x69 ;
  assign n3638 = n3583 & n3637 ;
  assign n3639 = n3638 ^ n3410 ;
  assign n3630 = n3400 ^ x68 ;
  assign n3631 = n3583 & n3630 ;
  assign n3632 = n3631 ^ n3403 ;
  assign n3623 = n3393 ^ x67 ;
  assign n3624 = n3583 & n3623 ;
  assign n3625 = n3624 ^ n3396 ;
  assign n3616 = n3386 ^ x66 ;
  assign n3617 = n3583 & n3616 ;
  assign n3618 = n3617 ^ n3389 ;
  assign n3610 = x64 & n3350 ;
  assign n3606 = ~x34 & x64 ;
  assign n3607 = n3606 ^ x65 ;
  assign n3608 = n3583 & n3607 ;
  assign n3609 = n3608 ^ x35 ;
  assign n3611 = n3610 ^ n3609 ;
  assign n3600 = x34 & x65 ;
  assign n3597 = x65 ^ x33 ;
  assign n3593 = x64 ^ x34 ;
  assign n3594 = n3593 ^ x65 ;
  assign n3598 = n3594 ^ n3583 ;
  assign n3599 = ~n3597 & n3598 ;
  assign n3601 = n3600 ^ n3599 ;
  assign n3602 = x64 & n3601 ;
  assign n3603 = n3602 ^ n3600 ;
  assign n3604 = n3603 ^ x65 ;
  assign n3612 = n3611 ^ n3604 ;
  assign n3613 = n3611 ^ x66 ;
  assign n3614 = n3612 & ~n3613 ;
  assign n3615 = n3614 ^ x66 ;
  assign n3619 = n3618 ^ n3615 ;
  assign n3620 = n3618 ^ x67 ;
  assign n3621 = n3619 & ~n3620 ;
  assign n3622 = n3621 ^ x67 ;
  assign n3626 = n3625 ^ n3622 ;
  assign n3627 = n3625 ^ x68 ;
  assign n3628 = n3626 & ~n3627 ;
  assign n3629 = n3628 ^ x68 ;
  assign n3633 = n3632 ^ n3629 ;
  assign n3634 = n3632 ^ x69 ;
  assign n3635 = n3633 & ~n3634 ;
  assign n3636 = n3635 ^ x69 ;
  assign n3640 = n3639 ^ n3636 ;
  assign n3641 = n3639 ^ x70 ;
  assign n3642 = n3640 & ~n3641 ;
  assign n3643 = n3642 ^ x70 ;
  assign n3647 = n3646 ^ n3643 ;
  assign n3648 = n3646 ^ x71 ;
  assign n3649 = n3647 & ~n3648 ;
  assign n3650 = n3649 ^ x71 ;
  assign n3654 = n3653 ^ n3650 ;
  assign n3655 = n3653 ^ x72 ;
  assign n3656 = n3654 & ~n3655 ;
  assign n3657 = n3656 ^ x72 ;
  assign n3661 = n3660 ^ n3657 ;
  assign n3662 = n3660 ^ x73 ;
  assign n3663 = n3661 & ~n3662 ;
  assign n3664 = n3663 ^ x73 ;
  assign n3668 = n3667 ^ n3664 ;
  assign n3669 = n3667 ^ x74 ;
  assign n3670 = n3668 & ~n3669 ;
  assign n3671 = n3670 ^ x74 ;
  assign n3675 = n3674 ^ n3671 ;
  assign n3676 = n3674 ^ x75 ;
  assign n3677 = n3675 & ~n3676 ;
  assign n3678 = n3677 ^ x75 ;
  assign n3682 = n3681 ^ n3678 ;
  assign n3683 = n3681 ^ x76 ;
  assign n3684 = n3682 & ~n3683 ;
  assign n3685 = n3684 ^ x76 ;
  assign n3689 = n3688 ^ n3685 ;
  assign n3690 = n3688 ^ x77 ;
  assign n3691 = n3689 & ~n3690 ;
  assign n3692 = n3691 ^ x77 ;
  assign n3704 = n3703 ^ n3692 ;
  assign n3705 = n3703 ^ x78 ;
  assign n3706 = n3704 & ~n3705 ;
  assign n3707 = n3706 ^ x78 ;
  assign n3711 = n3710 ^ n3707 ;
  assign n3712 = n3710 ^ x79 ;
  assign n3713 = n3711 & ~n3712 ;
  assign n3714 = n3713 ^ x79 ;
  assign n3718 = n3717 ^ n3714 ;
  assign n3719 = n3717 ^ x80 ;
  assign n3720 = n3718 & ~n3719 ;
  assign n3721 = n3720 ^ x80 ;
  assign n3725 = n3724 ^ n3721 ;
  assign n3726 = n3724 ^ x81 ;
  assign n3727 = n3725 & ~n3726 ;
  assign n3728 = n3727 ^ x81 ;
  assign n3732 = n3731 ^ n3728 ;
  assign n3733 = n3731 ^ x82 ;
  assign n3734 = n3732 & ~n3733 ;
  assign n3735 = n3734 ^ x82 ;
  assign n3736 = n3735 ^ n3585 ;
  assign n3737 = n3736 ^ n3591 ;
  assign n3738 = ~n3592 & n3737 ;
  assign n3739 = n3738 ^ n3591 ;
  assign n3740 = ~n3586 & n3739 ;
  assign n3741 = n3740 ^ x84 ;
  assign n3745 = n3744 ^ n3741 ;
  assign n3746 = n3744 ^ x85 ;
  assign n3747 = n3745 & ~n3746 ;
  assign n3748 = n3747 ^ x85 ;
  assign n3752 = n3751 ^ n3748 ;
  assign n3753 = n3751 ^ x86 ;
  assign n3754 = n3752 & ~n3753 ;
  assign n3755 = n3754 ^ x86 ;
  assign n3759 = n3758 ^ n3755 ;
  assign n3760 = n3758 ^ x87 ;
  assign n3761 = n3759 & ~n3760 ;
  assign n3762 = n3761 ^ x87 ;
  assign n3766 = n3765 ^ n3762 ;
  assign n3767 = n3765 ^ x88 ;
  assign n3768 = n3766 & ~n3767 ;
  assign n3769 = n3768 ^ x88 ;
  assign n3773 = n3772 ^ n3769 ;
  assign n3774 = n3772 ^ x89 ;
  assign n3775 = n3773 & ~n3774 ;
  assign n3776 = n3775 ^ x89 ;
  assign n3780 = n3779 ^ n3776 ;
  assign n3781 = n3779 ^ x90 ;
  assign n3782 = n3780 & ~n3781 ;
  assign n3783 = n3782 ^ x90 ;
  assign n3787 = n3786 ^ n3783 ;
  assign n3788 = n3786 ^ x91 ;
  assign n3789 = n3787 & ~n3788 ;
  assign n3790 = n3789 ^ x91 ;
  assign n3802 = n3801 ^ n3790 ;
  assign n4056 = n3790 ^ x92 ;
  assign n3806 = n3802 & n4056 ;
  assign n3803 = x93 ^ x92 ;
  assign n3807 = n3806 ^ n3803 ;
  assign n3812 = n3811 ^ n3807 ;
  assign n3816 = n3812 ^ n3811 ;
  assign n3813 = n3812 ^ x93 ;
  assign n3815 = n3813 ^ n3577 ;
  assign n3817 = n3816 ^ n3815 ;
  assign n3820 = n3817 ^ n3816 ;
  assign n3821 = n3820 ^ n3813 ;
  assign n3822 = x94 & n3821 ;
  assign n3808 = n3807 ^ n3577 ;
  assign n3814 = n3813 ^ n3808 ;
  assign n3823 = n3822 ^ n3814 ;
  assign n3825 = n3813 ^ n3811 ;
  assign n3827 = n3812 & n3825 ;
  assign n3828 = n3827 ^ n3811 ;
  assign n3829 = ~n3823 & ~n3828 ;
  assign n3830 = n3829 ^ n3811 ;
  assign n3831 = n162 & n3830 ;
  assign n3832 = x94 & ~n3353 ;
  assign n3833 = n3831 & n3832 ;
  assign n3834 = n3833 ^ n3831 ;
  assign n3835 = n3577 & ~n3834 ;
  assign n3836 = n3835 ^ n375 ;
  assign n3837 = n3836 ^ x95 ;
  assign n3841 = n3836 ^ x94 ;
  assign n3838 = n3807 & n3834 ;
  assign n3839 = n3838 ^ n3811 ;
  assign n3840 = n3839 ^ n3836 ;
  assign n3842 = n3841 ^ n3840 ;
  assign n4057 = n3834 & n4056 ;
  assign n4058 = n4057 ^ n3801 ;
  assign n4049 = n3783 ^ x91 ;
  assign n4050 = n3834 & n4049 ;
  assign n4051 = n4050 ^ n3786 ;
  assign n4042 = n3776 ^ x90 ;
  assign n4043 = n3834 & n4042 ;
  assign n4044 = n4043 ^ n3779 ;
  assign n4035 = n3769 ^ x89 ;
  assign n4036 = n3834 & n4035 ;
  assign n4037 = n4036 ^ n3772 ;
  assign n4028 = n3762 ^ x88 ;
  assign n4029 = n3834 & n4028 ;
  assign n4030 = n4029 ^ n3765 ;
  assign n4021 = n3755 ^ x87 ;
  assign n4022 = n3834 & n4021 ;
  assign n4023 = n4022 ^ n3758 ;
  assign n4014 = n3748 ^ x86 ;
  assign n4015 = n3834 & n4014 ;
  assign n4016 = n4015 ^ n3751 ;
  assign n3843 = n3741 ^ x85 ;
  assign n3844 = n3834 & n3843 ;
  assign n3845 = n3844 ^ n3744 ;
  assign n3846 = n3845 ^ x86 ;
  assign n3859 = n3845 ^ x85 ;
  assign n3847 = n3589 ^ x84 ;
  assign n3848 = n3847 ^ x83 ;
  assign n3849 = n3848 ^ n3735 ;
  assign n3850 = n3849 ^ n3847 ;
  assign n3852 = x84 ^ x83 ;
  assign n3853 = n3852 ^ n3847 ;
  assign n3854 = ~n3850 & ~n3853 ;
  assign n3855 = n3854 ^ n3847 ;
  assign n3856 = n3834 & ~n3855 ;
  assign n3857 = n3856 ^ n3585 ;
  assign n3858 = n3857 ^ n3845 ;
  assign n3860 = n3859 ^ n3858 ;
  assign n4001 = n3735 ^ x83 ;
  assign n4002 = n3834 & n4001 ;
  assign n4003 = n4002 ^ n3589 ;
  assign n3994 = n3728 ^ x82 ;
  assign n3995 = n3834 & n3994 ;
  assign n3996 = n3995 ^ n3731 ;
  assign n3987 = n3721 ^ x81 ;
  assign n3988 = n3834 & n3987 ;
  assign n3989 = n3988 ^ n3724 ;
  assign n3980 = n3714 ^ x80 ;
  assign n3981 = n3834 & n3980 ;
  assign n3982 = n3981 ^ n3717 ;
  assign n3973 = n3707 ^ x79 ;
  assign n3974 = n3834 & n3973 ;
  assign n3975 = n3974 ^ n3710 ;
  assign n3966 = n3692 ^ x78 ;
  assign n3967 = n3834 & n3966 ;
  assign n3968 = n3967 ^ n3703 ;
  assign n3959 = n3685 ^ x77 ;
  assign n3960 = n3834 & n3959 ;
  assign n3961 = n3960 ^ n3688 ;
  assign n3952 = n3678 ^ x76 ;
  assign n3953 = n3834 & n3952 ;
  assign n3954 = n3953 ^ n3681 ;
  assign n3945 = n3671 ^ x75 ;
  assign n3946 = n3834 & n3945 ;
  assign n3947 = n3946 ^ n3674 ;
  assign n3938 = n3664 ^ x74 ;
  assign n3939 = n3834 & n3938 ;
  assign n3940 = n3939 ^ n3667 ;
  assign n3931 = n3657 ^ x73 ;
  assign n3932 = n3834 & n3931 ;
  assign n3933 = n3932 ^ n3660 ;
  assign n3924 = n3650 ^ x72 ;
  assign n3925 = n3834 & n3924 ;
  assign n3926 = n3925 ^ n3653 ;
  assign n3917 = n3643 ^ x71 ;
  assign n3918 = n3834 & n3917 ;
  assign n3919 = n3918 ^ n3646 ;
  assign n3910 = n3636 ^ x70 ;
  assign n3911 = n3834 & n3910 ;
  assign n3912 = n3911 ^ n3639 ;
  assign n3903 = n3629 ^ x69 ;
  assign n3904 = n3834 & n3903 ;
  assign n3905 = n3904 ^ n3632 ;
  assign n3896 = n3622 ^ x68 ;
  assign n3897 = n3834 & n3896 ;
  assign n3898 = n3897 ^ n3625 ;
  assign n3889 = n3615 ^ x67 ;
  assign n3890 = n3834 & n3889 ;
  assign n3891 = n3890 ^ n3618 ;
  assign n3882 = n3604 ^ x66 ;
  assign n3883 = n3834 & n3882 ;
  assign n3884 = n3883 ^ n3611 ;
  assign n3876 = x64 & n3583 ;
  assign n3872 = ~x33 & x64 ;
  assign n3873 = n3872 ^ x65 ;
  assign n3874 = n3834 & n3873 ;
  assign n3875 = n3874 ^ x34 ;
  assign n3877 = n3876 ^ n3875 ;
  assign n3867 = ~x32 & x64 ;
  assign n3868 = n3867 ^ x65 ;
  assign n3869 = x33 & n3868 ;
  assign n3862 = x64 & ~x65 ;
  assign n3861 = x64 & n3834 ;
  assign n3863 = n3862 ^ n3861 ;
  assign n3864 = n3862 ^ x32 ;
  assign n3865 = n3863 & n3864 ;
  assign n3866 = n3865 ^ x65 ;
  assign n3870 = n3869 ^ n3866 ;
  assign n3878 = n3877 ^ n3870 ;
  assign n3879 = n3877 ^ x66 ;
  assign n3880 = n3878 & ~n3879 ;
  assign n3881 = n3880 ^ x66 ;
  assign n3885 = n3884 ^ n3881 ;
  assign n3886 = n3884 ^ x67 ;
  assign n3887 = n3885 & ~n3886 ;
  assign n3888 = n3887 ^ x67 ;
  assign n3892 = n3891 ^ n3888 ;
  assign n3893 = n3891 ^ x68 ;
  assign n3894 = n3892 & ~n3893 ;
  assign n3895 = n3894 ^ x68 ;
  assign n3899 = n3898 ^ n3895 ;
  assign n3900 = n3898 ^ x69 ;
  assign n3901 = n3899 & ~n3900 ;
  assign n3902 = n3901 ^ x69 ;
  assign n3906 = n3905 ^ n3902 ;
  assign n3907 = n3905 ^ x70 ;
  assign n3908 = n3906 & ~n3907 ;
  assign n3909 = n3908 ^ x70 ;
  assign n3913 = n3912 ^ n3909 ;
  assign n3914 = n3912 ^ x71 ;
  assign n3915 = n3913 & ~n3914 ;
  assign n3916 = n3915 ^ x71 ;
  assign n3920 = n3919 ^ n3916 ;
  assign n3921 = n3919 ^ x72 ;
  assign n3922 = n3920 & ~n3921 ;
  assign n3923 = n3922 ^ x72 ;
  assign n3927 = n3926 ^ n3923 ;
  assign n3928 = n3926 ^ x73 ;
  assign n3929 = n3927 & ~n3928 ;
  assign n3930 = n3929 ^ x73 ;
  assign n3934 = n3933 ^ n3930 ;
  assign n3935 = n3933 ^ x74 ;
  assign n3936 = n3934 & ~n3935 ;
  assign n3937 = n3936 ^ x74 ;
  assign n3941 = n3940 ^ n3937 ;
  assign n3942 = n3940 ^ x75 ;
  assign n3943 = n3941 & ~n3942 ;
  assign n3944 = n3943 ^ x75 ;
  assign n3948 = n3947 ^ n3944 ;
  assign n3949 = n3947 ^ x76 ;
  assign n3950 = n3948 & ~n3949 ;
  assign n3951 = n3950 ^ x76 ;
  assign n3955 = n3954 ^ n3951 ;
  assign n3956 = n3954 ^ x77 ;
  assign n3957 = n3955 & ~n3956 ;
  assign n3958 = n3957 ^ x77 ;
  assign n3962 = n3961 ^ n3958 ;
  assign n3963 = n3961 ^ x78 ;
  assign n3964 = n3962 & ~n3963 ;
  assign n3965 = n3964 ^ x78 ;
  assign n3969 = n3968 ^ n3965 ;
  assign n3970 = n3968 ^ x79 ;
  assign n3971 = n3969 & ~n3970 ;
  assign n3972 = n3971 ^ x79 ;
  assign n3976 = n3975 ^ n3972 ;
  assign n3977 = n3975 ^ x80 ;
  assign n3978 = n3976 & ~n3977 ;
  assign n3979 = n3978 ^ x80 ;
  assign n3983 = n3982 ^ n3979 ;
  assign n3984 = n3982 ^ x81 ;
  assign n3985 = n3983 & ~n3984 ;
  assign n3986 = n3985 ^ x81 ;
  assign n3990 = n3989 ^ n3986 ;
  assign n3991 = n3989 ^ x82 ;
  assign n3992 = n3990 & ~n3991 ;
  assign n3993 = n3992 ^ x82 ;
  assign n3997 = n3996 ^ n3993 ;
  assign n3998 = n3996 ^ x83 ;
  assign n3999 = n3997 & ~n3998 ;
  assign n4000 = n3999 ^ x83 ;
  assign n4004 = n4003 ^ n4000 ;
  assign n4005 = n4003 ^ x84 ;
  assign n4006 = n4004 & ~n4005 ;
  assign n4007 = n4006 ^ x84 ;
  assign n4008 = n4007 ^ n3845 ;
  assign n4009 = n4008 ^ n3859 ;
  assign n4010 = ~n3860 & n4009 ;
  assign n4011 = n4010 ^ n3859 ;
  assign n4012 = ~n3846 & n4011 ;
  assign n4013 = n4012 ^ x86 ;
  assign n4017 = n4016 ^ n4013 ;
  assign n4018 = n4016 ^ x87 ;
  assign n4019 = n4017 & ~n4018 ;
  assign n4020 = n4019 ^ x87 ;
  assign n4024 = n4023 ^ n4020 ;
  assign n4025 = n4023 ^ x88 ;
  assign n4026 = n4024 & ~n4025 ;
  assign n4027 = n4026 ^ x88 ;
  assign n4031 = n4030 ^ n4027 ;
  assign n4032 = n4030 ^ x89 ;
  assign n4033 = n4031 & ~n4032 ;
  assign n4034 = n4033 ^ x89 ;
  assign n4038 = n4037 ^ n4034 ;
  assign n4039 = n4037 ^ x90 ;
  assign n4040 = n4038 & ~n4039 ;
  assign n4041 = n4040 ^ x90 ;
  assign n4045 = n4044 ^ n4041 ;
  assign n4046 = n4044 ^ x91 ;
  assign n4047 = n4045 & ~n4046 ;
  assign n4048 = n4047 ^ x91 ;
  assign n4052 = n4051 ^ n4048 ;
  assign n4053 = n4051 ^ x92 ;
  assign n4054 = n4052 & ~n4053 ;
  assign n4055 = n4054 ^ x92 ;
  assign n4059 = n4058 ^ n4055 ;
  assign n4060 = n4058 ^ x93 ;
  assign n4061 = n4059 & ~n4060 ;
  assign n4062 = n4061 ^ x93 ;
  assign n4063 = n4062 ^ n3836 ;
  assign n4064 = n4063 ^ n3841 ;
  assign n4065 = ~n3842 & n4064 ;
  assign n4066 = n4065 ^ n3841 ;
  assign n4067 = ~n3837 & n4066 ;
  assign n4068 = n4067 ^ x95 ;
  assign n4069 = n161 & ~n4068 ;
  assign n4070 = n3836 & ~n4069 ;
  assign n4071 = n4070 ^ n375 ;
  assign n4072 = x96 & n160 ;
  assign n4291 = n4055 ^ x93 ;
  assign n4292 = n4069 & n4291 ;
  assign n4293 = n4292 ^ n4058 ;
  assign n4284 = n4048 ^ x92 ;
  assign n4285 = n4069 & n4284 ;
  assign n4286 = n4285 ^ n4051 ;
  assign n4277 = n4041 ^ x91 ;
  assign n4278 = n4069 & n4277 ;
  assign n4279 = n4278 ^ n4044 ;
  assign n4270 = n4034 ^ x90 ;
  assign n4271 = n4069 & n4270 ;
  assign n4272 = n4271 ^ n4037 ;
  assign n4263 = n4027 ^ x89 ;
  assign n4264 = n4069 & n4263 ;
  assign n4265 = n4264 ^ n4030 ;
  assign n4256 = n4020 ^ x88 ;
  assign n4257 = n4069 & n4256 ;
  assign n4258 = n4257 ^ n4023 ;
  assign n4249 = n4013 ^ x87 ;
  assign n4250 = n4069 & n4249 ;
  assign n4251 = n4250 ^ n4016 ;
  assign n4234 = n3857 ^ x86 ;
  assign n4235 = n4234 ^ x85 ;
  assign n4236 = n4235 ^ n4007 ;
  assign n4237 = n4236 ^ n4234 ;
  assign n4239 = x86 ^ x85 ;
  assign n4240 = n4239 ^ n4234 ;
  assign n4241 = ~n4237 & ~n4240 ;
  assign n4242 = n4241 ^ n4234 ;
  assign n4243 = n4069 & ~n4242 ;
  assign n4244 = n4243 ^ n3845 ;
  assign n4227 = n4007 ^ x85 ;
  assign n4228 = n4069 & n4227 ;
  assign n4229 = n4228 ^ n3857 ;
  assign n4220 = n4000 ^ x84 ;
  assign n4221 = n4069 & n4220 ;
  assign n4222 = n4221 ^ n4003 ;
  assign n4213 = n3993 ^ x83 ;
  assign n4214 = n4069 & n4213 ;
  assign n4215 = n4214 ^ n3996 ;
  assign n4206 = n3986 ^ x82 ;
  assign n4207 = n4069 & n4206 ;
  assign n4208 = n4207 ^ n3989 ;
  assign n4199 = n3979 ^ x81 ;
  assign n4200 = n4069 & n4199 ;
  assign n4201 = n4200 ^ n3982 ;
  assign n4192 = n3972 ^ x80 ;
  assign n4193 = n4069 & n4192 ;
  assign n4194 = n4193 ^ n3975 ;
  assign n4073 = n3965 ^ x79 ;
  assign n4074 = n4069 & n4073 ;
  assign n4075 = n4074 ^ n3968 ;
  assign n4076 = n4075 ^ x80 ;
  assign n4081 = n4075 ^ x79 ;
  assign n4077 = n3958 ^ x78 ;
  assign n4078 = n4069 & n4077 ;
  assign n4079 = n4078 ^ n3961 ;
  assign n4080 = n4079 ^ n4075 ;
  assign n4082 = n4081 ^ n4080 ;
  assign n4179 = n3951 ^ x77 ;
  assign n4180 = n4069 & n4179 ;
  assign n4181 = n4180 ^ n3954 ;
  assign n4172 = n3944 ^ x76 ;
  assign n4173 = n4069 & n4172 ;
  assign n4174 = n4173 ^ n3947 ;
  assign n4165 = n3937 ^ x75 ;
  assign n4166 = n4069 & n4165 ;
  assign n4167 = n4166 ^ n3940 ;
  assign n4158 = n3930 ^ x74 ;
  assign n4159 = n4069 & n4158 ;
  assign n4160 = n4159 ^ n3933 ;
  assign n4151 = n3923 ^ x73 ;
  assign n4152 = n4069 & n4151 ;
  assign n4153 = n4152 ^ n3926 ;
  assign n4144 = n3916 ^ x72 ;
  assign n4145 = n4069 & n4144 ;
  assign n4146 = n4145 ^ n3919 ;
  assign n4137 = n3909 ^ x71 ;
  assign n4138 = n4069 & n4137 ;
  assign n4139 = n4138 ^ n3912 ;
  assign n4130 = n3902 ^ x70 ;
  assign n4131 = n4069 & n4130 ;
  assign n4132 = n4131 ^ n3905 ;
  assign n4123 = n3895 ^ x69 ;
  assign n4124 = n4069 & n4123 ;
  assign n4125 = n4124 ^ n3898 ;
  assign n4116 = n3888 ^ x68 ;
  assign n4117 = n4069 & n4116 ;
  assign n4118 = n4117 ^ n3891 ;
  assign n4093 = x65 ^ x31 ;
  assign n4094 = x64 ^ x32 ;
  assign n4095 = n4094 ^ x65 ;
  assign n4096 = n4095 ^ n4069 ;
  assign n4097 = ~n4093 & n4096 ;
  assign n4092 = x32 & x65 ;
  assign n4098 = n4097 ^ n4092 ;
  assign n4101 = x64 & n4098 ;
  assign n4102 = n4101 ^ n4092 ;
  assign n4103 = n4102 ^ x65 ;
  assign n4090 = n3868 & n4069 ;
  assign n4089 = n3861 ^ x33 ;
  assign n4091 = n4090 ^ n4089 ;
  assign n4104 = n4103 ^ n4091 ;
  assign n4105 = n4103 ^ x66 ;
  assign n4106 = n4104 & n4105 ;
  assign n4107 = n4106 ^ x66 ;
  assign n4086 = n3870 ^ x66 ;
  assign n4087 = n4069 & n4086 ;
  assign n4088 = n4087 ^ n3877 ;
  assign n4108 = n4107 ^ n4088 ;
  assign n4109 = n4107 ^ x67 ;
  assign n4110 = n4108 & n4109 ;
  assign n4111 = n4110 ^ x67 ;
  assign n4083 = n3881 ^ x67 ;
  assign n4084 = n4069 & n4083 ;
  assign n4085 = n4084 ^ n3884 ;
  assign n4112 = n4111 ^ n4085 ;
  assign n4113 = n4111 ^ x68 ;
  assign n4114 = n4112 & n4113 ;
  assign n4115 = n4114 ^ x68 ;
  assign n4119 = n4118 ^ n4115 ;
  assign n4120 = n4118 ^ x69 ;
  assign n4121 = n4119 & ~n4120 ;
  assign n4122 = n4121 ^ x69 ;
  assign n4126 = n4125 ^ n4122 ;
  assign n4127 = n4125 ^ x70 ;
  assign n4128 = n4126 & ~n4127 ;
  assign n4129 = n4128 ^ x70 ;
  assign n4133 = n4132 ^ n4129 ;
  assign n4134 = n4132 ^ x71 ;
  assign n4135 = n4133 & ~n4134 ;
  assign n4136 = n4135 ^ x71 ;
  assign n4140 = n4139 ^ n4136 ;
  assign n4141 = n4139 ^ x72 ;
  assign n4142 = n4140 & ~n4141 ;
  assign n4143 = n4142 ^ x72 ;
  assign n4147 = n4146 ^ n4143 ;
  assign n4148 = n4146 ^ x73 ;
  assign n4149 = n4147 & ~n4148 ;
  assign n4150 = n4149 ^ x73 ;
  assign n4154 = n4153 ^ n4150 ;
  assign n4155 = n4153 ^ x74 ;
  assign n4156 = n4154 & ~n4155 ;
  assign n4157 = n4156 ^ x74 ;
  assign n4161 = n4160 ^ n4157 ;
  assign n4162 = n4160 ^ x75 ;
  assign n4163 = n4161 & ~n4162 ;
  assign n4164 = n4163 ^ x75 ;
  assign n4168 = n4167 ^ n4164 ;
  assign n4169 = n4167 ^ x76 ;
  assign n4170 = n4168 & ~n4169 ;
  assign n4171 = n4170 ^ x76 ;
  assign n4175 = n4174 ^ n4171 ;
  assign n4176 = n4174 ^ x77 ;
  assign n4177 = n4175 & ~n4176 ;
  assign n4178 = n4177 ^ x77 ;
  assign n4182 = n4181 ^ n4178 ;
  assign n4183 = n4181 ^ x78 ;
  assign n4184 = n4182 & ~n4183 ;
  assign n4185 = n4184 ^ x78 ;
  assign n4186 = n4185 ^ n4075 ;
  assign n4187 = n4186 ^ n4081 ;
  assign n4188 = ~n4082 & n4187 ;
  assign n4189 = n4188 ^ n4081 ;
  assign n4190 = ~n4076 & n4189 ;
  assign n4191 = n4190 ^ x80 ;
  assign n4195 = n4194 ^ n4191 ;
  assign n4196 = n4194 ^ x81 ;
  assign n4197 = n4195 & ~n4196 ;
  assign n4198 = n4197 ^ x81 ;
  assign n4202 = n4201 ^ n4198 ;
  assign n4203 = n4201 ^ x82 ;
  assign n4204 = n4202 & ~n4203 ;
  assign n4205 = n4204 ^ x82 ;
  assign n4209 = n4208 ^ n4205 ;
  assign n4210 = n4208 ^ x83 ;
  assign n4211 = n4209 & ~n4210 ;
  assign n4212 = n4211 ^ x83 ;
  assign n4216 = n4215 ^ n4212 ;
  assign n4217 = n4215 ^ x84 ;
  assign n4218 = n4216 & ~n4217 ;
  assign n4219 = n4218 ^ x84 ;
  assign n4223 = n4222 ^ n4219 ;
  assign n4224 = n4222 ^ x85 ;
  assign n4225 = n4223 & ~n4224 ;
  assign n4226 = n4225 ^ x85 ;
  assign n4230 = n4229 ^ n4226 ;
  assign n4231 = n4229 ^ x86 ;
  assign n4232 = n4230 & ~n4231 ;
  assign n4233 = n4232 ^ x86 ;
  assign n4245 = n4244 ^ n4233 ;
  assign n4246 = n4244 ^ x87 ;
  assign n4247 = n4245 & ~n4246 ;
  assign n4248 = n4247 ^ x87 ;
  assign n4252 = n4251 ^ n4248 ;
  assign n4253 = n4251 ^ x88 ;
  assign n4254 = n4252 & ~n4253 ;
  assign n4255 = n4254 ^ x88 ;
  assign n4259 = n4258 ^ n4255 ;
  assign n4260 = n4258 ^ x89 ;
  assign n4261 = n4259 & ~n4260 ;
  assign n4262 = n4261 ^ x89 ;
  assign n4266 = n4265 ^ n4262 ;
  assign n4267 = n4265 ^ x90 ;
  assign n4268 = n4266 & ~n4267 ;
  assign n4269 = n4268 ^ x90 ;
  assign n4273 = n4272 ^ n4269 ;
  assign n4274 = n4272 ^ x91 ;
  assign n4275 = n4273 & ~n4274 ;
  assign n4276 = n4275 ^ x91 ;
  assign n4280 = n4279 ^ n4276 ;
  assign n4281 = n4279 ^ x92 ;
  assign n4282 = n4280 & ~n4281 ;
  assign n4283 = n4282 ^ x92 ;
  assign n4287 = n4286 ^ n4283 ;
  assign n4288 = n4286 ^ x93 ;
  assign n4289 = n4287 & ~n4288 ;
  assign n4290 = n4289 ^ x93 ;
  assign n4294 = n4293 ^ n4290 ;
  assign n4295 = n4293 ^ x94 ;
  assign n4296 = n4294 & ~n4295 ;
  assign n4297 = n4296 ^ x94 ;
  assign n4298 = n4297 ^ x95 ;
  assign n4299 = n4062 ^ x94 ;
  assign n4300 = n4069 & n4299 ;
  assign n4301 = n4300 ^ n3839 ;
  assign n4302 = n4301 ^ x95 ;
  assign n4303 = n4298 & ~n4302 ;
  assign n4304 = n4303 ^ x95 ;
  assign n4305 = n4072 & n4304 ;
  assign n4306 = n4305 ^ n160 ;
  assign n4307 = n4071 & ~n4306 ;
  assign n4308 = x97 & ~n4071 ;
  assign n4309 = n159 & ~n4308 ;
  assign n4311 = n4308 ^ x97 ;
  assign n4310 = n4307 ^ n375 ;
  assign n4312 = n4311 ^ n4310 ;
  assign n4313 = x96 & ~n4071 ;
  assign n4314 = n160 & ~n4313 ;
  assign n4315 = n4071 ^ x96 ;
  assign n4316 = n4315 ^ n4313 ;
  assign n4317 = x95 & ~n4316 ;
  assign n4318 = ~n4301 & n4317 ;
  assign n4319 = n4314 & ~n4318 ;
  assign n4320 = n4297 & ~n4316 ;
  assign n4321 = ~x95 & n4301 ;
  assign n4322 = n4320 & n4321 ;
  assign n4323 = n4322 ^ n4320 ;
  assign n4324 = n4319 & ~n4323 ;
  assign n4325 = n4298 & n4324 ;
  assign n4326 = n4325 ^ n4301 ;
  assign n4327 = n4326 ^ x96 ;
  assign n4555 = n4290 ^ x94 ;
  assign n4556 = n4324 & n4555 ;
  assign n4557 = n4556 ^ n4293 ;
  assign n4548 = n4283 ^ x93 ;
  assign n4549 = n4324 & n4548 ;
  assign n4550 = n4549 ^ n4286 ;
  assign n4541 = n4276 ^ x92 ;
  assign n4542 = n4324 & n4541 ;
  assign n4543 = n4542 ^ n4279 ;
  assign n4534 = n4269 ^ x91 ;
  assign n4535 = n4324 & n4534 ;
  assign n4536 = n4535 ^ n4272 ;
  assign n4527 = n4262 ^ x90 ;
  assign n4528 = n4324 & n4527 ;
  assign n4529 = n4528 ^ n4265 ;
  assign n4520 = n4255 ^ x89 ;
  assign n4521 = n4324 & n4520 ;
  assign n4522 = n4521 ^ n4258 ;
  assign n4513 = n4248 ^ x88 ;
  assign n4514 = n4324 & n4513 ;
  assign n4515 = n4514 ^ n4251 ;
  assign n4506 = n4233 ^ x87 ;
  assign n4507 = n4324 & n4506 ;
  assign n4508 = n4507 ^ n4244 ;
  assign n4499 = n4226 ^ x86 ;
  assign n4500 = n4324 & n4499 ;
  assign n4501 = n4500 ^ n4229 ;
  assign n4492 = n4219 ^ x85 ;
  assign n4493 = n4324 & n4492 ;
  assign n4494 = n4493 ^ n4222 ;
  assign n4485 = n4212 ^ x84 ;
  assign n4486 = n4324 & n4485 ;
  assign n4487 = n4486 ^ n4215 ;
  assign n4478 = n4205 ^ x83 ;
  assign n4479 = n4324 & n4478 ;
  assign n4480 = n4479 ^ n4208 ;
  assign n4471 = n4198 ^ x82 ;
  assign n4472 = n4324 & n4471 ;
  assign n4473 = n4472 ^ n4201 ;
  assign n4464 = n4191 ^ x81 ;
  assign n4465 = n4324 & n4464 ;
  assign n4466 = n4465 ^ n4194 ;
  assign n4449 = n4079 ^ x80 ;
  assign n4450 = n4449 ^ x79 ;
  assign n4451 = n4450 ^ n4185 ;
  assign n4452 = n4451 ^ n4449 ;
  assign n4454 = x80 ^ x79 ;
  assign n4455 = n4454 ^ n4449 ;
  assign n4456 = ~n4452 & ~n4455 ;
  assign n4457 = n4456 ^ n4449 ;
  assign n4458 = n4324 & ~n4457 ;
  assign n4459 = n4458 ^ n4075 ;
  assign n4442 = n4185 ^ x79 ;
  assign n4443 = n4324 & n4442 ;
  assign n4444 = n4443 ^ n4079 ;
  assign n4435 = n4178 ^ x78 ;
  assign n4436 = n4324 & n4435 ;
  assign n4437 = n4436 ^ n4181 ;
  assign n4428 = n4171 ^ x77 ;
  assign n4429 = n4324 & n4428 ;
  assign n4430 = n4429 ^ n4174 ;
  assign n4421 = n4164 ^ x76 ;
  assign n4422 = n4324 & n4421 ;
  assign n4423 = n4422 ^ n4167 ;
  assign n4414 = n4157 ^ x75 ;
  assign n4415 = n4324 & n4414 ;
  assign n4416 = n4415 ^ n4160 ;
  assign n4407 = n4150 ^ x74 ;
  assign n4408 = n4324 & n4407 ;
  assign n4409 = n4408 ^ n4153 ;
  assign n4400 = n4143 ^ x73 ;
  assign n4401 = n4324 & n4400 ;
  assign n4402 = n4401 ^ n4146 ;
  assign n4393 = n4136 ^ x72 ;
  assign n4394 = n4324 & n4393 ;
  assign n4395 = n4394 ^ n4139 ;
  assign n4386 = n4129 ^ x71 ;
  assign n4387 = n4324 & n4386 ;
  assign n4388 = n4387 ^ n4132 ;
  assign n4379 = n4122 ^ x70 ;
  assign n4380 = n4324 & n4379 ;
  assign n4381 = n4380 ^ n4125 ;
  assign n4372 = n4115 ^ x69 ;
  assign n4373 = n4324 & n4372 ;
  assign n4374 = n4373 ^ n4118 ;
  assign n4366 = n4113 & n4324 ;
  assign n4367 = n4366 ^ n4085 ;
  assign n4360 = n4109 & n4324 ;
  assign n4361 = n4360 ^ n4088 ;
  assign n4354 = n4105 & n4324 ;
  assign n4355 = n4354 ^ n4091 ;
  assign n4331 = n4069 ^ x31 ;
  assign n4332 = n4331 ^ n4069 ;
  assign n4333 = n4324 & ~n4332 ;
  assign n4334 = n4333 ^ n4069 ;
  assign n4335 = x64 & n4334 ;
  assign n4336 = n4335 ^ x32 ;
  assign n4328 = x65 & n4324 ;
  assign n4337 = n4336 ^ n4328 ;
  assign n4338 = n4337 ^ x66 ;
  assign n4346 = x31 & x65 ;
  assign n4343 = x65 ^ x30 ;
  assign n4339 = x64 ^ x31 ;
  assign n4340 = n4339 ^ x65 ;
  assign n4344 = n4340 ^ n4324 ;
  assign n4345 = ~n4343 & n4344 ;
  assign n4347 = n4346 ^ n4345 ;
  assign n4348 = x64 & n4347 ;
  assign n4349 = n4348 ^ n4346 ;
  assign n4350 = n4349 ^ x65 ;
  assign n4351 = n4350 ^ n4337 ;
  assign n4352 = ~n4338 & n4351 ;
  assign n4353 = n4352 ^ x66 ;
  assign n4356 = n4355 ^ n4353 ;
  assign n4357 = n4355 ^ x67 ;
  assign n4358 = n4356 & ~n4357 ;
  assign n4359 = n4358 ^ x67 ;
  assign n4362 = n4361 ^ n4359 ;
  assign n4363 = n4361 ^ x68 ;
  assign n4364 = n4362 & ~n4363 ;
  assign n4365 = n4364 ^ x68 ;
  assign n4368 = n4367 ^ n4365 ;
  assign n4369 = n4367 ^ x69 ;
  assign n4370 = n4368 & ~n4369 ;
  assign n4371 = n4370 ^ x69 ;
  assign n4375 = n4374 ^ n4371 ;
  assign n4376 = n4374 ^ x70 ;
  assign n4377 = n4375 & ~n4376 ;
  assign n4378 = n4377 ^ x70 ;
  assign n4382 = n4381 ^ n4378 ;
  assign n4383 = n4381 ^ x71 ;
  assign n4384 = n4382 & ~n4383 ;
  assign n4385 = n4384 ^ x71 ;
  assign n4389 = n4388 ^ n4385 ;
  assign n4390 = n4388 ^ x72 ;
  assign n4391 = n4389 & ~n4390 ;
  assign n4392 = n4391 ^ x72 ;
  assign n4396 = n4395 ^ n4392 ;
  assign n4397 = n4395 ^ x73 ;
  assign n4398 = n4396 & ~n4397 ;
  assign n4399 = n4398 ^ x73 ;
  assign n4403 = n4402 ^ n4399 ;
  assign n4404 = n4402 ^ x74 ;
  assign n4405 = n4403 & ~n4404 ;
  assign n4406 = n4405 ^ x74 ;
  assign n4410 = n4409 ^ n4406 ;
  assign n4411 = n4409 ^ x75 ;
  assign n4412 = n4410 & ~n4411 ;
  assign n4413 = n4412 ^ x75 ;
  assign n4417 = n4416 ^ n4413 ;
  assign n4418 = n4416 ^ x76 ;
  assign n4419 = n4417 & ~n4418 ;
  assign n4420 = n4419 ^ x76 ;
  assign n4424 = n4423 ^ n4420 ;
  assign n4425 = n4423 ^ x77 ;
  assign n4426 = n4424 & ~n4425 ;
  assign n4427 = n4426 ^ x77 ;
  assign n4431 = n4430 ^ n4427 ;
  assign n4432 = n4430 ^ x78 ;
  assign n4433 = n4431 & ~n4432 ;
  assign n4434 = n4433 ^ x78 ;
  assign n4438 = n4437 ^ n4434 ;
  assign n4439 = n4437 ^ x79 ;
  assign n4440 = n4438 & ~n4439 ;
  assign n4441 = n4440 ^ x79 ;
  assign n4445 = n4444 ^ n4441 ;
  assign n4446 = n4444 ^ x80 ;
  assign n4447 = n4445 & ~n4446 ;
  assign n4448 = n4447 ^ x80 ;
  assign n4460 = n4459 ^ n4448 ;
  assign n4461 = n4459 ^ x81 ;
  assign n4462 = n4460 & ~n4461 ;
  assign n4463 = n4462 ^ x81 ;
  assign n4467 = n4466 ^ n4463 ;
  assign n4468 = n4466 ^ x82 ;
  assign n4469 = n4467 & ~n4468 ;
  assign n4470 = n4469 ^ x82 ;
  assign n4474 = n4473 ^ n4470 ;
  assign n4475 = n4473 ^ x83 ;
  assign n4476 = n4474 & ~n4475 ;
  assign n4477 = n4476 ^ x83 ;
  assign n4481 = n4480 ^ n4477 ;
  assign n4482 = n4480 ^ x84 ;
  assign n4483 = n4481 & ~n4482 ;
  assign n4484 = n4483 ^ x84 ;
  assign n4488 = n4487 ^ n4484 ;
  assign n4489 = n4487 ^ x85 ;
  assign n4490 = n4488 & ~n4489 ;
  assign n4491 = n4490 ^ x85 ;
  assign n4495 = n4494 ^ n4491 ;
  assign n4496 = n4494 ^ x86 ;
  assign n4497 = n4495 & ~n4496 ;
  assign n4498 = n4497 ^ x86 ;
  assign n4502 = n4501 ^ n4498 ;
  assign n4503 = n4501 ^ x87 ;
  assign n4504 = n4502 & ~n4503 ;
  assign n4505 = n4504 ^ x87 ;
  assign n4509 = n4508 ^ n4505 ;
  assign n4510 = n4508 ^ x88 ;
  assign n4511 = n4509 & ~n4510 ;
  assign n4512 = n4511 ^ x88 ;
  assign n4516 = n4515 ^ n4512 ;
  assign n4517 = n4515 ^ x89 ;
  assign n4518 = n4516 & ~n4517 ;
  assign n4519 = n4518 ^ x89 ;
  assign n4523 = n4522 ^ n4519 ;
  assign n4524 = n4522 ^ x90 ;
  assign n4525 = n4523 & ~n4524 ;
  assign n4526 = n4525 ^ x90 ;
  assign n4530 = n4529 ^ n4526 ;
  assign n4531 = n4529 ^ x91 ;
  assign n4532 = n4530 & ~n4531 ;
  assign n4533 = n4532 ^ x91 ;
  assign n4537 = n4536 ^ n4533 ;
  assign n4538 = n4536 ^ x92 ;
  assign n4539 = n4537 & ~n4538 ;
  assign n4540 = n4539 ^ x92 ;
  assign n4544 = n4543 ^ n4540 ;
  assign n4545 = n4543 ^ x93 ;
  assign n4546 = n4544 & ~n4545 ;
  assign n4547 = n4546 ^ x93 ;
  assign n4551 = n4550 ^ n4547 ;
  assign n4552 = n4550 ^ x94 ;
  assign n4553 = n4551 & ~n4552 ;
  assign n4554 = n4553 ^ x94 ;
  assign n4558 = n4557 ^ n4554 ;
  assign n4801 = n4554 ^ x95 ;
  assign n4562 = n4558 & n4801 ;
  assign n4559 = x96 ^ x95 ;
  assign n4563 = n4562 ^ n4559 ;
  assign n4566 = ~n4327 & n4563 ;
  assign n4567 = n4566 ^ x96 ;
  assign n4568 = ~n4312 & n4567 ;
  assign n4569 = n4309 & ~n4568 ;
  assign n4570 = n4307 & ~n4569 ;
  assign n4572 = n4310 ^ x98 ;
  assign n4571 = ~x98 & n4310 ;
  assign n4573 = n4572 ^ n4571 ;
  assign n4574 = n158 & ~n4573 ;
  assign n4814 = n4568 ^ n375 ;
  assign n4808 = n4563 & n4569 ;
  assign n4809 = n4808 ^ n4326 ;
  assign n4802 = n4569 & n4801 ;
  assign n4803 = n4802 ^ n4557 ;
  assign n4794 = n4547 ^ x94 ;
  assign n4795 = n4569 & n4794 ;
  assign n4796 = n4795 ^ n4550 ;
  assign n4787 = n4540 ^ x93 ;
  assign n4788 = n4569 & n4787 ;
  assign n4789 = n4788 ^ n4543 ;
  assign n4780 = n4533 ^ x92 ;
  assign n4781 = n4569 & n4780 ;
  assign n4782 = n4781 ^ n4536 ;
  assign n4773 = n4526 ^ x91 ;
  assign n4774 = n4569 & n4773 ;
  assign n4775 = n4774 ^ n4529 ;
  assign n4766 = n4519 ^ x90 ;
  assign n4767 = n4569 & n4766 ;
  assign n4768 = n4767 ^ n4522 ;
  assign n4759 = n4512 ^ x89 ;
  assign n4760 = n4569 & n4759 ;
  assign n4761 = n4760 ^ n4515 ;
  assign n4752 = n4505 ^ x88 ;
  assign n4753 = n4569 & n4752 ;
  assign n4754 = n4753 ^ n4508 ;
  assign n4745 = n4498 ^ x87 ;
  assign n4746 = n4569 & n4745 ;
  assign n4747 = n4746 ^ n4501 ;
  assign n4738 = n4491 ^ x86 ;
  assign n4739 = n4569 & n4738 ;
  assign n4740 = n4739 ^ n4494 ;
  assign n4731 = n4484 ^ x85 ;
  assign n4732 = n4569 & n4731 ;
  assign n4733 = n4732 ^ n4487 ;
  assign n4724 = n4477 ^ x84 ;
  assign n4725 = n4569 & n4724 ;
  assign n4726 = n4725 ^ n4480 ;
  assign n4717 = n4470 ^ x83 ;
  assign n4718 = n4569 & n4717 ;
  assign n4719 = n4718 ^ n4473 ;
  assign n4710 = n4463 ^ x82 ;
  assign n4711 = n4569 & n4710 ;
  assign n4712 = n4711 ^ n4466 ;
  assign n4703 = n4448 ^ x81 ;
  assign n4704 = n4569 & n4703 ;
  assign n4705 = n4704 ^ n4459 ;
  assign n4696 = n4441 ^ x80 ;
  assign n4697 = n4569 & n4696 ;
  assign n4698 = n4697 ^ n4444 ;
  assign n4689 = n4434 ^ x79 ;
  assign n4690 = n4569 & n4689 ;
  assign n4691 = n4690 ^ n4437 ;
  assign n4682 = n4427 ^ x78 ;
  assign n4683 = n4569 & n4682 ;
  assign n4684 = n4683 ^ n4430 ;
  assign n4675 = n4420 ^ x77 ;
  assign n4676 = n4569 & n4675 ;
  assign n4677 = n4676 ^ n4423 ;
  assign n4668 = n4413 ^ x76 ;
  assign n4669 = n4569 & n4668 ;
  assign n4670 = n4669 ^ n4416 ;
  assign n4661 = n4406 ^ x75 ;
  assign n4662 = n4569 & n4661 ;
  assign n4663 = n4662 ^ n4409 ;
  assign n4654 = n4399 ^ x74 ;
  assign n4655 = n4569 & n4654 ;
  assign n4656 = n4655 ^ n4402 ;
  assign n4647 = n4392 ^ x73 ;
  assign n4648 = n4569 & n4647 ;
  assign n4649 = n4648 ^ n4395 ;
  assign n4640 = n4385 ^ x72 ;
  assign n4641 = n4569 & n4640 ;
  assign n4642 = n4641 ^ n4388 ;
  assign n4633 = n4378 ^ x71 ;
  assign n4634 = n4569 & n4633 ;
  assign n4635 = n4634 ^ n4381 ;
  assign n4626 = n4371 ^ x70 ;
  assign n4627 = n4569 & n4626 ;
  assign n4628 = n4627 ^ n4374 ;
  assign n4619 = n4365 ^ x69 ;
  assign n4620 = n4569 & n4619 ;
  assign n4621 = n4620 ^ n4367 ;
  assign n4575 = n4359 ^ x68 ;
  assign n4576 = n4569 & n4575 ;
  assign n4577 = n4576 ^ n4361 ;
  assign n4578 = n4577 ^ x69 ;
  assign n4579 = n4353 ^ x67 ;
  assign n4580 = n4569 & n4579 ;
  assign n4581 = n4580 ^ n4355 ;
  assign n4582 = n4581 ^ x68 ;
  assign n4606 = n4350 ^ x66 ;
  assign n4607 = n4569 & n4606 ;
  assign n4608 = n4607 ^ n4337 ;
  assign n4600 = x64 & n4324 ;
  assign n4596 = ~x30 & x64 ;
  assign n4597 = n4596 ^ x65 ;
  assign n4598 = n4569 & n4597 ;
  assign n4599 = n4598 ^ x31 ;
  assign n4601 = n4600 ^ n4599 ;
  assign n4590 = x30 & x65 ;
  assign n4587 = x65 ^ x29 ;
  assign n4583 = x64 ^ x30 ;
  assign n4584 = n4583 ^ x65 ;
  assign n4588 = n4584 ^ n4569 ;
  assign n4589 = ~n4587 & n4588 ;
  assign n4591 = n4590 ^ n4589 ;
  assign n4592 = x64 & n4591 ;
  assign n4593 = n4592 ^ n4590 ;
  assign n4594 = n4593 ^ x65 ;
  assign n4602 = n4601 ^ n4594 ;
  assign n4603 = n4601 ^ x66 ;
  assign n4604 = n4602 & ~n4603 ;
  assign n4605 = n4604 ^ x66 ;
  assign n4609 = n4608 ^ n4605 ;
  assign n4610 = n4608 ^ x67 ;
  assign n4611 = n4609 & ~n4610 ;
  assign n4612 = n4611 ^ x67 ;
  assign n4613 = n4612 ^ n4581 ;
  assign n4614 = ~n4582 & n4613 ;
  assign n4615 = n4614 ^ x68 ;
  assign n4616 = n4615 ^ n4577 ;
  assign n4617 = ~n4578 & n4616 ;
  assign n4618 = n4617 ^ x69 ;
  assign n4622 = n4621 ^ n4618 ;
  assign n4623 = n4621 ^ x70 ;
  assign n4624 = n4622 & ~n4623 ;
  assign n4625 = n4624 ^ x70 ;
  assign n4629 = n4628 ^ n4625 ;
  assign n4630 = n4628 ^ x71 ;
  assign n4631 = n4629 & ~n4630 ;
  assign n4632 = n4631 ^ x71 ;
  assign n4636 = n4635 ^ n4632 ;
  assign n4637 = n4635 ^ x72 ;
  assign n4638 = n4636 & ~n4637 ;
  assign n4639 = n4638 ^ x72 ;
  assign n4643 = n4642 ^ n4639 ;
  assign n4644 = n4642 ^ x73 ;
  assign n4645 = n4643 & ~n4644 ;
  assign n4646 = n4645 ^ x73 ;
  assign n4650 = n4649 ^ n4646 ;
  assign n4651 = n4649 ^ x74 ;
  assign n4652 = n4650 & ~n4651 ;
  assign n4653 = n4652 ^ x74 ;
  assign n4657 = n4656 ^ n4653 ;
  assign n4658 = n4656 ^ x75 ;
  assign n4659 = n4657 & ~n4658 ;
  assign n4660 = n4659 ^ x75 ;
  assign n4664 = n4663 ^ n4660 ;
  assign n4665 = n4663 ^ x76 ;
  assign n4666 = n4664 & ~n4665 ;
  assign n4667 = n4666 ^ x76 ;
  assign n4671 = n4670 ^ n4667 ;
  assign n4672 = n4670 ^ x77 ;
  assign n4673 = n4671 & ~n4672 ;
  assign n4674 = n4673 ^ x77 ;
  assign n4678 = n4677 ^ n4674 ;
  assign n4679 = n4677 ^ x78 ;
  assign n4680 = n4678 & ~n4679 ;
  assign n4681 = n4680 ^ x78 ;
  assign n4685 = n4684 ^ n4681 ;
  assign n4686 = n4684 ^ x79 ;
  assign n4687 = n4685 & ~n4686 ;
  assign n4688 = n4687 ^ x79 ;
  assign n4692 = n4691 ^ n4688 ;
  assign n4693 = n4691 ^ x80 ;
  assign n4694 = n4692 & ~n4693 ;
  assign n4695 = n4694 ^ x80 ;
  assign n4699 = n4698 ^ n4695 ;
  assign n4700 = n4698 ^ x81 ;
  assign n4701 = n4699 & ~n4700 ;
  assign n4702 = n4701 ^ x81 ;
  assign n4706 = n4705 ^ n4702 ;
  assign n4707 = n4705 ^ x82 ;
  assign n4708 = n4706 & ~n4707 ;
  assign n4709 = n4708 ^ x82 ;
  assign n4713 = n4712 ^ n4709 ;
  assign n4714 = n4712 ^ x83 ;
  assign n4715 = n4713 & ~n4714 ;
  assign n4716 = n4715 ^ x83 ;
  assign n4720 = n4719 ^ n4716 ;
  assign n4721 = n4719 ^ x84 ;
  assign n4722 = n4720 & ~n4721 ;
  assign n4723 = n4722 ^ x84 ;
  assign n4727 = n4726 ^ n4723 ;
  assign n4728 = n4726 ^ x85 ;
  assign n4729 = n4727 & ~n4728 ;
  assign n4730 = n4729 ^ x85 ;
  assign n4734 = n4733 ^ n4730 ;
  assign n4735 = n4733 ^ x86 ;
  assign n4736 = n4734 & ~n4735 ;
  assign n4737 = n4736 ^ x86 ;
  assign n4741 = n4740 ^ n4737 ;
  assign n4742 = n4740 ^ x87 ;
  assign n4743 = n4741 & ~n4742 ;
  assign n4744 = n4743 ^ x87 ;
  assign n4748 = n4747 ^ n4744 ;
  assign n4749 = n4747 ^ x88 ;
  assign n4750 = n4748 & ~n4749 ;
  assign n4751 = n4750 ^ x88 ;
  assign n4755 = n4754 ^ n4751 ;
  assign n4756 = n4754 ^ x89 ;
  assign n4757 = n4755 & ~n4756 ;
  assign n4758 = n4757 ^ x89 ;
  assign n4762 = n4761 ^ n4758 ;
  assign n4763 = n4761 ^ x90 ;
  assign n4764 = n4762 & ~n4763 ;
  assign n4765 = n4764 ^ x90 ;
  assign n4769 = n4768 ^ n4765 ;
  assign n4770 = n4768 ^ x91 ;
  assign n4771 = n4769 & ~n4770 ;
  assign n4772 = n4771 ^ x91 ;
  assign n4776 = n4775 ^ n4772 ;
  assign n4777 = n4775 ^ x92 ;
  assign n4778 = n4776 & ~n4777 ;
  assign n4779 = n4778 ^ x92 ;
  assign n4783 = n4782 ^ n4779 ;
  assign n4784 = n4782 ^ x93 ;
  assign n4785 = n4783 & ~n4784 ;
  assign n4786 = n4785 ^ x93 ;
  assign n4790 = n4789 ^ n4786 ;
  assign n4791 = n4789 ^ x94 ;
  assign n4792 = n4790 & ~n4791 ;
  assign n4793 = n4792 ^ x94 ;
  assign n4797 = n4796 ^ n4793 ;
  assign n4798 = n4796 ^ x95 ;
  assign n4799 = n4797 & ~n4798 ;
  assign n4800 = n4799 ^ x95 ;
  assign n4804 = n4803 ^ n4800 ;
  assign n4805 = n4803 ^ x96 ;
  assign n4806 = n4804 & ~n4805 ;
  assign n4807 = n4806 ^ x96 ;
  assign n4810 = n4809 ^ n4807 ;
  assign n4811 = n4809 ^ x97 ;
  assign n4812 = n4810 & ~n4811 ;
  assign n4813 = n4812 ^ x97 ;
  assign n4815 = n4571 & n4813 ;
  assign n4816 = n4814 & n4815 ;
  assign n4817 = n4816 ^ n4813 ;
  assign n4818 = n4574 & ~n4817 ;
  assign n4819 = n4570 & ~n4818 ;
  assign n4820 = n4819 ^ n375 ;
  assign n4821 = n4820 ^ x99 ;
  assign n5059 = n4807 ^ x97 ;
  assign n5060 = n4818 & n5059 ;
  assign n5061 = n5060 ^ n4809 ;
  assign n5063 = n5061 ^ x97 ;
  assign n5052 = n4793 ^ x95 ;
  assign n5053 = n4818 & n5052 ;
  assign n5054 = n5053 ^ n4796 ;
  assign n5045 = n4786 ^ x94 ;
  assign n5046 = n4818 & n5045 ;
  assign n5047 = n5046 ^ n4789 ;
  assign n4822 = n4779 ^ x93 ;
  assign n4823 = n4818 & n4822 ;
  assign n4824 = n4823 ^ n4782 ;
  assign n4825 = n4824 ^ x94 ;
  assign n4830 = n4824 ^ x93 ;
  assign n4826 = n4772 ^ x92 ;
  assign n4827 = n4818 & n4826 ;
  assign n4828 = n4827 ^ n4775 ;
  assign n4829 = n4828 ^ n4824 ;
  assign n4831 = n4830 ^ n4829 ;
  assign n5032 = n4765 ^ x91 ;
  assign n5033 = n4818 & n5032 ;
  assign n5034 = n5033 ^ n4768 ;
  assign n5025 = n4758 ^ x90 ;
  assign n5026 = n4818 & n5025 ;
  assign n5027 = n5026 ^ n4761 ;
  assign n5018 = n4751 ^ x89 ;
  assign n5019 = n4818 & n5018 ;
  assign n5020 = n5019 ^ n4754 ;
  assign n5011 = n4744 ^ x88 ;
  assign n5012 = n4818 & n5011 ;
  assign n5013 = n5012 ^ n4747 ;
  assign n5004 = n4737 ^ x87 ;
  assign n5005 = n4818 & n5004 ;
  assign n5006 = n5005 ^ n4740 ;
  assign n4997 = n4730 ^ x86 ;
  assign n4998 = n4818 & n4997 ;
  assign n4999 = n4998 ^ n4733 ;
  assign n4990 = n4723 ^ x85 ;
  assign n4991 = n4818 & n4990 ;
  assign n4992 = n4991 ^ n4726 ;
  assign n4983 = n4716 ^ x84 ;
  assign n4984 = n4818 & n4983 ;
  assign n4985 = n4984 ^ n4719 ;
  assign n4976 = n4709 ^ x83 ;
  assign n4977 = n4818 & n4976 ;
  assign n4978 = n4977 ^ n4712 ;
  assign n4969 = n4702 ^ x82 ;
  assign n4970 = n4818 & n4969 ;
  assign n4971 = n4970 ^ n4705 ;
  assign n4962 = n4695 ^ x81 ;
  assign n4963 = n4818 & n4962 ;
  assign n4964 = n4963 ^ n4698 ;
  assign n4955 = n4688 ^ x80 ;
  assign n4956 = n4818 & n4955 ;
  assign n4957 = n4956 ^ n4691 ;
  assign n4948 = n4681 ^ x79 ;
  assign n4949 = n4818 & n4948 ;
  assign n4950 = n4949 ^ n4684 ;
  assign n4941 = n4674 ^ x78 ;
  assign n4942 = n4818 & n4941 ;
  assign n4943 = n4942 ^ n4677 ;
  assign n4934 = n4667 ^ x77 ;
  assign n4935 = n4818 & n4934 ;
  assign n4936 = n4935 ^ n4670 ;
  assign n4927 = n4660 ^ x76 ;
  assign n4928 = n4818 & n4927 ;
  assign n4929 = n4928 ^ n4663 ;
  assign n4920 = n4653 ^ x75 ;
  assign n4921 = n4818 & n4920 ;
  assign n4922 = n4921 ^ n4656 ;
  assign n4913 = n4646 ^ x74 ;
  assign n4914 = n4818 & n4913 ;
  assign n4915 = n4914 ^ n4649 ;
  assign n4906 = n4639 ^ x73 ;
  assign n4907 = n4818 & n4906 ;
  assign n4908 = n4907 ^ n4642 ;
  assign n4899 = n4632 ^ x72 ;
  assign n4900 = n4818 & n4899 ;
  assign n4901 = n4900 ^ n4635 ;
  assign n4892 = n4625 ^ x71 ;
  assign n4893 = n4818 & n4892 ;
  assign n4894 = n4893 ^ n4628 ;
  assign n4885 = n4618 ^ x70 ;
  assign n4886 = n4818 & n4885 ;
  assign n4887 = n4886 ^ n4621 ;
  assign n4832 = n4615 ^ x69 ;
  assign n4833 = n4818 & n4832 ;
  assign n4834 = n4833 ^ n4577 ;
  assign n4835 = n4834 ^ x70 ;
  assign n4840 = n4834 ^ x69 ;
  assign n4836 = n4612 ^ x68 ;
  assign n4837 = n4818 & n4836 ;
  assign n4838 = n4837 ^ n4581 ;
  assign n4839 = n4838 ^ n4834 ;
  assign n4841 = n4840 ^ n4839 ;
  assign n4872 = n4605 ^ x67 ;
  assign n4873 = n4818 & n4872 ;
  assign n4874 = n4873 ^ n4608 ;
  assign n4865 = n4594 ^ x66 ;
  assign n4866 = n4818 & n4865 ;
  assign n4867 = n4866 ^ n4601 ;
  assign n4859 = x64 & n4569 ;
  assign n4855 = ~x29 & x64 ;
  assign n4856 = n4855 ^ x65 ;
  assign n4857 = n4818 & n4856 ;
  assign n4858 = n4857 ^ x30 ;
  assign n4860 = n4859 ^ n4858 ;
  assign n4849 = x29 & x65 ;
  assign n4846 = x65 ^ x28 ;
  assign n4842 = x64 ^ x29 ;
  assign n4843 = n4842 ^ x65 ;
  assign n4847 = n4843 ^ n4818 ;
  assign n4848 = ~n4846 & n4847 ;
  assign n4850 = n4849 ^ n4848 ;
  assign n4851 = x64 & n4850 ;
  assign n4852 = n4851 ^ n4849 ;
  assign n4853 = n4852 ^ x65 ;
  assign n4861 = n4860 ^ n4853 ;
  assign n4862 = n4860 ^ x66 ;
  assign n4863 = n4861 & ~n4862 ;
  assign n4864 = n4863 ^ x66 ;
  assign n4868 = n4867 ^ n4864 ;
  assign n4869 = n4867 ^ x67 ;
  assign n4870 = n4868 & ~n4869 ;
  assign n4871 = n4870 ^ x67 ;
  assign n4875 = n4874 ^ n4871 ;
  assign n4876 = n4874 ^ x68 ;
  assign n4877 = n4875 & ~n4876 ;
  assign n4878 = n4877 ^ x68 ;
  assign n4879 = n4878 ^ n4834 ;
  assign n4880 = n4879 ^ n4840 ;
  assign n4881 = ~n4841 & n4880 ;
  assign n4882 = n4881 ^ n4840 ;
  assign n4883 = ~n4835 & n4882 ;
  assign n4884 = n4883 ^ x70 ;
  assign n4888 = n4887 ^ n4884 ;
  assign n4889 = n4887 ^ x71 ;
  assign n4890 = n4888 & ~n4889 ;
  assign n4891 = n4890 ^ x71 ;
  assign n4895 = n4894 ^ n4891 ;
  assign n4896 = n4894 ^ x72 ;
  assign n4897 = n4895 & ~n4896 ;
  assign n4898 = n4897 ^ x72 ;
  assign n4902 = n4901 ^ n4898 ;
  assign n4903 = n4901 ^ x73 ;
  assign n4904 = n4902 & ~n4903 ;
  assign n4905 = n4904 ^ x73 ;
  assign n4909 = n4908 ^ n4905 ;
  assign n4910 = n4908 ^ x74 ;
  assign n4911 = n4909 & ~n4910 ;
  assign n4912 = n4911 ^ x74 ;
  assign n4916 = n4915 ^ n4912 ;
  assign n4917 = n4915 ^ x75 ;
  assign n4918 = n4916 & ~n4917 ;
  assign n4919 = n4918 ^ x75 ;
  assign n4923 = n4922 ^ n4919 ;
  assign n4924 = n4922 ^ x76 ;
  assign n4925 = n4923 & ~n4924 ;
  assign n4926 = n4925 ^ x76 ;
  assign n4930 = n4929 ^ n4926 ;
  assign n4931 = n4929 ^ x77 ;
  assign n4932 = n4930 & ~n4931 ;
  assign n4933 = n4932 ^ x77 ;
  assign n4937 = n4936 ^ n4933 ;
  assign n4938 = n4936 ^ x78 ;
  assign n4939 = n4937 & ~n4938 ;
  assign n4940 = n4939 ^ x78 ;
  assign n4944 = n4943 ^ n4940 ;
  assign n4945 = n4943 ^ x79 ;
  assign n4946 = n4944 & ~n4945 ;
  assign n4947 = n4946 ^ x79 ;
  assign n4951 = n4950 ^ n4947 ;
  assign n4952 = n4950 ^ x80 ;
  assign n4953 = n4951 & ~n4952 ;
  assign n4954 = n4953 ^ x80 ;
  assign n4958 = n4957 ^ n4954 ;
  assign n4959 = n4957 ^ x81 ;
  assign n4960 = n4958 & ~n4959 ;
  assign n4961 = n4960 ^ x81 ;
  assign n4965 = n4964 ^ n4961 ;
  assign n4966 = n4964 ^ x82 ;
  assign n4967 = n4965 & ~n4966 ;
  assign n4968 = n4967 ^ x82 ;
  assign n4972 = n4971 ^ n4968 ;
  assign n4973 = n4971 ^ x83 ;
  assign n4974 = n4972 & ~n4973 ;
  assign n4975 = n4974 ^ x83 ;
  assign n4979 = n4978 ^ n4975 ;
  assign n4980 = n4978 ^ x84 ;
  assign n4981 = n4979 & ~n4980 ;
  assign n4982 = n4981 ^ x84 ;
  assign n4986 = n4985 ^ n4982 ;
  assign n4987 = n4985 ^ x85 ;
  assign n4988 = n4986 & ~n4987 ;
  assign n4989 = n4988 ^ x85 ;
  assign n4993 = n4992 ^ n4989 ;
  assign n4994 = n4992 ^ x86 ;
  assign n4995 = n4993 & ~n4994 ;
  assign n4996 = n4995 ^ x86 ;
  assign n5000 = n4999 ^ n4996 ;
  assign n5001 = n4999 ^ x87 ;
  assign n5002 = n5000 & ~n5001 ;
  assign n5003 = n5002 ^ x87 ;
  assign n5007 = n5006 ^ n5003 ;
  assign n5008 = n5006 ^ x88 ;
  assign n5009 = n5007 & ~n5008 ;
  assign n5010 = n5009 ^ x88 ;
  assign n5014 = n5013 ^ n5010 ;
  assign n5015 = n5013 ^ x89 ;
  assign n5016 = n5014 & ~n5015 ;
  assign n5017 = n5016 ^ x89 ;
  assign n5021 = n5020 ^ n5017 ;
  assign n5022 = n5020 ^ x90 ;
  assign n5023 = n5021 & ~n5022 ;
  assign n5024 = n5023 ^ x90 ;
  assign n5028 = n5027 ^ n5024 ;
  assign n5029 = n5027 ^ x91 ;
  assign n5030 = n5028 & ~n5029 ;
  assign n5031 = n5030 ^ x91 ;
  assign n5035 = n5034 ^ n5031 ;
  assign n5036 = n5034 ^ x92 ;
  assign n5037 = n5035 & ~n5036 ;
  assign n5038 = n5037 ^ x92 ;
  assign n5039 = n5038 ^ n4824 ;
  assign n5040 = n5039 ^ n4830 ;
  assign n5041 = ~n4831 & n5040 ;
  assign n5042 = n5041 ^ n4830 ;
  assign n5043 = ~n4825 & n5042 ;
  assign n5044 = n5043 ^ x94 ;
  assign n5048 = n5047 ^ n5044 ;
  assign n5049 = n5047 ^ x95 ;
  assign n5050 = n5048 & ~n5049 ;
  assign n5051 = n5050 ^ x95 ;
  assign n5055 = n5054 ^ n5051 ;
  assign n5056 = n5054 ^ x96 ;
  assign n5057 = n5055 & ~n5056 ;
  assign n5058 = n5057 ^ x96 ;
  assign n5062 = n5061 ^ n5058 ;
  assign n5064 = n5063 ^ n5062 ;
  assign n5065 = n4800 ^ x96 ;
  assign n5066 = n4818 & n5065 ;
  assign n5067 = n5066 ^ n4803 ;
  assign n5068 = n5067 ^ n5061 ;
  assign n5069 = n5068 ^ n5063 ;
  assign n5070 = n5064 & ~n5069 ;
  assign n5071 = n5070 ^ n5063 ;
  assign n5073 = n4820 ^ x98 ;
  assign n5072 = n5061 ^ n4820 ;
  assign n5074 = n5073 ^ n5072 ;
  assign n5075 = n5071 & ~n5074 ;
  assign n5076 = n5075 ^ n5073 ;
  assign n5077 = ~n4821 & n5076 ;
  assign n5078 = n5077 ^ x99 ;
  assign n5079 = n157 & ~n5078 ;
  assign n5080 = n4820 & ~n5079 ;
  assign n5352 = n5067 ^ x98 ;
  assign n5353 = n5352 ^ x97 ;
  assign n5354 = n5353 ^ n5058 ;
  assign n5355 = n5354 ^ n5352 ;
  assign n5357 = x98 ^ x97 ;
  assign n5358 = n5357 ^ n5352 ;
  assign n5359 = ~n5355 & ~n5358 ;
  assign n5360 = n5359 ^ n5352 ;
  assign n5361 = n5079 & ~n5360 ;
  assign n5362 = n5361 ^ n5061 ;
  assign n5345 = n5058 ^ x97 ;
  assign n5346 = n5079 & n5345 ;
  assign n5347 = n5346 ^ n5067 ;
  assign n5338 = n5051 ^ x96 ;
  assign n5339 = n5079 & n5338 ;
  assign n5340 = n5339 ^ n5054 ;
  assign n5331 = n5044 ^ x95 ;
  assign n5332 = n5079 & n5331 ;
  assign n5333 = n5332 ^ n5047 ;
  assign n5316 = n4828 ^ x94 ;
  assign n5317 = n5316 ^ x93 ;
  assign n5318 = n5317 ^ n5038 ;
  assign n5319 = n5318 ^ n5316 ;
  assign n5321 = x94 ^ x93 ;
  assign n5322 = n5321 ^ n5316 ;
  assign n5323 = ~n5319 & ~n5322 ;
  assign n5324 = n5323 ^ n5316 ;
  assign n5325 = n5079 & ~n5324 ;
  assign n5326 = n5325 ^ n4824 ;
  assign n5309 = n5038 ^ x93 ;
  assign n5310 = n5079 & n5309 ;
  assign n5311 = n5310 ^ n4828 ;
  assign n5081 = n5031 ^ x92 ;
  assign n5082 = n5079 & n5081 ;
  assign n5083 = n5082 ^ n5034 ;
  assign n5084 = n5083 ^ x93 ;
  assign n5089 = n5083 ^ x92 ;
  assign n5085 = n5024 ^ x91 ;
  assign n5086 = n5079 & n5085 ;
  assign n5087 = n5086 ^ n5027 ;
  assign n5088 = n5087 ^ n5083 ;
  assign n5090 = n5089 ^ n5088 ;
  assign n5296 = n5017 ^ x90 ;
  assign n5297 = n5079 & n5296 ;
  assign n5298 = n5297 ^ n5020 ;
  assign n5289 = n5010 ^ x89 ;
  assign n5290 = n5079 & n5289 ;
  assign n5291 = n5290 ^ n5013 ;
  assign n5282 = n5003 ^ x88 ;
  assign n5283 = n5079 & n5282 ;
  assign n5284 = n5283 ^ n5006 ;
  assign n5091 = n4996 ^ x87 ;
  assign n5092 = n5079 & n5091 ;
  assign n5093 = n5092 ^ n4999 ;
  assign n5094 = n5093 ^ x88 ;
  assign n5099 = n5093 ^ x87 ;
  assign n5095 = n4989 ^ x86 ;
  assign n5096 = n5079 & n5095 ;
  assign n5097 = n5096 ^ n4992 ;
  assign n5098 = n5097 ^ n5093 ;
  assign n5100 = n5099 ^ n5098 ;
  assign n5269 = n4982 ^ x85 ;
  assign n5270 = n5079 & n5269 ;
  assign n5271 = n5270 ^ n4985 ;
  assign n5262 = n4975 ^ x84 ;
  assign n5263 = n5079 & n5262 ;
  assign n5264 = n5263 ^ n4978 ;
  assign n5101 = n4968 ^ x83 ;
  assign n5102 = n5079 & n5101 ;
  assign n5103 = n5102 ^ n4971 ;
  assign n5104 = n5103 ^ x84 ;
  assign n5109 = n5103 ^ x83 ;
  assign n5105 = n4961 ^ x82 ;
  assign n5106 = n5079 & n5105 ;
  assign n5107 = n5106 ^ n4964 ;
  assign n5108 = n5107 ^ n5103 ;
  assign n5110 = n5109 ^ n5108 ;
  assign n5111 = n4954 ^ x81 ;
  assign n5112 = n5079 & n5111 ;
  assign n5113 = n5112 ^ n4957 ;
  assign n5114 = n5113 ^ x82 ;
  assign n5119 = n5113 ^ x81 ;
  assign n5115 = n4947 ^ x80 ;
  assign n5116 = n5079 & n5115 ;
  assign n5117 = n5116 ^ n4950 ;
  assign n5118 = n5117 ^ n5113 ;
  assign n5120 = n5119 ^ n5118 ;
  assign n5243 = n4940 ^ x79 ;
  assign n5244 = n5079 & n5243 ;
  assign n5245 = n5244 ^ n4943 ;
  assign n5236 = n4933 ^ x78 ;
  assign n5237 = n5079 & n5236 ;
  assign n5238 = n5237 ^ n4936 ;
  assign n5121 = n4926 ^ x77 ;
  assign n5122 = n5079 & n5121 ;
  assign n5123 = n5122 ^ n4929 ;
  assign n5124 = n5123 ^ x78 ;
  assign n5125 = n4919 ^ x76 ;
  assign n5126 = n5079 & n5125 ;
  assign n5127 = n5126 ^ n4922 ;
  assign n5128 = n5127 ^ x77 ;
  assign n5223 = n4912 ^ x75 ;
  assign n5224 = n5079 & n5223 ;
  assign n5225 = n5224 ^ n4915 ;
  assign n5216 = n4905 ^ x74 ;
  assign n5217 = n5079 & n5216 ;
  assign n5218 = n5217 ^ n4908 ;
  assign n5209 = n4898 ^ x73 ;
  assign n5210 = n5079 & n5209 ;
  assign n5211 = n5210 ^ n4901 ;
  assign n5202 = n4891 ^ x72 ;
  assign n5203 = n5079 & n5202 ;
  assign n5204 = n5203 ^ n4894 ;
  assign n5195 = n4884 ^ x71 ;
  assign n5196 = n5079 & n5195 ;
  assign n5197 = n5196 ^ n4887 ;
  assign n5180 = n4838 ^ x70 ;
  assign n5181 = n5180 ^ x69 ;
  assign n5182 = n5181 ^ n4878 ;
  assign n5183 = n5182 ^ n5180 ;
  assign n5185 = x70 ^ x69 ;
  assign n5186 = n5185 ^ n5180 ;
  assign n5187 = ~n5183 & ~n5186 ;
  assign n5188 = n5187 ^ n5180 ;
  assign n5189 = n5079 & ~n5188 ;
  assign n5190 = n5189 ^ n4834 ;
  assign n5173 = n4878 ^ x69 ;
  assign n5174 = n5079 & n5173 ;
  assign n5175 = n5174 ^ n4838 ;
  assign n5166 = n4871 ^ x68 ;
  assign n5167 = n5079 & n5166 ;
  assign n5168 = n5167 ^ n4874 ;
  assign n5159 = n4864 ^ x67 ;
  assign n5160 = n5079 & n5159 ;
  assign n5161 = n5160 ^ n4867 ;
  assign n5152 = n4853 ^ x66 ;
  assign n5153 = n5079 & n5152 ;
  assign n5154 = n5153 ^ n4860 ;
  assign n5146 = x64 & n4818 ;
  assign n5142 = ~x28 & x64 ;
  assign n5143 = n5142 ^ x65 ;
  assign n5144 = n5079 & n5143 ;
  assign n5145 = n5144 ^ x29 ;
  assign n5147 = n5146 ^ n5145 ;
  assign n5130 = x65 ^ x27 ;
  assign n5131 = x64 ^ x28 ;
  assign n5132 = n5131 ^ x65 ;
  assign n5133 = n5132 ^ n5079 ;
  assign n5134 = ~n5130 & n5133 ;
  assign n5129 = x28 & x65 ;
  assign n5135 = n5134 ^ n5129 ;
  assign n5138 = x64 & n5135 ;
  assign n5139 = n5138 ^ n5129 ;
  assign n5140 = n5139 ^ x65 ;
  assign n5148 = n5147 ^ n5140 ;
  assign n5149 = n5147 ^ x66 ;
  assign n5150 = n5148 & ~n5149 ;
  assign n5151 = n5150 ^ x66 ;
  assign n5155 = n5154 ^ n5151 ;
  assign n5156 = n5154 ^ x67 ;
  assign n5157 = n5155 & ~n5156 ;
  assign n5158 = n5157 ^ x67 ;
  assign n5162 = n5161 ^ n5158 ;
  assign n5163 = n5161 ^ x68 ;
  assign n5164 = n5162 & ~n5163 ;
  assign n5165 = n5164 ^ x68 ;
  assign n5169 = n5168 ^ n5165 ;
  assign n5170 = n5168 ^ x69 ;
  assign n5171 = n5169 & ~n5170 ;
  assign n5172 = n5171 ^ x69 ;
  assign n5176 = n5175 ^ n5172 ;
  assign n5177 = n5175 ^ x70 ;
  assign n5178 = n5176 & ~n5177 ;
  assign n5179 = n5178 ^ x70 ;
  assign n5191 = n5190 ^ n5179 ;
  assign n5192 = n5190 ^ x71 ;
  assign n5193 = n5191 & ~n5192 ;
  assign n5194 = n5193 ^ x71 ;
  assign n5198 = n5197 ^ n5194 ;
  assign n5199 = n5197 ^ x72 ;
  assign n5200 = n5198 & ~n5199 ;
  assign n5201 = n5200 ^ x72 ;
  assign n5205 = n5204 ^ n5201 ;
  assign n5206 = n5204 ^ x73 ;
  assign n5207 = n5205 & ~n5206 ;
  assign n5208 = n5207 ^ x73 ;
  assign n5212 = n5211 ^ n5208 ;
  assign n5213 = n5211 ^ x74 ;
  assign n5214 = n5212 & ~n5213 ;
  assign n5215 = n5214 ^ x74 ;
  assign n5219 = n5218 ^ n5215 ;
  assign n5220 = n5218 ^ x75 ;
  assign n5221 = n5219 & ~n5220 ;
  assign n5222 = n5221 ^ x75 ;
  assign n5226 = n5225 ^ n5222 ;
  assign n5227 = n5225 ^ x76 ;
  assign n5228 = n5226 & ~n5227 ;
  assign n5229 = n5228 ^ x76 ;
  assign n5230 = n5229 ^ n5127 ;
  assign n5231 = ~n5128 & n5230 ;
  assign n5232 = n5231 ^ x77 ;
  assign n5233 = n5232 ^ n5123 ;
  assign n5234 = ~n5124 & n5233 ;
  assign n5235 = n5234 ^ x78 ;
  assign n5239 = n5238 ^ n5235 ;
  assign n5240 = n5238 ^ x79 ;
  assign n5241 = n5239 & ~n5240 ;
  assign n5242 = n5241 ^ x79 ;
  assign n5246 = n5245 ^ n5242 ;
  assign n5247 = n5245 ^ x80 ;
  assign n5248 = n5246 & ~n5247 ;
  assign n5249 = n5248 ^ x80 ;
  assign n5250 = n5249 ^ n5113 ;
  assign n5251 = n5250 ^ n5119 ;
  assign n5252 = ~n5120 & n5251 ;
  assign n5253 = n5252 ^ n5119 ;
  assign n5254 = ~n5114 & n5253 ;
  assign n5255 = n5254 ^ x82 ;
  assign n5256 = n5255 ^ n5103 ;
  assign n5257 = n5256 ^ n5109 ;
  assign n5258 = ~n5110 & n5257 ;
  assign n5259 = n5258 ^ n5109 ;
  assign n5260 = ~n5104 & n5259 ;
  assign n5261 = n5260 ^ x84 ;
  assign n5265 = n5264 ^ n5261 ;
  assign n5266 = n5264 ^ x85 ;
  assign n5267 = n5265 & ~n5266 ;
  assign n5268 = n5267 ^ x85 ;
  assign n5272 = n5271 ^ n5268 ;
  assign n5273 = n5271 ^ x86 ;
  assign n5274 = n5272 & ~n5273 ;
  assign n5275 = n5274 ^ x86 ;
  assign n5276 = n5275 ^ n5093 ;
  assign n5277 = n5276 ^ n5099 ;
  assign n5278 = ~n5100 & n5277 ;
  assign n5279 = n5278 ^ n5099 ;
  assign n5280 = ~n5094 & n5279 ;
  assign n5281 = n5280 ^ x88 ;
  assign n5285 = n5284 ^ n5281 ;
  assign n5286 = n5284 ^ x89 ;
  assign n5287 = n5285 & ~n5286 ;
  assign n5288 = n5287 ^ x89 ;
  assign n5292 = n5291 ^ n5288 ;
  assign n5293 = n5291 ^ x90 ;
  assign n5294 = n5292 & ~n5293 ;
  assign n5295 = n5294 ^ x90 ;
  assign n5299 = n5298 ^ n5295 ;
  assign n5300 = n5298 ^ x91 ;
  assign n5301 = n5299 & ~n5300 ;
  assign n5302 = n5301 ^ x91 ;
  assign n5303 = n5302 ^ n5083 ;
  assign n5304 = n5303 ^ n5089 ;
  assign n5305 = ~n5090 & n5304 ;
  assign n5306 = n5305 ^ n5089 ;
  assign n5307 = ~n5084 & n5306 ;
  assign n5308 = n5307 ^ x93 ;
  assign n5312 = n5311 ^ n5308 ;
  assign n5313 = n5311 ^ x94 ;
  assign n5314 = n5312 & ~n5313 ;
  assign n5315 = n5314 ^ x94 ;
  assign n5327 = n5326 ^ n5315 ;
  assign n5328 = n5326 ^ x95 ;
  assign n5329 = n5327 & ~n5328 ;
  assign n5330 = n5329 ^ x95 ;
  assign n5334 = n5333 ^ n5330 ;
  assign n5335 = n5333 ^ x96 ;
  assign n5336 = n5334 & ~n5335 ;
  assign n5337 = n5336 ^ x96 ;
  assign n5341 = n5340 ^ n5337 ;
  assign n5342 = n5340 ^ x97 ;
  assign n5343 = n5341 & ~n5342 ;
  assign n5344 = n5343 ^ x97 ;
  assign n5348 = n5347 ^ n5344 ;
  assign n5349 = n5347 ^ x98 ;
  assign n5350 = n5348 & ~n5349 ;
  assign n5351 = n5350 ^ x98 ;
  assign n5363 = n5362 ^ n5351 ;
  assign n5614 = n5351 ^ x99 ;
  assign n5367 = n5363 & n5614 ;
  assign n5364 = x100 ^ x99 ;
  assign n5368 = n5367 ^ n5364 ;
  assign n5373 = ~n375 & ~n5080 ;
  assign n5374 = n5373 ^ x100 ;
  assign n5375 = n5368 & n5374 ;
  assign n5376 = n5375 ^ x100 ;
  assign n5377 = n156 & ~n5376 ;
  assign n5378 = n5080 & ~n5377 ;
  assign n5379 = ~n155 & n5378 ;
  assign n5610 = n5378 ^ n375 ;
  assign n5612 = x101 & ~n5610 ;
  assign n5613 = n155 & ~n5612 ;
  assign n5615 = n5377 & n5614 ;
  assign n5616 = n5615 ^ n5362 ;
  assign n5617 = n5610 ^ x101 ;
  assign n5618 = n5617 ^ n5612 ;
  assign n5619 = ~n5616 & ~n5618 ;
  assign n5620 = x100 & n5619 ;
  assign n5621 = n5613 & ~n5620 ;
  assign n5680 = n5344 ^ x98 ;
  assign n5681 = n5377 & n5680 ;
  assign n5682 = n5681 ^ n5347 ;
  assign n5673 = n5337 ^ x97 ;
  assign n5674 = n5377 & n5673 ;
  assign n5675 = n5674 ^ n5340 ;
  assign n5622 = n5330 ^ x96 ;
  assign n5623 = n5377 & n5622 ;
  assign n5624 = n5623 ^ n5333 ;
  assign n5625 = n5624 ^ x97 ;
  assign n5630 = n5624 ^ x96 ;
  assign n5626 = n5315 ^ x95 ;
  assign n5627 = n5377 & n5626 ;
  assign n5628 = n5627 ^ n5326 ;
  assign n5629 = n5628 ^ n5624 ;
  assign n5631 = n5630 ^ n5629 ;
  assign n5660 = n5308 ^ x94 ;
  assign n5661 = n5377 & n5660 ;
  assign n5662 = n5661 ^ n5311 ;
  assign n5632 = n5087 ^ x93 ;
  assign n5633 = n5632 ^ x92 ;
  assign n5634 = n5633 ^ n5302 ;
  assign n5635 = n5634 ^ n5632 ;
  assign n5638 = n5632 ^ n3803 ;
  assign n5639 = ~n5635 & ~n5638 ;
  assign n5640 = n5639 ^ n5632 ;
  assign n5641 = n5377 & ~n5640 ;
  assign n5642 = n5641 ^ n5083 ;
  assign n5643 = n5642 ^ x94 ;
  assign n5644 = n5302 ^ x92 ;
  assign n5645 = n5377 & n5644 ;
  assign n5646 = n5645 ^ n5087 ;
  assign n5647 = n5646 ^ x93 ;
  assign n5602 = n5288 ^ x90 ;
  assign n5603 = n5377 & n5602 ;
  assign n5604 = n5603 ^ n5291 ;
  assign n5380 = n5281 ^ x89 ;
  assign n5381 = n5377 & n5380 ;
  assign n5382 = n5381 ^ n5284 ;
  assign n5383 = n5382 ^ x90 ;
  assign n5396 = n5382 ^ x89 ;
  assign n5384 = n5097 ^ x88 ;
  assign n5385 = n5384 ^ x87 ;
  assign n5386 = n5385 ^ n5275 ;
  assign n5387 = n5386 ^ n5384 ;
  assign n5390 = n5384 ^ n3553 ;
  assign n5391 = ~n5387 & ~n5390 ;
  assign n5392 = n5391 ^ n5384 ;
  assign n5393 = n5377 & ~n5392 ;
  assign n5394 = n5393 ^ n5093 ;
  assign n5395 = n5394 ^ n5382 ;
  assign n5397 = n5396 ^ n5395 ;
  assign n5589 = n5275 ^ x87 ;
  assign n5590 = n5377 & n5589 ;
  assign n5591 = n5590 ^ n5097 ;
  assign n5582 = n5268 ^ x86 ;
  assign n5583 = n5377 & n5582 ;
  assign n5584 = n5583 ^ n5271 ;
  assign n5575 = n5261 ^ x85 ;
  assign n5576 = n5377 & n5575 ;
  assign n5577 = n5576 ^ n5264 ;
  assign n5560 = n5107 ^ x84 ;
  assign n5561 = n5560 ^ x83 ;
  assign n5562 = n5561 ^ n5255 ;
  assign n5563 = n5562 ^ n5560 ;
  assign n5566 = n5560 ^ n3852 ;
  assign n5567 = ~n5563 & ~n5566 ;
  assign n5568 = n5567 ^ n5560 ;
  assign n5569 = n5377 & ~n5568 ;
  assign n5570 = n5569 ^ n5103 ;
  assign n5553 = n5255 ^ x83 ;
  assign n5554 = n5377 & n5553 ;
  assign n5555 = n5554 ^ n5107 ;
  assign n5538 = n5117 ^ x82 ;
  assign n5539 = n5538 ^ x81 ;
  assign n5540 = n5539 ^ n5249 ;
  assign n5541 = n5540 ^ n5538 ;
  assign n5543 = x82 ^ x81 ;
  assign n5544 = n5543 ^ n5538 ;
  assign n5545 = ~n5541 & ~n5544 ;
  assign n5546 = n5545 ^ n5538 ;
  assign n5547 = n5377 & ~n5546 ;
  assign n5548 = n5547 ^ n5113 ;
  assign n5531 = n5249 ^ x81 ;
  assign n5532 = n5377 & n5531 ;
  assign n5533 = n5532 ^ n5117 ;
  assign n5524 = n5242 ^ x80 ;
  assign n5525 = n5377 & n5524 ;
  assign n5526 = n5525 ^ n5245 ;
  assign n5517 = n5235 ^ x79 ;
  assign n5518 = n5377 & n5517 ;
  assign n5519 = n5518 ^ n5238 ;
  assign n5510 = n5232 ^ x78 ;
  assign n5511 = n5377 & n5510 ;
  assign n5512 = n5511 ^ n5123 ;
  assign n5398 = n5229 ^ x77 ;
  assign n5399 = n5377 & n5398 ;
  assign n5400 = n5399 ^ n5127 ;
  assign n5401 = n5400 ^ x78 ;
  assign n5406 = n5400 ^ x77 ;
  assign n5402 = n5222 ^ x76 ;
  assign n5403 = n5377 & n5402 ;
  assign n5404 = n5403 ^ n5225 ;
  assign n5405 = n5404 ^ n5400 ;
  assign n5407 = n5406 ^ n5405 ;
  assign n5497 = n5215 ^ x75 ;
  assign n5498 = n5377 & n5497 ;
  assign n5499 = n5498 ^ n5218 ;
  assign n5490 = n5208 ^ x74 ;
  assign n5491 = n5377 & n5490 ;
  assign n5492 = n5491 ^ n5211 ;
  assign n5483 = n5201 ^ x73 ;
  assign n5484 = n5377 & n5483 ;
  assign n5485 = n5484 ^ n5204 ;
  assign n5476 = n5194 ^ x72 ;
  assign n5477 = n5377 & n5476 ;
  assign n5478 = n5477 ^ n5197 ;
  assign n5469 = n5179 ^ x71 ;
  assign n5470 = n5377 & n5469 ;
  assign n5471 = n5470 ^ n5190 ;
  assign n5462 = n5172 ^ x70 ;
  assign n5463 = n5377 & n5462 ;
  assign n5464 = n5463 ^ n5175 ;
  assign n5455 = n5165 ^ x69 ;
  assign n5456 = n5377 & n5455 ;
  assign n5457 = n5456 ^ n5168 ;
  assign n5448 = n5158 ^ x68 ;
  assign n5449 = n5377 & n5448 ;
  assign n5450 = n5449 ^ n5161 ;
  assign n5441 = n5151 ^ x67 ;
  assign n5442 = n5377 & n5441 ;
  assign n5443 = n5442 ^ n5154 ;
  assign n5434 = n5140 ^ x66 ;
  assign n5435 = n5377 & n5434 ;
  assign n5436 = n5435 ^ n5147 ;
  assign n5416 = x65 & n5377 ;
  assign n5410 = n5079 ^ x27 ;
  assign n5411 = n5410 ^ n5079 ;
  assign n5412 = n5377 & ~n5411 ;
  assign n5413 = n5412 ^ n5079 ;
  assign n5414 = x64 & n5413 ;
  assign n5415 = n5414 ^ x28 ;
  assign n5417 = n5416 ^ n5415 ;
  assign n5418 = n5417 ^ x66 ;
  assign n5420 = x65 ^ x26 ;
  assign n5421 = x64 ^ x27 ;
  assign n5422 = n5421 ^ x65 ;
  assign n5423 = n5422 ^ n5377 ;
  assign n5424 = ~n5420 & n5423 ;
  assign n5419 = x27 & x65 ;
  assign n5425 = n5424 ^ n5419 ;
  assign n5428 = x64 & n5425 ;
  assign n5429 = n5428 ^ n5419 ;
  assign n5430 = n5429 ^ x65 ;
  assign n5431 = n5430 ^ n5417 ;
  assign n5432 = ~n5418 & n5431 ;
  assign n5433 = n5432 ^ x66 ;
  assign n5437 = n5436 ^ n5433 ;
  assign n5438 = n5436 ^ x67 ;
  assign n5439 = n5437 & ~n5438 ;
  assign n5440 = n5439 ^ x67 ;
  assign n5444 = n5443 ^ n5440 ;
  assign n5445 = n5443 ^ x68 ;
  assign n5446 = n5444 & ~n5445 ;
  assign n5447 = n5446 ^ x68 ;
  assign n5451 = n5450 ^ n5447 ;
  assign n5452 = n5450 ^ x69 ;
  assign n5453 = n5451 & ~n5452 ;
  assign n5454 = n5453 ^ x69 ;
  assign n5458 = n5457 ^ n5454 ;
  assign n5459 = n5457 ^ x70 ;
  assign n5460 = n5458 & ~n5459 ;
  assign n5461 = n5460 ^ x70 ;
  assign n5465 = n5464 ^ n5461 ;
  assign n5466 = n5464 ^ x71 ;
  assign n5467 = n5465 & ~n5466 ;
  assign n5468 = n5467 ^ x71 ;
  assign n5472 = n5471 ^ n5468 ;
  assign n5473 = n5471 ^ x72 ;
  assign n5474 = n5472 & ~n5473 ;
  assign n5475 = n5474 ^ x72 ;
  assign n5479 = n5478 ^ n5475 ;
  assign n5480 = n5478 ^ x73 ;
  assign n5481 = n5479 & ~n5480 ;
  assign n5482 = n5481 ^ x73 ;
  assign n5486 = n5485 ^ n5482 ;
  assign n5487 = n5485 ^ x74 ;
  assign n5488 = n5486 & ~n5487 ;
  assign n5489 = n5488 ^ x74 ;
  assign n5493 = n5492 ^ n5489 ;
  assign n5494 = n5492 ^ x75 ;
  assign n5495 = n5493 & ~n5494 ;
  assign n5496 = n5495 ^ x75 ;
  assign n5500 = n5499 ^ n5496 ;
  assign n5501 = n5499 ^ x76 ;
  assign n5502 = n5500 & ~n5501 ;
  assign n5503 = n5502 ^ x76 ;
  assign n5504 = n5503 ^ n5400 ;
  assign n5505 = n5504 ^ n5406 ;
  assign n5506 = ~n5407 & n5505 ;
  assign n5507 = n5506 ^ n5406 ;
  assign n5508 = ~n5401 & n5507 ;
  assign n5509 = n5508 ^ x78 ;
  assign n5513 = n5512 ^ n5509 ;
  assign n5514 = n5512 ^ x79 ;
  assign n5515 = n5513 & ~n5514 ;
  assign n5516 = n5515 ^ x79 ;
  assign n5520 = n5519 ^ n5516 ;
  assign n5521 = n5519 ^ x80 ;
  assign n5522 = n5520 & ~n5521 ;
  assign n5523 = n5522 ^ x80 ;
  assign n5527 = n5526 ^ n5523 ;
  assign n5528 = n5526 ^ x81 ;
  assign n5529 = n5527 & ~n5528 ;
  assign n5530 = n5529 ^ x81 ;
  assign n5534 = n5533 ^ n5530 ;
  assign n5535 = n5533 ^ x82 ;
  assign n5536 = n5534 & ~n5535 ;
  assign n5537 = n5536 ^ x82 ;
  assign n5549 = n5548 ^ n5537 ;
  assign n5550 = n5548 ^ x83 ;
  assign n5551 = n5549 & ~n5550 ;
  assign n5552 = n5551 ^ x83 ;
  assign n5556 = n5555 ^ n5552 ;
  assign n5557 = n5555 ^ x84 ;
  assign n5558 = n5556 & ~n5557 ;
  assign n5559 = n5558 ^ x84 ;
  assign n5571 = n5570 ^ n5559 ;
  assign n5572 = n5570 ^ x85 ;
  assign n5573 = n5571 & ~n5572 ;
  assign n5574 = n5573 ^ x85 ;
  assign n5578 = n5577 ^ n5574 ;
  assign n5579 = n5577 ^ x86 ;
  assign n5580 = n5578 & ~n5579 ;
  assign n5581 = n5580 ^ x86 ;
  assign n5585 = n5584 ^ n5581 ;
  assign n5586 = n5584 ^ x87 ;
  assign n5587 = n5585 & ~n5586 ;
  assign n5588 = n5587 ^ x87 ;
  assign n5592 = n5591 ^ n5588 ;
  assign n5593 = n5591 ^ x88 ;
  assign n5594 = n5592 & ~n5593 ;
  assign n5595 = n5594 ^ x88 ;
  assign n5596 = n5595 ^ n5382 ;
  assign n5597 = n5596 ^ n5396 ;
  assign n5598 = ~n5397 & n5597 ;
  assign n5599 = n5598 ^ n5396 ;
  assign n5600 = ~n5383 & n5599 ;
  assign n5601 = n5600 ^ x90 ;
  assign n5605 = n5604 ^ n5601 ;
  assign n5606 = n5604 ^ x91 ;
  assign n5607 = n5605 & ~n5606 ;
  assign n5608 = n5607 ^ x91 ;
  assign n5609 = n5608 ^ x92 ;
  assign n5648 = n5295 ^ x91 ;
  assign n5649 = n5377 & n5648 ;
  assign n5650 = n5649 ^ n5298 ;
  assign n5651 = n5650 ^ n5608 ;
  assign n5652 = n5609 & n5651 ;
  assign n5653 = n5652 ^ x92 ;
  assign n5654 = n5653 ^ n5646 ;
  assign n5655 = ~n5647 & n5654 ;
  assign n5656 = n5655 ^ x93 ;
  assign n5657 = n5656 ^ n5642 ;
  assign n5658 = ~n5643 & n5657 ;
  assign n5659 = n5658 ^ x94 ;
  assign n5663 = n5662 ^ n5659 ;
  assign n5664 = n5662 ^ x95 ;
  assign n5665 = n5663 & ~n5664 ;
  assign n5666 = n5665 ^ x95 ;
  assign n5667 = n5666 ^ n5624 ;
  assign n5668 = n5667 ^ n5630 ;
  assign n5669 = ~n5631 & n5668 ;
  assign n5670 = n5669 ^ n5630 ;
  assign n5671 = ~n5625 & n5670 ;
  assign n5672 = n5671 ^ x97 ;
  assign n5676 = n5675 ^ n5672 ;
  assign n5677 = n5675 ^ x98 ;
  assign n5678 = n5676 & ~n5677 ;
  assign n5679 = n5678 ^ x98 ;
  assign n5683 = n5682 ^ n5679 ;
  assign n5684 = n5682 ^ x99 ;
  assign n5685 = n5683 & ~n5684 ;
  assign n5686 = n5685 ^ x99 ;
  assign n5691 = x100 & x101 ;
  assign n5692 = n5691 ^ n5619 ;
  assign n5693 = n5686 & n5692 ;
  assign n5694 = n5621 & ~n5693 ;
  assign n5989 = n5686 ^ x100 ;
  assign n5990 = n5694 & n5989 ;
  assign n5991 = n5990 ^ n5616 ;
  assign n5611 = x100 & ~n5610 ;
  assign n5695 = n5686 & n5694 ;
  assign n5696 = n5611 & n5695 ;
  assign n5697 = n5696 ^ n5694 ;
  assign n5982 = n5679 ^ x99 ;
  assign n5983 = n5697 & n5982 ;
  assign n5984 = n5983 ^ n5682 ;
  assign n5975 = n5672 ^ x98 ;
  assign n5976 = n5697 & n5975 ;
  assign n5977 = n5976 ^ n5675 ;
  assign n5960 = n5628 ^ x97 ;
  assign n5961 = n5960 ^ x96 ;
  assign n5962 = n5961 ^ n5666 ;
  assign n5963 = n5962 ^ n5960 ;
  assign n5965 = x97 ^ x96 ;
  assign n5966 = n5965 ^ n5960 ;
  assign n5967 = ~n5963 & ~n5966 ;
  assign n5968 = n5967 ^ n5960 ;
  assign n5969 = n5697 & ~n5968 ;
  assign n5970 = n5969 ^ n5624 ;
  assign n5953 = n5666 ^ x96 ;
  assign n5954 = n5697 & n5953 ;
  assign n5955 = n5954 ^ n5628 ;
  assign n5946 = n5659 ^ x95 ;
  assign n5947 = n5697 & n5946 ;
  assign n5948 = n5947 ^ n5662 ;
  assign n5939 = n5656 ^ x94 ;
  assign n5940 = n5697 & n5939 ;
  assign n5941 = n5940 ^ n5642 ;
  assign n5932 = n5653 ^ x93 ;
  assign n5933 = n5697 & n5932 ;
  assign n5934 = n5933 ^ n5646 ;
  assign n5698 = n5609 & n5697 ;
  assign n5699 = n5698 ^ n5650 ;
  assign n5700 = n5699 ^ x93 ;
  assign n5705 = n5699 ^ x92 ;
  assign n5701 = n5601 ^ x91 ;
  assign n5702 = n5697 & n5701 ;
  assign n5703 = n5702 ^ n5604 ;
  assign n5704 = n5703 ^ n5699 ;
  assign n5706 = n5705 ^ n5704 ;
  assign n5707 = n5394 ^ x90 ;
  assign n5708 = n5707 ^ x89 ;
  assign n5709 = n5708 ^ n5595 ;
  assign n5710 = n5709 ^ n5707 ;
  assign n5712 = x90 ^ x89 ;
  assign n5713 = n5712 ^ n5707 ;
  assign n5714 = ~n5710 & ~n5713 ;
  assign n5715 = n5714 ^ n5707 ;
  assign n5716 = n5697 & ~n5715 ;
  assign n5717 = n5716 ^ n5382 ;
  assign n5718 = n5717 ^ x91 ;
  assign n5723 = n5717 ^ x90 ;
  assign n5719 = n5595 ^ x89 ;
  assign n5720 = n5697 & n5719 ;
  assign n5721 = n5720 ^ n5394 ;
  assign n5722 = n5721 ^ n5717 ;
  assign n5724 = n5723 ^ n5722 ;
  assign n5913 = n5588 ^ x88 ;
  assign n5914 = n5697 & n5913 ;
  assign n5915 = n5914 ^ n5591 ;
  assign n5906 = n5581 ^ x87 ;
  assign n5907 = n5697 & n5906 ;
  assign n5908 = n5907 ^ n5584 ;
  assign n5899 = n5574 ^ x86 ;
  assign n5900 = n5697 & n5899 ;
  assign n5901 = n5900 ^ n5577 ;
  assign n5892 = n5559 ^ x85 ;
  assign n5893 = n5697 & n5892 ;
  assign n5894 = n5893 ^ n5570 ;
  assign n5885 = n5552 ^ x84 ;
  assign n5886 = n5697 & n5885 ;
  assign n5887 = n5886 ^ n5555 ;
  assign n5878 = n5537 ^ x83 ;
  assign n5879 = n5697 & n5878 ;
  assign n5880 = n5879 ^ n5548 ;
  assign n5871 = n5530 ^ x82 ;
  assign n5872 = n5697 & n5871 ;
  assign n5873 = n5872 ^ n5533 ;
  assign n5864 = n5523 ^ x81 ;
  assign n5865 = n5697 & n5864 ;
  assign n5866 = n5865 ^ n5526 ;
  assign n5857 = n5516 ^ x80 ;
  assign n5858 = n5697 & n5857 ;
  assign n5859 = n5858 ^ n5519 ;
  assign n5850 = n5509 ^ x79 ;
  assign n5851 = n5697 & n5850 ;
  assign n5852 = n5851 ^ n5512 ;
  assign n5835 = n5404 ^ x78 ;
  assign n5836 = n5835 ^ x77 ;
  assign n5837 = n5836 ^ n5503 ;
  assign n5838 = n5837 ^ n5835 ;
  assign n5840 = x78 ^ x77 ;
  assign n5841 = n5840 ^ n5835 ;
  assign n5842 = ~n5838 & ~n5841 ;
  assign n5843 = n5842 ^ n5835 ;
  assign n5844 = n5697 & ~n5843 ;
  assign n5845 = n5844 ^ n5400 ;
  assign n5828 = n5503 ^ x77 ;
  assign n5829 = n5697 & n5828 ;
  assign n5830 = n5829 ^ n5404 ;
  assign n5821 = n5496 ^ x76 ;
  assign n5822 = n5697 & n5821 ;
  assign n5823 = n5822 ^ n5499 ;
  assign n5814 = n5489 ^ x75 ;
  assign n5815 = n5697 & n5814 ;
  assign n5816 = n5815 ^ n5492 ;
  assign n5807 = n5482 ^ x74 ;
  assign n5808 = n5697 & n5807 ;
  assign n5809 = n5808 ^ n5485 ;
  assign n5800 = n5475 ^ x73 ;
  assign n5801 = n5697 & n5800 ;
  assign n5802 = n5801 ^ n5478 ;
  assign n5793 = n5468 ^ x72 ;
  assign n5794 = n5697 & n5793 ;
  assign n5795 = n5794 ^ n5471 ;
  assign n5786 = n5461 ^ x71 ;
  assign n5787 = n5697 & n5786 ;
  assign n5788 = n5787 ^ n5464 ;
  assign n5779 = n5454 ^ x70 ;
  assign n5780 = n5697 & n5779 ;
  assign n5781 = n5780 ^ n5457 ;
  assign n5772 = n5447 ^ x69 ;
  assign n5773 = n5697 & n5772 ;
  assign n5774 = n5773 ^ n5450 ;
  assign n5765 = n5440 ^ x68 ;
  assign n5766 = n5697 & n5765 ;
  assign n5767 = n5766 ^ n5443 ;
  assign n5758 = n5433 ^ x67 ;
  assign n5759 = n5697 & n5758 ;
  assign n5760 = n5759 ^ n5436 ;
  assign n5751 = n5430 ^ x66 ;
  assign n5752 = n5697 & n5751 ;
  assign n5753 = n5752 ^ n5417 ;
  assign n5740 = n5377 ^ x26 ;
  assign n5741 = n5740 ^ n5377 ;
  assign n5742 = n5697 & ~n5741 ;
  assign n5743 = n5742 ^ n5377 ;
  assign n5744 = x64 & n5743 ;
  assign n5745 = n5744 ^ x27 ;
  assign n5737 = x65 & n5697 ;
  assign n5746 = n5745 ^ n5737 ;
  assign n5732 = x26 & x65 ;
  assign n5729 = x65 ^ x25 ;
  assign n5725 = x64 ^ x26 ;
  assign n5726 = n5725 ^ x65 ;
  assign n5730 = n5726 ^ n5697 ;
  assign n5731 = ~n5729 & n5730 ;
  assign n5733 = n5732 ^ n5731 ;
  assign n5734 = x64 & n5733 ;
  assign n5735 = n5734 ^ n5732 ;
  assign n5736 = n5735 ^ x65 ;
  assign n5747 = n5746 ^ n5736 ;
  assign n5748 = n5746 ^ x66 ;
  assign n5749 = n5747 & ~n5748 ;
  assign n5750 = n5749 ^ x66 ;
  assign n5754 = n5753 ^ n5750 ;
  assign n5755 = n5753 ^ x67 ;
  assign n5756 = n5754 & ~n5755 ;
  assign n5757 = n5756 ^ x67 ;
  assign n5761 = n5760 ^ n5757 ;
  assign n5762 = n5760 ^ x68 ;
  assign n5763 = n5761 & ~n5762 ;
  assign n5764 = n5763 ^ x68 ;
  assign n5768 = n5767 ^ n5764 ;
  assign n5769 = n5767 ^ x69 ;
  assign n5770 = n5768 & ~n5769 ;
  assign n5771 = n5770 ^ x69 ;
  assign n5775 = n5774 ^ n5771 ;
  assign n5776 = n5774 ^ x70 ;
  assign n5777 = n5775 & ~n5776 ;
  assign n5778 = n5777 ^ x70 ;
  assign n5782 = n5781 ^ n5778 ;
  assign n5783 = n5781 ^ x71 ;
  assign n5784 = n5782 & ~n5783 ;
  assign n5785 = n5784 ^ x71 ;
  assign n5789 = n5788 ^ n5785 ;
  assign n5790 = n5788 ^ x72 ;
  assign n5791 = n5789 & ~n5790 ;
  assign n5792 = n5791 ^ x72 ;
  assign n5796 = n5795 ^ n5792 ;
  assign n5797 = n5795 ^ x73 ;
  assign n5798 = n5796 & ~n5797 ;
  assign n5799 = n5798 ^ x73 ;
  assign n5803 = n5802 ^ n5799 ;
  assign n5804 = n5802 ^ x74 ;
  assign n5805 = n5803 & ~n5804 ;
  assign n5806 = n5805 ^ x74 ;
  assign n5810 = n5809 ^ n5806 ;
  assign n5811 = n5809 ^ x75 ;
  assign n5812 = n5810 & ~n5811 ;
  assign n5813 = n5812 ^ x75 ;
  assign n5817 = n5816 ^ n5813 ;
  assign n5818 = n5816 ^ x76 ;
  assign n5819 = n5817 & ~n5818 ;
  assign n5820 = n5819 ^ x76 ;
  assign n5824 = n5823 ^ n5820 ;
  assign n5825 = n5823 ^ x77 ;
  assign n5826 = n5824 & ~n5825 ;
  assign n5827 = n5826 ^ x77 ;
  assign n5831 = n5830 ^ n5827 ;
  assign n5832 = n5830 ^ x78 ;
  assign n5833 = n5831 & ~n5832 ;
  assign n5834 = n5833 ^ x78 ;
  assign n5846 = n5845 ^ n5834 ;
  assign n5847 = n5845 ^ x79 ;
  assign n5848 = n5846 & ~n5847 ;
  assign n5849 = n5848 ^ x79 ;
  assign n5853 = n5852 ^ n5849 ;
  assign n5854 = n5852 ^ x80 ;
  assign n5855 = n5853 & ~n5854 ;
  assign n5856 = n5855 ^ x80 ;
  assign n5860 = n5859 ^ n5856 ;
  assign n5861 = n5859 ^ x81 ;
  assign n5862 = n5860 & ~n5861 ;
  assign n5863 = n5862 ^ x81 ;
  assign n5867 = n5866 ^ n5863 ;
  assign n5868 = n5866 ^ x82 ;
  assign n5869 = n5867 & ~n5868 ;
  assign n5870 = n5869 ^ x82 ;
  assign n5874 = n5873 ^ n5870 ;
  assign n5875 = n5873 ^ x83 ;
  assign n5876 = n5874 & ~n5875 ;
  assign n5877 = n5876 ^ x83 ;
  assign n5881 = n5880 ^ n5877 ;
  assign n5882 = n5880 ^ x84 ;
  assign n5883 = n5881 & ~n5882 ;
  assign n5884 = n5883 ^ x84 ;
  assign n5888 = n5887 ^ n5884 ;
  assign n5889 = n5887 ^ x85 ;
  assign n5890 = n5888 & ~n5889 ;
  assign n5891 = n5890 ^ x85 ;
  assign n5895 = n5894 ^ n5891 ;
  assign n5896 = n5894 ^ x86 ;
  assign n5897 = n5895 & ~n5896 ;
  assign n5898 = n5897 ^ x86 ;
  assign n5902 = n5901 ^ n5898 ;
  assign n5903 = n5901 ^ x87 ;
  assign n5904 = n5902 & ~n5903 ;
  assign n5905 = n5904 ^ x87 ;
  assign n5909 = n5908 ^ n5905 ;
  assign n5910 = n5908 ^ x88 ;
  assign n5911 = n5909 & ~n5910 ;
  assign n5912 = n5911 ^ x88 ;
  assign n5916 = n5915 ^ n5912 ;
  assign n5917 = n5915 ^ x89 ;
  assign n5918 = n5916 & ~n5917 ;
  assign n5919 = n5918 ^ x89 ;
  assign n5920 = n5919 ^ n5717 ;
  assign n5921 = n5920 ^ n5723 ;
  assign n5922 = ~n5724 & n5921 ;
  assign n5923 = n5922 ^ n5723 ;
  assign n5924 = ~n5718 & n5923 ;
  assign n5925 = n5924 ^ x91 ;
  assign n5926 = n5925 ^ n5699 ;
  assign n5927 = n5926 ^ n5705 ;
  assign n5928 = ~n5706 & n5927 ;
  assign n5929 = n5928 ^ n5705 ;
  assign n5930 = ~n5700 & n5929 ;
  assign n5931 = n5930 ^ x93 ;
  assign n5935 = n5934 ^ n5931 ;
  assign n5936 = n5934 ^ x94 ;
  assign n5937 = n5935 & ~n5936 ;
  assign n5938 = n5937 ^ x94 ;
  assign n5942 = n5941 ^ n5938 ;
  assign n5943 = n5941 ^ x95 ;
  assign n5944 = n5942 & ~n5943 ;
  assign n5945 = n5944 ^ x95 ;
  assign n5949 = n5948 ^ n5945 ;
  assign n5950 = n5948 ^ x96 ;
  assign n5951 = n5949 & ~n5950 ;
  assign n5952 = n5951 ^ x96 ;
  assign n5956 = n5955 ^ n5952 ;
  assign n5957 = n5955 ^ x97 ;
  assign n5958 = n5956 & ~n5957 ;
  assign n5959 = n5958 ^ x97 ;
  assign n5971 = n5970 ^ n5959 ;
  assign n5972 = n5970 ^ x98 ;
  assign n5973 = n5971 & ~n5972 ;
  assign n5974 = n5973 ^ x98 ;
  assign n5978 = n5977 ^ n5974 ;
  assign n5979 = n5977 ^ x99 ;
  assign n5980 = n5978 & ~n5979 ;
  assign n5981 = n5980 ^ x99 ;
  assign n5985 = n5984 ^ n5981 ;
  assign n5986 = n5984 ^ x100 ;
  assign n5987 = n5985 & ~n5986 ;
  assign n5988 = n5987 ^ x100 ;
  assign n5992 = n5991 ^ n5988 ;
  assign n5993 = n5991 ^ x101 ;
  assign n5994 = n5992 & ~n5993 ;
  assign n5995 = n5994 ^ x101 ;
  assign n5996 = n154 & ~n5995 ;
  assign n5997 = n5379 & ~n5996 ;
  assign n6313 = n5997 ^ n375 ;
  assign n5998 = n153 & ~n154 ;
  assign n5999 = n5610 & n5998 ;
  assign n6000 = n5999 ^ n154 ;
  assign n6001 = n5988 ^ x101 ;
  assign n6002 = n5995 ^ x102 ;
  assign n6009 = ~n375 & n5694 ;
  assign n6010 = n5610 & n6009 ;
  assign n6011 = n6010 ^ n5610 ;
  assign n6012 = n6011 ^ n5995 ;
  assign n6013 = n6002 & n6012 ;
  assign n6014 = n6013 ^ x102 ;
  assign n6015 = n154 & ~n6014 ;
  assign n6016 = n6001 & n6015 ;
  assign n6017 = n6016 ^ n5991 ;
  assign n6018 = n6017 ^ x102 ;
  assign n6298 = n5981 ^ x100 ;
  assign n6299 = n6015 & n6298 ;
  assign n6300 = n6299 ^ n5984 ;
  assign n6291 = n5974 ^ x99 ;
  assign n6292 = n6015 & n6291 ;
  assign n6293 = n6292 ^ n5977 ;
  assign n6284 = n5959 ^ x98 ;
  assign n6285 = n6015 & n6284 ;
  assign n6286 = n6285 ^ n5970 ;
  assign n6019 = n5952 ^ x97 ;
  assign n6020 = n6015 & n6019 ;
  assign n6021 = n6020 ^ n5955 ;
  assign n6022 = n6021 ^ x98 ;
  assign n6023 = n5945 ^ x96 ;
  assign n6024 = n6015 & n6023 ;
  assign n6025 = n6024 ^ n5948 ;
  assign n6026 = n6025 ^ x97 ;
  assign n6271 = n5938 ^ x95 ;
  assign n6272 = n6015 & n6271 ;
  assign n6273 = n6272 ^ n5941 ;
  assign n6264 = n5931 ^ x94 ;
  assign n6265 = n6015 & n6264 ;
  assign n6266 = n6265 ^ n5934 ;
  assign n6249 = n5703 ^ x93 ;
  assign n6250 = n6249 ^ x92 ;
  assign n6251 = n6250 ^ n5925 ;
  assign n6252 = n6251 ^ n6249 ;
  assign n6255 = n6249 ^ n3803 ;
  assign n6256 = ~n6252 & ~n6255 ;
  assign n6257 = n6256 ^ n6249 ;
  assign n6258 = n6015 & ~n6257 ;
  assign n6259 = n6258 ^ n5699 ;
  assign n6242 = n5925 ^ x92 ;
  assign n6243 = n6015 & n6242 ;
  assign n6244 = n6243 ^ n5703 ;
  assign n6227 = n5721 ^ x91 ;
  assign n6228 = n6227 ^ x90 ;
  assign n6229 = n6228 ^ n5919 ;
  assign n6230 = n6229 ^ n6227 ;
  assign n6232 = x91 ^ x90 ;
  assign n6233 = n6232 ^ n6227 ;
  assign n6234 = ~n6230 & ~n6233 ;
  assign n6235 = n6234 ^ n6227 ;
  assign n6236 = n6015 & ~n6235 ;
  assign n6237 = n6236 ^ n5717 ;
  assign n6220 = n5919 ^ x90 ;
  assign n6221 = n6015 & n6220 ;
  assign n6222 = n6221 ^ n5721 ;
  assign n6213 = n5912 ^ x89 ;
  assign n6214 = n6015 & n6213 ;
  assign n6215 = n6214 ^ n5915 ;
  assign n6206 = n5905 ^ x88 ;
  assign n6207 = n6015 & n6206 ;
  assign n6208 = n6207 ^ n5908 ;
  assign n6199 = n5898 ^ x87 ;
  assign n6200 = n6015 & n6199 ;
  assign n6201 = n6200 ^ n5901 ;
  assign n6192 = n5891 ^ x86 ;
  assign n6193 = n6015 & n6192 ;
  assign n6194 = n6193 ^ n5894 ;
  assign n6185 = n5884 ^ x85 ;
  assign n6186 = n6015 & n6185 ;
  assign n6187 = n6186 ^ n5887 ;
  assign n6178 = n5877 ^ x84 ;
  assign n6179 = n6015 & n6178 ;
  assign n6180 = n6179 ^ n5880 ;
  assign n6171 = n5870 ^ x83 ;
  assign n6172 = n6015 & n6171 ;
  assign n6173 = n6172 ^ n5873 ;
  assign n6164 = n5863 ^ x82 ;
  assign n6165 = n6015 & n6164 ;
  assign n6166 = n6165 ^ n5866 ;
  assign n6157 = n5856 ^ x81 ;
  assign n6158 = n6015 & n6157 ;
  assign n6159 = n6158 ^ n5859 ;
  assign n6150 = n5849 ^ x80 ;
  assign n6151 = n6015 & n6150 ;
  assign n6152 = n6151 ^ n5852 ;
  assign n6143 = n5834 ^ x79 ;
  assign n6144 = n6015 & n6143 ;
  assign n6145 = n6144 ^ n5845 ;
  assign n6136 = n5827 ^ x78 ;
  assign n6137 = n6015 & n6136 ;
  assign n6138 = n6137 ^ n5830 ;
  assign n6129 = n5820 ^ x77 ;
  assign n6130 = n6015 & n6129 ;
  assign n6131 = n6130 ^ n5823 ;
  assign n6122 = n5813 ^ x76 ;
  assign n6123 = n6015 & n6122 ;
  assign n6124 = n6123 ^ n5816 ;
  assign n6115 = n5806 ^ x75 ;
  assign n6116 = n6015 & n6115 ;
  assign n6117 = n6116 ^ n5809 ;
  assign n6108 = n5799 ^ x74 ;
  assign n6109 = n6015 & n6108 ;
  assign n6110 = n6109 ^ n5802 ;
  assign n6097 = n5785 ^ x72 ;
  assign n6098 = n6015 & n6097 ;
  assign n6099 = n6098 ^ n5788 ;
  assign n6030 = n5778 ^ x71 ;
  assign n6031 = n6015 & n6030 ;
  assign n6032 = n6031 ^ n5781 ;
  assign n6033 = n6032 ^ x72 ;
  assign n6038 = n6032 ^ x71 ;
  assign n6034 = n5771 ^ x70 ;
  assign n6035 = n6015 & n6034 ;
  assign n6036 = n6035 ^ n5774 ;
  assign n6037 = n6036 ^ n6032 ;
  assign n6039 = n6038 ^ n6037 ;
  assign n6084 = n5764 ^ x69 ;
  assign n6085 = n6015 & n6084 ;
  assign n6086 = n6085 ^ n5767 ;
  assign n6077 = n5757 ^ x68 ;
  assign n6078 = n6015 & n6077 ;
  assign n6079 = n6078 ^ n5760 ;
  assign n6070 = n5750 ^ x67 ;
  assign n6071 = n6015 & n6070 ;
  assign n6072 = n6071 ^ n5753 ;
  assign n6063 = n5736 ^ x66 ;
  assign n6064 = n6015 & n6063 ;
  assign n6065 = n6064 ^ n5746 ;
  assign n6045 = x64 & n5697 ;
  assign n6041 = ~x25 & x64 ;
  assign n6042 = n6041 ^ x65 ;
  assign n6043 = n6015 & n6042 ;
  assign n6044 = n6043 ^ x26 ;
  assign n6046 = n6045 ^ n6044 ;
  assign n6047 = n6046 ^ x66 ;
  assign n6055 = x25 & x65 ;
  assign n6052 = x65 ^ x24 ;
  assign n6048 = x64 ^ x25 ;
  assign n6049 = n6048 ^ x65 ;
  assign n6053 = n6049 ^ n6015 ;
  assign n6054 = ~n6052 & n6053 ;
  assign n6056 = n6055 ^ n6054 ;
  assign n6057 = x64 & n6056 ;
  assign n6058 = n6057 ^ n6055 ;
  assign n6059 = n6058 ^ x65 ;
  assign n6060 = n6059 ^ n6046 ;
  assign n6061 = ~n6047 & n6060 ;
  assign n6062 = n6061 ^ x66 ;
  assign n6066 = n6065 ^ n6062 ;
  assign n6067 = n6065 ^ x67 ;
  assign n6068 = n6066 & ~n6067 ;
  assign n6069 = n6068 ^ x67 ;
  assign n6073 = n6072 ^ n6069 ;
  assign n6074 = n6072 ^ x68 ;
  assign n6075 = n6073 & ~n6074 ;
  assign n6076 = n6075 ^ x68 ;
  assign n6080 = n6079 ^ n6076 ;
  assign n6081 = n6079 ^ x69 ;
  assign n6082 = n6080 & ~n6081 ;
  assign n6083 = n6082 ^ x69 ;
  assign n6087 = n6086 ^ n6083 ;
  assign n6088 = n6086 ^ x70 ;
  assign n6089 = n6087 & ~n6088 ;
  assign n6090 = n6089 ^ x70 ;
  assign n6091 = n6090 ^ n6032 ;
  assign n6092 = n6091 ^ n6038 ;
  assign n6093 = ~n6039 & n6092 ;
  assign n6094 = n6093 ^ n6038 ;
  assign n6095 = ~n6033 & n6094 ;
  assign n6096 = n6095 ^ x72 ;
  assign n6100 = n6099 ^ n6096 ;
  assign n6101 = n6099 ^ x73 ;
  assign n6102 = n6100 & ~n6101 ;
  assign n6103 = n6102 ^ x73 ;
  assign n6027 = n5792 ^ x73 ;
  assign n6028 = n6015 & n6027 ;
  assign n6029 = n6028 ^ n5795 ;
  assign n6104 = n6103 ^ n6029 ;
  assign n6105 = n6103 ^ x74 ;
  assign n6106 = n6104 & n6105 ;
  assign n6107 = n6106 ^ x74 ;
  assign n6111 = n6110 ^ n6107 ;
  assign n6112 = n6110 ^ x75 ;
  assign n6113 = n6111 & ~n6112 ;
  assign n6114 = n6113 ^ x75 ;
  assign n6118 = n6117 ^ n6114 ;
  assign n6119 = n6117 ^ x76 ;
  assign n6120 = n6118 & ~n6119 ;
  assign n6121 = n6120 ^ x76 ;
  assign n6125 = n6124 ^ n6121 ;
  assign n6126 = n6124 ^ x77 ;
  assign n6127 = n6125 & ~n6126 ;
  assign n6128 = n6127 ^ x77 ;
  assign n6132 = n6131 ^ n6128 ;
  assign n6133 = n6131 ^ x78 ;
  assign n6134 = n6132 & ~n6133 ;
  assign n6135 = n6134 ^ x78 ;
  assign n6139 = n6138 ^ n6135 ;
  assign n6140 = n6138 ^ x79 ;
  assign n6141 = n6139 & ~n6140 ;
  assign n6142 = n6141 ^ x79 ;
  assign n6146 = n6145 ^ n6142 ;
  assign n6147 = n6145 ^ x80 ;
  assign n6148 = n6146 & ~n6147 ;
  assign n6149 = n6148 ^ x80 ;
  assign n6153 = n6152 ^ n6149 ;
  assign n6154 = n6152 ^ x81 ;
  assign n6155 = n6153 & ~n6154 ;
  assign n6156 = n6155 ^ x81 ;
  assign n6160 = n6159 ^ n6156 ;
  assign n6161 = n6159 ^ x82 ;
  assign n6162 = n6160 & ~n6161 ;
  assign n6163 = n6162 ^ x82 ;
  assign n6167 = n6166 ^ n6163 ;
  assign n6168 = n6166 ^ x83 ;
  assign n6169 = n6167 & ~n6168 ;
  assign n6170 = n6169 ^ x83 ;
  assign n6174 = n6173 ^ n6170 ;
  assign n6175 = n6173 ^ x84 ;
  assign n6176 = n6174 & ~n6175 ;
  assign n6177 = n6176 ^ x84 ;
  assign n6181 = n6180 ^ n6177 ;
  assign n6182 = n6180 ^ x85 ;
  assign n6183 = n6181 & ~n6182 ;
  assign n6184 = n6183 ^ x85 ;
  assign n6188 = n6187 ^ n6184 ;
  assign n6189 = n6187 ^ x86 ;
  assign n6190 = n6188 & ~n6189 ;
  assign n6191 = n6190 ^ x86 ;
  assign n6195 = n6194 ^ n6191 ;
  assign n6196 = n6194 ^ x87 ;
  assign n6197 = n6195 & ~n6196 ;
  assign n6198 = n6197 ^ x87 ;
  assign n6202 = n6201 ^ n6198 ;
  assign n6203 = n6201 ^ x88 ;
  assign n6204 = n6202 & ~n6203 ;
  assign n6205 = n6204 ^ x88 ;
  assign n6209 = n6208 ^ n6205 ;
  assign n6210 = n6208 ^ x89 ;
  assign n6211 = n6209 & ~n6210 ;
  assign n6212 = n6211 ^ x89 ;
  assign n6216 = n6215 ^ n6212 ;
  assign n6217 = n6215 ^ x90 ;
  assign n6218 = n6216 & ~n6217 ;
  assign n6219 = n6218 ^ x90 ;
  assign n6223 = n6222 ^ n6219 ;
  assign n6224 = n6222 ^ x91 ;
  assign n6225 = n6223 & ~n6224 ;
  assign n6226 = n6225 ^ x91 ;
  assign n6238 = n6237 ^ n6226 ;
  assign n6239 = n6237 ^ x92 ;
  assign n6240 = n6238 & ~n6239 ;
  assign n6241 = n6240 ^ x92 ;
  assign n6245 = n6244 ^ n6241 ;
  assign n6246 = n6244 ^ x93 ;
  assign n6247 = n6245 & ~n6246 ;
  assign n6248 = n6247 ^ x93 ;
  assign n6260 = n6259 ^ n6248 ;
  assign n6261 = n6259 ^ x94 ;
  assign n6262 = n6260 & ~n6261 ;
  assign n6263 = n6262 ^ x94 ;
  assign n6267 = n6266 ^ n6263 ;
  assign n6268 = n6266 ^ x95 ;
  assign n6269 = n6267 & ~n6268 ;
  assign n6270 = n6269 ^ x95 ;
  assign n6274 = n6273 ^ n6270 ;
  assign n6275 = n6273 ^ x96 ;
  assign n6276 = n6274 & ~n6275 ;
  assign n6277 = n6276 ^ x96 ;
  assign n6278 = n6277 ^ n6025 ;
  assign n6279 = ~n6026 & n6278 ;
  assign n6280 = n6279 ^ x97 ;
  assign n6281 = n6280 ^ n6021 ;
  assign n6282 = ~n6022 & n6281 ;
  assign n6283 = n6282 ^ x98 ;
  assign n6287 = n6286 ^ n6283 ;
  assign n6288 = n6286 ^ x99 ;
  assign n6289 = n6287 & ~n6288 ;
  assign n6290 = n6289 ^ x99 ;
  assign n6294 = n6293 ^ n6290 ;
  assign n6295 = n6293 ^ x100 ;
  assign n6296 = n6294 & ~n6295 ;
  assign n6297 = n6296 ^ x100 ;
  assign n6301 = n6300 ^ n6297 ;
  assign n6605 = n6297 ^ x101 ;
  assign n6305 = n6301 & n6605 ;
  assign n6302 = x102 ^ x101 ;
  assign n6306 = n6305 ^ n6302 ;
  assign n6309 = ~n6018 & n6306 ;
  assign n6310 = n6309 ^ x102 ;
  assign n6311 = n6000 & n6310 ;
  assign n6314 = ~x103 & n6311 ;
  assign n6315 = n6313 & n6314 ;
  assign n6312 = n6311 ^ n6000 ;
  assign n6316 = n6315 ^ n6312 ;
  assign n6317 = n5997 & ~n6316 ;
  assign n6320 = ~x105 & n6319 ;
  assign n6321 = n6317 ^ n375 ;
  assign n6322 = n6321 ^ x104 ;
  assign n6326 = n6321 ^ x103 ;
  assign n6323 = n6306 & n6316 ;
  assign n6324 = n6323 ^ n6017 ;
  assign n6325 = n6324 ^ n6321 ;
  assign n6327 = n6326 ^ n6325 ;
  assign n6606 = n6316 & n6605 ;
  assign n6607 = n6606 ^ n6300 ;
  assign n6598 = n6290 ^ x100 ;
  assign n6599 = n6316 & n6598 ;
  assign n6600 = n6599 ^ n6293 ;
  assign n6591 = n6283 ^ x99 ;
  assign n6592 = n6316 & n6591 ;
  assign n6593 = n6592 ^ n6286 ;
  assign n6584 = n6280 ^ x98 ;
  assign n6585 = n6316 & n6584 ;
  assign n6586 = n6585 ^ n6021 ;
  assign n6577 = n6277 ^ x97 ;
  assign n6578 = n6316 & n6577 ;
  assign n6579 = n6578 ^ n6025 ;
  assign n6328 = n6270 ^ x96 ;
  assign n6329 = n6316 & n6328 ;
  assign n6330 = n6329 ^ n6273 ;
  assign n6331 = n6330 ^ x97 ;
  assign n6332 = n6263 ^ x95 ;
  assign n6333 = n6316 & n6332 ;
  assign n6334 = n6333 ^ n6266 ;
  assign n6335 = n6334 ^ x96 ;
  assign n6564 = n6248 ^ x94 ;
  assign n6565 = n6316 & n6564 ;
  assign n6566 = n6565 ^ n6259 ;
  assign n6557 = n6241 ^ x93 ;
  assign n6558 = n6316 & n6557 ;
  assign n6559 = n6558 ^ n6244 ;
  assign n6336 = n6226 ^ x92 ;
  assign n6337 = n6316 & n6336 ;
  assign n6338 = n6337 ^ n6237 ;
  assign n6339 = n6338 ^ x93 ;
  assign n6344 = n6338 ^ x92 ;
  assign n6340 = n6219 ^ x91 ;
  assign n6341 = n6316 & n6340 ;
  assign n6342 = n6341 ^ n6222 ;
  assign n6343 = n6342 ^ n6338 ;
  assign n6345 = n6344 ^ n6343 ;
  assign n6544 = n6212 ^ x90 ;
  assign n6545 = n6316 & n6544 ;
  assign n6546 = n6545 ^ n6215 ;
  assign n6537 = n6205 ^ x89 ;
  assign n6538 = n6316 & n6537 ;
  assign n6539 = n6538 ^ n6208 ;
  assign n6346 = n6198 ^ x88 ;
  assign n6347 = n6316 & n6346 ;
  assign n6348 = n6347 ^ n6201 ;
  assign n6349 = n6348 ^ x89 ;
  assign n6354 = n6348 ^ x88 ;
  assign n6350 = n6191 ^ x87 ;
  assign n6351 = n6316 & n6350 ;
  assign n6352 = n6351 ^ n6194 ;
  assign n6353 = n6352 ^ n6348 ;
  assign n6355 = n6354 ^ n6353 ;
  assign n6356 = n6184 ^ x86 ;
  assign n6357 = n6316 & n6356 ;
  assign n6358 = n6357 ^ n6187 ;
  assign n6359 = n6358 ^ x87 ;
  assign n6364 = n6358 ^ x86 ;
  assign n6360 = n6177 ^ x85 ;
  assign n6361 = n6316 & n6360 ;
  assign n6362 = n6361 ^ n6180 ;
  assign n6363 = n6362 ^ n6358 ;
  assign n6365 = n6364 ^ n6363 ;
  assign n6518 = n6170 ^ x84 ;
  assign n6519 = n6316 & n6518 ;
  assign n6520 = n6519 ^ n6173 ;
  assign n6511 = n6163 ^ x83 ;
  assign n6512 = n6316 & n6511 ;
  assign n6513 = n6512 ^ n6166 ;
  assign n6504 = n6156 ^ x82 ;
  assign n6505 = n6316 & n6504 ;
  assign n6506 = n6505 ^ n6159 ;
  assign n6497 = n6149 ^ x81 ;
  assign n6498 = n6316 & n6497 ;
  assign n6499 = n6498 ^ n6152 ;
  assign n6490 = n6142 ^ x80 ;
  assign n6491 = n6316 & n6490 ;
  assign n6492 = n6491 ^ n6145 ;
  assign n6483 = n6135 ^ x79 ;
  assign n6484 = n6316 & n6483 ;
  assign n6485 = n6484 ^ n6138 ;
  assign n6476 = n6128 ^ x78 ;
  assign n6477 = n6316 & n6476 ;
  assign n6478 = n6477 ^ n6131 ;
  assign n6469 = n6121 ^ x77 ;
  assign n6470 = n6316 & n6469 ;
  assign n6471 = n6470 ^ n6124 ;
  assign n6462 = n6114 ^ x76 ;
  assign n6463 = n6316 & n6462 ;
  assign n6464 = n6463 ^ n6117 ;
  assign n6455 = n6107 ^ x75 ;
  assign n6456 = n6316 & n6455 ;
  assign n6457 = n6456 ^ n6110 ;
  assign n6449 = n6105 & n6316 ;
  assign n6450 = n6449 ^ n6029 ;
  assign n6442 = n6096 ^ x73 ;
  assign n6443 = n6316 & n6442 ;
  assign n6444 = n6443 ^ n6099 ;
  assign n6427 = n6036 ^ x72 ;
  assign n6428 = n6427 ^ x71 ;
  assign n6429 = n6428 ^ n6090 ;
  assign n6430 = n6429 ^ n6427 ;
  assign n6433 = n6427 ^ n3023 ;
  assign n6434 = ~n6430 & ~n6433 ;
  assign n6435 = n6434 ^ n6427 ;
  assign n6436 = n6316 & ~n6435 ;
  assign n6437 = n6436 ^ n6032 ;
  assign n6420 = n6090 ^ x71 ;
  assign n6421 = n6316 & n6420 ;
  assign n6422 = n6421 ^ n6036 ;
  assign n6413 = n6083 ^ x70 ;
  assign n6414 = n6316 & n6413 ;
  assign n6415 = n6414 ^ n6086 ;
  assign n6406 = n6076 ^ x69 ;
  assign n6407 = n6316 & n6406 ;
  assign n6408 = n6407 ^ n6079 ;
  assign n6399 = n6069 ^ x68 ;
  assign n6400 = n6316 & n6399 ;
  assign n6401 = n6400 ^ n6072 ;
  assign n6392 = n6062 ^ x67 ;
  assign n6393 = n6316 & n6392 ;
  assign n6394 = n6393 ^ n6065 ;
  assign n6385 = n6059 ^ x66 ;
  assign n6386 = n6316 & n6385 ;
  assign n6387 = n6386 ^ n6046 ;
  assign n6371 = x64 & n6015 ;
  assign n6367 = ~x24 & x64 ;
  assign n6368 = n6367 ^ x65 ;
  assign n6369 = n6316 & n6368 ;
  assign n6370 = n6369 ^ x25 ;
  assign n6372 = n6371 ^ n6370 ;
  assign n6373 = n6372 ^ x66 ;
  assign n6376 = ~x23 & x64 ;
  assign n6379 = n6316 ^ x24 ;
  assign n6380 = n6376 & ~n6379 ;
  assign n6374 = x64 & n6316 ;
  assign n6375 = n6374 ^ x24 ;
  assign n6377 = n6376 ^ n6375 ;
  assign n6378 = x65 & ~n6377 ;
  assign n6381 = n6380 ^ n6378 ;
  assign n6382 = n6381 ^ n6372 ;
  assign n6383 = ~n6373 & n6382 ;
  assign n6384 = n6383 ^ x66 ;
  assign n6388 = n6387 ^ n6384 ;
  assign n6389 = n6387 ^ x67 ;
  assign n6390 = n6388 & ~n6389 ;
  assign n6391 = n6390 ^ x67 ;
  assign n6395 = n6394 ^ n6391 ;
  assign n6396 = n6394 ^ x68 ;
  assign n6397 = n6395 & ~n6396 ;
  assign n6398 = n6397 ^ x68 ;
  assign n6402 = n6401 ^ n6398 ;
  assign n6403 = n6401 ^ x69 ;
  assign n6404 = n6402 & ~n6403 ;
  assign n6405 = n6404 ^ x69 ;
  assign n6409 = n6408 ^ n6405 ;
  assign n6410 = n6408 ^ x70 ;
  assign n6411 = n6409 & ~n6410 ;
  assign n6412 = n6411 ^ x70 ;
  assign n6416 = n6415 ^ n6412 ;
  assign n6417 = n6415 ^ x71 ;
  assign n6418 = n6416 & ~n6417 ;
  assign n6419 = n6418 ^ x71 ;
  assign n6423 = n6422 ^ n6419 ;
  assign n6424 = n6422 ^ x72 ;
  assign n6425 = n6423 & ~n6424 ;
  assign n6426 = n6425 ^ x72 ;
  assign n6438 = n6437 ^ n6426 ;
  assign n6439 = n6437 ^ x73 ;
  assign n6440 = n6438 & ~n6439 ;
  assign n6441 = n6440 ^ x73 ;
  assign n6445 = n6444 ^ n6441 ;
  assign n6446 = n6444 ^ x74 ;
  assign n6447 = n6445 & ~n6446 ;
  assign n6448 = n6447 ^ x74 ;
  assign n6451 = n6450 ^ n6448 ;
  assign n6452 = n6450 ^ x75 ;
  assign n6453 = n6451 & ~n6452 ;
  assign n6454 = n6453 ^ x75 ;
  assign n6458 = n6457 ^ n6454 ;
  assign n6459 = n6457 ^ x76 ;
  assign n6460 = n6458 & ~n6459 ;
  assign n6461 = n6460 ^ x76 ;
  assign n6465 = n6464 ^ n6461 ;
  assign n6466 = n6464 ^ x77 ;
  assign n6467 = n6465 & ~n6466 ;
  assign n6468 = n6467 ^ x77 ;
  assign n6472 = n6471 ^ n6468 ;
  assign n6473 = n6471 ^ x78 ;
  assign n6474 = n6472 & ~n6473 ;
  assign n6475 = n6474 ^ x78 ;
  assign n6479 = n6478 ^ n6475 ;
  assign n6480 = n6478 ^ x79 ;
  assign n6481 = n6479 & ~n6480 ;
  assign n6482 = n6481 ^ x79 ;
  assign n6486 = n6485 ^ n6482 ;
  assign n6487 = n6485 ^ x80 ;
  assign n6488 = n6486 & ~n6487 ;
  assign n6489 = n6488 ^ x80 ;
  assign n6493 = n6492 ^ n6489 ;
  assign n6494 = n6492 ^ x81 ;
  assign n6495 = n6493 & ~n6494 ;
  assign n6496 = n6495 ^ x81 ;
  assign n6500 = n6499 ^ n6496 ;
  assign n6501 = n6499 ^ x82 ;
  assign n6502 = n6500 & ~n6501 ;
  assign n6503 = n6502 ^ x82 ;
  assign n6507 = n6506 ^ n6503 ;
  assign n6508 = n6506 ^ x83 ;
  assign n6509 = n6507 & ~n6508 ;
  assign n6510 = n6509 ^ x83 ;
  assign n6514 = n6513 ^ n6510 ;
  assign n6515 = n6513 ^ x84 ;
  assign n6516 = n6514 & ~n6515 ;
  assign n6517 = n6516 ^ x84 ;
  assign n6521 = n6520 ^ n6517 ;
  assign n6522 = n6520 ^ x85 ;
  assign n6523 = n6521 & ~n6522 ;
  assign n6524 = n6523 ^ x85 ;
  assign n6525 = n6524 ^ n6358 ;
  assign n6526 = n6525 ^ n6364 ;
  assign n6527 = ~n6365 & n6526 ;
  assign n6528 = n6527 ^ n6364 ;
  assign n6529 = ~n6359 & n6528 ;
  assign n6530 = n6529 ^ x87 ;
  assign n6531 = n6530 ^ n6348 ;
  assign n6532 = n6531 ^ n6354 ;
  assign n6533 = ~n6355 & n6532 ;
  assign n6534 = n6533 ^ n6354 ;
  assign n6535 = ~n6349 & n6534 ;
  assign n6536 = n6535 ^ x89 ;
  assign n6540 = n6539 ^ n6536 ;
  assign n6541 = n6539 ^ x90 ;
  assign n6542 = n6540 & ~n6541 ;
  assign n6543 = n6542 ^ x90 ;
  assign n6547 = n6546 ^ n6543 ;
  assign n6548 = n6546 ^ x91 ;
  assign n6549 = n6547 & ~n6548 ;
  assign n6550 = n6549 ^ x91 ;
  assign n6551 = n6550 ^ n6338 ;
  assign n6552 = n6551 ^ n6344 ;
  assign n6553 = ~n6345 & n6552 ;
  assign n6554 = n6553 ^ n6344 ;
  assign n6555 = ~n6339 & n6554 ;
  assign n6556 = n6555 ^ x93 ;
  assign n6560 = n6559 ^ n6556 ;
  assign n6561 = n6559 ^ x94 ;
  assign n6562 = n6560 & ~n6561 ;
  assign n6563 = n6562 ^ x94 ;
  assign n6567 = n6566 ^ n6563 ;
  assign n6568 = n6566 ^ x95 ;
  assign n6569 = n6567 & ~n6568 ;
  assign n6570 = n6569 ^ x95 ;
  assign n6571 = n6570 ^ n6334 ;
  assign n6572 = ~n6335 & n6571 ;
  assign n6573 = n6572 ^ x96 ;
  assign n6574 = n6573 ^ n6330 ;
  assign n6575 = ~n6331 & n6574 ;
  assign n6576 = n6575 ^ x97 ;
  assign n6580 = n6579 ^ n6576 ;
  assign n6581 = n6579 ^ x98 ;
  assign n6582 = n6580 & ~n6581 ;
  assign n6583 = n6582 ^ x98 ;
  assign n6587 = n6586 ^ n6583 ;
  assign n6588 = n6586 ^ x99 ;
  assign n6589 = n6587 & ~n6588 ;
  assign n6590 = n6589 ^ x99 ;
  assign n6594 = n6593 ^ n6590 ;
  assign n6595 = n6593 ^ x100 ;
  assign n6596 = n6594 & ~n6595 ;
  assign n6597 = n6596 ^ x100 ;
  assign n6601 = n6600 ^ n6597 ;
  assign n6602 = n6600 ^ x101 ;
  assign n6603 = n6601 & ~n6602 ;
  assign n6604 = n6603 ^ x101 ;
  assign n6608 = n6607 ^ n6604 ;
  assign n6609 = n6607 ^ x102 ;
  assign n6610 = n6608 & ~n6609 ;
  assign n6611 = n6610 ^ x102 ;
  assign n6612 = n6611 ^ n6321 ;
  assign n6613 = n6612 ^ n6326 ;
  assign n6614 = ~n6327 & n6613 ;
  assign n6615 = n6614 ^ n6326 ;
  assign n6616 = ~n6322 & n6615 ;
  assign n6617 = n6616 ^ x104 ;
  assign n6618 = n6320 & ~n6617 ;
  assign n6619 = n6317 & ~n6618 ;
  assign n6620 = n6619 ^ n375 ;
  assign n6900 = n6620 ^ x105 ;
  assign n6922 = n6611 ^ x103 ;
  assign n6923 = n6618 & n6922 ;
  assign n6924 = n6923 ^ n6324 ;
  assign n6915 = n6604 ^ x102 ;
  assign n6916 = n6618 & n6915 ;
  assign n6917 = n6916 ^ n6607 ;
  assign n6908 = n6597 ^ x101 ;
  assign n6909 = n6618 & n6908 ;
  assign n6910 = n6909 ^ n6600 ;
  assign n6901 = n6590 ^ x100 ;
  assign n6902 = n6618 & n6901 ;
  assign n6903 = n6902 ^ n6593 ;
  assign n6892 = n6583 ^ x99 ;
  assign n6893 = n6618 & n6892 ;
  assign n6894 = n6893 ^ n6586 ;
  assign n6621 = n6576 ^ x98 ;
  assign n6622 = n6618 & n6621 ;
  assign n6623 = n6622 ^ n6579 ;
  assign n6624 = n6623 ^ x99 ;
  assign n6888 = n6623 ^ x98 ;
  assign n6875 = n6570 ^ x96 ;
  assign n6876 = n6618 & n6875 ;
  assign n6877 = n6876 ^ n6334 ;
  assign n6868 = n6563 ^ x95 ;
  assign n6869 = n6618 & n6868 ;
  assign n6870 = n6869 ^ n6566 ;
  assign n6861 = n6556 ^ x94 ;
  assign n6862 = n6618 & n6861 ;
  assign n6863 = n6862 ^ n6559 ;
  assign n6846 = n6342 ^ x93 ;
  assign n6847 = n6846 ^ x92 ;
  assign n6848 = n6847 ^ n6550 ;
  assign n6849 = n6848 ^ n6846 ;
  assign n6852 = n6846 ^ n3803 ;
  assign n6853 = ~n6849 & ~n6852 ;
  assign n6854 = n6853 ^ n6846 ;
  assign n6855 = n6618 & ~n6854 ;
  assign n6856 = n6855 ^ n6338 ;
  assign n6839 = n6550 ^ x92 ;
  assign n6840 = n6618 & n6839 ;
  assign n6841 = n6840 ^ n6342 ;
  assign n6832 = n6543 ^ x91 ;
  assign n6833 = n6618 & n6832 ;
  assign n6834 = n6833 ^ n6546 ;
  assign n6825 = n6536 ^ x90 ;
  assign n6826 = n6618 & n6825 ;
  assign n6827 = n6826 ^ n6539 ;
  assign n6810 = n6352 ^ x89 ;
  assign n6811 = n6810 ^ x88 ;
  assign n6812 = n6811 ^ n6530 ;
  assign n6813 = n6812 ^ n6810 ;
  assign n6815 = x89 ^ x88 ;
  assign n6816 = n6815 ^ n6810 ;
  assign n6817 = ~n6813 & ~n6816 ;
  assign n6818 = n6817 ^ n6810 ;
  assign n6819 = n6618 & ~n6818 ;
  assign n6820 = n6819 ^ n6348 ;
  assign n6803 = n6530 ^ x88 ;
  assign n6804 = n6618 & n6803 ;
  assign n6805 = n6804 ^ n6352 ;
  assign n6788 = n6362 ^ x87 ;
  assign n6789 = n6788 ^ x86 ;
  assign n6790 = n6789 ^ n6524 ;
  assign n6791 = n6790 ^ n6788 ;
  assign n6794 = n6788 ^ n2532 ;
  assign n6795 = ~n6791 & ~n6794 ;
  assign n6796 = n6795 ^ n6788 ;
  assign n6797 = n6618 & ~n6796 ;
  assign n6798 = n6797 ^ n6358 ;
  assign n6781 = n6524 ^ x86 ;
  assign n6782 = n6618 & n6781 ;
  assign n6783 = n6782 ^ n6362 ;
  assign n6774 = n6517 ^ x85 ;
  assign n6775 = n6618 & n6774 ;
  assign n6776 = n6775 ^ n6520 ;
  assign n6767 = n6510 ^ x84 ;
  assign n6768 = n6618 & n6767 ;
  assign n6769 = n6768 ^ n6513 ;
  assign n6760 = n6503 ^ x83 ;
  assign n6761 = n6618 & n6760 ;
  assign n6762 = n6761 ^ n6506 ;
  assign n6753 = n6496 ^ x82 ;
  assign n6754 = n6618 & n6753 ;
  assign n6755 = n6754 ^ n6499 ;
  assign n6746 = n6489 ^ x81 ;
  assign n6747 = n6618 & n6746 ;
  assign n6748 = n6747 ^ n6492 ;
  assign n6739 = n6482 ^ x80 ;
  assign n6740 = n6618 & n6739 ;
  assign n6741 = n6740 ^ n6485 ;
  assign n6732 = n6475 ^ x79 ;
  assign n6733 = n6618 & n6732 ;
  assign n6734 = n6733 ^ n6478 ;
  assign n6725 = n6468 ^ x78 ;
  assign n6726 = n6618 & n6725 ;
  assign n6727 = n6726 ^ n6471 ;
  assign n6718 = n6461 ^ x77 ;
  assign n6719 = n6618 & n6718 ;
  assign n6720 = n6719 ^ n6464 ;
  assign n6711 = n6454 ^ x76 ;
  assign n6712 = n6618 & n6711 ;
  assign n6713 = n6712 ^ n6457 ;
  assign n6704 = n6448 ^ x75 ;
  assign n6705 = n6618 & n6704 ;
  assign n6706 = n6705 ^ n6450 ;
  assign n6697 = n6441 ^ x74 ;
  assign n6698 = n6618 & n6697 ;
  assign n6699 = n6698 ^ n6444 ;
  assign n6690 = n6426 ^ x73 ;
  assign n6691 = n6618 & n6690 ;
  assign n6692 = n6691 ^ n6437 ;
  assign n6683 = n6419 ^ x72 ;
  assign n6684 = n6618 & n6683 ;
  assign n6685 = n6684 ^ n6422 ;
  assign n6625 = n6412 ^ x71 ;
  assign n6626 = n6618 & n6625 ;
  assign n6627 = n6626 ^ n6415 ;
  assign n6628 = n6627 ^ x72 ;
  assign n6633 = n6627 ^ x71 ;
  assign n6629 = n6405 ^ x70 ;
  assign n6630 = n6618 & n6629 ;
  assign n6631 = n6630 ^ n6408 ;
  assign n6632 = n6631 ^ n6627 ;
  assign n6634 = n6633 ^ n6632 ;
  assign n6670 = n6398 ^ x69 ;
  assign n6671 = n6618 & n6670 ;
  assign n6672 = n6671 ^ n6401 ;
  assign n6663 = n6391 ^ x68 ;
  assign n6664 = n6618 & n6663 ;
  assign n6665 = n6664 ^ n6394 ;
  assign n6656 = n6384 ^ x67 ;
  assign n6657 = n6618 & n6656 ;
  assign n6658 = n6657 ^ n6387 ;
  assign n6649 = n6381 ^ x66 ;
  assign n6650 = n6618 & n6649 ;
  assign n6651 = n6650 ^ n6372 ;
  assign n6635 = n6376 ^ x65 ;
  assign n6636 = n6618 & n6635 ;
  assign n6637 = n6636 ^ n6375 ;
  assign n6638 = n6637 ^ x66 ;
  assign n6639 = ~x22 & x64 ;
  assign n6640 = n6639 ^ x65 ;
  assign n6641 = x64 & n6618 ;
  assign n6642 = n6641 ^ x23 ;
  assign n6643 = n6642 ^ n6639 ;
  assign n6644 = n6640 & n6643 ;
  assign n6645 = n6644 ^ x65 ;
  assign n6646 = n6645 ^ n6637 ;
  assign n6647 = ~n6638 & n6646 ;
  assign n6648 = n6647 ^ x66 ;
  assign n6652 = n6651 ^ n6648 ;
  assign n6653 = n6651 ^ x67 ;
  assign n6654 = n6652 & ~n6653 ;
  assign n6655 = n6654 ^ x67 ;
  assign n6659 = n6658 ^ n6655 ;
  assign n6660 = n6658 ^ x68 ;
  assign n6661 = n6659 & ~n6660 ;
  assign n6662 = n6661 ^ x68 ;
  assign n6666 = n6665 ^ n6662 ;
  assign n6667 = n6665 ^ x69 ;
  assign n6668 = n6666 & ~n6667 ;
  assign n6669 = n6668 ^ x69 ;
  assign n6673 = n6672 ^ n6669 ;
  assign n6674 = n6672 ^ x70 ;
  assign n6675 = n6673 & ~n6674 ;
  assign n6676 = n6675 ^ x70 ;
  assign n6677 = n6676 ^ n6627 ;
  assign n6678 = n6677 ^ n6633 ;
  assign n6679 = ~n6634 & n6678 ;
  assign n6680 = n6679 ^ n6633 ;
  assign n6681 = ~n6628 & n6680 ;
  assign n6682 = n6681 ^ x72 ;
  assign n6686 = n6685 ^ n6682 ;
  assign n6687 = n6685 ^ x73 ;
  assign n6688 = n6686 & ~n6687 ;
  assign n6689 = n6688 ^ x73 ;
  assign n6693 = n6692 ^ n6689 ;
  assign n6694 = n6692 ^ x74 ;
  assign n6695 = n6693 & ~n6694 ;
  assign n6696 = n6695 ^ x74 ;
  assign n6700 = n6699 ^ n6696 ;
  assign n6701 = n6699 ^ x75 ;
  assign n6702 = n6700 & ~n6701 ;
  assign n6703 = n6702 ^ x75 ;
  assign n6707 = n6706 ^ n6703 ;
  assign n6708 = n6706 ^ x76 ;
  assign n6709 = n6707 & ~n6708 ;
  assign n6710 = n6709 ^ x76 ;
  assign n6714 = n6713 ^ n6710 ;
  assign n6715 = n6713 ^ x77 ;
  assign n6716 = n6714 & ~n6715 ;
  assign n6717 = n6716 ^ x77 ;
  assign n6721 = n6720 ^ n6717 ;
  assign n6722 = n6720 ^ x78 ;
  assign n6723 = n6721 & ~n6722 ;
  assign n6724 = n6723 ^ x78 ;
  assign n6728 = n6727 ^ n6724 ;
  assign n6729 = n6727 ^ x79 ;
  assign n6730 = n6728 & ~n6729 ;
  assign n6731 = n6730 ^ x79 ;
  assign n6735 = n6734 ^ n6731 ;
  assign n6736 = n6734 ^ x80 ;
  assign n6737 = n6735 & ~n6736 ;
  assign n6738 = n6737 ^ x80 ;
  assign n6742 = n6741 ^ n6738 ;
  assign n6743 = n6741 ^ x81 ;
  assign n6744 = n6742 & ~n6743 ;
  assign n6745 = n6744 ^ x81 ;
  assign n6749 = n6748 ^ n6745 ;
  assign n6750 = n6748 ^ x82 ;
  assign n6751 = n6749 & ~n6750 ;
  assign n6752 = n6751 ^ x82 ;
  assign n6756 = n6755 ^ n6752 ;
  assign n6757 = n6755 ^ x83 ;
  assign n6758 = n6756 & ~n6757 ;
  assign n6759 = n6758 ^ x83 ;
  assign n6763 = n6762 ^ n6759 ;
  assign n6764 = n6762 ^ x84 ;
  assign n6765 = n6763 & ~n6764 ;
  assign n6766 = n6765 ^ x84 ;
  assign n6770 = n6769 ^ n6766 ;
  assign n6771 = n6769 ^ x85 ;
  assign n6772 = n6770 & ~n6771 ;
  assign n6773 = n6772 ^ x85 ;
  assign n6777 = n6776 ^ n6773 ;
  assign n6778 = n6776 ^ x86 ;
  assign n6779 = n6777 & ~n6778 ;
  assign n6780 = n6779 ^ x86 ;
  assign n6784 = n6783 ^ n6780 ;
  assign n6785 = n6783 ^ x87 ;
  assign n6786 = n6784 & ~n6785 ;
  assign n6787 = n6786 ^ x87 ;
  assign n6799 = n6798 ^ n6787 ;
  assign n6800 = n6798 ^ x88 ;
  assign n6801 = n6799 & ~n6800 ;
  assign n6802 = n6801 ^ x88 ;
  assign n6806 = n6805 ^ n6802 ;
  assign n6807 = n6805 ^ x89 ;
  assign n6808 = n6806 & ~n6807 ;
  assign n6809 = n6808 ^ x89 ;
  assign n6821 = n6820 ^ n6809 ;
  assign n6822 = n6820 ^ x90 ;
  assign n6823 = n6821 & ~n6822 ;
  assign n6824 = n6823 ^ x90 ;
  assign n6828 = n6827 ^ n6824 ;
  assign n6829 = n6827 ^ x91 ;
  assign n6830 = n6828 & ~n6829 ;
  assign n6831 = n6830 ^ x91 ;
  assign n6835 = n6834 ^ n6831 ;
  assign n6836 = n6834 ^ x92 ;
  assign n6837 = n6835 & ~n6836 ;
  assign n6838 = n6837 ^ x92 ;
  assign n6842 = n6841 ^ n6838 ;
  assign n6843 = n6841 ^ x93 ;
  assign n6844 = n6842 & ~n6843 ;
  assign n6845 = n6844 ^ x93 ;
  assign n6857 = n6856 ^ n6845 ;
  assign n6858 = n6856 ^ x94 ;
  assign n6859 = n6857 & ~n6858 ;
  assign n6860 = n6859 ^ x94 ;
  assign n6864 = n6863 ^ n6860 ;
  assign n6865 = n6863 ^ x95 ;
  assign n6866 = n6864 & ~n6865 ;
  assign n6867 = n6866 ^ x95 ;
  assign n6871 = n6870 ^ n6867 ;
  assign n6872 = n6870 ^ x96 ;
  assign n6873 = n6871 & ~n6872 ;
  assign n6874 = n6873 ^ x96 ;
  assign n6878 = n6877 ^ n6874 ;
  assign n6879 = n6877 ^ x97 ;
  assign n6880 = n6878 & ~n6879 ;
  assign n6881 = n6880 ^ x97 ;
  assign n6882 = n6881 ^ x98 ;
  assign n6883 = n6573 ^ x97 ;
  assign n6884 = n6618 & n6883 ;
  assign n6885 = n6884 ^ n6330 ;
  assign n6886 = n6885 ^ n6881 ;
  assign n6887 = n6882 & n6886 ;
  assign n6889 = n6888 ^ n6887 ;
  assign n6890 = ~n6624 & n6889 ;
  assign n6891 = n6890 ^ x99 ;
  assign n6895 = n6894 ^ n6891 ;
  assign n6896 = n6894 ^ x100 ;
  assign n6897 = n6895 & ~n6896 ;
  assign n6898 = n6897 ^ x100 ;
  assign n6904 = n6903 ^ n6898 ;
  assign n6905 = n6903 ^ x101 ;
  assign n6906 = n6904 & ~n6905 ;
  assign n6907 = n6906 ^ x101 ;
  assign n6911 = n6910 ^ n6907 ;
  assign n6912 = n6910 ^ x102 ;
  assign n6913 = n6911 & ~n6912 ;
  assign n6914 = n6913 ^ x102 ;
  assign n6918 = n6917 ^ n6914 ;
  assign n6919 = n6917 ^ x103 ;
  assign n6920 = n6918 & ~n6919 ;
  assign n6921 = n6920 ^ x103 ;
  assign n6925 = n6924 ^ n6921 ;
  assign n7271 = n6921 ^ x104 ;
  assign n6929 = n6925 & n7271 ;
  assign n6926 = x105 ^ x104 ;
  assign n6930 = n6929 ^ n6926 ;
  assign n6933 = ~n6900 & n6930 ;
  assign n6934 = n6933 ^ x105 ;
  assign n6935 = n6319 & ~n6934 ;
  assign n7257 = n6907 ^ x102 ;
  assign n7258 = n6935 & n7257 ;
  assign n7259 = n7258 ^ n6910 ;
  assign n6899 = n6898 ^ x101 ;
  assign n6936 = n6899 & n6935 ;
  assign n6937 = n6936 ^ n6903 ;
  assign n6938 = n6937 ^ x102 ;
  assign n6943 = n6937 ^ x101 ;
  assign n6939 = n6891 ^ x100 ;
  assign n6940 = n6935 & n6939 ;
  assign n6941 = n6940 ^ n6894 ;
  assign n6942 = n6941 ^ n6937 ;
  assign n6944 = n6943 ^ n6942 ;
  assign n6945 = n6887 ^ x99 ;
  assign n6946 = n6945 ^ x98 ;
  assign n6947 = n6935 & n6946 ;
  assign n6948 = n6947 ^ n6623 ;
  assign n6949 = n6948 ^ x100 ;
  assign n6953 = n6948 ^ x99 ;
  assign n6950 = n6882 & n6935 ;
  assign n6951 = n6950 ^ n6885 ;
  assign n6952 = n6951 ^ n6948 ;
  assign n6954 = n6953 ^ n6952 ;
  assign n7238 = n6874 ^ x97 ;
  assign n7239 = n6935 & n7238 ;
  assign n7240 = n7239 ^ n6877 ;
  assign n7231 = n6867 ^ x96 ;
  assign n7232 = n6935 & n7231 ;
  assign n7233 = n7232 ^ n6870 ;
  assign n7224 = n6860 ^ x95 ;
  assign n7225 = n6935 & n7224 ;
  assign n7226 = n7225 ^ n6863 ;
  assign n6955 = n6845 ^ x94 ;
  assign n6956 = n6935 & n6955 ;
  assign n6957 = n6956 ^ n6856 ;
  assign n6958 = n6957 ^ x95 ;
  assign n6963 = n6957 ^ x94 ;
  assign n6959 = n6838 ^ x93 ;
  assign n6960 = n6935 & n6959 ;
  assign n6961 = n6960 ^ n6841 ;
  assign n6962 = n6961 ^ n6957 ;
  assign n6964 = n6963 ^ n6962 ;
  assign n6965 = n6831 ^ x92 ;
  assign n6966 = n6935 & n6965 ;
  assign n6967 = n6966 ^ n6834 ;
  assign n6968 = n6967 ^ x93 ;
  assign n6973 = n6967 ^ x92 ;
  assign n6969 = n6824 ^ x91 ;
  assign n6970 = n6935 & n6969 ;
  assign n6971 = n6970 ^ n6827 ;
  assign n6972 = n6971 ^ n6967 ;
  assign n6974 = n6973 ^ n6972 ;
  assign n7205 = n6809 ^ x90 ;
  assign n7206 = n6935 & n7205 ;
  assign n7207 = n7206 ^ n6820 ;
  assign n7198 = n6802 ^ x89 ;
  assign n7199 = n6935 & n7198 ;
  assign n7200 = n7199 ^ n6805 ;
  assign n7191 = n6787 ^ x88 ;
  assign n7192 = n6935 & n7191 ;
  assign n7193 = n7192 ^ n6798 ;
  assign n7184 = n6780 ^ x87 ;
  assign n7185 = n6935 & n7184 ;
  assign n7186 = n7185 ^ n6783 ;
  assign n7177 = n6773 ^ x86 ;
  assign n7178 = n6935 & n7177 ;
  assign n7179 = n7178 ^ n6776 ;
  assign n7170 = n6766 ^ x85 ;
  assign n7171 = n6935 & n7170 ;
  assign n7172 = n7171 ^ n6769 ;
  assign n7163 = n6759 ^ x84 ;
  assign n7164 = n6935 & n7163 ;
  assign n7165 = n7164 ^ n6762 ;
  assign n7156 = n6752 ^ x83 ;
  assign n7157 = n6935 & n7156 ;
  assign n7158 = n7157 ^ n6755 ;
  assign n7149 = n6745 ^ x82 ;
  assign n7150 = n6935 & n7149 ;
  assign n7151 = n7150 ^ n6748 ;
  assign n7142 = n6738 ^ x81 ;
  assign n7143 = n6935 & n7142 ;
  assign n7144 = n7143 ^ n6741 ;
  assign n7135 = n6731 ^ x80 ;
  assign n7136 = n6935 & n7135 ;
  assign n7137 = n7136 ^ n6734 ;
  assign n7128 = n6724 ^ x79 ;
  assign n7129 = n6935 & n7128 ;
  assign n7130 = n7129 ^ n6727 ;
  assign n7121 = n6717 ^ x78 ;
  assign n7122 = n6935 & n7121 ;
  assign n7123 = n7122 ^ n6720 ;
  assign n7114 = n6710 ^ x77 ;
  assign n7115 = n6935 & n7114 ;
  assign n7116 = n7115 ^ n6713 ;
  assign n7107 = n6703 ^ x76 ;
  assign n7108 = n6935 & n7107 ;
  assign n7109 = n7108 ^ n6706 ;
  assign n7100 = n6696 ^ x75 ;
  assign n7101 = n6935 & n7100 ;
  assign n7102 = n7101 ^ n6699 ;
  assign n7093 = n6689 ^ x74 ;
  assign n7094 = n6935 & n7093 ;
  assign n7095 = n7094 ^ n6692 ;
  assign n7086 = n6682 ^ x73 ;
  assign n7087 = n6935 & n7086 ;
  assign n7088 = n7087 ^ n6685 ;
  assign n7071 = n6631 ^ x72 ;
  assign n7072 = n7071 ^ n6676 ;
  assign n7073 = n7072 ^ x71 ;
  assign n7074 = n7073 ^ n7071 ;
  assign n7076 = n6676 ^ x72 ;
  assign n7077 = n7076 ^ n7071 ;
  assign n7078 = ~n7074 & ~n7077 ;
  assign n7079 = n7078 ^ n7071 ;
  assign n7080 = n6935 & ~n7079 ;
  assign n7081 = n7080 ^ n6627 ;
  assign n7064 = n6676 ^ x71 ;
  assign n7065 = n6935 & n7064 ;
  assign n7066 = n7065 ^ n6631 ;
  assign n7057 = n6669 ^ x70 ;
  assign n7058 = n6935 & n7057 ;
  assign n7059 = n7058 ^ n6672 ;
  assign n7050 = n6662 ^ x69 ;
  assign n7051 = n6935 & n7050 ;
  assign n7052 = n7051 ^ n6665 ;
  assign n7043 = n6655 ^ x68 ;
  assign n7044 = n6935 & n7043 ;
  assign n7045 = n7044 ^ n6658 ;
  assign n7036 = n6648 ^ x67 ;
  assign n7037 = n6935 & n7036 ;
  assign n7038 = n7037 ^ n6651 ;
  assign n7029 = n6645 ^ x66 ;
  assign n7030 = n6935 & n7029 ;
  assign n7031 = n7030 ^ n6637 ;
  assign n6998 = x64 ^ x22 ;
  assign n6999 = n6642 ^ n196 ;
  assign n7000 = n6998 & n6999 ;
  assign n7001 = n6642 ^ x65 ;
  assign n6978 = ~x21 & x65 ;
  assign n7002 = n6978 ^ n6642 ;
  assign n7003 = ~n7001 & ~n7002 ;
  assign n7004 = n7003 ^ x65 ;
  assign n7005 = n7000 & n7004 ;
  assign n7006 = n6935 & n7005 ;
  assign n6977 = ~x22 & x65 ;
  assign n6979 = n6978 ^ x21 ;
  assign n6980 = x22 & ~n6979 ;
  assign n6981 = n6980 ^ x21 ;
  assign n6982 = x64 & ~n6981 ;
  assign n6983 = ~n6977 & ~n6982 ;
  assign n6975 = x64 & n6935 ;
  assign n6976 = ~x21 & n6975 ;
  assign n6984 = n6983 ^ n6976 ;
  assign n6985 = n6642 & n6935 ;
  assign n6986 = n6985 ^ n6642 ;
  assign n6987 = n6986 ^ n6639 ;
  assign n6988 = n6987 ^ n6986 ;
  assign n6993 = ~x65 & n6985 ;
  assign n6994 = ~n6988 & n6993 ;
  assign n6995 = n6994 ^ n6988 ;
  assign n6996 = n6995 ^ n6987 ;
  assign n6997 = n6984 & n6996 ;
  assign n7007 = n7006 ^ n6997 ;
  assign n7023 = ~n6975 & n6977 ;
  assign n7008 = ~n6642 & n6982 ;
  assign n7009 = ~x66 & n6975 ;
  assign n7011 = x65 ^ x21 ;
  assign n7010 = n6981 ^ n6977 ;
  assign n7012 = n7011 ^ n7010 ;
  assign n7013 = ~n7001 & n7012 ;
  assign n7014 = n7009 & n7013 ;
  assign n7015 = n7014 ^ x66 ;
  assign n7016 = n7008 & ~n7015 ;
  assign n7021 = n7016 ^ n7015 ;
  assign n7017 = n6935 & n7016 ;
  assign n7018 = ~x22 & n7017 ;
  assign n7019 = n6978 & n7018 ;
  assign n7020 = n7019 ^ n7017 ;
  assign n7022 = n7021 ^ n7020 ;
  assign n7024 = n6935 ^ n6642 ;
  assign n7025 = ~n7022 & ~n7024 ;
  assign n7026 = n7023 & n7025 ;
  assign n7027 = n7026 ^ n7022 ;
  assign n7028 = ~n7007 & n7027 ;
  assign n7032 = n7031 ^ n7028 ;
  assign n7033 = n7031 ^ x67 ;
  assign n7034 = n7032 & ~n7033 ;
  assign n7035 = n7034 ^ x67 ;
  assign n7039 = n7038 ^ n7035 ;
  assign n7040 = n7038 ^ x68 ;
  assign n7041 = n7039 & ~n7040 ;
  assign n7042 = n7041 ^ x68 ;
  assign n7046 = n7045 ^ n7042 ;
  assign n7047 = n7045 ^ x69 ;
  assign n7048 = n7046 & ~n7047 ;
  assign n7049 = n7048 ^ x69 ;
  assign n7053 = n7052 ^ n7049 ;
  assign n7054 = n7052 ^ x70 ;
  assign n7055 = n7053 & ~n7054 ;
  assign n7056 = n7055 ^ x70 ;
  assign n7060 = n7059 ^ n7056 ;
  assign n7061 = n7059 ^ x71 ;
  assign n7062 = n7060 & ~n7061 ;
  assign n7063 = n7062 ^ x71 ;
  assign n7067 = n7066 ^ n7063 ;
  assign n7068 = n7066 ^ x72 ;
  assign n7069 = n7067 & ~n7068 ;
  assign n7070 = n7069 ^ x72 ;
  assign n7082 = n7081 ^ n7070 ;
  assign n7083 = n7081 ^ x73 ;
  assign n7084 = n7082 & ~n7083 ;
  assign n7085 = n7084 ^ x73 ;
  assign n7089 = n7088 ^ n7085 ;
  assign n7090 = n7088 ^ x74 ;
  assign n7091 = n7089 & ~n7090 ;
  assign n7092 = n7091 ^ x74 ;
  assign n7096 = n7095 ^ n7092 ;
  assign n7097 = n7095 ^ x75 ;
  assign n7098 = n7096 & ~n7097 ;
  assign n7099 = n7098 ^ x75 ;
  assign n7103 = n7102 ^ n7099 ;
  assign n7104 = n7102 ^ x76 ;
  assign n7105 = n7103 & ~n7104 ;
  assign n7106 = n7105 ^ x76 ;
  assign n7110 = n7109 ^ n7106 ;
  assign n7111 = n7109 ^ x77 ;
  assign n7112 = n7110 & ~n7111 ;
  assign n7113 = n7112 ^ x77 ;
  assign n7117 = n7116 ^ n7113 ;
  assign n7118 = n7116 ^ x78 ;
  assign n7119 = n7117 & ~n7118 ;
  assign n7120 = n7119 ^ x78 ;
  assign n7124 = n7123 ^ n7120 ;
  assign n7125 = n7123 ^ x79 ;
  assign n7126 = n7124 & ~n7125 ;
  assign n7127 = n7126 ^ x79 ;
  assign n7131 = n7130 ^ n7127 ;
  assign n7132 = n7130 ^ x80 ;
  assign n7133 = n7131 & ~n7132 ;
  assign n7134 = n7133 ^ x80 ;
  assign n7138 = n7137 ^ n7134 ;
  assign n7139 = n7137 ^ x81 ;
  assign n7140 = n7138 & ~n7139 ;
  assign n7141 = n7140 ^ x81 ;
  assign n7145 = n7144 ^ n7141 ;
  assign n7146 = n7144 ^ x82 ;
  assign n7147 = n7145 & ~n7146 ;
  assign n7148 = n7147 ^ x82 ;
  assign n7152 = n7151 ^ n7148 ;
  assign n7153 = n7151 ^ x83 ;
  assign n7154 = n7152 & ~n7153 ;
  assign n7155 = n7154 ^ x83 ;
  assign n7159 = n7158 ^ n7155 ;
  assign n7160 = n7158 ^ x84 ;
  assign n7161 = n7159 & ~n7160 ;
  assign n7162 = n7161 ^ x84 ;
  assign n7166 = n7165 ^ n7162 ;
  assign n7167 = n7165 ^ x85 ;
  assign n7168 = n7166 & ~n7167 ;
  assign n7169 = n7168 ^ x85 ;
  assign n7173 = n7172 ^ n7169 ;
  assign n7174 = n7172 ^ x86 ;
  assign n7175 = n7173 & ~n7174 ;
  assign n7176 = n7175 ^ x86 ;
  assign n7180 = n7179 ^ n7176 ;
  assign n7181 = n7179 ^ x87 ;
  assign n7182 = n7180 & ~n7181 ;
  assign n7183 = n7182 ^ x87 ;
  assign n7187 = n7186 ^ n7183 ;
  assign n7188 = n7186 ^ x88 ;
  assign n7189 = n7187 & ~n7188 ;
  assign n7190 = n7189 ^ x88 ;
  assign n7194 = n7193 ^ n7190 ;
  assign n7195 = n7193 ^ x89 ;
  assign n7196 = n7194 & ~n7195 ;
  assign n7197 = n7196 ^ x89 ;
  assign n7201 = n7200 ^ n7197 ;
  assign n7202 = n7200 ^ x90 ;
  assign n7203 = n7201 & ~n7202 ;
  assign n7204 = n7203 ^ x90 ;
  assign n7208 = n7207 ^ n7204 ;
  assign n7209 = n7207 ^ x91 ;
  assign n7210 = n7208 & ~n7209 ;
  assign n7211 = n7210 ^ x91 ;
  assign n7212 = n7211 ^ n6967 ;
  assign n7213 = n7212 ^ n6973 ;
  assign n7214 = ~n6974 & n7213 ;
  assign n7215 = n7214 ^ n6973 ;
  assign n7216 = ~n6968 & n7215 ;
  assign n7217 = n7216 ^ x93 ;
  assign n7218 = n7217 ^ n6957 ;
  assign n7219 = n7218 ^ n6963 ;
  assign n7220 = ~n6964 & n7219 ;
  assign n7221 = n7220 ^ n6963 ;
  assign n7222 = ~n6958 & n7221 ;
  assign n7223 = n7222 ^ x95 ;
  assign n7227 = n7226 ^ n7223 ;
  assign n7228 = n7226 ^ x96 ;
  assign n7229 = n7227 & ~n7228 ;
  assign n7230 = n7229 ^ x96 ;
  assign n7234 = n7233 ^ n7230 ;
  assign n7235 = n7233 ^ x97 ;
  assign n7236 = n7234 & ~n7235 ;
  assign n7237 = n7236 ^ x97 ;
  assign n7241 = n7240 ^ n7237 ;
  assign n7242 = n7240 ^ x98 ;
  assign n7243 = n7241 & ~n7242 ;
  assign n7244 = n7243 ^ x98 ;
  assign n7245 = n7244 ^ n6948 ;
  assign n7246 = n7245 ^ n6953 ;
  assign n7247 = ~n6954 & n7246 ;
  assign n7248 = n7247 ^ n6953 ;
  assign n7249 = ~n6949 & n7248 ;
  assign n7250 = n7249 ^ x100 ;
  assign n7251 = n7250 ^ n6937 ;
  assign n7252 = n7251 ^ n6943 ;
  assign n7253 = ~n6944 & n7252 ;
  assign n7254 = n7253 ^ n6943 ;
  assign n7255 = ~n6938 & n7254 ;
  assign n7256 = n7255 ^ x102 ;
  assign n7260 = n7259 ^ n7256 ;
  assign n7261 = n7259 ^ x103 ;
  assign n7262 = n7260 & ~n7261 ;
  assign n7263 = n7262 ^ x103 ;
  assign n7287 = n7263 ^ x104 ;
  assign n7288 = n6620 ^ x106 ;
  assign n7272 = n6935 & n7271 ;
  assign n7273 = n7272 ^ n6924 ;
  assign n7264 = n6914 ^ x103 ;
  assign n7265 = n6935 & n7264 ;
  assign n7266 = n7265 ^ n6917 ;
  assign n7267 = n7266 ^ n7263 ;
  assign n7268 = n7266 ^ x104 ;
  assign n7269 = n7267 & ~n7268 ;
  assign n7270 = n7269 ^ x104 ;
  assign n7274 = n7273 ^ n7270 ;
  assign n7275 = n7273 ^ x105 ;
  assign n7276 = n7274 & ~n7275 ;
  assign n7277 = n7276 ^ x105 ;
  assign n7289 = n7277 ^ n6620 ;
  assign n7290 = n7288 & ~n7289 ;
  assign n7278 = ~x107 & n6318 ;
  assign n7291 = n7290 ^ n7277 ;
  assign n7292 = n7278 & ~n7291 ;
  assign n7293 = n7290 & n7292 ;
  assign n7294 = n6930 & n7293 ;
  assign n7295 = n7294 ^ n7292 ;
  assign n7296 = n7287 & n7295 ;
  assign n7297 = n7296 ^ n7266 ;
  assign n7298 = n7297 ^ x105 ;
  assign n7299 = n7256 ^ x103 ;
  assign n7300 = n7295 & n7299 ;
  assign n7301 = n7300 ^ n7259 ;
  assign n7302 = n7301 ^ x104 ;
  assign n7303 = n6941 ^ x102 ;
  assign n7304 = n7303 ^ x101 ;
  assign n7305 = n7304 ^ n7250 ;
  assign n7306 = n7305 ^ n7303 ;
  assign n7309 = n7303 ^ n6302 ;
  assign n7310 = ~n7306 & ~n7309 ;
  assign n7311 = n7310 ^ n7303 ;
  assign n7312 = n7295 & ~n7311 ;
  assign n7313 = n7312 ^ n6937 ;
  assign n7314 = n7313 ^ x103 ;
  assign n7315 = n7250 ^ x101 ;
  assign n7316 = n7295 & n7315 ;
  assign n7317 = n7316 ^ n6941 ;
  assign n7318 = n7317 ^ x102 ;
  assign n7607 = n6951 ^ x100 ;
  assign n7608 = n7607 ^ x99 ;
  assign n7609 = n7608 ^ n7244 ;
  assign n7610 = n7609 ^ n7607 ;
  assign n7613 = n7607 ^ n5364 ;
  assign n7614 = ~n7610 & ~n7613 ;
  assign n7615 = n7614 ^ n7607 ;
  assign n7616 = n7295 & ~n7615 ;
  assign n7617 = n7616 ^ n6948 ;
  assign n7600 = n7244 ^ x99 ;
  assign n7601 = n7295 & n7600 ;
  assign n7602 = n7601 ^ n6951 ;
  assign n7319 = n7237 ^ x98 ;
  assign n7320 = n7295 & n7319 ;
  assign n7321 = n7320 ^ n7240 ;
  assign n7322 = n7321 ^ x99 ;
  assign n7327 = n7321 ^ x98 ;
  assign n7323 = n7230 ^ x97 ;
  assign n7324 = n7295 & n7323 ;
  assign n7325 = n7324 ^ n7233 ;
  assign n7326 = n7325 ^ n7321 ;
  assign n7328 = n7327 ^ n7326 ;
  assign n7587 = n7223 ^ x96 ;
  assign n7588 = n7295 & n7587 ;
  assign n7589 = n7588 ^ n7226 ;
  assign n7572 = n6961 ^ x95 ;
  assign n7573 = n7572 ^ x94 ;
  assign n7574 = n7573 ^ n7217 ;
  assign n7575 = n7574 ^ n7572 ;
  assign n7577 = x95 ^ x94 ;
  assign n7578 = n7577 ^ n7572 ;
  assign n7579 = ~n7575 & ~n7578 ;
  assign n7580 = n7579 ^ n7572 ;
  assign n7581 = n7295 & ~n7580 ;
  assign n7582 = n7581 ^ n6957 ;
  assign n7565 = n7217 ^ x94 ;
  assign n7566 = n7295 & n7565 ;
  assign n7567 = n7566 ^ n6961 ;
  assign n7550 = n6971 ^ x93 ;
  assign n7551 = n7550 ^ x92 ;
  assign n7552 = n7551 ^ n7211 ;
  assign n7553 = n7552 ^ n7550 ;
  assign n7556 = n7550 ^ n3803 ;
  assign n7557 = ~n7553 & ~n7556 ;
  assign n7558 = n7557 ^ n7550 ;
  assign n7559 = n7295 & ~n7558 ;
  assign n7560 = n7559 ^ n6967 ;
  assign n7543 = n7211 ^ x92 ;
  assign n7544 = n7295 & n7543 ;
  assign n7545 = n7544 ^ n6971 ;
  assign n7536 = n7204 ^ x91 ;
  assign n7537 = n7295 & n7536 ;
  assign n7538 = n7537 ^ n7207 ;
  assign n7529 = n7197 ^ x90 ;
  assign n7530 = n7295 & n7529 ;
  assign n7531 = n7530 ^ n7200 ;
  assign n7522 = n7190 ^ x89 ;
  assign n7523 = n7295 & n7522 ;
  assign n7524 = n7523 ^ n7193 ;
  assign n7515 = n7183 ^ x88 ;
  assign n7516 = n7295 & n7515 ;
  assign n7517 = n7516 ^ n7186 ;
  assign n7508 = n7176 ^ x87 ;
  assign n7509 = n7295 & n7508 ;
  assign n7510 = n7509 ^ n7179 ;
  assign n7501 = n7169 ^ x86 ;
  assign n7502 = n7295 & n7501 ;
  assign n7503 = n7502 ^ n7172 ;
  assign n7494 = n7162 ^ x85 ;
  assign n7495 = n7295 & n7494 ;
  assign n7496 = n7495 ^ n7165 ;
  assign n7487 = n7155 ^ x84 ;
  assign n7488 = n7295 & n7487 ;
  assign n7489 = n7488 ^ n7158 ;
  assign n7480 = n7148 ^ x83 ;
  assign n7481 = n7295 & n7480 ;
  assign n7482 = n7481 ^ n7151 ;
  assign n7473 = n7141 ^ x82 ;
  assign n7474 = n7295 & n7473 ;
  assign n7475 = n7474 ^ n7144 ;
  assign n7329 = n7134 ^ x81 ;
  assign n7330 = n7295 & n7329 ;
  assign n7331 = n7330 ^ n7137 ;
  assign n7332 = n7331 ^ x82 ;
  assign n7337 = n7331 ^ x81 ;
  assign n7333 = n7127 ^ x80 ;
  assign n7334 = n7295 & n7333 ;
  assign n7335 = n7334 ^ n7130 ;
  assign n7336 = n7335 ^ n7331 ;
  assign n7338 = n7337 ^ n7336 ;
  assign n7460 = n7120 ^ x79 ;
  assign n7461 = n7295 & n7460 ;
  assign n7462 = n7461 ^ n7123 ;
  assign n7453 = n7113 ^ x78 ;
  assign n7454 = n7295 & n7453 ;
  assign n7455 = n7454 ^ n7116 ;
  assign n7446 = n7106 ^ x77 ;
  assign n7447 = n7295 & n7446 ;
  assign n7448 = n7447 ^ n7109 ;
  assign n7439 = n7099 ^ x76 ;
  assign n7440 = n7295 & n7439 ;
  assign n7441 = n7440 ^ n7102 ;
  assign n7432 = n7092 ^ x75 ;
  assign n7433 = n7295 & n7432 ;
  assign n7434 = n7433 ^ n7095 ;
  assign n7425 = n7085 ^ x74 ;
  assign n7426 = n7295 & n7425 ;
  assign n7427 = n7426 ^ n7088 ;
  assign n7418 = n7070 ^ x73 ;
  assign n7419 = n7295 & n7418 ;
  assign n7420 = n7419 ^ n7081 ;
  assign n7411 = n7063 ^ x72 ;
  assign n7412 = n7295 & n7411 ;
  assign n7413 = n7412 ^ n7066 ;
  assign n7404 = n7056 ^ x71 ;
  assign n7405 = n7295 & n7404 ;
  assign n7406 = n7405 ^ n7059 ;
  assign n7339 = n7049 ^ x70 ;
  assign n7340 = n7295 & n7339 ;
  assign n7341 = n7340 ^ n7052 ;
  assign n7342 = n7341 ^ x71 ;
  assign n7343 = n7042 ^ x69 ;
  assign n7344 = n7295 & n7343 ;
  assign n7345 = n7344 ^ n7045 ;
  assign n7346 = n7345 ^ x70 ;
  assign n7380 = x65 & n7295 ;
  assign n7370 = x64 & n7295 ;
  assign n7378 = ~x21 & n7370 ;
  assign n7377 = n6975 ^ x22 ;
  assign n7379 = n7378 ^ n7377 ;
  assign n7381 = n7380 ^ n7379 ;
  assign n7372 = ~x20 & x64 ;
  assign n7371 = n7370 ^ x21 ;
  assign n7373 = n7372 ^ n7371 ;
  assign n7374 = n7372 ^ x65 ;
  assign n7375 = n7373 & n7374 ;
  assign n7376 = n7375 ^ x65 ;
  assign n7382 = n7381 ^ n7376 ;
  assign n7383 = n7381 ^ x66 ;
  assign n7384 = n7382 & ~n7383 ;
  assign n7385 = n7384 ^ x66 ;
  assign n7368 = n6640 & n6935 ;
  assign n7362 = x22 & x65 ;
  assign n7353 = n6998 ^ x65 ;
  assign n7354 = n7353 ^ n6935 ;
  assign n7355 = ~n7011 & n7354 ;
  assign n7363 = n7362 ^ n7355 ;
  assign n7364 = ~x64 & n7363 ;
  assign n7358 = x66 ^ x65 ;
  assign n7359 = n7358 ^ n7355 ;
  assign n7365 = n7364 ^ n7359 ;
  assign n7366 = n7295 & n7365 ;
  assign n7367 = n7366 ^ n6642 ;
  assign n7369 = n7368 ^ n7367 ;
  assign n7386 = n7385 ^ n7369 ;
  assign n7387 = n7385 ^ x67 ;
  assign n7388 = n7386 & n7387 ;
  assign n7389 = n7388 ^ x67 ;
  assign n7350 = n7028 ^ x67 ;
  assign n7351 = n7295 & n7350 ;
  assign n7352 = n7351 ^ n7031 ;
  assign n7390 = n7389 ^ n7352 ;
  assign n7391 = n7389 ^ x68 ;
  assign n7392 = n7390 & n7391 ;
  assign n7393 = n7392 ^ x68 ;
  assign n7347 = n7035 ^ x68 ;
  assign n7348 = n7295 & n7347 ;
  assign n7349 = n7348 ^ n7038 ;
  assign n7394 = n7393 ^ n7349 ;
  assign n7395 = n7393 ^ x69 ;
  assign n7396 = n7394 & n7395 ;
  assign n7397 = n7396 ^ x69 ;
  assign n7398 = n7397 ^ n7345 ;
  assign n7399 = ~n7346 & n7398 ;
  assign n7400 = n7399 ^ x70 ;
  assign n7401 = n7400 ^ n7341 ;
  assign n7402 = ~n7342 & n7401 ;
  assign n7403 = n7402 ^ x71 ;
  assign n7407 = n7406 ^ n7403 ;
  assign n7408 = n7406 ^ x72 ;
  assign n7409 = n7407 & ~n7408 ;
  assign n7410 = n7409 ^ x72 ;
  assign n7414 = n7413 ^ n7410 ;
  assign n7415 = n7413 ^ x73 ;
  assign n7416 = n7414 & ~n7415 ;
  assign n7417 = n7416 ^ x73 ;
  assign n7421 = n7420 ^ n7417 ;
  assign n7422 = n7420 ^ x74 ;
  assign n7423 = n7421 & ~n7422 ;
  assign n7424 = n7423 ^ x74 ;
  assign n7428 = n7427 ^ n7424 ;
  assign n7429 = n7427 ^ x75 ;
  assign n7430 = n7428 & ~n7429 ;
  assign n7431 = n7430 ^ x75 ;
  assign n7435 = n7434 ^ n7431 ;
  assign n7436 = n7434 ^ x76 ;
  assign n7437 = n7435 & ~n7436 ;
  assign n7438 = n7437 ^ x76 ;
  assign n7442 = n7441 ^ n7438 ;
  assign n7443 = n7441 ^ x77 ;
  assign n7444 = n7442 & ~n7443 ;
  assign n7445 = n7444 ^ x77 ;
  assign n7449 = n7448 ^ n7445 ;
  assign n7450 = n7448 ^ x78 ;
  assign n7451 = n7449 & ~n7450 ;
  assign n7452 = n7451 ^ x78 ;
  assign n7456 = n7455 ^ n7452 ;
  assign n7457 = n7455 ^ x79 ;
  assign n7458 = n7456 & ~n7457 ;
  assign n7459 = n7458 ^ x79 ;
  assign n7463 = n7462 ^ n7459 ;
  assign n7464 = n7462 ^ x80 ;
  assign n7465 = n7463 & ~n7464 ;
  assign n7466 = n7465 ^ x80 ;
  assign n7467 = n7466 ^ n7331 ;
  assign n7468 = n7467 ^ n7337 ;
  assign n7469 = ~n7338 & n7468 ;
  assign n7470 = n7469 ^ n7337 ;
  assign n7471 = ~n7332 & n7470 ;
  assign n7472 = n7471 ^ x82 ;
  assign n7476 = n7475 ^ n7472 ;
  assign n7477 = n7475 ^ x83 ;
  assign n7478 = n7476 & ~n7477 ;
  assign n7479 = n7478 ^ x83 ;
  assign n7483 = n7482 ^ n7479 ;
  assign n7484 = n7482 ^ x84 ;
  assign n7485 = n7483 & ~n7484 ;
  assign n7486 = n7485 ^ x84 ;
  assign n7490 = n7489 ^ n7486 ;
  assign n7491 = n7489 ^ x85 ;
  assign n7492 = n7490 & ~n7491 ;
  assign n7493 = n7492 ^ x85 ;
  assign n7497 = n7496 ^ n7493 ;
  assign n7498 = n7496 ^ x86 ;
  assign n7499 = n7497 & ~n7498 ;
  assign n7500 = n7499 ^ x86 ;
  assign n7504 = n7503 ^ n7500 ;
  assign n7505 = n7503 ^ x87 ;
  assign n7506 = n7504 & ~n7505 ;
  assign n7507 = n7506 ^ x87 ;
  assign n7511 = n7510 ^ n7507 ;
  assign n7512 = n7510 ^ x88 ;
  assign n7513 = n7511 & ~n7512 ;
  assign n7514 = n7513 ^ x88 ;
  assign n7518 = n7517 ^ n7514 ;
  assign n7519 = n7517 ^ x89 ;
  assign n7520 = n7518 & ~n7519 ;
  assign n7521 = n7520 ^ x89 ;
  assign n7525 = n7524 ^ n7521 ;
  assign n7526 = n7524 ^ x90 ;
  assign n7527 = n7525 & ~n7526 ;
  assign n7528 = n7527 ^ x90 ;
  assign n7532 = n7531 ^ n7528 ;
  assign n7533 = n7531 ^ x91 ;
  assign n7534 = n7532 & ~n7533 ;
  assign n7535 = n7534 ^ x91 ;
  assign n7539 = n7538 ^ n7535 ;
  assign n7540 = n7538 ^ x92 ;
  assign n7541 = n7539 & ~n7540 ;
  assign n7542 = n7541 ^ x92 ;
  assign n7546 = n7545 ^ n7542 ;
  assign n7547 = n7545 ^ x93 ;
  assign n7548 = n7546 & ~n7547 ;
  assign n7549 = n7548 ^ x93 ;
  assign n7561 = n7560 ^ n7549 ;
  assign n7562 = n7560 ^ x94 ;
  assign n7563 = n7561 & ~n7562 ;
  assign n7564 = n7563 ^ x94 ;
  assign n7568 = n7567 ^ n7564 ;
  assign n7569 = n7567 ^ x95 ;
  assign n7570 = n7568 & ~n7569 ;
  assign n7571 = n7570 ^ x95 ;
  assign n7583 = n7582 ^ n7571 ;
  assign n7584 = n7582 ^ x96 ;
  assign n7585 = n7583 & ~n7584 ;
  assign n7586 = n7585 ^ x96 ;
  assign n7590 = n7589 ^ n7586 ;
  assign n7591 = n7589 ^ x97 ;
  assign n7592 = n7590 & ~n7591 ;
  assign n7593 = n7592 ^ x97 ;
  assign n7594 = n7593 ^ n7321 ;
  assign n7595 = n7594 ^ n7327 ;
  assign n7596 = ~n7328 & n7595 ;
  assign n7597 = n7596 ^ n7327 ;
  assign n7598 = ~n7322 & n7597 ;
  assign n7599 = n7598 ^ x99 ;
  assign n7603 = n7602 ^ n7599 ;
  assign n7604 = n7602 ^ x100 ;
  assign n7605 = n7603 & ~n7604 ;
  assign n7606 = n7605 ^ x100 ;
  assign n7618 = n7617 ^ n7606 ;
  assign n7619 = n7617 ^ x101 ;
  assign n7620 = n7618 & ~n7619 ;
  assign n7621 = n7620 ^ x101 ;
  assign n7622 = n7621 ^ n7317 ;
  assign n7623 = ~n7318 & n7622 ;
  assign n7624 = n7623 ^ x102 ;
  assign n7625 = n7624 ^ n7313 ;
  assign n7626 = ~n7314 & n7625 ;
  assign n7627 = n7626 ^ x103 ;
  assign n7628 = n7627 ^ n7301 ;
  assign n7629 = ~n7302 & n7628 ;
  assign n7630 = n7629 ^ x104 ;
  assign n7631 = n7630 ^ n7297 ;
  assign n7632 = ~n7298 & n7631 ;
  assign n7633 = n7632 ^ x105 ;
  assign n7644 = n7633 ^ x106 ;
  assign n7645 = x107 & ~n6620 ;
  assign n7646 = n6318 & ~n7645 ;
  assign n7634 = n7270 ^ x105 ;
  assign n7635 = n7295 & n7634 ;
  assign n7636 = n7635 ^ n7273 ;
  assign n7637 = n7636 ^ n7633 ;
  assign n7638 = n7636 ^ x106 ;
  assign n7639 = n7637 & ~n7638 ;
  assign n7640 = n7639 ^ x106 ;
  assign n7279 = n7277 ^ x106 ;
  assign n7280 = n7278 & ~n7279 ;
  assign n7281 = n6930 & n7280 ;
  assign n7282 = ~n7277 & n7281 ;
  assign n7283 = n7282 ^ n7280 ;
  assign n7284 = n7283 ^ n7278 ;
  assign n7285 = n6620 & ~n7284 ;
  assign n7647 = n7645 ^ n7285 ;
  assign n7648 = n7647 ^ x107 ;
  assign n7649 = n7640 & ~n7648 ;
  assign n7650 = n7646 & ~n7649 ;
  assign n7651 = n7644 & n7650 ;
  assign n7652 = n7651 ^ n7636 ;
  assign n7653 = ~x107 & n7652 ;
  assign n7654 = n7652 ^ x107 ;
  assign n7655 = n7654 ^ n7653 ;
  assign n7984 = n7630 ^ x105 ;
  assign n7985 = n7650 & n7984 ;
  assign n7986 = n7985 ^ n7297 ;
  assign n7977 = n7627 ^ x104 ;
  assign n7978 = n7650 & n7977 ;
  assign n7979 = n7978 ^ n7301 ;
  assign n7970 = n7624 ^ x103 ;
  assign n7971 = n7650 & n7970 ;
  assign n7972 = n7971 ^ n7313 ;
  assign n7963 = n7621 ^ x102 ;
  assign n7964 = n7650 & n7963 ;
  assign n7965 = n7964 ^ n7317 ;
  assign n7956 = n7606 ^ x101 ;
  assign n7957 = n7650 & n7956 ;
  assign n7958 = n7957 ^ n7617 ;
  assign n7949 = n7599 ^ x100 ;
  assign n7950 = n7650 & n7949 ;
  assign n7951 = n7950 ^ n7602 ;
  assign n7934 = n7325 ^ x99 ;
  assign n7935 = n7934 ^ x98 ;
  assign n7936 = n7935 ^ n7593 ;
  assign n7937 = n7936 ^ n7934 ;
  assign n7939 = x99 ^ x98 ;
  assign n7940 = n7939 ^ n7934 ;
  assign n7941 = ~n7937 & ~n7940 ;
  assign n7942 = n7941 ^ n7934 ;
  assign n7943 = n7650 & ~n7942 ;
  assign n7944 = n7943 ^ n7321 ;
  assign n7927 = n7593 ^ x98 ;
  assign n7928 = n7650 & n7927 ;
  assign n7929 = n7928 ^ n7325 ;
  assign n7920 = n7586 ^ x97 ;
  assign n7921 = n7650 & n7920 ;
  assign n7922 = n7921 ^ n7589 ;
  assign n7913 = n7571 ^ x96 ;
  assign n7914 = n7650 & n7913 ;
  assign n7915 = n7914 ^ n7582 ;
  assign n7906 = n7564 ^ x95 ;
  assign n7907 = n7650 & n7906 ;
  assign n7908 = n7907 ^ n7567 ;
  assign n7899 = n7549 ^ x94 ;
  assign n7900 = n7650 & n7899 ;
  assign n7901 = n7900 ^ n7560 ;
  assign n7892 = n7542 ^ x93 ;
  assign n7893 = n7650 & n7892 ;
  assign n7894 = n7893 ^ n7545 ;
  assign n7885 = n7535 ^ x92 ;
  assign n7886 = n7650 & n7885 ;
  assign n7887 = n7886 ^ n7538 ;
  assign n7878 = n7528 ^ x91 ;
  assign n7879 = n7650 & n7878 ;
  assign n7880 = n7879 ^ n7531 ;
  assign n7871 = n7521 ^ x90 ;
  assign n7872 = n7650 & n7871 ;
  assign n7873 = n7872 ^ n7524 ;
  assign n7864 = n7514 ^ x89 ;
  assign n7865 = n7650 & n7864 ;
  assign n7866 = n7865 ^ n7517 ;
  assign n7857 = n7507 ^ x88 ;
  assign n7858 = n7650 & n7857 ;
  assign n7859 = n7858 ^ n7510 ;
  assign n7850 = n7500 ^ x87 ;
  assign n7851 = n7650 & n7850 ;
  assign n7852 = n7851 ^ n7503 ;
  assign n7843 = n7493 ^ x86 ;
  assign n7844 = n7650 & n7843 ;
  assign n7845 = n7844 ^ n7496 ;
  assign n7836 = n7486 ^ x85 ;
  assign n7837 = n7650 & n7836 ;
  assign n7838 = n7837 ^ n7489 ;
  assign n7829 = n7479 ^ x84 ;
  assign n7830 = n7650 & n7829 ;
  assign n7831 = n7830 ^ n7482 ;
  assign n7822 = n7472 ^ x83 ;
  assign n7823 = n7650 & n7822 ;
  assign n7824 = n7823 ^ n7475 ;
  assign n7807 = n7335 ^ x82 ;
  assign n7808 = n7807 ^ x81 ;
  assign n7809 = n7808 ^ n7466 ;
  assign n7810 = n7809 ^ n7807 ;
  assign n7813 = n7807 ^ n5543 ;
  assign n7814 = ~n7810 & ~n7813 ;
  assign n7815 = n7814 ^ n7807 ;
  assign n7816 = n7650 & ~n7815 ;
  assign n7817 = n7816 ^ n7331 ;
  assign n7800 = n7466 ^ x81 ;
  assign n7801 = n7650 & n7800 ;
  assign n7802 = n7801 ^ n7335 ;
  assign n7793 = n7459 ^ x80 ;
  assign n7794 = n7650 & n7793 ;
  assign n7795 = n7794 ^ n7462 ;
  assign n7786 = n7452 ^ x79 ;
  assign n7787 = n7650 & n7786 ;
  assign n7788 = n7787 ^ n7455 ;
  assign n7779 = n7445 ^ x78 ;
  assign n7780 = n7650 & n7779 ;
  assign n7781 = n7780 ^ n7448 ;
  assign n7772 = n7438 ^ x77 ;
  assign n7773 = n7650 & n7772 ;
  assign n7774 = n7773 ^ n7441 ;
  assign n7765 = n7431 ^ x76 ;
  assign n7766 = n7650 & n7765 ;
  assign n7767 = n7766 ^ n7434 ;
  assign n7758 = n7424 ^ x75 ;
  assign n7759 = n7650 & n7758 ;
  assign n7760 = n7759 ^ n7427 ;
  assign n7751 = n7417 ^ x74 ;
  assign n7752 = n7650 & n7751 ;
  assign n7753 = n7752 ^ n7420 ;
  assign n7744 = n7410 ^ x73 ;
  assign n7745 = n7650 & n7744 ;
  assign n7746 = n7745 ^ n7413 ;
  assign n7737 = n7403 ^ x72 ;
  assign n7738 = n7650 & n7737 ;
  assign n7739 = n7738 ^ n7406 ;
  assign n7730 = n7400 ^ x71 ;
  assign n7731 = n7650 & n7730 ;
  assign n7732 = n7731 ^ n7341 ;
  assign n7723 = n7397 ^ x70 ;
  assign n7724 = n7650 & n7723 ;
  assign n7725 = n7724 ^ n7345 ;
  assign n7717 = n7395 & n7650 ;
  assign n7718 = n7717 ^ n7349 ;
  assign n7711 = n7391 & n7650 ;
  assign n7712 = n7711 ^ n7352 ;
  assign n7705 = n7387 & n7650 ;
  assign n7706 = n7705 ^ n7369 ;
  assign n7698 = n7376 ^ x66 ;
  assign n7699 = n7650 & n7698 ;
  assign n7700 = n7699 ^ n7381 ;
  assign n7667 = x64 & n7650 ;
  assign n7668 = n7371 ^ x65 ;
  assign n7669 = n7372 & ~n7668 ;
  assign n7670 = n7667 & n7669 ;
  assign n7672 = ~x19 & x65 ;
  assign n7673 = n7670 & n7672 ;
  assign n7664 = x20 & ~x21 ;
  assign n7665 = n926 & n7650 ;
  assign n7666 = n7664 & n7665 ;
  assign n7671 = n7670 ^ n7666 ;
  assign n7674 = n7673 ^ n7671 ;
  assign n7656 = ~x20 & x65 ;
  assign n7657 = n7371 & ~n7656 ;
  assign n7658 = ~x19 & x64 ;
  assign n7659 = n7658 ^ n7650 ;
  assign n7660 = n7658 ^ n7374 ;
  assign n7661 = n7659 & ~n7660 ;
  assign n7662 = n7661 ^ n7650 ;
  assign n7663 = n7657 & ~n7662 ;
  assign n7675 = n7674 ^ n7663 ;
  assign n7676 = n7371 ^ x19 ;
  assign n7677 = n7676 ^ x65 ;
  assign n7678 = n7677 ^ n7650 ;
  assign n7679 = n7678 ^ x20 ;
  assign n7680 = ~x19 & ~n7679 ;
  assign n7681 = n7680 ^ n7676 ;
  assign n7682 = n7650 ^ x20 ;
  assign n7683 = n7676 ^ x20 ;
  assign n7684 = n7683 ^ x19 ;
  assign n7685 = ~n7682 & ~n7684 ;
  assign n7686 = n7685 ^ n7676 ;
  assign n7687 = ~n7681 & ~n7686 ;
  assign n7688 = n7687 ^ n7676 ;
  assign n7689 = ~x66 & ~n7667 ;
  assign n7690 = n7650 ^ n7371 ;
  assign n7691 = n7656 & ~n7690 ;
  assign n7692 = n7689 & n7691 ;
  assign n7693 = n7692 ^ x66 ;
  assign n7694 = x64 & ~n7693 ;
  assign n7695 = ~n7688 & n7694 ;
  assign n7696 = n7695 ^ n7693 ;
  assign n7697 = ~n7675 & n7696 ;
  assign n7701 = n7700 ^ n7697 ;
  assign n7702 = n7700 ^ x67 ;
  assign n7703 = n7701 & ~n7702 ;
  assign n7704 = n7703 ^ x67 ;
  assign n7707 = n7706 ^ n7704 ;
  assign n7708 = n7706 ^ x68 ;
  assign n7709 = n7707 & ~n7708 ;
  assign n7710 = n7709 ^ x68 ;
  assign n7713 = n7712 ^ n7710 ;
  assign n7714 = n7712 ^ x69 ;
  assign n7715 = n7713 & ~n7714 ;
  assign n7716 = n7715 ^ x69 ;
  assign n7719 = n7718 ^ n7716 ;
  assign n7720 = n7718 ^ x70 ;
  assign n7721 = n7719 & ~n7720 ;
  assign n7722 = n7721 ^ x70 ;
  assign n7726 = n7725 ^ n7722 ;
  assign n7727 = n7725 ^ x71 ;
  assign n7728 = n7726 & ~n7727 ;
  assign n7729 = n7728 ^ x71 ;
  assign n7733 = n7732 ^ n7729 ;
  assign n7734 = n7732 ^ x72 ;
  assign n7735 = n7733 & ~n7734 ;
  assign n7736 = n7735 ^ x72 ;
  assign n7740 = n7739 ^ n7736 ;
  assign n7741 = n7739 ^ x73 ;
  assign n7742 = n7740 & ~n7741 ;
  assign n7743 = n7742 ^ x73 ;
  assign n7747 = n7746 ^ n7743 ;
  assign n7748 = n7746 ^ x74 ;
  assign n7749 = n7747 & ~n7748 ;
  assign n7750 = n7749 ^ x74 ;
  assign n7754 = n7753 ^ n7750 ;
  assign n7755 = n7753 ^ x75 ;
  assign n7756 = n7754 & ~n7755 ;
  assign n7757 = n7756 ^ x75 ;
  assign n7761 = n7760 ^ n7757 ;
  assign n7762 = n7760 ^ x76 ;
  assign n7763 = n7761 & ~n7762 ;
  assign n7764 = n7763 ^ x76 ;
  assign n7768 = n7767 ^ n7764 ;
  assign n7769 = n7767 ^ x77 ;
  assign n7770 = n7768 & ~n7769 ;
  assign n7771 = n7770 ^ x77 ;
  assign n7775 = n7774 ^ n7771 ;
  assign n7776 = n7774 ^ x78 ;
  assign n7777 = n7775 & ~n7776 ;
  assign n7778 = n7777 ^ x78 ;
  assign n7782 = n7781 ^ n7778 ;
  assign n7783 = n7781 ^ x79 ;
  assign n7784 = n7782 & ~n7783 ;
  assign n7785 = n7784 ^ x79 ;
  assign n7789 = n7788 ^ n7785 ;
  assign n7790 = n7788 ^ x80 ;
  assign n7791 = n7789 & ~n7790 ;
  assign n7792 = n7791 ^ x80 ;
  assign n7796 = n7795 ^ n7792 ;
  assign n7797 = n7795 ^ x81 ;
  assign n7798 = n7796 & ~n7797 ;
  assign n7799 = n7798 ^ x81 ;
  assign n7803 = n7802 ^ n7799 ;
  assign n7804 = n7802 ^ x82 ;
  assign n7805 = n7803 & ~n7804 ;
  assign n7806 = n7805 ^ x82 ;
  assign n7818 = n7817 ^ n7806 ;
  assign n7819 = n7817 ^ x83 ;
  assign n7820 = n7818 & ~n7819 ;
  assign n7821 = n7820 ^ x83 ;
  assign n7825 = n7824 ^ n7821 ;
  assign n7826 = n7824 ^ x84 ;
  assign n7827 = n7825 & ~n7826 ;
  assign n7828 = n7827 ^ x84 ;
  assign n7832 = n7831 ^ n7828 ;
  assign n7833 = n7831 ^ x85 ;
  assign n7834 = n7832 & ~n7833 ;
  assign n7835 = n7834 ^ x85 ;
  assign n7839 = n7838 ^ n7835 ;
  assign n7840 = n7838 ^ x86 ;
  assign n7841 = n7839 & ~n7840 ;
  assign n7842 = n7841 ^ x86 ;
  assign n7846 = n7845 ^ n7842 ;
  assign n7847 = n7845 ^ x87 ;
  assign n7848 = n7846 & ~n7847 ;
  assign n7849 = n7848 ^ x87 ;
  assign n7853 = n7852 ^ n7849 ;
  assign n7854 = n7852 ^ x88 ;
  assign n7855 = n7853 & ~n7854 ;
  assign n7856 = n7855 ^ x88 ;
  assign n7860 = n7859 ^ n7856 ;
  assign n7861 = n7859 ^ x89 ;
  assign n7862 = n7860 & ~n7861 ;
  assign n7863 = n7862 ^ x89 ;
  assign n7867 = n7866 ^ n7863 ;
  assign n7868 = n7866 ^ x90 ;
  assign n7869 = n7867 & ~n7868 ;
  assign n7870 = n7869 ^ x90 ;
  assign n7874 = n7873 ^ n7870 ;
  assign n7875 = n7873 ^ x91 ;
  assign n7876 = n7874 & ~n7875 ;
  assign n7877 = n7876 ^ x91 ;
  assign n7881 = n7880 ^ n7877 ;
  assign n7882 = n7880 ^ x92 ;
  assign n7883 = n7881 & ~n7882 ;
  assign n7884 = n7883 ^ x92 ;
  assign n7888 = n7887 ^ n7884 ;
  assign n7889 = n7887 ^ x93 ;
  assign n7890 = n7888 & ~n7889 ;
  assign n7891 = n7890 ^ x93 ;
  assign n7895 = n7894 ^ n7891 ;
  assign n7896 = n7894 ^ x94 ;
  assign n7897 = n7895 & ~n7896 ;
  assign n7898 = n7897 ^ x94 ;
  assign n7902 = n7901 ^ n7898 ;
  assign n7903 = n7901 ^ x95 ;
  assign n7904 = n7902 & ~n7903 ;
  assign n7905 = n7904 ^ x95 ;
  assign n7909 = n7908 ^ n7905 ;
  assign n7910 = n7908 ^ x96 ;
  assign n7911 = n7909 & ~n7910 ;
  assign n7912 = n7911 ^ x96 ;
  assign n7916 = n7915 ^ n7912 ;
  assign n7917 = n7915 ^ x97 ;
  assign n7918 = n7916 & ~n7917 ;
  assign n7919 = n7918 ^ x97 ;
  assign n7923 = n7922 ^ n7919 ;
  assign n7924 = n7922 ^ x98 ;
  assign n7925 = n7923 & ~n7924 ;
  assign n7926 = n7925 ^ x98 ;
  assign n7930 = n7929 ^ n7926 ;
  assign n7931 = n7929 ^ x99 ;
  assign n7932 = n7930 & ~n7931 ;
  assign n7933 = n7932 ^ x99 ;
  assign n7945 = n7944 ^ n7933 ;
  assign n7946 = n7944 ^ x100 ;
  assign n7947 = n7945 & ~n7946 ;
  assign n7948 = n7947 ^ x100 ;
  assign n7952 = n7951 ^ n7948 ;
  assign n7953 = n7951 ^ x101 ;
  assign n7954 = n7952 & ~n7953 ;
  assign n7955 = n7954 ^ x101 ;
  assign n7959 = n7958 ^ n7955 ;
  assign n7960 = n7958 ^ x102 ;
  assign n7961 = n7959 & ~n7960 ;
  assign n7962 = n7961 ^ x102 ;
  assign n7966 = n7965 ^ n7962 ;
  assign n7967 = n7965 ^ x103 ;
  assign n7968 = n7966 & ~n7967 ;
  assign n7969 = n7968 ^ x103 ;
  assign n7973 = n7972 ^ n7969 ;
  assign n7974 = n7972 ^ x104 ;
  assign n7975 = n7973 & ~n7974 ;
  assign n7976 = n7975 ^ x104 ;
  assign n7980 = n7979 ^ n7976 ;
  assign n7981 = n7979 ^ x105 ;
  assign n7982 = n7980 & ~n7981 ;
  assign n7983 = n7982 ^ x105 ;
  assign n7987 = n7986 ^ n7983 ;
  assign n7988 = n7986 ^ x106 ;
  assign n7989 = n7987 & ~n7988 ;
  assign n7990 = n7989 ^ x106 ;
  assign n7991 = ~n7655 & ~n7990 ;
  assign n7992 = ~n7653 & ~n7991 ;
  assign n8000 = n6318 & ~n7992 ;
  assign n8001 = n148 & n6620 ;
  assign n8002 = n7653 ^ n7284 ;
  assign n8003 = n8002 ^ n7653 ;
  assign n7641 = n7640 ^ x107 ;
  assign n7642 = ~x108 & ~n7641 ;
  assign n8004 = n7653 ^ n7642 ;
  assign n8005 = n8004 ^ n7653 ;
  assign n8006 = ~n8003 & n8005 ;
  assign n8007 = n8006 ^ n7653 ;
  assign n8008 = ~n7991 & ~n8007 ;
  assign n8009 = n8001 & ~n8008 ;
  assign n8010 = ~n8000 & ~n8009 ;
  assign n8340 = n7990 ^ x107 ;
  assign n8341 = ~n8010 & n8340 ;
  assign n8342 = n8341 ^ n7652 ;
  assign n7999 = n7983 ^ x106 ;
  assign n8011 = n7999 & ~n8010 ;
  assign n8012 = n8011 ^ n7986 ;
  assign n8013 = n8012 ^ x107 ;
  assign n8018 = n8012 ^ x106 ;
  assign n8014 = n7976 ^ x105 ;
  assign n8015 = ~n8010 & n8014 ;
  assign n8016 = n8015 ^ n7979 ;
  assign n8017 = n8016 ^ n8012 ;
  assign n8019 = n8018 ^ n8017 ;
  assign n8327 = n7969 ^ x104 ;
  assign n8328 = ~n8010 & n8327 ;
  assign n8329 = n8328 ^ n7972 ;
  assign n8320 = n7962 ^ x103 ;
  assign n8321 = ~n8010 & n8320 ;
  assign n8322 = n8321 ^ n7965 ;
  assign n8313 = n7955 ^ x102 ;
  assign n8314 = ~n8010 & n8313 ;
  assign n8315 = n8314 ^ n7958 ;
  assign n8306 = n7948 ^ x101 ;
  assign n8307 = ~n8010 & n8306 ;
  assign n8308 = n8307 ^ n7951 ;
  assign n8299 = n7933 ^ x100 ;
  assign n8300 = ~n8010 & n8299 ;
  assign n8301 = n8300 ^ n7944 ;
  assign n8020 = n7926 ^ x99 ;
  assign n8021 = ~n8010 & n8020 ;
  assign n8022 = n8021 ^ n7929 ;
  assign n8023 = n8022 ^ x100 ;
  assign n8028 = n8022 ^ x99 ;
  assign n8024 = n7919 ^ x98 ;
  assign n8025 = ~n8010 & n8024 ;
  assign n8026 = n8025 ^ n7922 ;
  assign n8027 = n8026 ^ n8022 ;
  assign n8029 = n8028 ^ n8027 ;
  assign n8030 = n7912 ^ x97 ;
  assign n8031 = ~n8010 & n8030 ;
  assign n8032 = n8031 ^ n7915 ;
  assign n8033 = n8032 ^ x98 ;
  assign n8038 = n8032 ^ x97 ;
  assign n8034 = n7905 ^ x96 ;
  assign n8035 = ~n8010 & n8034 ;
  assign n8036 = n8035 ^ n7908 ;
  assign n8037 = n8036 ^ n8032 ;
  assign n8039 = n8038 ^ n8037 ;
  assign n8280 = n7898 ^ x95 ;
  assign n8281 = ~n8010 & n8280 ;
  assign n8282 = n8281 ^ n7901 ;
  assign n8273 = n7891 ^ x94 ;
  assign n8274 = ~n8010 & n8273 ;
  assign n8275 = n8274 ^ n7894 ;
  assign n8266 = n7884 ^ x93 ;
  assign n8267 = ~n8010 & n8266 ;
  assign n8268 = n8267 ^ n7887 ;
  assign n8259 = n7877 ^ x92 ;
  assign n8260 = ~n8010 & n8259 ;
  assign n8261 = n8260 ^ n7880 ;
  assign n8252 = n7870 ^ x91 ;
  assign n8253 = ~n8010 & n8252 ;
  assign n8254 = n8253 ^ n7873 ;
  assign n8245 = n7863 ^ x90 ;
  assign n8246 = ~n8010 & n8245 ;
  assign n8247 = n8246 ^ n7866 ;
  assign n8238 = n7856 ^ x89 ;
  assign n8239 = ~n8010 & n8238 ;
  assign n8240 = n8239 ^ n7859 ;
  assign n8231 = n7849 ^ x88 ;
  assign n8232 = ~n8010 & n8231 ;
  assign n8233 = n8232 ^ n7852 ;
  assign n8224 = n7842 ^ x87 ;
  assign n8225 = ~n8010 & n8224 ;
  assign n8226 = n8225 ^ n7845 ;
  assign n8217 = n7835 ^ x86 ;
  assign n8218 = ~n8010 & n8217 ;
  assign n8219 = n8218 ^ n7838 ;
  assign n8210 = n7828 ^ x85 ;
  assign n8211 = ~n8010 & n8210 ;
  assign n8212 = n8211 ^ n7831 ;
  assign n8203 = n7821 ^ x84 ;
  assign n8204 = ~n8010 & n8203 ;
  assign n8205 = n8204 ^ n7824 ;
  assign n8196 = n7806 ^ x83 ;
  assign n8197 = ~n8010 & n8196 ;
  assign n8198 = n8197 ^ n7817 ;
  assign n8189 = n7799 ^ x82 ;
  assign n8190 = ~n8010 & n8189 ;
  assign n8191 = n8190 ^ n7802 ;
  assign n8182 = n7792 ^ x81 ;
  assign n8183 = ~n8010 & n8182 ;
  assign n8184 = n8183 ^ n7795 ;
  assign n8040 = n7785 ^ x80 ;
  assign n8041 = ~n8010 & n8040 ;
  assign n8042 = n8041 ^ n7788 ;
  assign n8043 = n8042 ^ x81 ;
  assign n8048 = n8042 ^ x80 ;
  assign n8044 = n7778 ^ x79 ;
  assign n8045 = ~n8010 & n8044 ;
  assign n8046 = n8045 ^ n7781 ;
  assign n8047 = n8046 ^ n8042 ;
  assign n8049 = n8048 ^ n8047 ;
  assign n8169 = n7771 ^ x78 ;
  assign n8170 = ~n8010 & n8169 ;
  assign n8171 = n8170 ^ n7774 ;
  assign n8162 = n7764 ^ x77 ;
  assign n8163 = ~n8010 & n8162 ;
  assign n8164 = n8163 ^ n7767 ;
  assign n8155 = n7757 ^ x76 ;
  assign n8156 = ~n8010 & n8155 ;
  assign n8157 = n8156 ^ n7760 ;
  assign n8148 = n7750 ^ x75 ;
  assign n8149 = ~n8010 & n8148 ;
  assign n8150 = n8149 ^ n7753 ;
  assign n8141 = n7743 ^ x74 ;
  assign n8142 = ~n8010 & n8141 ;
  assign n8143 = n8142 ^ n7746 ;
  assign n8134 = n7736 ^ x73 ;
  assign n8135 = ~n8010 & n8134 ;
  assign n8136 = n8135 ^ n7739 ;
  assign n8127 = n7729 ^ x72 ;
  assign n8128 = ~n8010 & n8127 ;
  assign n8129 = n8128 ^ n7732 ;
  assign n8120 = n7722 ^ x71 ;
  assign n8121 = ~n8010 & n8120 ;
  assign n8122 = n8121 ^ n7725 ;
  assign n8113 = n7716 ^ x70 ;
  assign n8114 = ~n8010 & n8113 ;
  assign n8115 = n8114 ^ n7718 ;
  assign n8106 = n7710 ^ x69 ;
  assign n8107 = ~n8010 & n8106 ;
  assign n8108 = n8107 ^ n7712 ;
  assign n8099 = n7704 ^ x68 ;
  assign n8100 = ~n8010 & n8099 ;
  assign n8101 = n8100 ^ n7706 ;
  assign n8092 = n7697 ^ x67 ;
  assign n8093 = ~n8010 & n8092 ;
  assign n8094 = n8093 ^ n7700 ;
  assign n8051 = n7658 ^ x65 ;
  assign n8052 = ~n8010 & n8051 ;
  assign n8050 = n7667 ^ x20 ;
  assign n8053 = n8052 ^ n8050 ;
  assign n8054 = n8053 ^ x66 ;
  assign n8062 = x19 & x65 ;
  assign n8059 = x65 ^ x18 ;
  assign n8055 = x64 ^ x19 ;
  assign n8056 = n8055 ^ x65 ;
  assign n8060 = n8056 ^ n8010 ;
  assign n8061 = ~n8059 & ~n8060 ;
  assign n8063 = n8062 ^ n8061 ;
  assign n8064 = x64 & n8063 ;
  assign n8065 = n8064 ^ n8062 ;
  assign n8066 = n8065 ^ x65 ;
  assign n8067 = n8066 ^ n8053 ;
  assign n8068 = ~n8054 & n8067 ;
  assign n8069 = n8068 ^ x66 ;
  assign n8070 = n8069 ^ x67 ;
  assign n8087 = n7374 & n7650 ;
  assign n8081 = x20 & x65 ;
  assign n8071 = x65 ^ x19 ;
  assign n8072 = x64 ^ x20 ;
  assign n8073 = n8072 ^ x65 ;
  assign n8074 = n8073 ^ n7650 ;
  assign n8075 = ~n8071 & n8074 ;
  assign n8082 = n8081 ^ n8075 ;
  assign n8083 = ~x64 & n8082 ;
  assign n8078 = n8075 ^ n7358 ;
  assign n8084 = n8083 ^ n8078 ;
  assign n8085 = ~n8010 & n8084 ;
  assign n8086 = n8085 ^ n7371 ;
  assign n8088 = n8087 ^ n8086 ;
  assign n8089 = n8088 ^ n8069 ;
  assign n8090 = n8070 & n8089 ;
  assign n8091 = n8090 ^ x67 ;
  assign n8095 = n8094 ^ n8091 ;
  assign n8096 = n8094 ^ x68 ;
  assign n8097 = n8095 & ~n8096 ;
  assign n8098 = n8097 ^ x68 ;
  assign n8102 = n8101 ^ n8098 ;
  assign n8103 = n8101 ^ x69 ;
  assign n8104 = n8102 & ~n8103 ;
  assign n8105 = n8104 ^ x69 ;
  assign n8109 = n8108 ^ n8105 ;
  assign n8110 = n8108 ^ x70 ;
  assign n8111 = n8109 & ~n8110 ;
  assign n8112 = n8111 ^ x70 ;
  assign n8116 = n8115 ^ n8112 ;
  assign n8117 = n8115 ^ x71 ;
  assign n8118 = n8116 & ~n8117 ;
  assign n8119 = n8118 ^ x71 ;
  assign n8123 = n8122 ^ n8119 ;
  assign n8124 = n8122 ^ x72 ;
  assign n8125 = n8123 & ~n8124 ;
  assign n8126 = n8125 ^ x72 ;
  assign n8130 = n8129 ^ n8126 ;
  assign n8131 = n8129 ^ x73 ;
  assign n8132 = n8130 & ~n8131 ;
  assign n8133 = n8132 ^ x73 ;
  assign n8137 = n8136 ^ n8133 ;
  assign n8138 = n8136 ^ x74 ;
  assign n8139 = n8137 & ~n8138 ;
  assign n8140 = n8139 ^ x74 ;
  assign n8144 = n8143 ^ n8140 ;
  assign n8145 = n8143 ^ x75 ;
  assign n8146 = n8144 & ~n8145 ;
  assign n8147 = n8146 ^ x75 ;
  assign n8151 = n8150 ^ n8147 ;
  assign n8152 = n8150 ^ x76 ;
  assign n8153 = n8151 & ~n8152 ;
  assign n8154 = n8153 ^ x76 ;
  assign n8158 = n8157 ^ n8154 ;
  assign n8159 = n8157 ^ x77 ;
  assign n8160 = n8158 & ~n8159 ;
  assign n8161 = n8160 ^ x77 ;
  assign n8165 = n8164 ^ n8161 ;
  assign n8166 = n8164 ^ x78 ;
  assign n8167 = n8165 & ~n8166 ;
  assign n8168 = n8167 ^ x78 ;
  assign n8172 = n8171 ^ n8168 ;
  assign n8173 = n8171 ^ x79 ;
  assign n8174 = n8172 & ~n8173 ;
  assign n8175 = n8174 ^ x79 ;
  assign n8176 = n8175 ^ n8042 ;
  assign n8177 = n8176 ^ n8048 ;
  assign n8178 = ~n8049 & n8177 ;
  assign n8179 = n8178 ^ n8048 ;
  assign n8180 = ~n8043 & n8179 ;
  assign n8181 = n8180 ^ x81 ;
  assign n8185 = n8184 ^ n8181 ;
  assign n8186 = n8184 ^ x82 ;
  assign n8187 = n8185 & ~n8186 ;
  assign n8188 = n8187 ^ x82 ;
  assign n8192 = n8191 ^ n8188 ;
  assign n8193 = n8191 ^ x83 ;
  assign n8194 = n8192 & ~n8193 ;
  assign n8195 = n8194 ^ x83 ;
  assign n8199 = n8198 ^ n8195 ;
  assign n8200 = n8198 ^ x84 ;
  assign n8201 = n8199 & ~n8200 ;
  assign n8202 = n8201 ^ x84 ;
  assign n8206 = n8205 ^ n8202 ;
  assign n8207 = n8205 ^ x85 ;
  assign n8208 = n8206 & ~n8207 ;
  assign n8209 = n8208 ^ x85 ;
  assign n8213 = n8212 ^ n8209 ;
  assign n8214 = n8212 ^ x86 ;
  assign n8215 = n8213 & ~n8214 ;
  assign n8216 = n8215 ^ x86 ;
  assign n8220 = n8219 ^ n8216 ;
  assign n8221 = n8219 ^ x87 ;
  assign n8222 = n8220 & ~n8221 ;
  assign n8223 = n8222 ^ x87 ;
  assign n8227 = n8226 ^ n8223 ;
  assign n8228 = n8226 ^ x88 ;
  assign n8229 = n8227 & ~n8228 ;
  assign n8230 = n8229 ^ x88 ;
  assign n8234 = n8233 ^ n8230 ;
  assign n8235 = n8233 ^ x89 ;
  assign n8236 = n8234 & ~n8235 ;
  assign n8237 = n8236 ^ x89 ;
  assign n8241 = n8240 ^ n8237 ;
  assign n8242 = n8240 ^ x90 ;
  assign n8243 = n8241 & ~n8242 ;
  assign n8244 = n8243 ^ x90 ;
  assign n8248 = n8247 ^ n8244 ;
  assign n8249 = n8247 ^ x91 ;
  assign n8250 = n8248 & ~n8249 ;
  assign n8251 = n8250 ^ x91 ;
  assign n8255 = n8254 ^ n8251 ;
  assign n8256 = n8254 ^ x92 ;
  assign n8257 = n8255 & ~n8256 ;
  assign n8258 = n8257 ^ x92 ;
  assign n8262 = n8261 ^ n8258 ;
  assign n8263 = n8261 ^ x93 ;
  assign n8264 = n8262 & ~n8263 ;
  assign n8265 = n8264 ^ x93 ;
  assign n8269 = n8268 ^ n8265 ;
  assign n8270 = n8268 ^ x94 ;
  assign n8271 = n8269 & ~n8270 ;
  assign n8272 = n8271 ^ x94 ;
  assign n8276 = n8275 ^ n8272 ;
  assign n8277 = n8275 ^ x95 ;
  assign n8278 = n8276 & ~n8277 ;
  assign n8279 = n8278 ^ x95 ;
  assign n8283 = n8282 ^ n8279 ;
  assign n8284 = n8282 ^ x96 ;
  assign n8285 = n8283 & ~n8284 ;
  assign n8286 = n8285 ^ x96 ;
  assign n8287 = n8286 ^ n8032 ;
  assign n8288 = n8287 ^ n8038 ;
  assign n8289 = ~n8039 & n8288 ;
  assign n8290 = n8289 ^ n8038 ;
  assign n8291 = ~n8033 & n8290 ;
  assign n8292 = n8291 ^ x98 ;
  assign n8293 = n8292 ^ n8022 ;
  assign n8294 = n8293 ^ n8028 ;
  assign n8295 = ~n8029 & n8294 ;
  assign n8296 = n8295 ^ n8028 ;
  assign n8297 = ~n8023 & n8296 ;
  assign n8298 = n8297 ^ x100 ;
  assign n8302 = n8301 ^ n8298 ;
  assign n8303 = n8301 ^ x101 ;
  assign n8304 = n8302 & ~n8303 ;
  assign n8305 = n8304 ^ x101 ;
  assign n8309 = n8308 ^ n8305 ;
  assign n8310 = n8308 ^ x102 ;
  assign n8311 = n8309 & ~n8310 ;
  assign n8312 = n8311 ^ x102 ;
  assign n8316 = n8315 ^ n8312 ;
  assign n8317 = n8315 ^ x103 ;
  assign n8318 = n8316 & ~n8317 ;
  assign n8319 = n8318 ^ x103 ;
  assign n8323 = n8322 ^ n8319 ;
  assign n8324 = n8322 ^ x104 ;
  assign n8325 = n8323 & ~n8324 ;
  assign n8326 = n8325 ^ x104 ;
  assign n8330 = n8329 ^ n8326 ;
  assign n8331 = n8329 ^ x105 ;
  assign n8332 = n8330 & ~n8331 ;
  assign n8333 = n8332 ^ x105 ;
  assign n8334 = n8333 ^ n8012 ;
  assign n8335 = n8334 ^ n8018 ;
  assign n8336 = ~n8019 & n8335 ;
  assign n8337 = n8336 ^ n8018 ;
  assign n8338 = ~n8013 & n8337 ;
  assign n8339 = n8338 ^ x107 ;
  assign n8343 = n8342 ^ n8339 ;
  assign n8344 = n8342 ^ x108 ;
  assign n8345 = n8343 & ~n8344 ;
  assign n8346 = n8345 ^ x108 ;
  assign n8347 = n8346 ^ x109 ;
  assign n7286 = n148 & n7285 ;
  assign n7643 = n7642 ^ x108 ;
  assign n7995 = n7643 & ~n7992 ;
  assign n7996 = n7995 ^ x108 ;
  assign n7997 = n7286 & ~n7996 ;
  assign n7998 = n7997 ^ n7285 ;
  assign n8348 = n147 & n7998 ;
  assign n8349 = n8347 & n8348 ;
  assign n8350 = n8349 ^ n7998 ;
  assign n8351 = n146 & n8350 ;
  assign n8353 = x109 & n147 ;
  assign n8354 = ~n6620 & n8353 ;
  assign n8355 = n8354 ^ n147 ;
  assign n8356 = n8346 & n8355 ;
  assign n8357 = n8354 ^ x109 ;
  assign n8358 = n8357 ^ n7998 ;
  assign n8359 = n8356 & ~n8358 ;
  assign n8360 = n8359 ^ n8355 ;
  assign n8705 = n8339 ^ x108 ;
  assign n8706 = n8360 & n8705 ;
  assign n8707 = n8706 ^ n8342 ;
  assign n8690 = n8016 ^ x107 ;
  assign n8691 = n8690 ^ x106 ;
  assign n8692 = n8691 ^ n8333 ;
  assign n8693 = n8692 ^ n8690 ;
  assign n8695 = x107 ^ x106 ;
  assign n8696 = n8695 ^ n8690 ;
  assign n8697 = ~n8693 & ~n8696 ;
  assign n8698 = n8697 ^ n8690 ;
  assign n8699 = n8360 & ~n8698 ;
  assign n8700 = n8699 ^ n8012 ;
  assign n8683 = n8333 ^ x106 ;
  assign n8684 = n8360 & n8683 ;
  assign n8685 = n8684 ^ n8016 ;
  assign n8676 = n8326 ^ x105 ;
  assign n8677 = n8360 & n8676 ;
  assign n8678 = n8677 ^ n8329 ;
  assign n8669 = n8319 ^ x104 ;
  assign n8670 = n8360 & n8669 ;
  assign n8671 = n8670 ^ n8322 ;
  assign n8662 = n8312 ^ x103 ;
  assign n8663 = n8360 & n8662 ;
  assign n8664 = n8663 ^ n8315 ;
  assign n8655 = n8305 ^ x102 ;
  assign n8656 = n8360 & n8655 ;
  assign n8657 = n8656 ^ n8308 ;
  assign n8648 = n8298 ^ x101 ;
  assign n8649 = n8360 & n8648 ;
  assign n8650 = n8649 ^ n8301 ;
  assign n8633 = n8026 ^ x100 ;
  assign n8634 = n8633 ^ x99 ;
  assign n8635 = n8634 ^ n8292 ;
  assign n8636 = n8635 ^ n8633 ;
  assign n8639 = n8633 ^ n5364 ;
  assign n8640 = ~n8636 & ~n8639 ;
  assign n8641 = n8640 ^ n8633 ;
  assign n8642 = n8360 & ~n8641 ;
  assign n8643 = n8642 ^ n8022 ;
  assign n8626 = n8292 ^ x99 ;
  assign n8627 = n8360 & n8626 ;
  assign n8628 = n8627 ^ n8026 ;
  assign n8611 = n8036 ^ x98 ;
  assign n8612 = n8611 ^ x97 ;
  assign n8613 = n8612 ^ n8286 ;
  assign n8614 = n8613 ^ n8611 ;
  assign n8617 = n8611 ^ n5357 ;
  assign n8618 = ~n8614 & ~n8617 ;
  assign n8619 = n8618 ^ n8611 ;
  assign n8620 = n8360 & ~n8619 ;
  assign n8621 = n8620 ^ n8032 ;
  assign n8604 = n8286 ^ x97 ;
  assign n8605 = n8360 & n8604 ;
  assign n8606 = n8605 ^ n8036 ;
  assign n8597 = n8279 ^ x96 ;
  assign n8598 = n8360 & n8597 ;
  assign n8599 = n8598 ^ n8282 ;
  assign n8590 = n8272 ^ x95 ;
  assign n8591 = n8360 & n8590 ;
  assign n8592 = n8591 ^ n8275 ;
  assign n8583 = n8265 ^ x94 ;
  assign n8584 = n8360 & n8583 ;
  assign n8585 = n8584 ^ n8268 ;
  assign n8576 = n8258 ^ x93 ;
  assign n8577 = n8360 & n8576 ;
  assign n8578 = n8577 ^ n8261 ;
  assign n8569 = n8251 ^ x92 ;
  assign n8570 = n8360 & n8569 ;
  assign n8571 = n8570 ^ n8254 ;
  assign n8562 = n8244 ^ x91 ;
  assign n8563 = n8360 & n8562 ;
  assign n8564 = n8563 ^ n8247 ;
  assign n8555 = n8237 ^ x90 ;
  assign n8556 = n8360 & n8555 ;
  assign n8557 = n8556 ^ n8240 ;
  assign n8548 = n8230 ^ x89 ;
  assign n8549 = n8360 & n8548 ;
  assign n8550 = n8549 ^ n8233 ;
  assign n8541 = n8223 ^ x88 ;
  assign n8542 = n8360 & n8541 ;
  assign n8543 = n8542 ^ n8226 ;
  assign n8534 = n8216 ^ x87 ;
  assign n8535 = n8360 & n8534 ;
  assign n8536 = n8535 ^ n8219 ;
  assign n8527 = n8209 ^ x86 ;
  assign n8528 = n8360 & n8527 ;
  assign n8529 = n8528 ^ n8212 ;
  assign n8352 = n8202 ^ x85 ;
  assign n8361 = n8352 & n8360 ;
  assign n8362 = n8361 ^ n8205 ;
  assign n8363 = n8362 ^ x86 ;
  assign n8368 = n8362 ^ x85 ;
  assign n8364 = n8195 ^ x84 ;
  assign n8365 = n8360 & n8364 ;
  assign n8366 = n8365 ^ n8198 ;
  assign n8367 = n8366 ^ n8362 ;
  assign n8369 = n8368 ^ n8367 ;
  assign n8514 = n8188 ^ x83 ;
  assign n8515 = n8360 & n8514 ;
  assign n8516 = n8515 ^ n8191 ;
  assign n8507 = n8181 ^ x82 ;
  assign n8508 = n8360 & n8507 ;
  assign n8509 = n8508 ^ n8184 ;
  assign n8492 = n8046 ^ x81 ;
  assign n8493 = n8492 ^ x80 ;
  assign n8494 = n8493 ^ n8175 ;
  assign n8495 = n8494 ^ n8492 ;
  assign n8497 = x81 ^ x80 ;
  assign n8498 = n8497 ^ n8492 ;
  assign n8499 = ~n8495 & ~n8498 ;
  assign n8500 = n8499 ^ n8492 ;
  assign n8501 = n8360 & ~n8500 ;
  assign n8502 = n8501 ^ n8042 ;
  assign n8485 = n8175 ^ x80 ;
  assign n8486 = n8360 & n8485 ;
  assign n8487 = n8486 ^ n8046 ;
  assign n8478 = n8168 ^ x79 ;
  assign n8479 = n8360 & n8478 ;
  assign n8480 = n8479 ^ n8171 ;
  assign n8471 = n8161 ^ x78 ;
  assign n8472 = n8360 & n8471 ;
  assign n8473 = n8472 ^ n8164 ;
  assign n8464 = n8154 ^ x77 ;
  assign n8465 = n8360 & n8464 ;
  assign n8466 = n8465 ^ n8157 ;
  assign n8457 = n8147 ^ x76 ;
  assign n8458 = n8360 & n8457 ;
  assign n8459 = n8458 ^ n8150 ;
  assign n8450 = n8140 ^ x75 ;
  assign n8451 = n8360 & n8450 ;
  assign n8452 = n8451 ^ n8143 ;
  assign n8443 = n8133 ^ x74 ;
  assign n8444 = n8360 & n8443 ;
  assign n8445 = n8444 ^ n8136 ;
  assign n8436 = n8126 ^ x73 ;
  assign n8437 = n8360 & n8436 ;
  assign n8438 = n8437 ^ n8129 ;
  assign n8429 = n8119 ^ x72 ;
  assign n8430 = n8360 & n8429 ;
  assign n8431 = n8430 ^ n8122 ;
  assign n8422 = n8112 ^ x71 ;
  assign n8423 = n8360 & n8422 ;
  assign n8424 = n8423 ^ n8115 ;
  assign n8415 = n8105 ^ x70 ;
  assign n8416 = n8360 & n8415 ;
  assign n8417 = n8416 ^ n8108 ;
  assign n8408 = n8098 ^ x69 ;
  assign n8409 = n8360 & n8408 ;
  assign n8410 = n8409 ^ n8101 ;
  assign n8401 = n8091 ^ x68 ;
  assign n8402 = n8360 & n8401 ;
  assign n8403 = n8402 ^ n8094 ;
  assign n8395 = n8070 & n8360 ;
  assign n8396 = n8395 ^ n8088 ;
  assign n8388 = n8066 ^ x66 ;
  assign n8389 = n8360 & n8388 ;
  assign n8390 = n8389 ^ n8053 ;
  assign n8370 = ~x17 & x64 ;
  assign n8371 = n8370 ^ x65 ;
  assign n8372 = x64 & n8360 ;
  assign n8373 = n8372 ^ x18 ;
  assign n8374 = n8373 ^ n8370 ;
  assign n8375 = n8371 & n8374 ;
  assign n8376 = n8375 ^ x65 ;
  assign n8377 = n8376 ^ x66 ;
  assign n8383 = x64 & ~n8010 ;
  assign n8379 = ~x18 & x64 ;
  assign n8380 = n8379 ^ x65 ;
  assign n8381 = n8360 & n8380 ;
  assign n8382 = n8381 ^ x19 ;
  assign n8384 = n8383 ^ n8382 ;
  assign n8385 = n8384 ^ n8376 ;
  assign n8386 = n8377 & n8385 ;
  assign n8387 = n8386 ^ x66 ;
  assign n8391 = n8390 ^ n8387 ;
  assign n8392 = n8390 ^ x67 ;
  assign n8393 = n8391 & ~n8392 ;
  assign n8394 = n8393 ^ x67 ;
  assign n8397 = n8396 ^ n8394 ;
  assign n8398 = n8396 ^ x68 ;
  assign n8399 = n8397 & ~n8398 ;
  assign n8400 = n8399 ^ x68 ;
  assign n8404 = n8403 ^ n8400 ;
  assign n8405 = n8403 ^ x69 ;
  assign n8406 = n8404 & ~n8405 ;
  assign n8407 = n8406 ^ x69 ;
  assign n8411 = n8410 ^ n8407 ;
  assign n8412 = n8410 ^ x70 ;
  assign n8413 = n8411 & ~n8412 ;
  assign n8414 = n8413 ^ x70 ;
  assign n8418 = n8417 ^ n8414 ;
  assign n8419 = n8417 ^ x71 ;
  assign n8420 = n8418 & ~n8419 ;
  assign n8421 = n8420 ^ x71 ;
  assign n8425 = n8424 ^ n8421 ;
  assign n8426 = n8424 ^ x72 ;
  assign n8427 = n8425 & ~n8426 ;
  assign n8428 = n8427 ^ x72 ;
  assign n8432 = n8431 ^ n8428 ;
  assign n8433 = n8431 ^ x73 ;
  assign n8434 = n8432 & ~n8433 ;
  assign n8435 = n8434 ^ x73 ;
  assign n8439 = n8438 ^ n8435 ;
  assign n8440 = n8438 ^ x74 ;
  assign n8441 = n8439 & ~n8440 ;
  assign n8442 = n8441 ^ x74 ;
  assign n8446 = n8445 ^ n8442 ;
  assign n8447 = n8445 ^ x75 ;
  assign n8448 = n8446 & ~n8447 ;
  assign n8449 = n8448 ^ x75 ;
  assign n8453 = n8452 ^ n8449 ;
  assign n8454 = n8452 ^ x76 ;
  assign n8455 = n8453 & ~n8454 ;
  assign n8456 = n8455 ^ x76 ;
  assign n8460 = n8459 ^ n8456 ;
  assign n8461 = n8459 ^ x77 ;
  assign n8462 = n8460 & ~n8461 ;
  assign n8463 = n8462 ^ x77 ;
  assign n8467 = n8466 ^ n8463 ;
  assign n8468 = n8466 ^ x78 ;
  assign n8469 = n8467 & ~n8468 ;
  assign n8470 = n8469 ^ x78 ;
  assign n8474 = n8473 ^ n8470 ;
  assign n8475 = n8473 ^ x79 ;
  assign n8476 = n8474 & ~n8475 ;
  assign n8477 = n8476 ^ x79 ;
  assign n8481 = n8480 ^ n8477 ;
  assign n8482 = n8480 ^ x80 ;
  assign n8483 = n8481 & ~n8482 ;
  assign n8484 = n8483 ^ x80 ;
  assign n8488 = n8487 ^ n8484 ;
  assign n8489 = n8487 ^ x81 ;
  assign n8490 = n8488 & ~n8489 ;
  assign n8491 = n8490 ^ x81 ;
  assign n8503 = n8502 ^ n8491 ;
  assign n8504 = n8502 ^ x82 ;
  assign n8505 = n8503 & ~n8504 ;
  assign n8506 = n8505 ^ x82 ;
  assign n8510 = n8509 ^ n8506 ;
  assign n8511 = n8509 ^ x83 ;
  assign n8512 = n8510 & ~n8511 ;
  assign n8513 = n8512 ^ x83 ;
  assign n8517 = n8516 ^ n8513 ;
  assign n8518 = n8516 ^ x84 ;
  assign n8519 = n8517 & ~n8518 ;
  assign n8520 = n8519 ^ x84 ;
  assign n8521 = n8520 ^ n8362 ;
  assign n8522 = n8521 ^ n8368 ;
  assign n8523 = ~n8369 & n8522 ;
  assign n8524 = n8523 ^ n8368 ;
  assign n8525 = ~n8363 & n8524 ;
  assign n8526 = n8525 ^ x86 ;
  assign n8530 = n8529 ^ n8526 ;
  assign n8531 = n8529 ^ x87 ;
  assign n8532 = n8530 & ~n8531 ;
  assign n8533 = n8532 ^ x87 ;
  assign n8537 = n8536 ^ n8533 ;
  assign n8538 = n8536 ^ x88 ;
  assign n8539 = n8537 & ~n8538 ;
  assign n8540 = n8539 ^ x88 ;
  assign n8544 = n8543 ^ n8540 ;
  assign n8545 = n8543 ^ x89 ;
  assign n8546 = n8544 & ~n8545 ;
  assign n8547 = n8546 ^ x89 ;
  assign n8551 = n8550 ^ n8547 ;
  assign n8552 = n8550 ^ x90 ;
  assign n8553 = n8551 & ~n8552 ;
  assign n8554 = n8553 ^ x90 ;
  assign n8558 = n8557 ^ n8554 ;
  assign n8559 = n8557 ^ x91 ;
  assign n8560 = n8558 & ~n8559 ;
  assign n8561 = n8560 ^ x91 ;
  assign n8565 = n8564 ^ n8561 ;
  assign n8566 = n8564 ^ x92 ;
  assign n8567 = n8565 & ~n8566 ;
  assign n8568 = n8567 ^ x92 ;
  assign n8572 = n8571 ^ n8568 ;
  assign n8573 = n8571 ^ x93 ;
  assign n8574 = n8572 & ~n8573 ;
  assign n8575 = n8574 ^ x93 ;
  assign n8579 = n8578 ^ n8575 ;
  assign n8580 = n8578 ^ x94 ;
  assign n8581 = n8579 & ~n8580 ;
  assign n8582 = n8581 ^ x94 ;
  assign n8586 = n8585 ^ n8582 ;
  assign n8587 = n8585 ^ x95 ;
  assign n8588 = n8586 & ~n8587 ;
  assign n8589 = n8588 ^ x95 ;
  assign n8593 = n8592 ^ n8589 ;
  assign n8594 = n8592 ^ x96 ;
  assign n8595 = n8593 & ~n8594 ;
  assign n8596 = n8595 ^ x96 ;
  assign n8600 = n8599 ^ n8596 ;
  assign n8601 = n8599 ^ x97 ;
  assign n8602 = n8600 & ~n8601 ;
  assign n8603 = n8602 ^ x97 ;
  assign n8607 = n8606 ^ n8603 ;
  assign n8608 = n8606 ^ x98 ;
  assign n8609 = n8607 & ~n8608 ;
  assign n8610 = n8609 ^ x98 ;
  assign n8622 = n8621 ^ n8610 ;
  assign n8623 = n8621 ^ x99 ;
  assign n8624 = n8622 & ~n8623 ;
  assign n8625 = n8624 ^ x99 ;
  assign n8629 = n8628 ^ n8625 ;
  assign n8630 = n8628 ^ x100 ;
  assign n8631 = n8629 & ~n8630 ;
  assign n8632 = n8631 ^ x100 ;
  assign n8644 = n8643 ^ n8632 ;
  assign n8645 = n8643 ^ x101 ;
  assign n8646 = n8644 & ~n8645 ;
  assign n8647 = n8646 ^ x101 ;
  assign n8651 = n8650 ^ n8647 ;
  assign n8652 = n8650 ^ x102 ;
  assign n8653 = n8651 & ~n8652 ;
  assign n8654 = n8653 ^ x102 ;
  assign n8658 = n8657 ^ n8654 ;
  assign n8659 = n8657 ^ x103 ;
  assign n8660 = n8658 & ~n8659 ;
  assign n8661 = n8660 ^ x103 ;
  assign n8665 = n8664 ^ n8661 ;
  assign n8666 = n8664 ^ x104 ;
  assign n8667 = n8665 & ~n8666 ;
  assign n8668 = n8667 ^ x104 ;
  assign n8672 = n8671 ^ n8668 ;
  assign n8673 = n8671 ^ x105 ;
  assign n8674 = n8672 & ~n8673 ;
  assign n8675 = n8674 ^ x105 ;
  assign n8679 = n8678 ^ n8675 ;
  assign n8680 = n8678 ^ x106 ;
  assign n8681 = n8679 & ~n8680 ;
  assign n8682 = n8681 ^ x106 ;
  assign n8686 = n8685 ^ n8682 ;
  assign n8687 = n8685 ^ x107 ;
  assign n8688 = n8686 & ~n8687 ;
  assign n8689 = n8688 ^ x107 ;
  assign n8701 = n8700 ^ n8689 ;
  assign n8702 = n8700 ^ x108 ;
  assign n8703 = n8701 & ~n8702 ;
  assign n8704 = n8703 ^ x108 ;
  assign n8708 = n8707 ^ n8704 ;
  assign n9090 = n8704 ^ x109 ;
  assign n8712 = n8708 & n9090 ;
  assign n8709 = x110 ^ x109 ;
  assign n8713 = n8712 ^ n8709 ;
  assign n8714 = n8351 & n8713 ;
  assign n8715 = n8714 ^ n8350 ;
  assign n8716 = n141 & n144 ;
  assign n8718 = n8350 ^ x110 ;
  assign n8721 = n8713 & ~n8718 ;
  assign n8722 = n8721 ^ x110 ;
  assign n8723 = n146 & ~n8722 ;
  assign n9080 = n8689 ^ x108 ;
  assign n9081 = n8723 & n9080 ;
  assign n9082 = n9081 ^ n8700 ;
  assign n9073 = n8682 ^ x107 ;
  assign n9074 = n8723 & n9073 ;
  assign n9075 = n9074 ^ n8685 ;
  assign n8717 = n8675 ^ x106 ;
  assign n8724 = n8717 & n8723 ;
  assign n8725 = n8724 ^ n8678 ;
  assign n8726 = n8725 ^ x107 ;
  assign n8727 = n8668 ^ x105 ;
  assign n8728 = n8723 & n8727 ;
  assign n8729 = n8728 ^ n8671 ;
  assign n8730 = n8729 ^ x106 ;
  assign n9060 = n8661 ^ x104 ;
  assign n9061 = n8723 & n9060 ;
  assign n9062 = n9061 ^ n8664 ;
  assign n9053 = n8654 ^ x103 ;
  assign n9054 = n8723 & n9053 ;
  assign n9055 = n9054 ^ n8657 ;
  assign n9046 = n8647 ^ x102 ;
  assign n9047 = n8723 & n9046 ;
  assign n9048 = n9047 ^ n8650 ;
  assign n9039 = n8632 ^ x101 ;
  assign n9040 = n8723 & n9039 ;
  assign n9041 = n9040 ^ n8643 ;
  assign n8731 = n8625 ^ x100 ;
  assign n8732 = n8723 & n8731 ;
  assign n8733 = n8732 ^ n8628 ;
  assign n8734 = n8733 ^ x101 ;
  assign n8735 = n8610 ^ x99 ;
  assign n8736 = n8723 & n8735 ;
  assign n8737 = n8736 ^ n8621 ;
  assign n8738 = n8737 ^ x100 ;
  assign n9026 = n8603 ^ x98 ;
  assign n9027 = n8723 & n9026 ;
  assign n9028 = n9027 ^ n8606 ;
  assign n9019 = n8596 ^ x97 ;
  assign n9020 = n8723 & n9019 ;
  assign n9021 = n9020 ^ n8599 ;
  assign n9012 = n8589 ^ x96 ;
  assign n9013 = n8723 & n9012 ;
  assign n9014 = n9013 ^ n8592 ;
  assign n9005 = n8582 ^ x95 ;
  assign n9006 = n8723 & n9005 ;
  assign n9007 = n9006 ^ n8585 ;
  assign n8739 = n8575 ^ x94 ;
  assign n8740 = n8723 & n8739 ;
  assign n8741 = n8740 ^ n8578 ;
  assign n8742 = n8741 ^ x95 ;
  assign n8743 = n8568 ^ x93 ;
  assign n8744 = n8723 & n8743 ;
  assign n8745 = n8744 ^ n8571 ;
  assign n8746 = n8745 ^ x94 ;
  assign n8992 = n8561 ^ x92 ;
  assign n8993 = n8723 & n8992 ;
  assign n8994 = n8993 ^ n8564 ;
  assign n8985 = n8554 ^ x91 ;
  assign n8986 = n8723 & n8985 ;
  assign n8987 = n8986 ^ n8557 ;
  assign n8978 = n8547 ^ x90 ;
  assign n8979 = n8723 & n8978 ;
  assign n8980 = n8979 ^ n8550 ;
  assign n8971 = n8540 ^ x89 ;
  assign n8972 = n8723 & n8971 ;
  assign n8973 = n8972 ^ n8543 ;
  assign n8964 = n8533 ^ x88 ;
  assign n8965 = n8723 & n8964 ;
  assign n8966 = n8965 ^ n8536 ;
  assign n8957 = n8526 ^ x87 ;
  assign n8958 = n8723 & n8957 ;
  assign n8959 = n8958 ^ n8529 ;
  assign n8942 = n8366 ^ x86 ;
  assign n8943 = n8942 ^ n8520 ;
  assign n8944 = n8943 ^ x85 ;
  assign n8945 = n8944 ^ n8942 ;
  assign n8947 = n8520 ^ x86 ;
  assign n8948 = n8947 ^ n8942 ;
  assign n8949 = ~n8945 & ~n8948 ;
  assign n8950 = n8949 ^ n8942 ;
  assign n8951 = n8723 & ~n8950 ;
  assign n8952 = n8951 ^ n8362 ;
  assign n8935 = n8520 ^ x85 ;
  assign n8936 = n8723 & n8935 ;
  assign n8937 = n8936 ^ n8366 ;
  assign n8928 = n8513 ^ x84 ;
  assign n8929 = n8723 & n8928 ;
  assign n8930 = n8929 ^ n8516 ;
  assign n8921 = n8506 ^ x83 ;
  assign n8922 = n8723 & n8921 ;
  assign n8923 = n8922 ^ n8509 ;
  assign n8914 = n8491 ^ x82 ;
  assign n8915 = n8723 & n8914 ;
  assign n8916 = n8915 ^ n8502 ;
  assign n8907 = n8484 ^ x81 ;
  assign n8908 = n8723 & n8907 ;
  assign n8909 = n8908 ^ n8487 ;
  assign n8900 = n8477 ^ x80 ;
  assign n8901 = n8723 & n8900 ;
  assign n8902 = n8901 ^ n8480 ;
  assign n8893 = n8470 ^ x79 ;
  assign n8894 = n8723 & n8893 ;
  assign n8895 = n8894 ^ n8473 ;
  assign n8886 = n8463 ^ x78 ;
  assign n8887 = n8723 & n8886 ;
  assign n8888 = n8887 ^ n8466 ;
  assign n8879 = n8456 ^ x77 ;
  assign n8880 = n8723 & n8879 ;
  assign n8881 = n8880 ^ n8459 ;
  assign n8872 = n8449 ^ x76 ;
  assign n8873 = n8723 & n8872 ;
  assign n8874 = n8873 ^ n8452 ;
  assign n8865 = n8442 ^ x75 ;
  assign n8866 = n8723 & n8865 ;
  assign n8867 = n8866 ^ n8445 ;
  assign n8858 = n8435 ^ x74 ;
  assign n8859 = n8723 & n8858 ;
  assign n8860 = n8859 ^ n8438 ;
  assign n8851 = n8428 ^ x73 ;
  assign n8852 = n8723 & n8851 ;
  assign n8853 = n8852 ^ n8431 ;
  assign n8844 = n8421 ^ x72 ;
  assign n8845 = n8723 & n8844 ;
  assign n8846 = n8845 ^ n8424 ;
  assign n8837 = n8414 ^ x71 ;
  assign n8838 = n8723 & n8837 ;
  assign n8839 = n8838 ^ n8417 ;
  assign n8830 = n8407 ^ x70 ;
  assign n8831 = n8723 & n8830 ;
  assign n8832 = n8831 ^ n8410 ;
  assign n8747 = n8400 ^ x69 ;
  assign n8748 = n8723 & n8747 ;
  assign n8749 = n8748 ^ n8403 ;
  assign n8750 = n8749 ^ x70 ;
  assign n8751 = n8394 ^ x68 ;
  assign n8752 = n8723 & n8751 ;
  assign n8753 = n8752 ^ n8396 ;
  assign n8754 = n8753 ^ x69 ;
  assign n8817 = n8387 ^ x67 ;
  assign n8818 = n8723 & n8817 ;
  assign n8819 = n8818 ^ n8390 ;
  assign n8811 = n8377 & n8723 ;
  assign n8812 = n8811 ^ n8384 ;
  assign n8765 = ~x16 & x64 ;
  assign n8766 = x17 & ~x65 ;
  assign n8767 = n8766 ^ n8723 ;
  assign n8768 = n8765 & ~n8767 ;
  assign n8769 = x65 ^ x17 ;
  assign n8770 = n8769 ^ n8766 ;
  assign n8771 = n8373 & ~n8770 ;
  assign n8772 = n8371 & n8723 ;
  assign n8773 = n8771 & ~n8772 ;
  assign n8774 = ~n8768 & n8773 ;
  assign n8755 = x64 ^ x17 ;
  assign n8756 = n8723 & n8755 ;
  assign n8757 = x16 & x65 ;
  assign n8760 = x64 & ~n8757 ;
  assign n8761 = n8760 ^ x65 ;
  assign n8762 = n8373 & n8761 ;
  assign n8763 = n8762 ^ n196 ;
  assign n8764 = n8756 & n8763 ;
  assign n8775 = n8774 ^ n8764 ;
  assign n8776 = n8723 ^ n8373 ;
  assign n8777 = n8770 & ~n8776 ;
  assign n8778 = x64 & n8723 ;
  assign n8779 = ~x17 & ~x66 ;
  assign n8780 = ~n8373 & n8765 ;
  assign n8781 = n8779 & n8780 ;
  assign n8782 = n8781 ^ x66 ;
  assign n8783 = ~n8778 & ~n8782 ;
  assign n8784 = n8777 & n8783 ;
  assign n8785 = n8784 ^ n8782 ;
  assign n8786 = n8373 ^ x65 ;
  assign n8787 = n8786 ^ n8723 ;
  assign n8788 = x17 ^ x16 ;
  assign n8789 = n8788 ^ n8776 ;
  assign n8790 = n8373 ^ x16 ;
  assign n8791 = n8790 ^ n8788 ;
  assign n8792 = ~n8789 & ~n8791 ;
  assign n8793 = n8792 ^ n8788 ;
  assign n8794 = n8787 & n8793 ;
  assign n8795 = x64 & n8794 ;
  assign n8796 = ~n8785 & n8795 ;
  assign n8797 = n8796 ^ n8785 ;
  assign n8800 = n8797 ^ x16 ;
  assign n8801 = n8800 ^ n8797 ;
  assign n8806 = ~x17 & n8796 ;
  assign n8807 = n8801 & n8806 ;
  assign n8808 = n8807 ^ n8801 ;
  assign n8809 = n8808 ^ n8800 ;
  assign n8810 = ~n8775 & n8809 ;
  assign n8813 = n8812 ^ n8810 ;
  assign n8814 = n8812 ^ x67 ;
  assign n8815 = n8813 & ~n8814 ;
  assign n8816 = n8815 ^ x67 ;
  assign n8820 = n8819 ^ n8816 ;
  assign n8821 = n8819 ^ x68 ;
  assign n8822 = n8820 & ~n8821 ;
  assign n8823 = n8822 ^ x68 ;
  assign n8824 = n8823 ^ n8753 ;
  assign n8825 = ~n8754 & n8824 ;
  assign n8826 = n8825 ^ x69 ;
  assign n8827 = n8826 ^ n8749 ;
  assign n8828 = ~n8750 & n8827 ;
  assign n8829 = n8828 ^ x70 ;
  assign n8833 = n8832 ^ n8829 ;
  assign n8834 = n8832 ^ x71 ;
  assign n8835 = n8833 & ~n8834 ;
  assign n8836 = n8835 ^ x71 ;
  assign n8840 = n8839 ^ n8836 ;
  assign n8841 = n8839 ^ x72 ;
  assign n8842 = n8840 & ~n8841 ;
  assign n8843 = n8842 ^ x72 ;
  assign n8847 = n8846 ^ n8843 ;
  assign n8848 = n8846 ^ x73 ;
  assign n8849 = n8847 & ~n8848 ;
  assign n8850 = n8849 ^ x73 ;
  assign n8854 = n8853 ^ n8850 ;
  assign n8855 = n8853 ^ x74 ;
  assign n8856 = n8854 & ~n8855 ;
  assign n8857 = n8856 ^ x74 ;
  assign n8861 = n8860 ^ n8857 ;
  assign n8862 = n8860 ^ x75 ;
  assign n8863 = n8861 & ~n8862 ;
  assign n8864 = n8863 ^ x75 ;
  assign n8868 = n8867 ^ n8864 ;
  assign n8869 = n8867 ^ x76 ;
  assign n8870 = n8868 & ~n8869 ;
  assign n8871 = n8870 ^ x76 ;
  assign n8875 = n8874 ^ n8871 ;
  assign n8876 = n8874 ^ x77 ;
  assign n8877 = n8875 & ~n8876 ;
  assign n8878 = n8877 ^ x77 ;
  assign n8882 = n8881 ^ n8878 ;
  assign n8883 = n8881 ^ x78 ;
  assign n8884 = n8882 & ~n8883 ;
  assign n8885 = n8884 ^ x78 ;
  assign n8889 = n8888 ^ n8885 ;
  assign n8890 = n8888 ^ x79 ;
  assign n8891 = n8889 & ~n8890 ;
  assign n8892 = n8891 ^ x79 ;
  assign n8896 = n8895 ^ n8892 ;
  assign n8897 = n8895 ^ x80 ;
  assign n8898 = n8896 & ~n8897 ;
  assign n8899 = n8898 ^ x80 ;
  assign n8903 = n8902 ^ n8899 ;
  assign n8904 = n8902 ^ x81 ;
  assign n8905 = n8903 & ~n8904 ;
  assign n8906 = n8905 ^ x81 ;
  assign n8910 = n8909 ^ n8906 ;
  assign n8911 = n8909 ^ x82 ;
  assign n8912 = n8910 & ~n8911 ;
  assign n8913 = n8912 ^ x82 ;
  assign n8917 = n8916 ^ n8913 ;
  assign n8918 = n8916 ^ x83 ;
  assign n8919 = n8917 & ~n8918 ;
  assign n8920 = n8919 ^ x83 ;
  assign n8924 = n8923 ^ n8920 ;
  assign n8925 = n8923 ^ x84 ;
  assign n8926 = n8924 & ~n8925 ;
  assign n8927 = n8926 ^ x84 ;
  assign n8931 = n8930 ^ n8927 ;
  assign n8932 = n8930 ^ x85 ;
  assign n8933 = n8931 & ~n8932 ;
  assign n8934 = n8933 ^ x85 ;
  assign n8938 = n8937 ^ n8934 ;
  assign n8939 = n8937 ^ x86 ;
  assign n8940 = n8938 & ~n8939 ;
  assign n8941 = n8940 ^ x86 ;
  assign n8953 = n8952 ^ n8941 ;
  assign n8954 = n8952 ^ x87 ;
  assign n8955 = n8953 & ~n8954 ;
  assign n8956 = n8955 ^ x87 ;
  assign n8960 = n8959 ^ n8956 ;
  assign n8961 = n8959 ^ x88 ;
  assign n8962 = n8960 & ~n8961 ;
  assign n8963 = n8962 ^ x88 ;
  assign n8967 = n8966 ^ n8963 ;
  assign n8968 = n8966 ^ x89 ;
  assign n8969 = n8967 & ~n8968 ;
  assign n8970 = n8969 ^ x89 ;
  assign n8974 = n8973 ^ n8970 ;
  assign n8975 = n8973 ^ x90 ;
  assign n8976 = n8974 & ~n8975 ;
  assign n8977 = n8976 ^ x90 ;
  assign n8981 = n8980 ^ n8977 ;
  assign n8982 = n8980 ^ x91 ;
  assign n8983 = n8981 & ~n8982 ;
  assign n8984 = n8983 ^ x91 ;
  assign n8988 = n8987 ^ n8984 ;
  assign n8989 = n8987 ^ x92 ;
  assign n8990 = n8988 & ~n8989 ;
  assign n8991 = n8990 ^ x92 ;
  assign n8995 = n8994 ^ n8991 ;
  assign n8996 = n8994 ^ x93 ;
  assign n8997 = n8995 & ~n8996 ;
  assign n8998 = n8997 ^ x93 ;
  assign n8999 = n8998 ^ n8745 ;
  assign n9000 = ~n8746 & n8999 ;
  assign n9001 = n9000 ^ x94 ;
  assign n9002 = n9001 ^ n8741 ;
  assign n9003 = ~n8742 & n9002 ;
  assign n9004 = n9003 ^ x95 ;
  assign n9008 = n9007 ^ n9004 ;
  assign n9009 = n9007 ^ x96 ;
  assign n9010 = n9008 & ~n9009 ;
  assign n9011 = n9010 ^ x96 ;
  assign n9015 = n9014 ^ n9011 ;
  assign n9016 = n9014 ^ x97 ;
  assign n9017 = n9015 & ~n9016 ;
  assign n9018 = n9017 ^ x97 ;
  assign n9022 = n9021 ^ n9018 ;
  assign n9023 = n9021 ^ x98 ;
  assign n9024 = n9022 & ~n9023 ;
  assign n9025 = n9024 ^ x98 ;
  assign n9029 = n9028 ^ n9025 ;
  assign n9030 = n9028 ^ x99 ;
  assign n9031 = n9029 & ~n9030 ;
  assign n9032 = n9031 ^ x99 ;
  assign n9033 = n9032 ^ n8737 ;
  assign n9034 = ~n8738 & n9033 ;
  assign n9035 = n9034 ^ x100 ;
  assign n9036 = n9035 ^ n8733 ;
  assign n9037 = ~n8734 & n9036 ;
  assign n9038 = n9037 ^ x101 ;
  assign n9042 = n9041 ^ n9038 ;
  assign n9043 = n9041 ^ x102 ;
  assign n9044 = n9042 & ~n9043 ;
  assign n9045 = n9044 ^ x102 ;
  assign n9049 = n9048 ^ n9045 ;
  assign n9050 = n9048 ^ x103 ;
  assign n9051 = n9049 & ~n9050 ;
  assign n9052 = n9051 ^ x103 ;
  assign n9056 = n9055 ^ n9052 ;
  assign n9057 = n9055 ^ x104 ;
  assign n9058 = n9056 & ~n9057 ;
  assign n9059 = n9058 ^ x104 ;
  assign n9063 = n9062 ^ n9059 ;
  assign n9064 = n9062 ^ x105 ;
  assign n9065 = n9063 & ~n9064 ;
  assign n9066 = n9065 ^ x105 ;
  assign n9067 = n9066 ^ n8729 ;
  assign n9068 = ~n8730 & n9067 ;
  assign n9069 = n9068 ^ x106 ;
  assign n9070 = n9069 ^ n8725 ;
  assign n9071 = ~n8726 & n9070 ;
  assign n9072 = n9071 ^ x107 ;
  assign n9076 = n9075 ^ n9072 ;
  assign n9077 = n9075 ^ x108 ;
  assign n9078 = n9076 & ~n9077 ;
  assign n9079 = n9078 ^ x108 ;
  assign n9083 = n9082 ^ n9079 ;
  assign n9084 = n9082 ^ x109 ;
  assign n9085 = n9083 & ~n9084 ;
  assign n9086 = n9085 ^ x109 ;
  assign n9087 = n9086 ^ x110 ;
  assign n9088 = ~x112 & n8716 ;
  assign n9089 = n8715 ^ x111 ;
  assign n9091 = n8723 & n9090 ;
  assign n9092 = n9091 ^ n8707 ;
  assign n9093 = n9092 ^ x110 ;
  assign n9094 = n9092 ^ n9086 ;
  assign n9095 = ~n9093 & n9094 ;
  assign n9096 = n9095 ^ x110 ;
  assign n9097 = n9096 ^ n8715 ;
  assign n9098 = ~n9089 & ~n9097 ;
  assign n9099 = n9098 ^ n8715 ;
  assign n9100 = n9088 & n9099 ;
  assign n9101 = n9087 & n9100 ;
  assign n9102 = n9101 ^ n9092 ;
  assign n9103 = n9079 ^ x109 ;
  assign n9104 = n9100 & n9103 ;
  assign n9105 = n9104 ^ n9082 ;
  assign n9106 = n9105 ^ x110 ;
  assign n9107 = n9072 ^ x108 ;
  assign n9108 = n9100 & n9107 ;
  assign n9109 = n9108 ^ n9075 ;
  assign n9110 = n9109 ^ x109 ;
  assign n9431 = n9069 ^ x107 ;
  assign n9432 = n9100 & n9431 ;
  assign n9433 = n9432 ^ n8725 ;
  assign n9424 = n9066 ^ x106 ;
  assign n9425 = n9100 & n9424 ;
  assign n9426 = n9425 ^ n8729 ;
  assign n9417 = n9059 ^ x105 ;
  assign n9418 = n9100 & n9417 ;
  assign n9419 = n9418 ^ n9062 ;
  assign n9111 = n9052 ^ x104 ;
  assign n9112 = n9100 & n9111 ;
  assign n9113 = n9112 ^ n9055 ;
  assign n9114 = n9113 ^ x105 ;
  assign n9119 = n9113 ^ x104 ;
  assign n9115 = n9045 ^ x103 ;
  assign n9116 = n9100 & n9115 ;
  assign n9117 = n9116 ^ n9048 ;
  assign n9118 = n9117 ^ n9113 ;
  assign n9120 = n9119 ^ n9118 ;
  assign n9404 = n9038 ^ x102 ;
  assign n9405 = n9100 & n9404 ;
  assign n9406 = n9405 ^ n9041 ;
  assign n9397 = n9035 ^ x101 ;
  assign n9398 = n9100 & n9397 ;
  assign n9399 = n9398 ^ n8733 ;
  assign n9390 = n9032 ^ x100 ;
  assign n9391 = n9100 & n9390 ;
  assign n9392 = n9391 ^ n8737 ;
  assign n9383 = n9025 ^ x99 ;
  assign n9384 = n9100 & n9383 ;
  assign n9385 = n9384 ^ n9028 ;
  assign n9376 = n9018 ^ x98 ;
  assign n9377 = n9100 & n9376 ;
  assign n9378 = n9377 ^ n9021 ;
  assign n9369 = n9011 ^ x97 ;
  assign n9370 = n9100 & n9369 ;
  assign n9371 = n9370 ^ n9014 ;
  assign n9362 = n9004 ^ x96 ;
  assign n9363 = n9100 & n9362 ;
  assign n9364 = n9363 ^ n9007 ;
  assign n9355 = n9001 ^ x95 ;
  assign n9356 = n9100 & n9355 ;
  assign n9357 = n9356 ^ n8741 ;
  assign n9348 = n8998 ^ x94 ;
  assign n9349 = n9100 & n9348 ;
  assign n9350 = n9349 ^ n8745 ;
  assign n9341 = n8991 ^ x93 ;
  assign n9342 = n9100 & n9341 ;
  assign n9343 = n9342 ^ n8994 ;
  assign n9334 = n8984 ^ x92 ;
  assign n9335 = n9100 & n9334 ;
  assign n9336 = n9335 ^ n8987 ;
  assign n9327 = n8977 ^ x91 ;
  assign n9328 = n9100 & n9327 ;
  assign n9329 = n9328 ^ n8980 ;
  assign n9320 = n8970 ^ x90 ;
  assign n9321 = n9100 & n9320 ;
  assign n9322 = n9321 ^ n8973 ;
  assign n9313 = n8963 ^ x89 ;
  assign n9314 = n9100 & n9313 ;
  assign n9315 = n9314 ^ n8966 ;
  assign n9306 = n8956 ^ x88 ;
  assign n9307 = n9100 & n9306 ;
  assign n9308 = n9307 ^ n8959 ;
  assign n9299 = n8941 ^ x87 ;
  assign n9300 = n9100 & n9299 ;
  assign n9301 = n9300 ^ n8952 ;
  assign n9292 = n8934 ^ x86 ;
  assign n9293 = n9100 & n9292 ;
  assign n9294 = n9293 ^ n8937 ;
  assign n9285 = n8927 ^ x85 ;
  assign n9286 = n9100 & n9285 ;
  assign n9287 = n9286 ^ n8930 ;
  assign n9278 = n8920 ^ x84 ;
  assign n9279 = n9100 & n9278 ;
  assign n9280 = n9279 ^ n8923 ;
  assign n9271 = n8913 ^ x83 ;
  assign n9272 = n9100 & n9271 ;
  assign n9273 = n9272 ^ n8916 ;
  assign n9264 = n8906 ^ x82 ;
  assign n9265 = n9100 & n9264 ;
  assign n9266 = n9265 ^ n8909 ;
  assign n9121 = n8899 ^ x81 ;
  assign n9122 = n9100 & n9121 ;
  assign n9123 = n9122 ^ n8902 ;
  assign n9124 = n9123 ^ x82 ;
  assign n9129 = n9123 ^ x81 ;
  assign n9125 = n8892 ^ x80 ;
  assign n9126 = n9100 & n9125 ;
  assign n9127 = n9126 ^ n8895 ;
  assign n9128 = n9127 ^ n9123 ;
  assign n9130 = n9129 ^ n9128 ;
  assign n9251 = n8885 ^ x79 ;
  assign n9252 = n9100 & n9251 ;
  assign n9253 = n9252 ^ n8888 ;
  assign n9244 = n8878 ^ x78 ;
  assign n9245 = n9100 & n9244 ;
  assign n9246 = n9245 ^ n8881 ;
  assign n9237 = n8871 ^ x77 ;
  assign n9238 = n9100 & n9237 ;
  assign n9239 = n9238 ^ n8874 ;
  assign n9230 = n8864 ^ x76 ;
  assign n9231 = n9100 & n9230 ;
  assign n9232 = n9231 ^ n8867 ;
  assign n9223 = n8857 ^ x75 ;
  assign n9224 = n9100 & n9223 ;
  assign n9225 = n9224 ^ n8860 ;
  assign n9216 = n8850 ^ x74 ;
  assign n9217 = n9100 & n9216 ;
  assign n9218 = n9217 ^ n8853 ;
  assign n9209 = n8843 ^ x73 ;
  assign n9210 = n9100 & n9209 ;
  assign n9211 = n9210 ^ n8846 ;
  assign n9202 = n8836 ^ x72 ;
  assign n9203 = n9100 & n9202 ;
  assign n9204 = n9203 ^ n8839 ;
  assign n9195 = n8829 ^ x71 ;
  assign n9196 = n9100 & n9195 ;
  assign n9197 = n9196 ^ n8832 ;
  assign n9188 = n8826 ^ x70 ;
  assign n9189 = n9100 & n9188 ;
  assign n9190 = n9189 ^ n8749 ;
  assign n9181 = n8823 ^ x69 ;
  assign n9182 = n9100 & n9181 ;
  assign n9183 = n9182 ^ n8753 ;
  assign n9174 = n8816 ^ x68 ;
  assign n9175 = n9100 & n9174 ;
  assign n9176 = n9175 ^ n8819 ;
  assign n9167 = n8810 ^ x67 ;
  assign n9168 = n9100 & n9167 ;
  assign n9169 = n9168 ^ n8812 ;
  assign n9161 = n8772 ^ n8373 ;
  assign n9156 = x17 & x65 ;
  assign n9147 = x65 ^ x16 ;
  assign n9148 = n8755 ^ x65 ;
  assign n9149 = n9148 ^ n8723 ;
  assign n9150 = ~n9147 & n9149 ;
  assign n9157 = n9156 ^ n9150 ;
  assign n9158 = ~x64 & n9157 ;
  assign n9153 = n9150 ^ n7358 ;
  assign n9159 = n9158 ^ n9153 ;
  assign n9160 = n9100 & n9159 ;
  assign n9162 = n9161 ^ n9160 ;
  assign n9132 = n8765 ^ x65 ;
  assign n9133 = n9100 & n9132 ;
  assign n9131 = n8778 ^ x17 ;
  assign n9134 = n9133 ^ n9131 ;
  assign n9135 = n9134 ^ x66 ;
  assign n9136 = x65 ^ x15 ;
  assign n9137 = x64 ^ x16 ;
  assign n9138 = n9137 ^ x65 ;
  assign n9139 = n9138 ^ n9100 ;
  assign n9140 = ~n9136 & n9139 ;
  assign n9141 = n9140 ^ n8757 ;
  assign n9142 = x64 & n9141 ;
  assign n8758 = n8757 ^ x65 ;
  assign n9143 = n9142 ^ n8758 ;
  assign n9144 = n9143 ^ n9134 ;
  assign n9145 = ~n9135 & n9144 ;
  assign n9146 = n9145 ^ x66 ;
  assign n9163 = n9162 ^ n9146 ;
  assign n9164 = n9162 ^ x67 ;
  assign n9165 = n9163 & ~n9164 ;
  assign n9166 = n9165 ^ x67 ;
  assign n9170 = n9169 ^ n9166 ;
  assign n9171 = n9169 ^ x68 ;
  assign n9172 = n9170 & ~n9171 ;
  assign n9173 = n9172 ^ x68 ;
  assign n9177 = n9176 ^ n9173 ;
  assign n9178 = n9176 ^ x69 ;
  assign n9179 = n9177 & ~n9178 ;
  assign n9180 = n9179 ^ x69 ;
  assign n9184 = n9183 ^ n9180 ;
  assign n9185 = n9183 ^ x70 ;
  assign n9186 = n9184 & ~n9185 ;
  assign n9187 = n9186 ^ x70 ;
  assign n9191 = n9190 ^ n9187 ;
  assign n9192 = n9190 ^ x71 ;
  assign n9193 = n9191 & ~n9192 ;
  assign n9194 = n9193 ^ x71 ;
  assign n9198 = n9197 ^ n9194 ;
  assign n9199 = n9197 ^ x72 ;
  assign n9200 = n9198 & ~n9199 ;
  assign n9201 = n9200 ^ x72 ;
  assign n9205 = n9204 ^ n9201 ;
  assign n9206 = n9204 ^ x73 ;
  assign n9207 = n9205 & ~n9206 ;
  assign n9208 = n9207 ^ x73 ;
  assign n9212 = n9211 ^ n9208 ;
  assign n9213 = n9211 ^ x74 ;
  assign n9214 = n9212 & ~n9213 ;
  assign n9215 = n9214 ^ x74 ;
  assign n9219 = n9218 ^ n9215 ;
  assign n9220 = n9218 ^ x75 ;
  assign n9221 = n9219 & ~n9220 ;
  assign n9222 = n9221 ^ x75 ;
  assign n9226 = n9225 ^ n9222 ;
  assign n9227 = n9225 ^ x76 ;
  assign n9228 = n9226 & ~n9227 ;
  assign n9229 = n9228 ^ x76 ;
  assign n9233 = n9232 ^ n9229 ;
  assign n9234 = n9232 ^ x77 ;
  assign n9235 = n9233 & ~n9234 ;
  assign n9236 = n9235 ^ x77 ;
  assign n9240 = n9239 ^ n9236 ;
  assign n9241 = n9239 ^ x78 ;
  assign n9242 = n9240 & ~n9241 ;
  assign n9243 = n9242 ^ x78 ;
  assign n9247 = n9246 ^ n9243 ;
  assign n9248 = n9246 ^ x79 ;
  assign n9249 = n9247 & ~n9248 ;
  assign n9250 = n9249 ^ x79 ;
  assign n9254 = n9253 ^ n9250 ;
  assign n9255 = n9253 ^ x80 ;
  assign n9256 = n9254 & ~n9255 ;
  assign n9257 = n9256 ^ x80 ;
  assign n9258 = n9257 ^ n9123 ;
  assign n9259 = n9258 ^ n9129 ;
  assign n9260 = ~n9130 & n9259 ;
  assign n9261 = n9260 ^ n9129 ;
  assign n9262 = ~n9124 & n9261 ;
  assign n9263 = n9262 ^ x82 ;
  assign n9267 = n9266 ^ n9263 ;
  assign n9268 = n9266 ^ x83 ;
  assign n9269 = n9267 & ~n9268 ;
  assign n9270 = n9269 ^ x83 ;
  assign n9274 = n9273 ^ n9270 ;
  assign n9275 = n9273 ^ x84 ;
  assign n9276 = n9274 & ~n9275 ;
  assign n9277 = n9276 ^ x84 ;
  assign n9281 = n9280 ^ n9277 ;
  assign n9282 = n9280 ^ x85 ;
  assign n9283 = n9281 & ~n9282 ;
  assign n9284 = n9283 ^ x85 ;
  assign n9288 = n9287 ^ n9284 ;
  assign n9289 = n9287 ^ x86 ;
  assign n9290 = n9288 & ~n9289 ;
  assign n9291 = n9290 ^ x86 ;
  assign n9295 = n9294 ^ n9291 ;
  assign n9296 = n9294 ^ x87 ;
  assign n9297 = n9295 & ~n9296 ;
  assign n9298 = n9297 ^ x87 ;
  assign n9302 = n9301 ^ n9298 ;
  assign n9303 = n9301 ^ x88 ;
  assign n9304 = n9302 & ~n9303 ;
  assign n9305 = n9304 ^ x88 ;
  assign n9309 = n9308 ^ n9305 ;
  assign n9310 = n9308 ^ x89 ;
  assign n9311 = n9309 & ~n9310 ;
  assign n9312 = n9311 ^ x89 ;
  assign n9316 = n9315 ^ n9312 ;
  assign n9317 = n9315 ^ x90 ;
  assign n9318 = n9316 & ~n9317 ;
  assign n9319 = n9318 ^ x90 ;
  assign n9323 = n9322 ^ n9319 ;
  assign n9324 = n9322 ^ x91 ;
  assign n9325 = n9323 & ~n9324 ;
  assign n9326 = n9325 ^ x91 ;
  assign n9330 = n9329 ^ n9326 ;
  assign n9331 = n9329 ^ x92 ;
  assign n9332 = n9330 & ~n9331 ;
  assign n9333 = n9332 ^ x92 ;
  assign n9337 = n9336 ^ n9333 ;
  assign n9338 = n9336 ^ x93 ;
  assign n9339 = n9337 & ~n9338 ;
  assign n9340 = n9339 ^ x93 ;
  assign n9344 = n9343 ^ n9340 ;
  assign n9345 = n9343 ^ x94 ;
  assign n9346 = n9344 & ~n9345 ;
  assign n9347 = n9346 ^ x94 ;
  assign n9351 = n9350 ^ n9347 ;
  assign n9352 = n9350 ^ x95 ;
  assign n9353 = n9351 & ~n9352 ;
  assign n9354 = n9353 ^ x95 ;
  assign n9358 = n9357 ^ n9354 ;
  assign n9359 = n9357 ^ x96 ;
  assign n9360 = n9358 & ~n9359 ;
  assign n9361 = n9360 ^ x96 ;
  assign n9365 = n9364 ^ n9361 ;
  assign n9366 = n9364 ^ x97 ;
  assign n9367 = n9365 & ~n9366 ;
  assign n9368 = n9367 ^ x97 ;
  assign n9372 = n9371 ^ n9368 ;
  assign n9373 = n9371 ^ x98 ;
  assign n9374 = n9372 & ~n9373 ;
  assign n9375 = n9374 ^ x98 ;
  assign n9379 = n9378 ^ n9375 ;
  assign n9380 = n9378 ^ x99 ;
  assign n9381 = n9379 & ~n9380 ;
  assign n9382 = n9381 ^ x99 ;
  assign n9386 = n9385 ^ n9382 ;
  assign n9387 = n9385 ^ x100 ;
  assign n9388 = n9386 & ~n9387 ;
  assign n9389 = n9388 ^ x100 ;
  assign n9393 = n9392 ^ n9389 ;
  assign n9394 = n9392 ^ x101 ;
  assign n9395 = n9393 & ~n9394 ;
  assign n9396 = n9395 ^ x101 ;
  assign n9400 = n9399 ^ n9396 ;
  assign n9401 = n9399 ^ x102 ;
  assign n9402 = n9400 & ~n9401 ;
  assign n9403 = n9402 ^ x102 ;
  assign n9407 = n9406 ^ n9403 ;
  assign n9408 = n9406 ^ x103 ;
  assign n9409 = n9407 & ~n9408 ;
  assign n9410 = n9409 ^ x103 ;
  assign n9411 = n9410 ^ n9113 ;
  assign n9412 = n9411 ^ n9119 ;
  assign n9413 = ~n9120 & n9412 ;
  assign n9414 = n9413 ^ n9119 ;
  assign n9415 = ~n9114 & n9414 ;
  assign n9416 = n9415 ^ x105 ;
  assign n9420 = n9419 ^ n9416 ;
  assign n9421 = n9419 ^ x106 ;
  assign n9422 = n9420 & ~n9421 ;
  assign n9423 = n9422 ^ x106 ;
  assign n9427 = n9426 ^ n9423 ;
  assign n9428 = n9426 ^ x107 ;
  assign n9429 = n9427 & ~n9428 ;
  assign n9430 = n9429 ^ x107 ;
  assign n9434 = n9433 ^ n9430 ;
  assign n9435 = n9433 ^ x108 ;
  assign n9436 = n9434 & ~n9435 ;
  assign n9437 = n9436 ^ x108 ;
  assign n9438 = n9437 ^ n9109 ;
  assign n9439 = ~n9110 & n9438 ;
  assign n9440 = n9439 ^ x109 ;
  assign n9441 = n9440 ^ n9105 ;
  assign n9442 = ~n9106 & n9441 ;
  assign n9443 = n9442 ^ x110 ;
  assign n9445 = n9102 & ~n9443 ;
  assign n9444 = n9443 ^ n9102 ;
  assign n9446 = n9445 ^ n9444 ;
  assign n9447 = ~x111 & ~n9446 ;
  assign n9448 = n9447 ^ x112 ;
  assign n9449 = n8716 & n9448 ;
  assign n9450 = n9445 ^ n9096 ;
  assign n9453 = ~n9447 & n9450 ;
  assign n9454 = n9453 ^ n9096 ;
  assign n9455 = n9449 & ~n9454 ;
  assign n9456 = n9455 ^ n8716 ;
  assign n9457 = n8715 & ~n9456 ;
  assign n9458 = n142 & n9457 ;
  assign n9469 = n9447 ^ x111 ;
  assign n9460 = ~n9445 & ~n9447 ;
  assign n9470 = n9469 ^ n9460 ;
  assign n9471 = n9470 ^ n9469 ;
  assign n9472 = n9469 ^ n9096 ;
  assign n9473 = n9472 ^ n9469 ;
  assign n9474 = n9471 & ~n9473 ;
  assign n9475 = n9474 ^ n9469 ;
  assign n9476 = n9100 & ~n9475 ;
  assign n9477 = n9476 ^ n9088 ;
  assign n9468 = ~n8715 & n9460 ;
  assign n9478 = n9477 ^ n9468 ;
  assign n9461 = n9460 ^ n7998 ;
  assign n9462 = n7998 ^ x112 ;
  assign n9465 = ~n8716 & ~n9462 ;
  assign n9466 = n9465 ^ x112 ;
  assign n9467 = n9461 & n9466 ;
  assign n9479 = n9478 ^ n9467 ;
  assign n9834 = n9443 ^ x111 ;
  assign n9835 = n9479 & n9834 ;
  assign n9836 = n9835 ^ n9102 ;
  assign n9827 = n9440 ^ x110 ;
  assign n9828 = n9479 & n9827 ;
  assign n9829 = n9828 ^ n9105 ;
  assign n9820 = n9437 ^ x109 ;
  assign n9821 = n9479 & n9820 ;
  assign n9822 = n9821 ^ n9109 ;
  assign n9813 = n9430 ^ x108 ;
  assign n9814 = n9479 & n9813 ;
  assign n9815 = n9814 ^ n9433 ;
  assign n9806 = n9423 ^ x107 ;
  assign n9807 = n9479 & n9806 ;
  assign n9808 = n9807 ^ n9426 ;
  assign n9799 = n9416 ^ x106 ;
  assign n9800 = n9479 & n9799 ;
  assign n9801 = n9800 ^ n9419 ;
  assign n9784 = n9117 ^ x105 ;
  assign n9785 = n9784 ^ x104 ;
  assign n9786 = n9785 ^ n9410 ;
  assign n9787 = n9786 ^ n9784 ;
  assign n9790 = n9784 ^ n6926 ;
  assign n9791 = ~n9787 & ~n9790 ;
  assign n9792 = n9791 ^ n9784 ;
  assign n9793 = n9479 & ~n9792 ;
  assign n9794 = n9793 ^ n9113 ;
  assign n9777 = n9410 ^ x104 ;
  assign n9778 = n9479 & n9777 ;
  assign n9779 = n9778 ^ n9117 ;
  assign n9770 = n9403 ^ x103 ;
  assign n9771 = n9479 & n9770 ;
  assign n9772 = n9771 ^ n9406 ;
  assign n9763 = n9396 ^ x102 ;
  assign n9764 = n9479 & n9763 ;
  assign n9765 = n9764 ^ n9399 ;
  assign n9756 = n9389 ^ x101 ;
  assign n9757 = n9479 & n9756 ;
  assign n9758 = n9757 ^ n9392 ;
  assign n9749 = n9382 ^ x100 ;
  assign n9750 = n9479 & n9749 ;
  assign n9751 = n9750 ^ n9385 ;
  assign n9742 = n9375 ^ x99 ;
  assign n9743 = n9479 & n9742 ;
  assign n9744 = n9743 ^ n9378 ;
  assign n9735 = n9368 ^ x98 ;
  assign n9736 = n9479 & n9735 ;
  assign n9737 = n9736 ^ n9371 ;
  assign n9728 = n9361 ^ x97 ;
  assign n9729 = n9479 & n9728 ;
  assign n9730 = n9729 ^ n9364 ;
  assign n9721 = n9354 ^ x96 ;
  assign n9722 = n9479 & n9721 ;
  assign n9723 = n9722 ^ n9357 ;
  assign n9714 = n9347 ^ x95 ;
  assign n9715 = n9479 & n9714 ;
  assign n9716 = n9715 ^ n9350 ;
  assign n9707 = n9340 ^ x94 ;
  assign n9708 = n9479 & n9707 ;
  assign n9709 = n9708 ^ n9343 ;
  assign n9700 = n9333 ^ x93 ;
  assign n9701 = n9479 & n9700 ;
  assign n9702 = n9701 ^ n9336 ;
  assign n9693 = n9326 ^ x92 ;
  assign n9694 = n9479 & n9693 ;
  assign n9695 = n9694 ^ n9329 ;
  assign n9686 = n9319 ^ x91 ;
  assign n9687 = n9479 & n9686 ;
  assign n9688 = n9687 ^ n9322 ;
  assign n9459 = n9312 ^ x90 ;
  assign n9480 = n9459 & n9479 ;
  assign n9481 = n9480 ^ n9315 ;
  assign n9482 = n9481 ^ x91 ;
  assign n9487 = n9481 ^ x90 ;
  assign n9483 = n9305 ^ x89 ;
  assign n9484 = n9479 & n9483 ;
  assign n9485 = n9484 ^ n9308 ;
  assign n9486 = n9485 ^ n9481 ;
  assign n9488 = n9487 ^ n9486 ;
  assign n9489 = n9298 ^ x88 ;
  assign n9490 = n9479 & n9489 ;
  assign n9491 = n9490 ^ n9301 ;
  assign n9492 = n9491 ^ x89 ;
  assign n9497 = n9491 ^ x88 ;
  assign n9493 = n9291 ^ x87 ;
  assign n9494 = n9479 & n9493 ;
  assign n9495 = n9494 ^ n9294 ;
  assign n9496 = n9495 ^ n9491 ;
  assign n9498 = n9497 ^ n9496 ;
  assign n9667 = n9284 ^ x86 ;
  assign n9668 = n9479 & n9667 ;
  assign n9669 = n9668 ^ n9287 ;
  assign n9499 = n9277 ^ x85 ;
  assign n9500 = n9479 & n9499 ;
  assign n9501 = n9500 ^ n9280 ;
  assign n9502 = n9501 ^ x86 ;
  assign n9503 = n9270 ^ x84 ;
  assign n9504 = n9479 & n9503 ;
  assign n9505 = n9504 ^ n9273 ;
  assign n9506 = n9505 ^ x85 ;
  assign n9654 = n9263 ^ x83 ;
  assign n9655 = n9479 & n9654 ;
  assign n9656 = n9655 ^ n9266 ;
  assign n9639 = n9127 ^ x82 ;
  assign n9640 = n9639 ^ x81 ;
  assign n9641 = n9640 ^ n9257 ;
  assign n9642 = n9641 ^ n9639 ;
  assign n9645 = n9639 ^ n5543 ;
  assign n9646 = ~n9642 & ~n9645 ;
  assign n9647 = n9646 ^ n9639 ;
  assign n9648 = n9479 & ~n9647 ;
  assign n9649 = n9648 ^ n9123 ;
  assign n9632 = n9257 ^ x81 ;
  assign n9633 = n9479 & n9632 ;
  assign n9634 = n9633 ^ n9127 ;
  assign n9625 = n9250 ^ x80 ;
  assign n9626 = n9479 & n9625 ;
  assign n9627 = n9626 ^ n9253 ;
  assign n9618 = n9243 ^ x79 ;
  assign n9619 = n9479 & n9618 ;
  assign n9620 = n9619 ^ n9246 ;
  assign n9611 = n9236 ^ x78 ;
  assign n9612 = n9479 & n9611 ;
  assign n9613 = n9612 ^ n9239 ;
  assign n9604 = n9229 ^ x77 ;
  assign n9605 = n9479 & n9604 ;
  assign n9606 = n9605 ^ n9232 ;
  assign n9507 = n9222 ^ x76 ;
  assign n9508 = n9479 & n9507 ;
  assign n9509 = n9508 ^ n9225 ;
  assign n9510 = n9509 ^ x77 ;
  assign n9515 = n9509 ^ x76 ;
  assign n9511 = n9215 ^ x75 ;
  assign n9512 = n9479 & n9511 ;
  assign n9513 = n9512 ^ n9218 ;
  assign n9514 = n9513 ^ n9509 ;
  assign n9516 = n9515 ^ n9514 ;
  assign n9591 = n9208 ^ x74 ;
  assign n9592 = n9479 & n9591 ;
  assign n9593 = n9592 ^ n9211 ;
  assign n9584 = n9201 ^ x73 ;
  assign n9585 = n9479 & n9584 ;
  assign n9586 = n9585 ^ n9204 ;
  assign n9577 = n9194 ^ x72 ;
  assign n9578 = n9479 & n9577 ;
  assign n9579 = n9578 ^ n9197 ;
  assign n9570 = n9187 ^ x71 ;
  assign n9571 = n9479 & n9570 ;
  assign n9572 = n9571 ^ n9190 ;
  assign n9563 = n9180 ^ x70 ;
  assign n9564 = n9479 & n9563 ;
  assign n9565 = n9564 ^ n9183 ;
  assign n9556 = n9173 ^ x69 ;
  assign n9557 = n9479 & n9556 ;
  assign n9558 = n9557 ^ n9176 ;
  assign n9549 = n9166 ^ x68 ;
  assign n9550 = n9479 & n9549 ;
  assign n9551 = n9550 ^ n9169 ;
  assign n9542 = n9146 ^ x67 ;
  assign n9543 = n9479 & n9542 ;
  assign n9544 = n9543 ^ n9162 ;
  assign n9535 = n9143 ^ x66 ;
  assign n9536 = n9479 & n9535 ;
  assign n9537 = n9536 ^ n9134 ;
  assign n9517 = ~x14 & x64 ;
  assign n9518 = n9517 ^ x65 ;
  assign n9519 = x64 & n9479 ;
  assign n9520 = n9519 ^ x15 ;
  assign n9521 = n9520 ^ n9517 ;
  assign n9522 = n9518 & n9521 ;
  assign n9523 = n9522 ^ x65 ;
  assign n9524 = n9523 ^ x66 ;
  assign n9530 = x64 & n9100 ;
  assign n9526 = ~x15 & x64 ;
  assign n9527 = n9526 ^ x65 ;
  assign n9528 = n9479 & n9527 ;
  assign n9529 = n9528 ^ x16 ;
  assign n9531 = n9530 ^ n9529 ;
  assign n9532 = n9531 ^ n9523 ;
  assign n9533 = n9524 & n9532 ;
  assign n9534 = n9533 ^ x66 ;
  assign n9538 = n9537 ^ n9534 ;
  assign n9539 = n9537 ^ x67 ;
  assign n9540 = n9538 & ~n9539 ;
  assign n9541 = n9540 ^ x67 ;
  assign n9545 = n9544 ^ n9541 ;
  assign n9546 = n9544 ^ x68 ;
  assign n9547 = n9545 & ~n9546 ;
  assign n9548 = n9547 ^ x68 ;
  assign n9552 = n9551 ^ n9548 ;
  assign n9553 = n9551 ^ x69 ;
  assign n9554 = n9552 & ~n9553 ;
  assign n9555 = n9554 ^ x69 ;
  assign n9559 = n9558 ^ n9555 ;
  assign n9560 = n9558 ^ x70 ;
  assign n9561 = n9559 & ~n9560 ;
  assign n9562 = n9561 ^ x70 ;
  assign n9566 = n9565 ^ n9562 ;
  assign n9567 = n9565 ^ x71 ;
  assign n9568 = n9566 & ~n9567 ;
  assign n9569 = n9568 ^ x71 ;
  assign n9573 = n9572 ^ n9569 ;
  assign n9574 = n9572 ^ x72 ;
  assign n9575 = n9573 & ~n9574 ;
  assign n9576 = n9575 ^ x72 ;
  assign n9580 = n9579 ^ n9576 ;
  assign n9581 = n9579 ^ x73 ;
  assign n9582 = n9580 & ~n9581 ;
  assign n9583 = n9582 ^ x73 ;
  assign n9587 = n9586 ^ n9583 ;
  assign n9588 = n9586 ^ x74 ;
  assign n9589 = n9587 & ~n9588 ;
  assign n9590 = n9589 ^ x74 ;
  assign n9594 = n9593 ^ n9590 ;
  assign n9595 = n9593 ^ x75 ;
  assign n9596 = n9594 & ~n9595 ;
  assign n9597 = n9596 ^ x75 ;
  assign n9598 = n9597 ^ n9509 ;
  assign n9599 = n9598 ^ n9515 ;
  assign n9600 = ~n9516 & n9599 ;
  assign n9601 = n9600 ^ n9515 ;
  assign n9602 = ~n9510 & n9601 ;
  assign n9603 = n9602 ^ x77 ;
  assign n9607 = n9606 ^ n9603 ;
  assign n9608 = n9606 ^ x78 ;
  assign n9609 = n9607 & ~n9608 ;
  assign n9610 = n9609 ^ x78 ;
  assign n9614 = n9613 ^ n9610 ;
  assign n9615 = n9613 ^ x79 ;
  assign n9616 = n9614 & ~n9615 ;
  assign n9617 = n9616 ^ x79 ;
  assign n9621 = n9620 ^ n9617 ;
  assign n9622 = n9620 ^ x80 ;
  assign n9623 = n9621 & ~n9622 ;
  assign n9624 = n9623 ^ x80 ;
  assign n9628 = n9627 ^ n9624 ;
  assign n9629 = n9627 ^ x81 ;
  assign n9630 = n9628 & ~n9629 ;
  assign n9631 = n9630 ^ x81 ;
  assign n9635 = n9634 ^ n9631 ;
  assign n9636 = n9634 ^ x82 ;
  assign n9637 = n9635 & ~n9636 ;
  assign n9638 = n9637 ^ x82 ;
  assign n9650 = n9649 ^ n9638 ;
  assign n9651 = n9649 ^ x83 ;
  assign n9652 = n9650 & ~n9651 ;
  assign n9653 = n9652 ^ x83 ;
  assign n9657 = n9656 ^ n9653 ;
  assign n9658 = n9656 ^ x84 ;
  assign n9659 = n9657 & ~n9658 ;
  assign n9660 = n9659 ^ x84 ;
  assign n9661 = n9660 ^ n9505 ;
  assign n9662 = ~n9506 & n9661 ;
  assign n9663 = n9662 ^ x85 ;
  assign n9664 = n9663 ^ n9501 ;
  assign n9665 = ~n9502 & n9664 ;
  assign n9666 = n9665 ^ x86 ;
  assign n9670 = n9669 ^ n9666 ;
  assign n9671 = n9669 ^ x87 ;
  assign n9672 = n9670 & ~n9671 ;
  assign n9673 = n9672 ^ x87 ;
  assign n9674 = n9673 ^ n9491 ;
  assign n9675 = n9674 ^ n9497 ;
  assign n9676 = ~n9498 & n9675 ;
  assign n9677 = n9676 ^ n9497 ;
  assign n9678 = ~n9492 & n9677 ;
  assign n9679 = n9678 ^ x89 ;
  assign n9680 = n9679 ^ n9481 ;
  assign n9681 = n9680 ^ n9487 ;
  assign n9682 = ~n9488 & n9681 ;
  assign n9683 = n9682 ^ n9487 ;
  assign n9684 = ~n9482 & n9683 ;
  assign n9685 = n9684 ^ x91 ;
  assign n9689 = n9688 ^ n9685 ;
  assign n9690 = n9688 ^ x92 ;
  assign n9691 = n9689 & ~n9690 ;
  assign n9692 = n9691 ^ x92 ;
  assign n9696 = n9695 ^ n9692 ;
  assign n9697 = n9695 ^ x93 ;
  assign n9698 = n9696 & ~n9697 ;
  assign n9699 = n9698 ^ x93 ;
  assign n9703 = n9702 ^ n9699 ;
  assign n9704 = n9702 ^ x94 ;
  assign n9705 = n9703 & ~n9704 ;
  assign n9706 = n9705 ^ x94 ;
  assign n9710 = n9709 ^ n9706 ;
  assign n9711 = n9709 ^ x95 ;
  assign n9712 = n9710 & ~n9711 ;
  assign n9713 = n9712 ^ x95 ;
  assign n9717 = n9716 ^ n9713 ;
  assign n9718 = n9716 ^ x96 ;
  assign n9719 = n9717 & ~n9718 ;
  assign n9720 = n9719 ^ x96 ;
  assign n9724 = n9723 ^ n9720 ;
  assign n9725 = n9723 ^ x97 ;
  assign n9726 = n9724 & ~n9725 ;
  assign n9727 = n9726 ^ x97 ;
  assign n9731 = n9730 ^ n9727 ;
  assign n9732 = n9730 ^ x98 ;
  assign n9733 = n9731 & ~n9732 ;
  assign n9734 = n9733 ^ x98 ;
  assign n9738 = n9737 ^ n9734 ;
  assign n9739 = n9737 ^ x99 ;
  assign n9740 = n9738 & ~n9739 ;
  assign n9741 = n9740 ^ x99 ;
  assign n9745 = n9744 ^ n9741 ;
  assign n9746 = n9744 ^ x100 ;
  assign n9747 = n9745 & ~n9746 ;
  assign n9748 = n9747 ^ x100 ;
  assign n9752 = n9751 ^ n9748 ;
  assign n9753 = n9751 ^ x101 ;
  assign n9754 = n9752 & ~n9753 ;
  assign n9755 = n9754 ^ x101 ;
  assign n9759 = n9758 ^ n9755 ;
  assign n9760 = n9758 ^ x102 ;
  assign n9761 = n9759 & ~n9760 ;
  assign n9762 = n9761 ^ x102 ;
  assign n9766 = n9765 ^ n9762 ;
  assign n9767 = n9765 ^ x103 ;
  assign n9768 = n9766 & ~n9767 ;
  assign n9769 = n9768 ^ x103 ;
  assign n9773 = n9772 ^ n9769 ;
  assign n9774 = n9772 ^ x104 ;
  assign n9775 = n9773 & ~n9774 ;
  assign n9776 = n9775 ^ x104 ;
  assign n9780 = n9779 ^ n9776 ;
  assign n9781 = n9779 ^ x105 ;
  assign n9782 = n9780 & ~n9781 ;
  assign n9783 = n9782 ^ x105 ;
  assign n9795 = n9794 ^ n9783 ;
  assign n9796 = n9794 ^ x106 ;
  assign n9797 = n9795 & ~n9796 ;
  assign n9798 = n9797 ^ x106 ;
  assign n9802 = n9801 ^ n9798 ;
  assign n9803 = n9801 ^ x107 ;
  assign n9804 = n9802 & ~n9803 ;
  assign n9805 = n9804 ^ x107 ;
  assign n9809 = n9808 ^ n9805 ;
  assign n9810 = n9808 ^ x108 ;
  assign n9811 = n9809 & ~n9810 ;
  assign n9812 = n9811 ^ x108 ;
  assign n9816 = n9815 ^ n9812 ;
  assign n9817 = n9815 ^ x109 ;
  assign n9818 = n9816 & ~n9817 ;
  assign n9819 = n9818 ^ x109 ;
  assign n9823 = n9822 ^ n9819 ;
  assign n9824 = n9822 ^ x110 ;
  assign n9825 = n9823 & ~n9824 ;
  assign n9826 = n9825 ^ x110 ;
  assign n9830 = n9829 ^ n9826 ;
  assign n9831 = n9829 ^ x111 ;
  assign n9832 = n9830 & ~n9831 ;
  assign n9833 = n9832 ^ x111 ;
  assign n9837 = n9836 ^ n9833 ;
  assign n10255 = n9833 ^ x112 ;
  assign n9841 = n9837 & n10255 ;
  assign n9838 = x113 ^ x112 ;
  assign n9842 = n9841 ^ n9838 ;
  assign n9843 = n9458 & n9842 ;
  assign n9844 = n9843 ^ n9457 ;
  assign n9845 = n141 & n9844 ;
  assign n9847 = n9457 ^ x113 ;
  assign n9850 = n9842 & ~n9847 ;
  assign n9851 = n9850 ^ x113 ;
  assign n9852 = n142 & ~n9851 ;
  assign n10256 = n9852 & n10255 ;
  assign n10257 = n10256 ^ n9836 ;
  assign n10248 = n9826 ^ x111 ;
  assign n10249 = n9852 & n10248 ;
  assign n10250 = n10249 ^ n9829 ;
  assign n10241 = n9819 ^ x110 ;
  assign n10242 = n9852 & n10241 ;
  assign n10243 = n10242 ^ n9822 ;
  assign n10234 = n9812 ^ x109 ;
  assign n10235 = n9852 & n10234 ;
  assign n10236 = n10235 ^ n9815 ;
  assign n10227 = n9805 ^ x108 ;
  assign n10228 = n9852 & n10227 ;
  assign n10229 = n10228 ^ n9808 ;
  assign n10220 = n9798 ^ x107 ;
  assign n10221 = n9852 & n10220 ;
  assign n10222 = n10221 ^ n9801 ;
  assign n9846 = n9783 ^ x106 ;
  assign n9853 = n9846 & n9852 ;
  assign n9854 = n9853 ^ n9794 ;
  assign n9855 = n9854 ^ x107 ;
  assign n9860 = n9854 ^ x106 ;
  assign n9856 = n9776 ^ x105 ;
  assign n9857 = n9852 & n9856 ;
  assign n9858 = n9857 ^ n9779 ;
  assign n9859 = n9858 ^ n9854 ;
  assign n9861 = n9860 ^ n9859 ;
  assign n10207 = n9769 ^ x104 ;
  assign n10208 = n9852 & n10207 ;
  assign n10209 = n10208 ^ n9772 ;
  assign n10200 = n9762 ^ x103 ;
  assign n10201 = n9852 & n10200 ;
  assign n10202 = n10201 ^ n9765 ;
  assign n10193 = n9755 ^ x102 ;
  assign n10194 = n9852 & n10193 ;
  assign n10195 = n10194 ^ n9758 ;
  assign n10186 = n9748 ^ x101 ;
  assign n10187 = n9852 & n10186 ;
  assign n10188 = n10187 ^ n9751 ;
  assign n10179 = n9741 ^ x100 ;
  assign n10180 = n9852 & n10179 ;
  assign n10181 = n10180 ^ n9744 ;
  assign n10172 = n9734 ^ x99 ;
  assign n10173 = n9852 & n10172 ;
  assign n10174 = n10173 ^ n9737 ;
  assign n10165 = n9727 ^ x98 ;
  assign n10166 = n9852 & n10165 ;
  assign n10167 = n10166 ^ n9730 ;
  assign n10158 = n9720 ^ x97 ;
  assign n10159 = n9852 & n10158 ;
  assign n10160 = n10159 ^ n9723 ;
  assign n9862 = n9713 ^ x96 ;
  assign n9863 = n9852 & n9862 ;
  assign n9864 = n9863 ^ n9716 ;
  assign n9865 = n9864 ^ x97 ;
  assign n9866 = n9706 ^ x95 ;
  assign n9867 = n9852 & n9866 ;
  assign n9868 = n9867 ^ n9709 ;
  assign n9869 = n9868 ^ x96 ;
  assign n10145 = n9699 ^ x94 ;
  assign n10146 = n9852 & n10145 ;
  assign n10147 = n10146 ^ n9702 ;
  assign n10138 = n9692 ^ x93 ;
  assign n10139 = n9852 & n10138 ;
  assign n10140 = n10139 ^ n9695 ;
  assign n10131 = n9685 ^ x92 ;
  assign n10132 = n9852 & n10131 ;
  assign n10133 = n10132 ^ n9688 ;
  assign n10116 = n9485 ^ x91 ;
  assign n10117 = n10116 ^ n9679 ;
  assign n10118 = n10117 ^ x90 ;
  assign n10119 = n10118 ^ n10116 ;
  assign n10121 = n9679 ^ x91 ;
  assign n10122 = n10121 ^ n10116 ;
  assign n10123 = ~n10119 & ~n10122 ;
  assign n10124 = n10123 ^ n10116 ;
  assign n10125 = n9852 & ~n10124 ;
  assign n10126 = n10125 ^ n9481 ;
  assign n10109 = n9679 ^ x90 ;
  assign n10110 = n9852 & n10109 ;
  assign n10111 = n10110 ^ n9485 ;
  assign n10094 = n9495 ^ x89 ;
  assign n10095 = n10094 ^ n9673 ;
  assign n10096 = n10095 ^ x88 ;
  assign n10097 = n10096 ^ n10094 ;
  assign n10099 = n9673 ^ x89 ;
  assign n10100 = n10099 ^ n10094 ;
  assign n10101 = ~n10097 & ~n10100 ;
  assign n10102 = n10101 ^ n10094 ;
  assign n10103 = n9852 & ~n10102 ;
  assign n10104 = n10103 ^ n9491 ;
  assign n10087 = n9673 ^ x88 ;
  assign n10088 = n9852 & n10087 ;
  assign n10089 = n10088 ^ n9495 ;
  assign n10080 = n9666 ^ x87 ;
  assign n10081 = n9852 & n10080 ;
  assign n10082 = n10081 ^ n9669 ;
  assign n10073 = n9663 ^ x86 ;
  assign n10074 = n9852 & n10073 ;
  assign n10075 = n10074 ^ n9501 ;
  assign n10066 = n9660 ^ x85 ;
  assign n10067 = n9852 & n10066 ;
  assign n10068 = n10067 ^ n9505 ;
  assign n9870 = n9653 ^ x84 ;
  assign n9871 = n9852 & n9870 ;
  assign n9872 = n9871 ^ n9656 ;
  assign n9873 = n9872 ^ x85 ;
  assign n9878 = n9872 ^ x84 ;
  assign n9874 = n9638 ^ x83 ;
  assign n9875 = n9852 & n9874 ;
  assign n9876 = n9875 ^ n9649 ;
  assign n9877 = n9876 ^ n9872 ;
  assign n9879 = n9878 ^ n9877 ;
  assign n10053 = n9631 ^ x82 ;
  assign n10054 = n9852 & n10053 ;
  assign n10055 = n10054 ^ n9634 ;
  assign n10046 = n9624 ^ x81 ;
  assign n10047 = n9852 & n10046 ;
  assign n10048 = n10047 ^ n9627 ;
  assign n10039 = n9617 ^ x80 ;
  assign n10040 = n9852 & n10039 ;
  assign n10041 = n10040 ^ n9620 ;
  assign n10032 = n9610 ^ x79 ;
  assign n10033 = n9852 & n10032 ;
  assign n10034 = n10033 ^ n9613 ;
  assign n10025 = n9603 ^ x78 ;
  assign n10026 = n9852 & n10025 ;
  assign n10027 = n10026 ^ n9606 ;
  assign n10010 = n9513 ^ x77 ;
  assign n10011 = n10010 ^ n9597 ;
  assign n10012 = n10011 ^ x76 ;
  assign n10013 = n10012 ^ n10010 ;
  assign n10015 = n9597 ^ x77 ;
  assign n10016 = n10015 ^ n10010 ;
  assign n10017 = ~n10013 & ~n10016 ;
  assign n10018 = n10017 ^ n10010 ;
  assign n10019 = n9852 & ~n10018 ;
  assign n10020 = n10019 ^ n9509 ;
  assign n10003 = n9597 ^ x76 ;
  assign n10004 = n9852 & n10003 ;
  assign n10005 = n10004 ^ n9513 ;
  assign n9996 = n9590 ^ x75 ;
  assign n9997 = n9852 & n9996 ;
  assign n9998 = n9997 ^ n9593 ;
  assign n9989 = n9583 ^ x74 ;
  assign n9990 = n9852 & n9989 ;
  assign n9991 = n9990 ^ n9586 ;
  assign n9982 = n9576 ^ x73 ;
  assign n9983 = n9852 & n9982 ;
  assign n9984 = n9983 ^ n9579 ;
  assign n9975 = n9569 ^ x72 ;
  assign n9976 = n9852 & n9975 ;
  assign n9977 = n9976 ^ n9572 ;
  assign n9968 = n9562 ^ x71 ;
  assign n9969 = n9852 & n9968 ;
  assign n9970 = n9969 ^ n9565 ;
  assign n9961 = n9555 ^ x70 ;
  assign n9962 = n9852 & n9961 ;
  assign n9963 = n9962 ^ n9558 ;
  assign n9954 = n9548 ^ x69 ;
  assign n9955 = n9852 & n9954 ;
  assign n9956 = n9955 ^ n9551 ;
  assign n9947 = n9541 ^ x68 ;
  assign n9948 = n9852 & n9947 ;
  assign n9949 = n9948 ^ n9544 ;
  assign n9940 = n9534 ^ x67 ;
  assign n9941 = n9852 & n9940 ;
  assign n9942 = n9941 ^ n9537 ;
  assign n9934 = n9524 & n9852 ;
  assign n9935 = n9934 ^ n9531 ;
  assign n9887 = n9520 ^ n196 ;
  assign n9888 = x64 ^ x14 ;
  assign n9889 = n9520 ^ x65 ;
  assign n9890 = ~x13 & x65 ;
  assign n9891 = n9890 ^ n9520 ;
  assign n9892 = ~n9889 & n9891 ;
  assign n9893 = n9892 ^ n9520 ;
  assign n9894 = n9888 & ~n9893 ;
  assign n9895 = n9887 & n9894 ;
  assign n9881 = x65 ^ x14 ;
  assign n9880 = x14 & ~x65 ;
  assign n9882 = n9881 ^ n9880 ;
  assign n9883 = ~x13 & x64 ;
  assign n9884 = ~n9880 & n9883 ;
  assign n9885 = ~n9882 & ~n9884 ;
  assign n9886 = n9520 & n9885 ;
  assign n9896 = n9895 ^ n9886 ;
  assign n9897 = n9852 & n9896 ;
  assign n9898 = ~x65 & ~n9517 ;
  assign n9899 = ~n9883 & n9898 ;
  assign n9900 = n9897 & ~n9899 ;
  assign n9901 = n9900 ^ n9886 ;
  assign n9902 = ~x66 & ~n9520 ;
  assign n9903 = ~n9852 & n9884 ;
  assign n9904 = n9902 & n9903 ;
  assign n9905 = n9904 ^ x66 ;
  assign n9906 = n9882 & ~n9905 ;
  assign n9907 = x64 & n9852 ;
  assign n9908 = n9852 ^ n9520 ;
  assign n9909 = ~n9907 & ~n9908 ;
  assign n9910 = n9906 & n9909 ;
  assign n9911 = n9910 ^ n9905 ;
  assign n9912 = x64 & ~n9911 ;
  assign n9913 = n9881 ^ n9520 ;
  assign n9914 = n9520 ^ x13 ;
  assign n9915 = n9914 ^ n9852 ;
  assign n9916 = x65 ^ x13 ;
  assign n9917 = n9916 ^ n9852 ;
  assign n9918 = ~n9915 & n9917 ;
  assign n9919 = n9918 ^ n9852 ;
  assign n9920 = n9913 & n9919 ;
  assign n9921 = n9912 & n9920 ;
  assign n9922 = n9921 ^ n9911 ;
  assign n9923 = n9922 ^ x13 ;
  assign n9924 = n9923 ^ n9922 ;
  assign n9929 = ~x65 & n9921 ;
  assign n9930 = n9924 & n9929 ;
  assign n9931 = n9930 ^ n9924 ;
  assign n9932 = n9931 ^ n9923 ;
  assign n9933 = ~n9901 & n9932 ;
  assign n9936 = n9935 ^ n9933 ;
  assign n9937 = n9935 ^ x67 ;
  assign n9938 = n9936 & ~n9937 ;
  assign n9939 = n9938 ^ x67 ;
  assign n9943 = n9942 ^ n9939 ;
  assign n9944 = n9942 ^ x68 ;
  assign n9945 = n9943 & ~n9944 ;
  assign n9946 = n9945 ^ x68 ;
  assign n9950 = n9949 ^ n9946 ;
  assign n9951 = n9949 ^ x69 ;
  assign n9952 = n9950 & ~n9951 ;
  assign n9953 = n9952 ^ x69 ;
  assign n9957 = n9956 ^ n9953 ;
  assign n9958 = n9956 ^ x70 ;
  assign n9959 = n9957 & ~n9958 ;
  assign n9960 = n9959 ^ x70 ;
  assign n9964 = n9963 ^ n9960 ;
  assign n9965 = n9963 ^ x71 ;
  assign n9966 = n9964 & ~n9965 ;
  assign n9967 = n9966 ^ x71 ;
  assign n9971 = n9970 ^ n9967 ;
  assign n9972 = n9970 ^ x72 ;
  assign n9973 = n9971 & ~n9972 ;
  assign n9974 = n9973 ^ x72 ;
  assign n9978 = n9977 ^ n9974 ;
  assign n9979 = n9977 ^ x73 ;
  assign n9980 = n9978 & ~n9979 ;
  assign n9981 = n9980 ^ x73 ;
  assign n9985 = n9984 ^ n9981 ;
  assign n9986 = n9984 ^ x74 ;
  assign n9987 = n9985 & ~n9986 ;
  assign n9988 = n9987 ^ x74 ;
  assign n9992 = n9991 ^ n9988 ;
  assign n9993 = n9991 ^ x75 ;
  assign n9994 = n9992 & ~n9993 ;
  assign n9995 = n9994 ^ x75 ;
  assign n9999 = n9998 ^ n9995 ;
  assign n10000 = n9998 ^ x76 ;
  assign n10001 = n9999 & ~n10000 ;
  assign n10002 = n10001 ^ x76 ;
  assign n10006 = n10005 ^ n10002 ;
  assign n10007 = n10005 ^ x77 ;
  assign n10008 = n10006 & ~n10007 ;
  assign n10009 = n10008 ^ x77 ;
  assign n10021 = n10020 ^ n10009 ;
  assign n10022 = n10020 ^ x78 ;
  assign n10023 = n10021 & ~n10022 ;
  assign n10024 = n10023 ^ x78 ;
  assign n10028 = n10027 ^ n10024 ;
  assign n10029 = n10027 ^ x79 ;
  assign n10030 = n10028 & ~n10029 ;
  assign n10031 = n10030 ^ x79 ;
  assign n10035 = n10034 ^ n10031 ;
  assign n10036 = n10034 ^ x80 ;
  assign n10037 = n10035 & ~n10036 ;
  assign n10038 = n10037 ^ x80 ;
  assign n10042 = n10041 ^ n10038 ;
  assign n10043 = n10041 ^ x81 ;
  assign n10044 = n10042 & ~n10043 ;
  assign n10045 = n10044 ^ x81 ;
  assign n10049 = n10048 ^ n10045 ;
  assign n10050 = n10048 ^ x82 ;
  assign n10051 = n10049 & ~n10050 ;
  assign n10052 = n10051 ^ x82 ;
  assign n10056 = n10055 ^ n10052 ;
  assign n10057 = n10055 ^ x83 ;
  assign n10058 = n10056 & ~n10057 ;
  assign n10059 = n10058 ^ x83 ;
  assign n10060 = n10059 ^ n9872 ;
  assign n10061 = n10060 ^ n9878 ;
  assign n10062 = ~n9879 & n10061 ;
  assign n10063 = n10062 ^ n9878 ;
  assign n10064 = ~n9873 & n10063 ;
  assign n10065 = n10064 ^ x85 ;
  assign n10069 = n10068 ^ n10065 ;
  assign n10070 = n10068 ^ x86 ;
  assign n10071 = n10069 & ~n10070 ;
  assign n10072 = n10071 ^ x86 ;
  assign n10076 = n10075 ^ n10072 ;
  assign n10077 = n10075 ^ x87 ;
  assign n10078 = n10076 & ~n10077 ;
  assign n10079 = n10078 ^ x87 ;
  assign n10083 = n10082 ^ n10079 ;
  assign n10084 = n10082 ^ x88 ;
  assign n10085 = n10083 & ~n10084 ;
  assign n10086 = n10085 ^ x88 ;
  assign n10090 = n10089 ^ n10086 ;
  assign n10091 = n10089 ^ x89 ;
  assign n10092 = n10090 & ~n10091 ;
  assign n10093 = n10092 ^ x89 ;
  assign n10105 = n10104 ^ n10093 ;
  assign n10106 = n10104 ^ x90 ;
  assign n10107 = n10105 & ~n10106 ;
  assign n10108 = n10107 ^ x90 ;
  assign n10112 = n10111 ^ n10108 ;
  assign n10113 = n10111 ^ x91 ;
  assign n10114 = n10112 & ~n10113 ;
  assign n10115 = n10114 ^ x91 ;
  assign n10127 = n10126 ^ n10115 ;
  assign n10128 = n10126 ^ x92 ;
  assign n10129 = n10127 & ~n10128 ;
  assign n10130 = n10129 ^ x92 ;
  assign n10134 = n10133 ^ n10130 ;
  assign n10135 = n10133 ^ x93 ;
  assign n10136 = n10134 & ~n10135 ;
  assign n10137 = n10136 ^ x93 ;
  assign n10141 = n10140 ^ n10137 ;
  assign n10142 = n10140 ^ x94 ;
  assign n10143 = n10141 & ~n10142 ;
  assign n10144 = n10143 ^ x94 ;
  assign n10148 = n10147 ^ n10144 ;
  assign n10149 = n10147 ^ x95 ;
  assign n10150 = n10148 & ~n10149 ;
  assign n10151 = n10150 ^ x95 ;
  assign n10152 = n10151 ^ n9868 ;
  assign n10153 = ~n9869 & n10152 ;
  assign n10154 = n10153 ^ x96 ;
  assign n10155 = n10154 ^ n9864 ;
  assign n10156 = ~n9865 & n10155 ;
  assign n10157 = n10156 ^ x97 ;
  assign n10161 = n10160 ^ n10157 ;
  assign n10162 = n10160 ^ x98 ;
  assign n10163 = n10161 & ~n10162 ;
  assign n10164 = n10163 ^ x98 ;
  assign n10168 = n10167 ^ n10164 ;
  assign n10169 = n10167 ^ x99 ;
  assign n10170 = n10168 & ~n10169 ;
  assign n10171 = n10170 ^ x99 ;
  assign n10175 = n10174 ^ n10171 ;
  assign n10176 = n10174 ^ x100 ;
  assign n10177 = n10175 & ~n10176 ;
  assign n10178 = n10177 ^ x100 ;
  assign n10182 = n10181 ^ n10178 ;
  assign n10183 = n10181 ^ x101 ;
  assign n10184 = n10182 & ~n10183 ;
  assign n10185 = n10184 ^ x101 ;
  assign n10189 = n10188 ^ n10185 ;
  assign n10190 = n10188 ^ x102 ;
  assign n10191 = n10189 & ~n10190 ;
  assign n10192 = n10191 ^ x102 ;
  assign n10196 = n10195 ^ n10192 ;
  assign n10197 = n10195 ^ x103 ;
  assign n10198 = n10196 & ~n10197 ;
  assign n10199 = n10198 ^ x103 ;
  assign n10203 = n10202 ^ n10199 ;
  assign n10204 = n10202 ^ x104 ;
  assign n10205 = n10203 & ~n10204 ;
  assign n10206 = n10205 ^ x104 ;
  assign n10210 = n10209 ^ n10206 ;
  assign n10211 = n10209 ^ x105 ;
  assign n10212 = n10210 & ~n10211 ;
  assign n10213 = n10212 ^ x105 ;
  assign n10214 = n10213 ^ n9854 ;
  assign n10215 = n10214 ^ n9860 ;
  assign n10216 = ~n9861 & n10215 ;
  assign n10217 = n10216 ^ n9860 ;
  assign n10218 = ~n9855 & n10217 ;
  assign n10219 = n10218 ^ x107 ;
  assign n10223 = n10222 ^ n10219 ;
  assign n10224 = n10222 ^ x108 ;
  assign n10225 = n10223 & ~n10224 ;
  assign n10226 = n10225 ^ x108 ;
  assign n10230 = n10229 ^ n10226 ;
  assign n10231 = n10229 ^ x109 ;
  assign n10232 = n10230 & ~n10231 ;
  assign n10233 = n10232 ^ x109 ;
  assign n10237 = n10236 ^ n10233 ;
  assign n10238 = n10236 ^ x110 ;
  assign n10239 = n10237 & ~n10238 ;
  assign n10240 = n10239 ^ x110 ;
  assign n10244 = n10243 ^ n10240 ;
  assign n10245 = n10243 ^ x111 ;
  assign n10246 = n10244 & ~n10245 ;
  assign n10247 = n10246 ^ x111 ;
  assign n10251 = n10250 ^ n10247 ;
  assign n10252 = n10250 ^ x112 ;
  assign n10253 = n10251 & ~n10252 ;
  assign n10254 = n10253 ^ x112 ;
  assign n10258 = n10257 ^ n10254 ;
  assign n10267 = n10254 ^ x113 ;
  assign n10262 = n10258 & n10267 ;
  assign n10259 = x114 ^ x113 ;
  assign n10263 = n10262 ^ n10259 ;
  assign n10264 = n9845 & n10263 ;
  assign n10265 = n10264 ^ n9844 ;
  assign n11070 = n10265 ^ x116 ;
  assign n10266 = n10265 ^ x115 ;
  assign n10268 = n9844 ^ x114 ;
  assign n10271 = n10263 & ~n10268 ;
  assign n10272 = n10271 ^ x114 ;
  assign n10273 = n141 & ~n10272 ;
  assign n10274 = n10267 & n10273 ;
  assign n10275 = n10274 ^ n10257 ;
  assign n10277 = n10275 ^ x114 ;
  assign n10276 = x114 & ~n10275 ;
  assign n10278 = n10277 ^ n10276 ;
  assign n10279 = ~n10266 & ~n10278 ;
  assign n10650 = n10247 ^ x112 ;
  assign n10651 = n10273 & n10650 ;
  assign n10652 = n10651 ^ n10250 ;
  assign n10643 = n10240 ^ x111 ;
  assign n10644 = n10273 & n10643 ;
  assign n10645 = n10644 ^ n10243 ;
  assign n10636 = n10233 ^ x110 ;
  assign n10637 = n10273 & n10636 ;
  assign n10638 = n10637 ^ n10236 ;
  assign n10629 = n10226 ^ x109 ;
  assign n10630 = n10273 & n10629 ;
  assign n10631 = n10630 ^ n10229 ;
  assign n10622 = n10219 ^ x108 ;
  assign n10623 = n10273 & n10622 ;
  assign n10624 = n10623 ^ n10222 ;
  assign n10607 = n9858 ^ x107 ;
  assign n10608 = n10607 ^ n10213 ;
  assign n10609 = n10608 ^ x106 ;
  assign n10610 = n10609 ^ n10607 ;
  assign n10612 = n10213 ^ x107 ;
  assign n10613 = n10612 ^ n10607 ;
  assign n10614 = ~n10610 & ~n10613 ;
  assign n10615 = n10614 ^ n10607 ;
  assign n10616 = n10273 & ~n10615 ;
  assign n10617 = n10616 ^ n9854 ;
  assign n10600 = n10213 ^ x106 ;
  assign n10601 = n10273 & n10600 ;
  assign n10602 = n10601 ^ n9858 ;
  assign n10593 = n10206 ^ x105 ;
  assign n10594 = n10273 & n10593 ;
  assign n10595 = n10594 ^ n10209 ;
  assign n10586 = n10199 ^ x104 ;
  assign n10587 = n10273 & n10586 ;
  assign n10588 = n10587 ^ n10202 ;
  assign n10579 = n10192 ^ x103 ;
  assign n10580 = n10273 & n10579 ;
  assign n10581 = n10580 ^ n10195 ;
  assign n10572 = n10185 ^ x102 ;
  assign n10573 = n10273 & n10572 ;
  assign n10574 = n10573 ^ n10188 ;
  assign n10565 = n10178 ^ x101 ;
  assign n10566 = n10273 & n10565 ;
  assign n10567 = n10566 ^ n10181 ;
  assign n10280 = n10171 ^ x100 ;
  assign n10281 = n10273 & n10280 ;
  assign n10282 = n10281 ^ n10174 ;
  assign n10283 = n10282 ^ x101 ;
  assign n10288 = n10282 ^ x100 ;
  assign n10284 = n10164 ^ x99 ;
  assign n10285 = n10273 & n10284 ;
  assign n10286 = n10285 ^ n10167 ;
  assign n10287 = n10286 ^ n10282 ;
  assign n10289 = n10288 ^ n10287 ;
  assign n10552 = n10157 ^ x98 ;
  assign n10553 = n10273 & n10552 ;
  assign n10554 = n10553 ^ n10160 ;
  assign n10545 = n10154 ^ x97 ;
  assign n10546 = n10273 & n10545 ;
  assign n10547 = n10546 ^ n9864 ;
  assign n10538 = n10151 ^ x96 ;
  assign n10539 = n10273 & n10538 ;
  assign n10540 = n10539 ^ n9868 ;
  assign n10531 = n10144 ^ x95 ;
  assign n10532 = n10273 & n10531 ;
  assign n10533 = n10532 ^ n10147 ;
  assign n10524 = n10137 ^ x94 ;
  assign n10525 = n10273 & n10524 ;
  assign n10526 = n10525 ^ n10140 ;
  assign n10517 = n10130 ^ x93 ;
  assign n10518 = n10273 & n10517 ;
  assign n10519 = n10518 ^ n10133 ;
  assign n10510 = n10115 ^ x92 ;
  assign n10511 = n10273 & n10510 ;
  assign n10512 = n10511 ^ n10126 ;
  assign n10503 = n10108 ^ x91 ;
  assign n10504 = n10273 & n10503 ;
  assign n10505 = n10504 ^ n10111 ;
  assign n10496 = n10093 ^ x90 ;
  assign n10497 = n10273 & n10496 ;
  assign n10498 = n10497 ^ n10104 ;
  assign n10489 = n10086 ^ x89 ;
  assign n10490 = n10273 & n10489 ;
  assign n10491 = n10490 ^ n10089 ;
  assign n10482 = n10079 ^ x88 ;
  assign n10483 = n10273 & n10482 ;
  assign n10484 = n10483 ^ n10082 ;
  assign n10475 = n10072 ^ x87 ;
  assign n10476 = n10273 & n10475 ;
  assign n10477 = n10476 ^ n10075 ;
  assign n10468 = n10065 ^ x86 ;
  assign n10469 = n10273 & n10468 ;
  assign n10470 = n10469 ^ n10068 ;
  assign n10453 = n9876 ^ x85 ;
  assign n10454 = n10453 ^ n10059 ;
  assign n10455 = n10454 ^ x84 ;
  assign n10456 = n10455 ^ n10453 ;
  assign n10458 = n10059 ^ x85 ;
  assign n10459 = n10458 ^ n10453 ;
  assign n10460 = ~n10456 & ~n10459 ;
  assign n10461 = n10460 ^ n10453 ;
  assign n10462 = n10273 & ~n10461 ;
  assign n10463 = n10462 ^ n9872 ;
  assign n10446 = n10059 ^ x84 ;
  assign n10447 = n10273 & n10446 ;
  assign n10448 = n10447 ^ n9876 ;
  assign n10439 = n10052 ^ x83 ;
  assign n10440 = n10273 & n10439 ;
  assign n10441 = n10440 ^ n10055 ;
  assign n10432 = n10045 ^ x82 ;
  assign n10433 = n10273 & n10432 ;
  assign n10434 = n10433 ^ n10048 ;
  assign n10425 = n10038 ^ x81 ;
  assign n10426 = n10273 & n10425 ;
  assign n10427 = n10426 ^ n10041 ;
  assign n10418 = n10031 ^ x80 ;
  assign n10419 = n10273 & n10418 ;
  assign n10420 = n10419 ^ n10034 ;
  assign n10411 = n10024 ^ x79 ;
  assign n10412 = n10273 & n10411 ;
  assign n10413 = n10412 ^ n10027 ;
  assign n10404 = n10009 ^ x78 ;
  assign n10405 = n10273 & n10404 ;
  assign n10406 = n10405 ^ n10020 ;
  assign n10397 = n10002 ^ x77 ;
  assign n10398 = n10273 & n10397 ;
  assign n10399 = n10398 ^ n10005 ;
  assign n10390 = n9995 ^ x76 ;
  assign n10391 = n10273 & n10390 ;
  assign n10392 = n10391 ^ n9998 ;
  assign n10290 = n9988 ^ x75 ;
  assign n10291 = n10273 & n10290 ;
  assign n10292 = n10291 ^ n9991 ;
  assign n10293 = n10292 ^ x76 ;
  assign n10298 = n10292 ^ x75 ;
  assign n10294 = n9981 ^ x74 ;
  assign n10295 = n10273 & n10294 ;
  assign n10296 = n10295 ^ n9984 ;
  assign n10297 = n10296 ^ n10292 ;
  assign n10299 = n10298 ^ n10297 ;
  assign n10377 = n9974 ^ x73 ;
  assign n10378 = n10273 & n10377 ;
  assign n10379 = n10378 ^ n9977 ;
  assign n10370 = n9967 ^ x72 ;
  assign n10371 = n10273 & n10370 ;
  assign n10372 = n10371 ^ n9970 ;
  assign n10363 = n9960 ^ x71 ;
  assign n10364 = n10273 & n10363 ;
  assign n10365 = n10364 ^ n9963 ;
  assign n10356 = n9953 ^ x70 ;
  assign n10357 = n10273 & n10356 ;
  assign n10358 = n10357 ^ n9956 ;
  assign n10349 = n9946 ^ x69 ;
  assign n10350 = n10273 & n10349 ;
  assign n10351 = n10350 ^ n9949 ;
  assign n10342 = n9939 ^ x68 ;
  assign n10343 = n10273 & n10342 ;
  assign n10344 = n10343 ^ n9942 ;
  assign n10335 = n9933 ^ x67 ;
  assign n10336 = n10273 & n10335 ;
  assign n10337 = n10336 ^ n9935 ;
  assign n10302 = n9907 ^ x14 ;
  assign n10300 = n9883 ^ x65 ;
  assign n10301 = n10273 & n10300 ;
  assign n10303 = n10302 ^ n10301 ;
  assign n10304 = n10303 ^ x66 ;
  assign n10310 = n1228 & n10273 ;
  assign n10306 = n9883 ^ n1228 ;
  assign n10305 = x64 & n10273 ;
  assign n10307 = n10306 ^ n10305 ;
  assign n10308 = ~x12 & n10307 ;
  assign n10309 = n10308 ^ n9890 ;
  assign n10311 = n10310 ^ n10309 ;
  assign n10312 = n10311 ^ n10303 ;
  assign n10313 = ~n10304 & n10312 ;
  assign n10314 = n10313 ^ x66 ;
  assign n10315 = n10314 ^ x67 ;
  assign n10330 = n9518 & n9852 ;
  assign n10324 = x14 & x65 ;
  assign n10316 = n9888 ^ x65 ;
  assign n10317 = n10316 ^ n9852 ;
  assign n10318 = ~n9916 & n10317 ;
  assign n10325 = n10324 ^ n10318 ;
  assign n10326 = ~x64 & n10325 ;
  assign n10321 = n10318 ^ n7358 ;
  assign n10327 = n10326 ^ n10321 ;
  assign n10328 = n10273 & n10327 ;
  assign n10329 = n10328 ^ n9520 ;
  assign n10331 = n10330 ^ n10329 ;
  assign n10332 = n10331 ^ n10314 ;
  assign n10333 = n10315 & n10332 ;
  assign n10334 = n10333 ^ x67 ;
  assign n10338 = n10337 ^ n10334 ;
  assign n10339 = n10337 ^ x68 ;
  assign n10340 = n10338 & ~n10339 ;
  assign n10341 = n10340 ^ x68 ;
  assign n10345 = n10344 ^ n10341 ;
  assign n10346 = n10344 ^ x69 ;
  assign n10347 = n10345 & ~n10346 ;
  assign n10348 = n10347 ^ x69 ;
  assign n10352 = n10351 ^ n10348 ;
  assign n10353 = n10351 ^ x70 ;
  assign n10354 = n10352 & ~n10353 ;
  assign n10355 = n10354 ^ x70 ;
  assign n10359 = n10358 ^ n10355 ;
  assign n10360 = n10358 ^ x71 ;
  assign n10361 = n10359 & ~n10360 ;
  assign n10362 = n10361 ^ x71 ;
  assign n10366 = n10365 ^ n10362 ;
  assign n10367 = n10365 ^ x72 ;
  assign n10368 = n10366 & ~n10367 ;
  assign n10369 = n10368 ^ x72 ;
  assign n10373 = n10372 ^ n10369 ;
  assign n10374 = n10372 ^ x73 ;
  assign n10375 = n10373 & ~n10374 ;
  assign n10376 = n10375 ^ x73 ;
  assign n10380 = n10379 ^ n10376 ;
  assign n10381 = n10379 ^ x74 ;
  assign n10382 = n10380 & ~n10381 ;
  assign n10383 = n10382 ^ x74 ;
  assign n10384 = n10383 ^ n10292 ;
  assign n10385 = n10384 ^ n10298 ;
  assign n10386 = ~n10299 & n10385 ;
  assign n10387 = n10386 ^ n10298 ;
  assign n10388 = ~n10293 & n10387 ;
  assign n10389 = n10388 ^ x76 ;
  assign n10393 = n10392 ^ n10389 ;
  assign n10394 = n10392 ^ x77 ;
  assign n10395 = n10393 & ~n10394 ;
  assign n10396 = n10395 ^ x77 ;
  assign n10400 = n10399 ^ n10396 ;
  assign n10401 = n10399 ^ x78 ;
  assign n10402 = n10400 & ~n10401 ;
  assign n10403 = n10402 ^ x78 ;
  assign n10407 = n10406 ^ n10403 ;
  assign n10408 = n10406 ^ x79 ;
  assign n10409 = n10407 & ~n10408 ;
  assign n10410 = n10409 ^ x79 ;
  assign n10414 = n10413 ^ n10410 ;
  assign n10415 = n10413 ^ x80 ;
  assign n10416 = n10414 & ~n10415 ;
  assign n10417 = n10416 ^ x80 ;
  assign n10421 = n10420 ^ n10417 ;
  assign n10422 = n10420 ^ x81 ;
  assign n10423 = n10421 & ~n10422 ;
  assign n10424 = n10423 ^ x81 ;
  assign n10428 = n10427 ^ n10424 ;
  assign n10429 = n10427 ^ x82 ;
  assign n10430 = n10428 & ~n10429 ;
  assign n10431 = n10430 ^ x82 ;
  assign n10435 = n10434 ^ n10431 ;
  assign n10436 = n10434 ^ x83 ;
  assign n10437 = n10435 & ~n10436 ;
  assign n10438 = n10437 ^ x83 ;
  assign n10442 = n10441 ^ n10438 ;
  assign n10443 = n10441 ^ x84 ;
  assign n10444 = n10442 & ~n10443 ;
  assign n10445 = n10444 ^ x84 ;
  assign n10449 = n10448 ^ n10445 ;
  assign n10450 = n10448 ^ x85 ;
  assign n10451 = n10449 & ~n10450 ;
  assign n10452 = n10451 ^ x85 ;
  assign n10464 = n10463 ^ n10452 ;
  assign n10465 = n10463 ^ x86 ;
  assign n10466 = n10464 & ~n10465 ;
  assign n10467 = n10466 ^ x86 ;
  assign n10471 = n10470 ^ n10467 ;
  assign n10472 = n10470 ^ x87 ;
  assign n10473 = n10471 & ~n10472 ;
  assign n10474 = n10473 ^ x87 ;
  assign n10478 = n10477 ^ n10474 ;
  assign n10479 = n10477 ^ x88 ;
  assign n10480 = n10478 & ~n10479 ;
  assign n10481 = n10480 ^ x88 ;
  assign n10485 = n10484 ^ n10481 ;
  assign n10486 = n10484 ^ x89 ;
  assign n10487 = n10485 & ~n10486 ;
  assign n10488 = n10487 ^ x89 ;
  assign n10492 = n10491 ^ n10488 ;
  assign n10493 = n10491 ^ x90 ;
  assign n10494 = n10492 & ~n10493 ;
  assign n10495 = n10494 ^ x90 ;
  assign n10499 = n10498 ^ n10495 ;
  assign n10500 = n10498 ^ x91 ;
  assign n10501 = n10499 & ~n10500 ;
  assign n10502 = n10501 ^ x91 ;
  assign n10506 = n10505 ^ n10502 ;
  assign n10507 = n10505 ^ x92 ;
  assign n10508 = n10506 & ~n10507 ;
  assign n10509 = n10508 ^ x92 ;
  assign n10513 = n10512 ^ n10509 ;
  assign n10514 = n10512 ^ x93 ;
  assign n10515 = n10513 & ~n10514 ;
  assign n10516 = n10515 ^ x93 ;
  assign n10520 = n10519 ^ n10516 ;
  assign n10521 = n10519 ^ x94 ;
  assign n10522 = n10520 & ~n10521 ;
  assign n10523 = n10522 ^ x94 ;
  assign n10527 = n10526 ^ n10523 ;
  assign n10528 = n10526 ^ x95 ;
  assign n10529 = n10527 & ~n10528 ;
  assign n10530 = n10529 ^ x95 ;
  assign n10534 = n10533 ^ n10530 ;
  assign n10535 = n10533 ^ x96 ;
  assign n10536 = n10534 & ~n10535 ;
  assign n10537 = n10536 ^ x96 ;
  assign n10541 = n10540 ^ n10537 ;
  assign n10542 = n10540 ^ x97 ;
  assign n10543 = n10541 & ~n10542 ;
  assign n10544 = n10543 ^ x97 ;
  assign n10548 = n10547 ^ n10544 ;
  assign n10549 = n10547 ^ x98 ;
  assign n10550 = n10548 & ~n10549 ;
  assign n10551 = n10550 ^ x98 ;
  assign n10555 = n10554 ^ n10551 ;
  assign n10556 = n10554 ^ x99 ;
  assign n10557 = n10555 & ~n10556 ;
  assign n10558 = n10557 ^ x99 ;
  assign n10559 = n10558 ^ n10282 ;
  assign n10560 = n10559 ^ n10288 ;
  assign n10561 = ~n10289 & n10560 ;
  assign n10562 = n10561 ^ n10288 ;
  assign n10563 = ~n10283 & n10562 ;
  assign n10564 = n10563 ^ x101 ;
  assign n10568 = n10567 ^ n10564 ;
  assign n10569 = n10567 ^ x102 ;
  assign n10570 = n10568 & ~n10569 ;
  assign n10571 = n10570 ^ x102 ;
  assign n10575 = n10574 ^ n10571 ;
  assign n10576 = n10574 ^ x103 ;
  assign n10577 = n10575 & ~n10576 ;
  assign n10578 = n10577 ^ x103 ;
  assign n10582 = n10581 ^ n10578 ;
  assign n10583 = n10581 ^ x104 ;
  assign n10584 = n10582 & ~n10583 ;
  assign n10585 = n10584 ^ x104 ;
  assign n10589 = n10588 ^ n10585 ;
  assign n10590 = n10588 ^ x105 ;
  assign n10591 = n10589 & ~n10590 ;
  assign n10592 = n10591 ^ x105 ;
  assign n10596 = n10595 ^ n10592 ;
  assign n10597 = n10595 ^ x106 ;
  assign n10598 = n10596 & ~n10597 ;
  assign n10599 = n10598 ^ x106 ;
  assign n10603 = n10602 ^ n10599 ;
  assign n10604 = n10602 ^ x107 ;
  assign n10605 = n10603 & ~n10604 ;
  assign n10606 = n10605 ^ x107 ;
  assign n10618 = n10617 ^ n10606 ;
  assign n10619 = n10617 ^ x108 ;
  assign n10620 = n10618 & ~n10619 ;
  assign n10621 = n10620 ^ x108 ;
  assign n10625 = n10624 ^ n10621 ;
  assign n10626 = n10624 ^ x109 ;
  assign n10627 = n10625 & ~n10626 ;
  assign n10628 = n10627 ^ x109 ;
  assign n10632 = n10631 ^ n10628 ;
  assign n10633 = n10631 ^ x110 ;
  assign n10634 = n10632 & ~n10633 ;
  assign n10635 = n10634 ^ x110 ;
  assign n10639 = n10638 ^ n10635 ;
  assign n10640 = n10638 ^ x111 ;
  assign n10641 = n10639 & ~n10640 ;
  assign n10642 = n10641 ^ x111 ;
  assign n10646 = n10645 ^ n10642 ;
  assign n10647 = n10645 ^ x112 ;
  assign n10648 = n10646 & ~n10647 ;
  assign n10649 = n10648 ^ x112 ;
  assign n10653 = n10652 ^ n10649 ;
  assign n10654 = n10652 ^ x113 ;
  assign n10655 = n10653 & ~n10654 ;
  assign n10656 = n10655 ^ x113 ;
  assign n10657 = n10279 & n10656 ;
  assign n10658 = n10276 ^ x115 ;
  assign n10659 = ~n10266 & n10658 ;
  assign n10660 = n10659 ^ x115 ;
  assign n10661 = n140 & ~n10660 ;
  assign n10662 = ~n10657 & n10661 ;
  assign n10663 = n10656 ^ x114 ;
  assign n10664 = n10662 & n10663 ;
  assign n10665 = n10664 ^ n10275 ;
  assign n10667 = n10665 ^ x115 ;
  assign n10666 = ~x115 & n10665 ;
  assign n10668 = n10667 ^ n10666 ;
  assign n11040 = n10649 ^ x113 ;
  assign n11041 = n10662 & n11040 ;
  assign n11042 = n11041 ^ n10652 ;
  assign n11033 = n10642 ^ x112 ;
  assign n11034 = n10662 & n11033 ;
  assign n11035 = n11034 ^ n10645 ;
  assign n11026 = n10635 ^ x111 ;
  assign n11027 = n10662 & n11026 ;
  assign n11028 = n11027 ^ n10638 ;
  assign n11019 = n10628 ^ x110 ;
  assign n11020 = n10662 & n11019 ;
  assign n11021 = n11020 ^ n10631 ;
  assign n11012 = n10621 ^ x109 ;
  assign n11013 = n10662 & n11012 ;
  assign n11014 = n11013 ^ n10624 ;
  assign n11005 = n10606 ^ x108 ;
  assign n11006 = n10662 & n11005 ;
  assign n11007 = n11006 ^ n10617 ;
  assign n10998 = n10599 ^ x107 ;
  assign n10999 = n10662 & n10998 ;
  assign n11000 = n10999 ^ n10602 ;
  assign n10991 = n10592 ^ x106 ;
  assign n10992 = n10662 & n10991 ;
  assign n10993 = n10992 ^ n10595 ;
  assign n10984 = n10585 ^ x105 ;
  assign n10985 = n10662 & n10984 ;
  assign n10986 = n10985 ^ n10588 ;
  assign n10977 = n10578 ^ x104 ;
  assign n10978 = n10662 & n10977 ;
  assign n10979 = n10978 ^ n10581 ;
  assign n10970 = n10571 ^ x103 ;
  assign n10971 = n10662 & n10970 ;
  assign n10972 = n10971 ^ n10574 ;
  assign n10963 = n10564 ^ x102 ;
  assign n10964 = n10662 & n10963 ;
  assign n10965 = n10964 ^ n10567 ;
  assign n10948 = n10286 ^ x101 ;
  assign n10949 = n10948 ^ x100 ;
  assign n10950 = n10949 ^ n10558 ;
  assign n10951 = n10950 ^ n10948 ;
  assign n10953 = x101 ^ x100 ;
  assign n10954 = n10953 ^ n10948 ;
  assign n10955 = ~n10951 & ~n10954 ;
  assign n10956 = n10955 ^ n10948 ;
  assign n10957 = n10662 & ~n10956 ;
  assign n10958 = n10957 ^ n10282 ;
  assign n10669 = n10558 ^ x100 ;
  assign n10670 = n10662 & n10669 ;
  assign n10671 = n10670 ^ n10286 ;
  assign n10672 = n10671 ^ x101 ;
  assign n10677 = n10671 ^ x100 ;
  assign n10673 = n10551 ^ x99 ;
  assign n10674 = n10662 & n10673 ;
  assign n10675 = n10674 ^ n10554 ;
  assign n10676 = n10675 ^ n10671 ;
  assign n10678 = n10677 ^ n10676 ;
  assign n10935 = n10544 ^ x98 ;
  assign n10936 = n10662 & n10935 ;
  assign n10937 = n10936 ^ n10547 ;
  assign n10928 = n10537 ^ x97 ;
  assign n10929 = n10662 & n10928 ;
  assign n10930 = n10929 ^ n10540 ;
  assign n10921 = n10530 ^ x96 ;
  assign n10922 = n10662 & n10921 ;
  assign n10923 = n10922 ^ n10533 ;
  assign n10914 = n10523 ^ x95 ;
  assign n10915 = n10662 & n10914 ;
  assign n10916 = n10915 ^ n10526 ;
  assign n10907 = n10516 ^ x94 ;
  assign n10908 = n10662 & n10907 ;
  assign n10909 = n10908 ^ n10519 ;
  assign n10900 = n10509 ^ x93 ;
  assign n10901 = n10662 & n10900 ;
  assign n10902 = n10901 ^ n10512 ;
  assign n10893 = n10502 ^ x92 ;
  assign n10894 = n10662 & n10893 ;
  assign n10895 = n10894 ^ n10505 ;
  assign n10886 = n10495 ^ x91 ;
  assign n10887 = n10662 & n10886 ;
  assign n10888 = n10887 ^ n10498 ;
  assign n10879 = n10488 ^ x90 ;
  assign n10880 = n10662 & n10879 ;
  assign n10881 = n10880 ^ n10491 ;
  assign n10872 = n10481 ^ x89 ;
  assign n10873 = n10662 & n10872 ;
  assign n10874 = n10873 ^ n10484 ;
  assign n10865 = n10474 ^ x88 ;
  assign n10866 = n10662 & n10865 ;
  assign n10867 = n10866 ^ n10477 ;
  assign n10858 = n10467 ^ x87 ;
  assign n10859 = n10662 & n10858 ;
  assign n10860 = n10859 ^ n10470 ;
  assign n10851 = n10452 ^ x86 ;
  assign n10852 = n10662 & n10851 ;
  assign n10853 = n10852 ^ n10463 ;
  assign n10844 = n10445 ^ x85 ;
  assign n10845 = n10662 & n10844 ;
  assign n10846 = n10845 ^ n10448 ;
  assign n10837 = n10438 ^ x84 ;
  assign n10838 = n10662 & n10837 ;
  assign n10839 = n10838 ^ n10441 ;
  assign n10830 = n10431 ^ x83 ;
  assign n10831 = n10662 & n10830 ;
  assign n10832 = n10831 ^ n10434 ;
  assign n10823 = n10424 ^ x82 ;
  assign n10824 = n10662 & n10823 ;
  assign n10825 = n10824 ^ n10427 ;
  assign n10816 = n10417 ^ x81 ;
  assign n10817 = n10662 & n10816 ;
  assign n10818 = n10817 ^ n10420 ;
  assign n10809 = n10410 ^ x80 ;
  assign n10810 = n10662 & n10809 ;
  assign n10811 = n10810 ^ n10413 ;
  assign n10802 = n10403 ^ x79 ;
  assign n10803 = n10662 & n10802 ;
  assign n10804 = n10803 ^ n10406 ;
  assign n10679 = n10396 ^ x78 ;
  assign n10680 = n10662 & n10679 ;
  assign n10681 = n10680 ^ n10399 ;
  assign n10682 = n10681 ^ x79 ;
  assign n10687 = n10681 ^ x78 ;
  assign n10683 = n10389 ^ x77 ;
  assign n10684 = n10662 & n10683 ;
  assign n10685 = n10684 ^ n10392 ;
  assign n10686 = n10685 ^ n10681 ;
  assign n10688 = n10687 ^ n10686 ;
  assign n10689 = n10296 ^ x76 ;
  assign n10690 = n10689 ^ x75 ;
  assign n10691 = n10690 ^ n10383 ;
  assign n10692 = n10691 ^ n10689 ;
  assign n10695 = n10689 ^ n888 ;
  assign n10696 = ~n10692 & ~n10695 ;
  assign n10697 = n10696 ^ n10689 ;
  assign n10698 = n10662 & ~n10697 ;
  assign n10699 = n10698 ^ n10292 ;
  assign n10700 = n10699 ^ x77 ;
  assign n10786 = n10383 ^ x75 ;
  assign n10787 = n10662 & n10786 ;
  assign n10788 = n10787 ^ n10296 ;
  assign n10779 = n10376 ^ x74 ;
  assign n10780 = n10662 & n10779 ;
  assign n10781 = n10780 ^ n10379 ;
  assign n10772 = n10369 ^ x73 ;
  assign n10773 = n10662 & n10772 ;
  assign n10774 = n10773 ^ n10372 ;
  assign n10701 = n10362 ^ x72 ;
  assign n10702 = n10662 & n10701 ;
  assign n10703 = n10702 ^ n10365 ;
  assign n10704 = n10703 ^ x73 ;
  assign n10705 = n10355 ^ x71 ;
  assign n10706 = n10662 & n10705 ;
  assign n10707 = n10706 ^ n10358 ;
  assign n10708 = n10707 ^ x72 ;
  assign n10759 = n10348 ^ x70 ;
  assign n10760 = n10662 & n10759 ;
  assign n10761 = n10760 ^ n10351 ;
  assign n10752 = n10341 ^ x69 ;
  assign n10753 = n10662 & n10752 ;
  assign n10754 = n10753 ^ n10344 ;
  assign n10745 = n10334 ^ x68 ;
  assign n10746 = n10662 & n10745 ;
  assign n10747 = n10746 ^ n10337 ;
  assign n10739 = n10315 & n10662 ;
  assign n10740 = n10739 ^ n10331 ;
  assign n10732 = n10311 ^ x66 ;
  assign n10733 = n10662 & n10732 ;
  assign n10734 = n10733 ^ n10303 ;
  assign n10714 = n10305 ^ x13 ;
  assign n10711 = ~x12 & x64 ;
  assign n10712 = n10711 ^ x65 ;
  assign n10713 = n10662 & n10712 ;
  assign n10715 = n10714 ^ n10713 ;
  assign n10716 = n10715 ^ x66 ;
  assign n10724 = x12 & x65 ;
  assign n10721 = x65 ^ x11 ;
  assign n10717 = x64 ^ x12 ;
  assign n10718 = n10717 ^ x65 ;
  assign n10722 = n10718 ^ n10662 ;
  assign n10723 = ~n10721 & n10722 ;
  assign n10725 = n10724 ^ n10723 ;
  assign n10726 = x64 & n10725 ;
  assign n10727 = n10726 ^ n10724 ;
  assign n10728 = n10727 ^ x65 ;
  assign n10729 = n10728 ^ n10715 ;
  assign n10730 = ~n10716 & n10729 ;
  assign n10731 = n10730 ^ x66 ;
  assign n10735 = n10734 ^ n10731 ;
  assign n10736 = n10734 ^ x67 ;
  assign n10737 = n10735 & ~n10736 ;
  assign n10738 = n10737 ^ x67 ;
  assign n10741 = n10740 ^ n10738 ;
  assign n10742 = n10740 ^ x68 ;
  assign n10743 = n10741 & ~n10742 ;
  assign n10744 = n10743 ^ x68 ;
  assign n10748 = n10747 ^ n10744 ;
  assign n10749 = n10747 ^ x69 ;
  assign n10750 = n10748 & ~n10749 ;
  assign n10751 = n10750 ^ x69 ;
  assign n10755 = n10754 ^ n10751 ;
  assign n10756 = n10754 ^ x70 ;
  assign n10757 = n10755 & ~n10756 ;
  assign n10758 = n10757 ^ x70 ;
  assign n10762 = n10761 ^ n10758 ;
  assign n10763 = n10761 ^ x71 ;
  assign n10764 = n10762 & ~n10763 ;
  assign n10765 = n10764 ^ x71 ;
  assign n10766 = n10765 ^ n10707 ;
  assign n10767 = ~n10708 & n10766 ;
  assign n10768 = n10767 ^ x72 ;
  assign n10769 = n10768 ^ n10703 ;
  assign n10770 = ~n10704 & n10769 ;
  assign n10771 = n10770 ^ x73 ;
  assign n10775 = n10774 ^ n10771 ;
  assign n10776 = n10774 ^ x74 ;
  assign n10777 = n10775 & ~n10776 ;
  assign n10778 = n10777 ^ x74 ;
  assign n10782 = n10781 ^ n10778 ;
  assign n10783 = n10781 ^ x75 ;
  assign n10784 = n10782 & ~n10783 ;
  assign n10785 = n10784 ^ x75 ;
  assign n10789 = n10788 ^ n10785 ;
  assign n10790 = n10788 ^ x76 ;
  assign n10791 = n10789 & ~n10790 ;
  assign n10792 = n10791 ^ x76 ;
  assign n10793 = n10792 ^ n10699 ;
  assign n10794 = ~n10700 & n10793 ;
  assign n10795 = n10794 ^ x77 ;
  assign n10796 = n10795 ^ n10681 ;
  assign n10797 = n10796 ^ n10687 ;
  assign n10798 = ~n10688 & n10797 ;
  assign n10799 = n10798 ^ n10687 ;
  assign n10800 = ~n10682 & n10799 ;
  assign n10801 = n10800 ^ x79 ;
  assign n10805 = n10804 ^ n10801 ;
  assign n10806 = n10804 ^ x80 ;
  assign n10807 = n10805 & ~n10806 ;
  assign n10808 = n10807 ^ x80 ;
  assign n10812 = n10811 ^ n10808 ;
  assign n10813 = n10811 ^ x81 ;
  assign n10814 = n10812 & ~n10813 ;
  assign n10815 = n10814 ^ x81 ;
  assign n10819 = n10818 ^ n10815 ;
  assign n10820 = n10818 ^ x82 ;
  assign n10821 = n10819 & ~n10820 ;
  assign n10822 = n10821 ^ x82 ;
  assign n10826 = n10825 ^ n10822 ;
  assign n10827 = n10825 ^ x83 ;
  assign n10828 = n10826 & ~n10827 ;
  assign n10829 = n10828 ^ x83 ;
  assign n10833 = n10832 ^ n10829 ;
  assign n10834 = n10832 ^ x84 ;
  assign n10835 = n10833 & ~n10834 ;
  assign n10836 = n10835 ^ x84 ;
  assign n10840 = n10839 ^ n10836 ;
  assign n10841 = n10839 ^ x85 ;
  assign n10842 = n10840 & ~n10841 ;
  assign n10843 = n10842 ^ x85 ;
  assign n10847 = n10846 ^ n10843 ;
  assign n10848 = n10846 ^ x86 ;
  assign n10849 = n10847 & ~n10848 ;
  assign n10850 = n10849 ^ x86 ;
  assign n10854 = n10853 ^ n10850 ;
  assign n10855 = n10853 ^ x87 ;
  assign n10856 = n10854 & ~n10855 ;
  assign n10857 = n10856 ^ x87 ;
  assign n10861 = n10860 ^ n10857 ;
  assign n10862 = n10860 ^ x88 ;
  assign n10863 = n10861 & ~n10862 ;
  assign n10864 = n10863 ^ x88 ;
  assign n10868 = n10867 ^ n10864 ;
  assign n10869 = n10867 ^ x89 ;
  assign n10870 = n10868 & ~n10869 ;
  assign n10871 = n10870 ^ x89 ;
  assign n10875 = n10874 ^ n10871 ;
  assign n10876 = n10874 ^ x90 ;
  assign n10877 = n10875 & ~n10876 ;
  assign n10878 = n10877 ^ x90 ;
  assign n10882 = n10881 ^ n10878 ;
  assign n10883 = n10881 ^ x91 ;
  assign n10884 = n10882 & ~n10883 ;
  assign n10885 = n10884 ^ x91 ;
  assign n10889 = n10888 ^ n10885 ;
  assign n10890 = n10888 ^ x92 ;
  assign n10891 = n10889 & ~n10890 ;
  assign n10892 = n10891 ^ x92 ;
  assign n10896 = n10895 ^ n10892 ;
  assign n10897 = n10895 ^ x93 ;
  assign n10898 = n10896 & ~n10897 ;
  assign n10899 = n10898 ^ x93 ;
  assign n10903 = n10902 ^ n10899 ;
  assign n10904 = n10902 ^ x94 ;
  assign n10905 = n10903 & ~n10904 ;
  assign n10906 = n10905 ^ x94 ;
  assign n10910 = n10909 ^ n10906 ;
  assign n10911 = n10909 ^ x95 ;
  assign n10912 = n10910 & ~n10911 ;
  assign n10913 = n10912 ^ x95 ;
  assign n10917 = n10916 ^ n10913 ;
  assign n10918 = n10916 ^ x96 ;
  assign n10919 = n10917 & ~n10918 ;
  assign n10920 = n10919 ^ x96 ;
  assign n10924 = n10923 ^ n10920 ;
  assign n10925 = n10923 ^ x97 ;
  assign n10926 = n10924 & ~n10925 ;
  assign n10927 = n10926 ^ x97 ;
  assign n10931 = n10930 ^ n10927 ;
  assign n10932 = n10930 ^ x98 ;
  assign n10933 = n10931 & ~n10932 ;
  assign n10934 = n10933 ^ x98 ;
  assign n10938 = n10937 ^ n10934 ;
  assign n10939 = n10937 ^ x99 ;
  assign n10940 = n10938 & ~n10939 ;
  assign n10941 = n10940 ^ x99 ;
  assign n10942 = n10941 ^ n10671 ;
  assign n10943 = n10942 ^ n10677 ;
  assign n10944 = ~n10678 & n10943 ;
  assign n10945 = n10944 ^ n10677 ;
  assign n10946 = ~n10672 & n10945 ;
  assign n10947 = n10946 ^ x101 ;
  assign n10959 = n10958 ^ n10947 ;
  assign n10960 = n10958 ^ x102 ;
  assign n10961 = n10959 & ~n10960 ;
  assign n10962 = n10961 ^ x102 ;
  assign n10966 = n10965 ^ n10962 ;
  assign n10967 = n10965 ^ x103 ;
  assign n10968 = n10966 & ~n10967 ;
  assign n10969 = n10968 ^ x103 ;
  assign n10973 = n10972 ^ n10969 ;
  assign n10974 = n10972 ^ x104 ;
  assign n10975 = n10973 & ~n10974 ;
  assign n10976 = n10975 ^ x104 ;
  assign n10980 = n10979 ^ n10976 ;
  assign n10981 = n10979 ^ x105 ;
  assign n10982 = n10980 & ~n10981 ;
  assign n10983 = n10982 ^ x105 ;
  assign n10987 = n10986 ^ n10983 ;
  assign n10988 = n10986 ^ x106 ;
  assign n10989 = n10987 & ~n10988 ;
  assign n10990 = n10989 ^ x106 ;
  assign n10994 = n10993 ^ n10990 ;
  assign n10995 = n10993 ^ x107 ;
  assign n10996 = n10994 & ~n10995 ;
  assign n10997 = n10996 ^ x107 ;
  assign n11001 = n11000 ^ n10997 ;
  assign n11002 = n11000 ^ x108 ;
  assign n11003 = n11001 & ~n11002 ;
  assign n11004 = n11003 ^ x108 ;
  assign n11008 = n11007 ^ n11004 ;
  assign n11009 = n11007 ^ x109 ;
  assign n11010 = n11008 & ~n11009 ;
  assign n11011 = n11010 ^ x109 ;
  assign n11015 = n11014 ^ n11011 ;
  assign n11016 = n11014 ^ x110 ;
  assign n11017 = n11015 & ~n11016 ;
  assign n11018 = n11017 ^ x110 ;
  assign n11022 = n11021 ^ n11018 ;
  assign n11023 = n11021 ^ x111 ;
  assign n11024 = n11022 & ~n11023 ;
  assign n11025 = n11024 ^ x111 ;
  assign n11029 = n11028 ^ n11025 ;
  assign n11030 = n11028 ^ x112 ;
  assign n11031 = n11029 & ~n11030 ;
  assign n11032 = n11031 ^ x112 ;
  assign n11036 = n11035 ^ n11032 ;
  assign n11037 = n11035 ^ x113 ;
  assign n11038 = n11036 & ~n11037 ;
  assign n11039 = n11038 ^ x113 ;
  assign n11043 = n11042 ^ n11039 ;
  assign n11044 = n11042 ^ x114 ;
  assign n11045 = n11043 & ~n11044 ;
  assign n11046 = n11045 ^ x114 ;
  assign n11047 = ~n10668 & ~n11046 ;
  assign n11071 = n11070 ^ n11047 ;
  assign n11072 = n11071 ^ n10265 ;
  assign n11083 = n11072 ^ x116 ;
  assign n11073 = n11072 ^ n11070 ;
  assign n11074 = n11073 ^ n10666 ;
  assign n11075 = n11074 ^ n11073 ;
  assign n11084 = n11083 ^ n11075 ;
  assign n11085 = n11084 ^ n11070 ;
  assign n11087 = n11083 & ~n11085 ;
  assign n11054 = n10656 ^ n10275 ;
  assign n11058 = n10663 & n11054 ;
  assign n11055 = x115 ^ x114 ;
  assign n11059 = n11058 ^ n11055 ;
  assign n11076 = n11075 ^ n11059 ;
  assign n11079 = n11075 ^ n11070 ;
  assign n11078 = n11072 ^ n11059 ;
  assign n11080 = n11079 ^ n11078 ;
  assign n11081 = ~n11076 & n11080 ;
  assign n11088 = n11087 ^ n11081 ;
  assign n11089 = n11088 ^ n11079 ;
  assign n11090 = n11087 ^ n11072 ;
  assign n11091 = n11090 ^ n11079 ;
  assign n11092 = ~n11089 & n11091 ;
  assign n11093 = n11070 & n11092 ;
  assign n11094 = n11093 ^ n11087 ;
  assign n11095 = n11094 ^ n11085 ;
  assign n11096 = n11095 ^ x116 ;
  assign n11105 = n11096 ^ n10265 ;
  assign n11106 = n139 & n11105 ;
  assign n11494 = n11046 ^ x115 ;
  assign n11495 = n11106 & n11494 ;
  assign n11496 = n11495 ^ n10665 ;
  assign n11487 = n11039 ^ x114 ;
  assign n11488 = n11106 & n11487 ;
  assign n11489 = n11488 ^ n11042 ;
  assign n11480 = n11032 ^ x113 ;
  assign n11481 = n11106 & n11480 ;
  assign n11482 = n11481 ^ n11035 ;
  assign n11069 = n11025 ^ x112 ;
  assign n11107 = n11069 & n11106 ;
  assign n11108 = n11107 ^ n11028 ;
  assign n11109 = n11108 ^ x113 ;
  assign n11114 = n11108 ^ x112 ;
  assign n11110 = n11018 ^ x111 ;
  assign n11111 = n11106 & n11110 ;
  assign n11112 = n11111 ^ n11021 ;
  assign n11113 = n11112 ^ n11108 ;
  assign n11115 = n11114 ^ n11113 ;
  assign n11467 = n11011 ^ x110 ;
  assign n11468 = n11106 & n11467 ;
  assign n11469 = n11468 ^ n11014 ;
  assign n11460 = n11004 ^ x109 ;
  assign n11461 = n11106 & n11460 ;
  assign n11462 = n11461 ^ n11007 ;
  assign n11453 = n10997 ^ x108 ;
  assign n11454 = n11106 & n11453 ;
  assign n11455 = n11454 ^ n11000 ;
  assign n11446 = n10990 ^ x107 ;
  assign n11447 = n11106 & n11446 ;
  assign n11448 = n11447 ^ n10993 ;
  assign n11439 = n10983 ^ x106 ;
  assign n11440 = n11106 & n11439 ;
  assign n11441 = n11440 ^ n10986 ;
  assign n11432 = n10976 ^ x105 ;
  assign n11433 = n11106 & n11432 ;
  assign n11434 = n11433 ^ n10979 ;
  assign n11425 = n10969 ^ x104 ;
  assign n11426 = n11106 & n11425 ;
  assign n11427 = n11426 ^ n10972 ;
  assign n11418 = n10962 ^ x103 ;
  assign n11419 = n11106 & n11418 ;
  assign n11420 = n11419 ^ n10965 ;
  assign n11411 = n10947 ^ x102 ;
  assign n11412 = n11106 & n11411 ;
  assign n11413 = n11412 ^ n10958 ;
  assign n11396 = n10675 ^ x101 ;
  assign n11397 = n11396 ^ x100 ;
  assign n11398 = n11397 ^ n10941 ;
  assign n11399 = n11398 ^ n11396 ;
  assign n11402 = n11396 ^ n10953 ;
  assign n11403 = ~n11399 & ~n11402 ;
  assign n11404 = n11403 ^ n11396 ;
  assign n11405 = n11106 & ~n11404 ;
  assign n11406 = n11405 ^ n10671 ;
  assign n11389 = n10941 ^ x100 ;
  assign n11390 = n11106 & n11389 ;
  assign n11391 = n11390 ^ n10675 ;
  assign n11382 = n10934 ^ x99 ;
  assign n11383 = n11106 & n11382 ;
  assign n11384 = n11383 ^ n10937 ;
  assign n11375 = n10927 ^ x98 ;
  assign n11376 = n11106 & n11375 ;
  assign n11377 = n11376 ^ n10930 ;
  assign n11368 = n10920 ^ x97 ;
  assign n11369 = n11106 & n11368 ;
  assign n11370 = n11369 ^ n10923 ;
  assign n11361 = n10913 ^ x96 ;
  assign n11362 = n11106 & n11361 ;
  assign n11363 = n11362 ^ n10916 ;
  assign n11354 = n10906 ^ x95 ;
  assign n11355 = n11106 & n11354 ;
  assign n11356 = n11355 ^ n10909 ;
  assign n11347 = n10899 ^ x94 ;
  assign n11348 = n11106 & n11347 ;
  assign n11349 = n11348 ^ n10902 ;
  assign n11340 = n10892 ^ x93 ;
  assign n11341 = n11106 & n11340 ;
  assign n11342 = n11341 ^ n10895 ;
  assign n11333 = n10885 ^ x92 ;
  assign n11334 = n11106 & n11333 ;
  assign n11335 = n11334 ^ n10888 ;
  assign n11326 = n10878 ^ x91 ;
  assign n11327 = n11106 & n11326 ;
  assign n11328 = n11327 ^ n10881 ;
  assign n11319 = n10871 ^ x90 ;
  assign n11320 = n11106 & n11319 ;
  assign n11321 = n11320 ^ n10874 ;
  assign n11312 = n10864 ^ x89 ;
  assign n11313 = n11106 & n11312 ;
  assign n11314 = n11313 ^ n10867 ;
  assign n11305 = n10857 ^ x88 ;
  assign n11306 = n11106 & n11305 ;
  assign n11307 = n11306 ^ n10860 ;
  assign n11298 = n10850 ^ x87 ;
  assign n11299 = n11106 & n11298 ;
  assign n11300 = n11299 ^ n10853 ;
  assign n11291 = n10843 ^ x86 ;
  assign n11292 = n11106 & n11291 ;
  assign n11293 = n11292 ^ n10846 ;
  assign n11284 = n10836 ^ x85 ;
  assign n11285 = n11106 & n11284 ;
  assign n11286 = n11285 ^ n10839 ;
  assign n11277 = n10829 ^ x84 ;
  assign n11278 = n11106 & n11277 ;
  assign n11279 = n11278 ^ n10832 ;
  assign n11270 = n10822 ^ x83 ;
  assign n11271 = n11106 & n11270 ;
  assign n11272 = n11271 ^ n10825 ;
  assign n11263 = n10815 ^ x82 ;
  assign n11264 = n11106 & n11263 ;
  assign n11265 = n11264 ^ n10818 ;
  assign n11256 = n10808 ^ x81 ;
  assign n11257 = n11106 & n11256 ;
  assign n11258 = n11257 ^ n10811 ;
  assign n11249 = n10801 ^ x80 ;
  assign n11250 = n11106 & n11249 ;
  assign n11251 = n11250 ^ n10804 ;
  assign n11234 = n10685 ^ x79 ;
  assign n11235 = n11234 ^ n10795 ;
  assign n11236 = n11235 ^ x78 ;
  assign n11237 = n11236 ^ n11234 ;
  assign n11239 = n10795 ^ x79 ;
  assign n11240 = n11239 ^ n11234 ;
  assign n11241 = ~n11237 & ~n11240 ;
  assign n11242 = n11241 ^ n11234 ;
  assign n11243 = n11106 & ~n11242 ;
  assign n11244 = n11243 ^ n10681 ;
  assign n11227 = n10795 ^ x78 ;
  assign n11228 = n11106 & n11227 ;
  assign n11229 = n11228 ^ n10685 ;
  assign n11220 = n10792 ^ x77 ;
  assign n11221 = n11106 & n11220 ;
  assign n11222 = n11221 ^ n10699 ;
  assign n11116 = n10785 ^ x76 ;
  assign n11117 = n11106 & n11116 ;
  assign n11118 = n11117 ^ n10788 ;
  assign n11119 = n11118 ^ x77 ;
  assign n11124 = n11118 ^ x76 ;
  assign n11120 = n10778 ^ x75 ;
  assign n11121 = n11106 & n11120 ;
  assign n11122 = n11121 ^ n10781 ;
  assign n11123 = n11122 ^ n11118 ;
  assign n11125 = n11124 ^ n11123 ;
  assign n11207 = n10771 ^ x74 ;
  assign n11208 = n11106 & n11207 ;
  assign n11209 = n11208 ^ n10774 ;
  assign n11200 = n10768 ^ x73 ;
  assign n11201 = n11106 & n11200 ;
  assign n11202 = n11201 ^ n10703 ;
  assign n11193 = n10765 ^ x72 ;
  assign n11194 = n11106 & n11193 ;
  assign n11195 = n11194 ^ n10707 ;
  assign n11186 = n10758 ^ x71 ;
  assign n11187 = n11106 & n11186 ;
  assign n11188 = n11187 ^ n10761 ;
  assign n11179 = n10751 ^ x70 ;
  assign n11180 = n11106 & n11179 ;
  assign n11181 = n11180 ^ n10754 ;
  assign n11126 = n10738 ^ x68 ;
  assign n11127 = n11106 & n11126 ;
  assign n11128 = n11127 ^ n10740 ;
  assign n11129 = n11128 ^ x69 ;
  assign n11162 = n10731 ^ x67 ;
  assign n11163 = n11106 & n11162 ;
  assign n11164 = n11163 ^ n10734 ;
  assign n11155 = n10728 ^ x66 ;
  assign n11156 = n11106 & n11155 ;
  assign n11157 = n11156 ^ n10715 ;
  assign n11135 = x64 & n10662 ;
  assign n11131 = ~x11 & x64 ;
  assign n11132 = n11131 ^ x65 ;
  assign n11133 = n11106 & n11132 ;
  assign n11134 = n11133 ^ x12 ;
  assign n11136 = n11135 ^ n11134 ;
  assign n11137 = n11136 ^ x66 ;
  assign n11145 = x64 & n11106 ;
  assign n11146 = n11145 ^ x11 ;
  assign n11147 = ~x10 & x64 ;
  assign n11148 = n11147 ^ x65 ;
  assign n11141 = ~x10 & x65 ;
  assign n11142 = ~x64 & n11141 ;
  assign n11149 = n11148 ^ n11142 ;
  assign n11150 = ~n11146 & n11149 ;
  assign n11138 = ~x11 & n926 ;
  assign n11139 = x10 & n11138 ;
  assign n11140 = n11139 ^ n11138 ;
  assign n11143 = n11142 ^ n11140 ;
  assign n11144 = n11143 ^ n11141 ;
  assign n11151 = n11150 ^ n11144 ;
  assign n11152 = n11151 ^ n11136 ;
  assign n11153 = ~n11137 & n11152 ;
  assign n11154 = n11153 ^ x66 ;
  assign n11158 = n11157 ^ n11154 ;
  assign n11159 = n11157 ^ x67 ;
  assign n11160 = n11158 & ~n11159 ;
  assign n11161 = n11160 ^ x67 ;
  assign n11165 = n11164 ^ n11161 ;
  assign n11166 = n11164 ^ x68 ;
  assign n11167 = n11165 & ~n11166 ;
  assign n11168 = n11167 ^ x68 ;
  assign n11169 = n11168 ^ n11128 ;
  assign n11170 = ~n11129 & n11169 ;
  assign n11171 = n11170 ^ x69 ;
  assign n11172 = n11171 ^ x70 ;
  assign n11173 = n10744 ^ x69 ;
  assign n11174 = n11106 & n11173 ;
  assign n11175 = n11174 ^ n10747 ;
  assign n11176 = n11175 ^ n11171 ;
  assign n11177 = n11172 & n11176 ;
  assign n11178 = n11177 ^ x70 ;
  assign n11182 = n11181 ^ n11178 ;
  assign n11183 = n11181 ^ x71 ;
  assign n11184 = n11182 & ~n11183 ;
  assign n11185 = n11184 ^ x71 ;
  assign n11189 = n11188 ^ n11185 ;
  assign n11190 = n11188 ^ x72 ;
  assign n11191 = n11189 & ~n11190 ;
  assign n11192 = n11191 ^ x72 ;
  assign n11196 = n11195 ^ n11192 ;
  assign n11197 = n11195 ^ x73 ;
  assign n11198 = n11196 & ~n11197 ;
  assign n11199 = n11198 ^ x73 ;
  assign n11203 = n11202 ^ n11199 ;
  assign n11204 = n11202 ^ x74 ;
  assign n11205 = n11203 & ~n11204 ;
  assign n11206 = n11205 ^ x74 ;
  assign n11210 = n11209 ^ n11206 ;
  assign n11211 = n11209 ^ x75 ;
  assign n11212 = n11210 & ~n11211 ;
  assign n11213 = n11212 ^ x75 ;
  assign n11214 = n11213 ^ n11118 ;
  assign n11215 = n11214 ^ n11124 ;
  assign n11216 = ~n11125 & n11215 ;
  assign n11217 = n11216 ^ n11124 ;
  assign n11218 = ~n11119 & n11217 ;
  assign n11219 = n11218 ^ x77 ;
  assign n11223 = n11222 ^ n11219 ;
  assign n11224 = n11222 ^ x78 ;
  assign n11225 = n11223 & ~n11224 ;
  assign n11226 = n11225 ^ x78 ;
  assign n11230 = n11229 ^ n11226 ;
  assign n11231 = n11229 ^ x79 ;
  assign n11232 = n11230 & ~n11231 ;
  assign n11233 = n11232 ^ x79 ;
  assign n11245 = n11244 ^ n11233 ;
  assign n11246 = n11244 ^ x80 ;
  assign n11247 = n11245 & ~n11246 ;
  assign n11248 = n11247 ^ x80 ;
  assign n11252 = n11251 ^ n11248 ;
  assign n11253 = n11251 ^ x81 ;
  assign n11254 = n11252 & ~n11253 ;
  assign n11255 = n11254 ^ x81 ;
  assign n11259 = n11258 ^ n11255 ;
  assign n11260 = n11258 ^ x82 ;
  assign n11261 = n11259 & ~n11260 ;
  assign n11262 = n11261 ^ x82 ;
  assign n11266 = n11265 ^ n11262 ;
  assign n11267 = n11265 ^ x83 ;
  assign n11268 = n11266 & ~n11267 ;
  assign n11269 = n11268 ^ x83 ;
  assign n11273 = n11272 ^ n11269 ;
  assign n11274 = n11272 ^ x84 ;
  assign n11275 = n11273 & ~n11274 ;
  assign n11276 = n11275 ^ x84 ;
  assign n11280 = n11279 ^ n11276 ;
  assign n11281 = n11279 ^ x85 ;
  assign n11282 = n11280 & ~n11281 ;
  assign n11283 = n11282 ^ x85 ;
  assign n11287 = n11286 ^ n11283 ;
  assign n11288 = n11286 ^ x86 ;
  assign n11289 = n11287 & ~n11288 ;
  assign n11290 = n11289 ^ x86 ;
  assign n11294 = n11293 ^ n11290 ;
  assign n11295 = n11293 ^ x87 ;
  assign n11296 = n11294 & ~n11295 ;
  assign n11297 = n11296 ^ x87 ;
  assign n11301 = n11300 ^ n11297 ;
  assign n11302 = n11300 ^ x88 ;
  assign n11303 = n11301 & ~n11302 ;
  assign n11304 = n11303 ^ x88 ;
  assign n11308 = n11307 ^ n11304 ;
  assign n11309 = n11307 ^ x89 ;
  assign n11310 = n11308 & ~n11309 ;
  assign n11311 = n11310 ^ x89 ;
  assign n11315 = n11314 ^ n11311 ;
  assign n11316 = n11314 ^ x90 ;
  assign n11317 = n11315 & ~n11316 ;
  assign n11318 = n11317 ^ x90 ;
  assign n11322 = n11321 ^ n11318 ;
  assign n11323 = n11321 ^ x91 ;
  assign n11324 = n11322 & ~n11323 ;
  assign n11325 = n11324 ^ x91 ;
  assign n11329 = n11328 ^ n11325 ;
  assign n11330 = n11328 ^ x92 ;
  assign n11331 = n11329 & ~n11330 ;
  assign n11332 = n11331 ^ x92 ;
  assign n11336 = n11335 ^ n11332 ;
  assign n11337 = n11335 ^ x93 ;
  assign n11338 = n11336 & ~n11337 ;
  assign n11339 = n11338 ^ x93 ;
  assign n11343 = n11342 ^ n11339 ;
  assign n11344 = n11342 ^ x94 ;
  assign n11345 = n11343 & ~n11344 ;
  assign n11346 = n11345 ^ x94 ;
  assign n11350 = n11349 ^ n11346 ;
  assign n11351 = n11349 ^ x95 ;
  assign n11352 = n11350 & ~n11351 ;
  assign n11353 = n11352 ^ x95 ;
  assign n11357 = n11356 ^ n11353 ;
  assign n11358 = n11356 ^ x96 ;
  assign n11359 = n11357 & ~n11358 ;
  assign n11360 = n11359 ^ x96 ;
  assign n11364 = n11363 ^ n11360 ;
  assign n11365 = n11363 ^ x97 ;
  assign n11366 = n11364 & ~n11365 ;
  assign n11367 = n11366 ^ x97 ;
  assign n11371 = n11370 ^ n11367 ;
  assign n11372 = n11370 ^ x98 ;
  assign n11373 = n11371 & ~n11372 ;
  assign n11374 = n11373 ^ x98 ;
  assign n11378 = n11377 ^ n11374 ;
  assign n11379 = n11377 ^ x99 ;
  assign n11380 = n11378 & ~n11379 ;
  assign n11381 = n11380 ^ x99 ;
  assign n11385 = n11384 ^ n11381 ;
  assign n11386 = n11384 ^ x100 ;
  assign n11387 = n11385 & ~n11386 ;
  assign n11388 = n11387 ^ x100 ;
  assign n11392 = n11391 ^ n11388 ;
  assign n11393 = n11391 ^ x101 ;
  assign n11394 = n11392 & ~n11393 ;
  assign n11395 = n11394 ^ x101 ;
  assign n11407 = n11406 ^ n11395 ;
  assign n11408 = n11406 ^ x102 ;
  assign n11409 = n11407 & ~n11408 ;
  assign n11410 = n11409 ^ x102 ;
  assign n11414 = n11413 ^ n11410 ;
  assign n11415 = n11413 ^ x103 ;
  assign n11416 = n11414 & ~n11415 ;
  assign n11417 = n11416 ^ x103 ;
  assign n11421 = n11420 ^ n11417 ;
  assign n11422 = n11420 ^ x104 ;
  assign n11423 = n11421 & ~n11422 ;
  assign n11424 = n11423 ^ x104 ;
  assign n11428 = n11427 ^ n11424 ;
  assign n11429 = n11427 ^ x105 ;
  assign n11430 = n11428 & ~n11429 ;
  assign n11431 = n11430 ^ x105 ;
  assign n11435 = n11434 ^ n11431 ;
  assign n11436 = n11434 ^ x106 ;
  assign n11437 = n11435 & ~n11436 ;
  assign n11438 = n11437 ^ x106 ;
  assign n11442 = n11441 ^ n11438 ;
  assign n11443 = n11441 ^ x107 ;
  assign n11444 = n11442 & ~n11443 ;
  assign n11445 = n11444 ^ x107 ;
  assign n11449 = n11448 ^ n11445 ;
  assign n11450 = n11448 ^ x108 ;
  assign n11451 = n11449 & ~n11450 ;
  assign n11452 = n11451 ^ x108 ;
  assign n11456 = n11455 ^ n11452 ;
  assign n11457 = n11455 ^ x109 ;
  assign n11458 = n11456 & ~n11457 ;
  assign n11459 = n11458 ^ x109 ;
  assign n11463 = n11462 ^ n11459 ;
  assign n11464 = n11462 ^ x110 ;
  assign n11465 = n11463 & ~n11464 ;
  assign n11466 = n11465 ^ x110 ;
  assign n11470 = n11469 ^ n11466 ;
  assign n11471 = n11469 ^ x111 ;
  assign n11472 = n11470 & ~n11471 ;
  assign n11473 = n11472 ^ x111 ;
  assign n11474 = n11473 ^ n11108 ;
  assign n11475 = n11474 ^ n11114 ;
  assign n11476 = ~n11115 & n11475 ;
  assign n11477 = n11476 ^ n11114 ;
  assign n11478 = ~n11109 & n11477 ;
  assign n11479 = n11478 ^ x113 ;
  assign n11483 = n11482 ^ n11479 ;
  assign n11484 = n11482 ^ x114 ;
  assign n11485 = n11483 & ~n11484 ;
  assign n11486 = n11485 ^ x114 ;
  assign n11490 = n11489 ^ n11486 ;
  assign n11491 = n11489 ^ x115 ;
  assign n11492 = n11490 & ~n11491 ;
  assign n11493 = n11492 ^ x115 ;
  assign n11497 = n11496 ^ n11493 ;
  assign n11940 = n11493 ^ x116 ;
  assign n11501 = n11497 & n11940 ;
  assign n11498 = x117 ^ x116 ;
  assign n11502 = n11501 ^ n11498 ;
  assign n11048 = ~n10666 & ~n11047 ;
  assign n11049 = n11048 ^ x116 ;
  assign n11050 = n139 & ~n11049 ;
  assign n11064 = n11050 & n11059 ;
  assign n11065 = ~n11048 & n11064 ;
  assign n11066 = n11065 ^ n11048 ;
  assign n11051 = n11050 ^ n139 ;
  assign n11052 = n11051 ^ n11048 ;
  assign n11067 = n11066 ^ n11052 ;
  assign n11068 = n10265 & ~n11067 ;
  assign n11503 = n11068 ^ x117 ;
  assign n11506 = n11502 & ~n11503 ;
  assign n11507 = n11506 ^ x117 ;
  assign n11508 = n138 & ~n11507 ;
  assign n11509 = n11502 & n11508 ;
  assign n11510 = n11509 ^ n11068 ;
  assign n11511 = n137 & n11510 ;
  assign n11941 = n11508 & n11940 ;
  assign n11942 = n11941 ^ n11496 ;
  assign n11512 = n11486 ^ x115 ;
  assign n11513 = n11508 & n11512 ;
  assign n11514 = n11513 ^ n11489 ;
  assign n11515 = n11514 ^ x116 ;
  assign n11520 = n11514 ^ x115 ;
  assign n11516 = n11479 ^ x114 ;
  assign n11517 = n11508 & n11516 ;
  assign n11518 = n11517 ^ n11482 ;
  assign n11519 = n11518 ^ n11514 ;
  assign n11521 = n11520 ^ n11519 ;
  assign n11522 = n11112 ^ x113 ;
  assign n11523 = n11522 ^ n11473 ;
  assign n11524 = n11523 ^ x112 ;
  assign n11525 = n11524 ^ n11522 ;
  assign n11527 = n11473 ^ x113 ;
  assign n11528 = n11527 ^ n11522 ;
  assign n11529 = ~n11525 & ~n11528 ;
  assign n11530 = n11529 ^ n11522 ;
  assign n11531 = n11508 & ~n11530 ;
  assign n11532 = n11531 ^ n11108 ;
  assign n11533 = n11532 ^ x114 ;
  assign n11538 = n11532 ^ x113 ;
  assign n11534 = n11473 ^ x112 ;
  assign n11535 = n11508 & n11534 ;
  assign n11536 = n11535 ^ n11112 ;
  assign n11537 = n11536 ^ n11532 ;
  assign n11539 = n11538 ^ n11537 ;
  assign n11921 = n11466 ^ x111 ;
  assign n11922 = n11508 & n11921 ;
  assign n11923 = n11922 ^ n11469 ;
  assign n11914 = n11459 ^ x110 ;
  assign n11915 = n11508 & n11914 ;
  assign n11916 = n11915 ^ n11462 ;
  assign n11907 = n11452 ^ x109 ;
  assign n11908 = n11508 & n11907 ;
  assign n11909 = n11908 ^ n11455 ;
  assign n11900 = n11445 ^ x108 ;
  assign n11901 = n11508 & n11900 ;
  assign n11902 = n11901 ^ n11448 ;
  assign n11540 = n11438 ^ x107 ;
  assign n11541 = n11508 & n11540 ;
  assign n11542 = n11541 ^ n11441 ;
  assign n11543 = n11542 ^ x108 ;
  assign n11548 = n11542 ^ x107 ;
  assign n11544 = n11431 ^ x106 ;
  assign n11545 = n11508 & n11544 ;
  assign n11546 = n11545 ^ n11434 ;
  assign n11547 = n11546 ^ n11542 ;
  assign n11549 = n11548 ^ n11547 ;
  assign n11887 = n11424 ^ x105 ;
  assign n11888 = n11508 & n11887 ;
  assign n11889 = n11888 ^ n11427 ;
  assign n11880 = n11417 ^ x104 ;
  assign n11881 = n11508 & n11880 ;
  assign n11882 = n11881 ^ n11420 ;
  assign n11873 = n11410 ^ x103 ;
  assign n11874 = n11508 & n11873 ;
  assign n11875 = n11874 ^ n11413 ;
  assign n11866 = n11395 ^ x102 ;
  assign n11867 = n11508 & n11866 ;
  assign n11868 = n11867 ^ n11406 ;
  assign n11859 = n11388 ^ x101 ;
  assign n11860 = n11508 & n11859 ;
  assign n11861 = n11860 ^ n11391 ;
  assign n11852 = n11381 ^ x100 ;
  assign n11853 = n11508 & n11852 ;
  assign n11854 = n11853 ^ n11384 ;
  assign n11845 = n11374 ^ x99 ;
  assign n11846 = n11508 & n11845 ;
  assign n11847 = n11846 ^ n11377 ;
  assign n11838 = n11367 ^ x98 ;
  assign n11839 = n11508 & n11838 ;
  assign n11840 = n11839 ^ n11370 ;
  assign n11831 = n11360 ^ x97 ;
  assign n11832 = n11508 & n11831 ;
  assign n11833 = n11832 ^ n11363 ;
  assign n11824 = n11353 ^ x96 ;
  assign n11825 = n11508 & n11824 ;
  assign n11826 = n11825 ^ n11356 ;
  assign n11817 = n11346 ^ x95 ;
  assign n11818 = n11508 & n11817 ;
  assign n11819 = n11818 ^ n11349 ;
  assign n11810 = n11339 ^ x94 ;
  assign n11811 = n11508 & n11810 ;
  assign n11812 = n11811 ^ n11342 ;
  assign n11803 = n11332 ^ x93 ;
  assign n11804 = n11508 & n11803 ;
  assign n11805 = n11804 ^ n11335 ;
  assign n11796 = n11325 ^ x92 ;
  assign n11797 = n11508 & n11796 ;
  assign n11798 = n11797 ^ n11328 ;
  assign n11789 = n11318 ^ x91 ;
  assign n11790 = n11508 & n11789 ;
  assign n11791 = n11790 ^ n11321 ;
  assign n11782 = n11311 ^ x90 ;
  assign n11783 = n11508 & n11782 ;
  assign n11784 = n11783 ^ n11314 ;
  assign n11775 = n11304 ^ x89 ;
  assign n11776 = n11508 & n11775 ;
  assign n11777 = n11776 ^ n11307 ;
  assign n11768 = n11297 ^ x88 ;
  assign n11769 = n11508 & n11768 ;
  assign n11770 = n11769 ^ n11300 ;
  assign n11761 = n11290 ^ x87 ;
  assign n11762 = n11508 & n11761 ;
  assign n11763 = n11762 ^ n11293 ;
  assign n11754 = n11283 ^ x86 ;
  assign n11755 = n11508 & n11754 ;
  assign n11756 = n11755 ^ n11286 ;
  assign n11747 = n11276 ^ x85 ;
  assign n11748 = n11508 & n11747 ;
  assign n11749 = n11748 ^ n11279 ;
  assign n11740 = n11269 ^ x84 ;
  assign n11741 = n11508 & n11740 ;
  assign n11742 = n11741 ^ n11272 ;
  assign n11733 = n11262 ^ x83 ;
  assign n11734 = n11508 & n11733 ;
  assign n11735 = n11734 ^ n11265 ;
  assign n11726 = n11255 ^ x82 ;
  assign n11727 = n11508 & n11726 ;
  assign n11728 = n11727 ^ n11258 ;
  assign n11719 = n11248 ^ x81 ;
  assign n11720 = n11508 & n11719 ;
  assign n11721 = n11720 ^ n11251 ;
  assign n11712 = n11233 ^ x80 ;
  assign n11713 = n11508 & n11712 ;
  assign n11714 = n11713 ^ n11244 ;
  assign n11705 = n11226 ^ x79 ;
  assign n11706 = n11508 & n11705 ;
  assign n11707 = n11706 ^ n11229 ;
  assign n11698 = n11219 ^ x78 ;
  assign n11699 = n11508 & n11698 ;
  assign n11700 = n11699 ^ n11222 ;
  assign n11683 = n11122 ^ x77 ;
  assign n11684 = n11683 ^ n11213 ;
  assign n11685 = n11684 ^ x76 ;
  assign n11686 = n11685 ^ n11683 ;
  assign n11687 = n11683 ^ n11122 ;
  assign n11688 = n11687 ^ n11213 ;
  assign n11689 = n11688 ^ n11683 ;
  assign n11690 = ~n11686 & ~n11689 ;
  assign n11691 = n11690 ^ n11683 ;
  assign n11692 = n11508 & ~n11691 ;
  assign n11693 = n11692 ^ n11118 ;
  assign n11676 = n11213 ^ x76 ;
  assign n11677 = n11508 & n11676 ;
  assign n11678 = n11677 ^ n11122 ;
  assign n11669 = n11206 ^ x75 ;
  assign n11670 = n11508 & n11669 ;
  assign n11671 = n11670 ^ n11209 ;
  assign n11662 = n11199 ^ x74 ;
  assign n11663 = n11508 & n11662 ;
  assign n11664 = n11663 ^ n11202 ;
  assign n11655 = n11192 ^ x73 ;
  assign n11656 = n11508 & n11655 ;
  assign n11657 = n11656 ^ n11195 ;
  assign n11648 = n11185 ^ x72 ;
  assign n11649 = n11508 & n11648 ;
  assign n11650 = n11649 ^ n11188 ;
  assign n11641 = n11178 ^ x71 ;
  assign n11642 = n11508 & n11641 ;
  assign n11643 = n11642 ^ n11181 ;
  assign n11550 = n11172 & n11508 ;
  assign n11551 = n11550 ^ n11175 ;
  assign n11552 = n11551 ^ x71 ;
  assign n11557 = n11551 ^ x70 ;
  assign n11553 = n11168 ^ x69 ;
  assign n11554 = n11508 & n11553 ;
  assign n11555 = n11554 ^ n11128 ;
  assign n11556 = n11555 ^ n11551 ;
  assign n11558 = n11557 ^ n11556 ;
  assign n11628 = n11161 ^ x68 ;
  assign n11629 = n11508 & n11628 ;
  assign n11630 = n11629 ^ n11164 ;
  assign n11621 = n11154 ^ x67 ;
  assign n11622 = n11508 & n11621 ;
  assign n11623 = n11622 ^ n11157 ;
  assign n11614 = n11151 ^ x66 ;
  assign n11615 = n11508 & n11614 ;
  assign n11616 = n11615 ^ n11136 ;
  assign n11559 = n11142 ^ n11141 ;
  assign n11560 = n11559 ^ n11148 ;
  assign n11561 = ~x9 & x64 ;
  assign n11562 = ~n11560 & ~n11561 ;
  assign n11564 = n11561 ^ n11560 ;
  assign n11565 = n11564 ^ n11562 ;
  assign n11566 = ~n11141 & n11565 ;
  assign n11571 = n11146 & n11566 ;
  assign n11572 = n11571 ^ n11139 ;
  assign n11563 = n11146 ^ x65 ;
  assign n11568 = n11565 ^ n11141 ;
  assign n11567 = n11566 ^ n11147 ;
  assign n11569 = n11568 ^ n11567 ;
  assign n11570 = ~n11563 & n11569 ;
  assign n11573 = n11572 ^ n11570 ;
  assign n11574 = ~n11562 & n11573 ;
  assign n11575 = n11508 & n11574 ;
  assign n11576 = n11575 ^ n11571 ;
  assign n11588 = x65 ^ x9 ;
  assign n11579 = n11146 ^ x9 ;
  assign n11589 = n11588 ^ n11579 ;
  assign n11590 = n11589 ^ x10 ;
  assign n11591 = n11590 ^ n11508 ;
  assign n11592 = n11591 ^ x9 ;
  assign n11577 = x65 ^ x10 ;
  assign n11578 = n11577 ^ n11508 ;
  assign n11580 = n11579 ^ n11146 ;
  assign n11581 = n11580 ^ n11508 ;
  assign n11582 = n11581 ^ n11579 ;
  assign n11585 = x65 & ~n11582 ;
  assign n11586 = n11585 ^ n11579 ;
  assign n11587 = n11578 & n11586 ;
  assign n11593 = n11592 ^ n11587 ;
  assign n11594 = ~x66 & n11141 ;
  assign n11595 = x64 & n11508 ;
  assign n11596 = n11508 ^ n11146 ;
  assign n11597 = ~n11595 & ~n11596 ;
  assign n11598 = n11594 & n11597 ;
  assign n11599 = n11598 ^ x66 ;
  assign n11600 = x64 & ~n11599 ;
  assign n11601 = ~n11593 & n11600 ;
  assign n11602 = n11601 ^ n11599 ;
  assign n11605 = n11602 ^ n11587 ;
  assign n11606 = n11605 ^ n11602 ;
  assign n11609 = n11601 & ~n11606 ;
  assign n11610 = n11591 & n11609 ;
  assign n11611 = n11610 ^ n11591 ;
  assign n11603 = n11602 ^ n11591 ;
  assign n11612 = n11611 ^ n11603 ;
  assign n11613 = ~n11576 & n11612 ;
  assign n11617 = n11616 ^ n11613 ;
  assign n11618 = n11616 ^ x67 ;
  assign n11619 = n11617 & ~n11618 ;
  assign n11620 = n11619 ^ x67 ;
  assign n11624 = n11623 ^ n11620 ;
  assign n11625 = n11623 ^ x68 ;
  assign n11626 = n11624 & ~n11625 ;
  assign n11627 = n11626 ^ x68 ;
  assign n11631 = n11630 ^ n11627 ;
  assign n11632 = n11630 ^ x69 ;
  assign n11633 = n11631 & ~n11632 ;
  assign n11634 = n11633 ^ x69 ;
  assign n11635 = n11634 ^ n11551 ;
  assign n11636 = n11635 ^ n11557 ;
  assign n11637 = ~n11558 & n11636 ;
  assign n11638 = n11637 ^ n11557 ;
  assign n11639 = ~n11552 & n11638 ;
  assign n11640 = n11639 ^ x71 ;
  assign n11644 = n11643 ^ n11640 ;
  assign n11645 = n11643 ^ x72 ;
  assign n11646 = n11644 & ~n11645 ;
  assign n11647 = n11646 ^ x72 ;
  assign n11651 = n11650 ^ n11647 ;
  assign n11652 = n11650 ^ x73 ;
  assign n11653 = n11651 & ~n11652 ;
  assign n11654 = n11653 ^ x73 ;
  assign n11658 = n11657 ^ n11654 ;
  assign n11659 = n11657 ^ x74 ;
  assign n11660 = n11658 & ~n11659 ;
  assign n11661 = n11660 ^ x74 ;
  assign n11665 = n11664 ^ n11661 ;
  assign n11666 = n11664 ^ x75 ;
  assign n11667 = n11665 & ~n11666 ;
  assign n11668 = n11667 ^ x75 ;
  assign n11672 = n11671 ^ n11668 ;
  assign n11673 = n11671 ^ x76 ;
  assign n11674 = n11672 & ~n11673 ;
  assign n11675 = n11674 ^ x76 ;
  assign n11679 = n11678 ^ n11675 ;
  assign n11680 = n11678 ^ x77 ;
  assign n11681 = n11679 & ~n11680 ;
  assign n11682 = n11681 ^ x77 ;
  assign n11694 = n11693 ^ n11682 ;
  assign n11695 = n11693 ^ x78 ;
  assign n11696 = n11694 & ~n11695 ;
  assign n11697 = n11696 ^ x78 ;
  assign n11701 = n11700 ^ n11697 ;
  assign n11702 = n11700 ^ x79 ;
  assign n11703 = n11701 & ~n11702 ;
  assign n11704 = n11703 ^ x79 ;
  assign n11708 = n11707 ^ n11704 ;
  assign n11709 = n11707 ^ x80 ;
  assign n11710 = n11708 & ~n11709 ;
  assign n11711 = n11710 ^ x80 ;
  assign n11715 = n11714 ^ n11711 ;
  assign n11716 = n11714 ^ x81 ;
  assign n11717 = n11715 & ~n11716 ;
  assign n11718 = n11717 ^ x81 ;
  assign n11722 = n11721 ^ n11718 ;
  assign n11723 = n11721 ^ x82 ;
  assign n11724 = n11722 & ~n11723 ;
  assign n11725 = n11724 ^ x82 ;
  assign n11729 = n11728 ^ n11725 ;
  assign n11730 = n11728 ^ x83 ;
  assign n11731 = n11729 & ~n11730 ;
  assign n11732 = n11731 ^ x83 ;
  assign n11736 = n11735 ^ n11732 ;
  assign n11737 = n11735 ^ x84 ;
  assign n11738 = n11736 & ~n11737 ;
  assign n11739 = n11738 ^ x84 ;
  assign n11743 = n11742 ^ n11739 ;
  assign n11744 = n11742 ^ x85 ;
  assign n11745 = n11743 & ~n11744 ;
  assign n11746 = n11745 ^ x85 ;
  assign n11750 = n11749 ^ n11746 ;
  assign n11751 = n11749 ^ x86 ;
  assign n11752 = n11750 & ~n11751 ;
  assign n11753 = n11752 ^ x86 ;
  assign n11757 = n11756 ^ n11753 ;
  assign n11758 = n11756 ^ x87 ;
  assign n11759 = n11757 & ~n11758 ;
  assign n11760 = n11759 ^ x87 ;
  assign n11764 = n11763 ^ n11760 ;
  assign n11765 = n11763 ^ x88 ;
  assign n11766 = n11764 & ~n11765 ;
  assign n11767 = n11766 ^ x88 ;
  assign n11771 = n11770 ^ n11767 ;
  assign n11772 = n11770 ^ x89 ;
  assign n11773 = n11771 & ~n11772 ;
  assign n11774 = n11773 ^ x89 ;
  assign n11778 = n11777 ^ n11774 ;
  assign n11779 = n11777 ^ x90 ;
  assign n11780 = n11778 & ~n11779 ;
  assign n11781 = n11780 ^ x90 ;
  assign n11785 = n11784 ^ n11781 ;
  assign n11786 = n11784 ^ x91 ;
  assign n11787 = n11785 & ~n11786 ;
  assign n11788 = n11787 ^ x91 ;
  assign n11792 = n11791 ^ n11788 ;
  assign n11793 = n11791 ^ x92 ;
  assign n11794 = n11792 & ~n11793 ;
  assign n11795 = n11794 ^ x92 ;
  assign n11799 = n11798 ^ n11795 ;
  assign n11800 = n11798 ^ x93 ;
  assign n11801 = n11799 & ~n11800 ;
  assign n11802 = n11801 ^ x93 ;
  assign n11806 = n11805 ^ n11802 ;
  assign n11807 = n11805 ^ x94 ;
  assign n11808 = n11806 & ~n11807 ;
  assign n11809 = n11808 ^ x94 ;
  assign n11813 = n11812 ^ n11809 ;
  assign n11814 = n11812 ^ x95 ;
  assign n11815 = n11813 & ~n11814 ;
  assign n11816 = n11815 ^ x95 ;
  assign n11820 = n11819 ^ n11816 ;
  assign n11821 = n11819 ^ x96 ;
  assign n11822 = n11820 & ~n11821 ;
  assign n11823 = n11822 ^ x96 ;
  assign n11827 = n11826 ^ n11823 ;
  assign n11828 = n11826 ^ x97 ;
  assign n11829 = n11827 & ~n11828 ;
  assign n11830 = n11829 ^ x97 ;
  assign n11834 = n11833 ^ n11830 ;
  assign n11835 = n11833 ^ x98 ;
  assign n11836 = n11834 & ~n11835 ;
  assign n11837 = n11836 ^ x98 ;
  assign n11841 = n11840 ^ n11837 ;
  assign n11842 = n11840 ^ x99 ;
  assign n11843 = n11841 & ~n11842 ;
  assign n11844 = n11843 ^ x99 ;
  assign n11848 = n11847 ^ n11844 ;
  assign n11849 = n11847 ^ x100 ;
  assign n11850 = n11848 & ~n11849 ;
  assign n11851 = n11850 ^ x100 ;
  assign n11855 = n11854 ^ n11851 ;
  assign n11856 = n11854 ^ x101 ;
  assign n11857 = n11855 & ~n11856 ;
  assign n11858 = n11857 ^ x101 ;
  assign n11862 = n11861 ^ n11858 ;
  assign n11863 = n11861 ^ x102 ;
  assign n11864 = n11862 & ~n11863 ;
  assign n11865 = n11864 ^ x102 ;
  assign n11869 = n11868 ^ n11865 ;
  assign n11870 = n11868 ^ x103 ;
  assign n11871 = n11869 & ~n11870 ;
  assign n11872 = n11871 ^ x103 ;
  assign n11876 = n11875 ^ n11872 ;
  assign n11877 = n11875 ^ x104 ;
  assign n11878 = n11876 & ~n11877 ;
  assign n11879 = n11878 ^ x104 ;
  assign n11883 = n11882 ^ n11879 ;
  assign n11884 = n11882 ^ x105 ;
  assign n11885 = n11883 & ~n11884 ;
  assign n11886 = n11885 ^ x105 ;
  assign n11890 = n11889 ^ n11886 ;
  assign n11891 = n11889 ^ x106 ;
  assign n11892 = n11890 & ~n11891 ;
  assign n11893 = n11892 ^ x106 ;
  assign n11894 = n11893 ^ n11542 ;
  assign n11895 = n11894 ^ n11548 ;
  assign n11896 = ~n11549 & n11895 ;
  assign n11897 = n11896 ^ n11548 ;
  assign n11898 = ~n11543 & n11897 ;
  assign n11899 = n11898 ^ x108 ;
  assign n11903 = n11902 ^ n11899 ;
  assign n11904 = n11902 ^ x109 ;
  assign n11905 = n11903 & ~n11904 ;
  assign n11906 = n11905 ^ x109 ;
  assign n11910 = n11909 ^ n11906 ;
  assign n11911 = n11909 ^ x110 ;
  assign n11912 = n11910 & ~n11911 ;
  assign n11913 = n11912 ^ x110 ;
  assign n11917 = n11916 ^ n11913 ;
  assign n11918 = n11916 ^ x111 ;
  assign n11919 = n11917 & ~n11918 ;
  assign n11920 = n11919 ^ x111 ;
  assign n11924 = n11923 ^ n11920 ;
  assign n11925 = n11923 ^ x112 ;
  assign n11926 = n11924 & ~n11925 ;
  assign n11927 = n11926 ^ x112 ;
  assign n11928 = n11927 ^ n11532 ;
  assign n11929 = n11928 ^ n11538 ;
  assign n11930 = ~n11539 & n11929 ;
  assign n11931 = n11930 ^ n11538 ;
  assign n11932 = ~n11533 & n11931 ;
  assign n11933 = n11932 ^ x114 ;
  assign n11934 = n11933 ^ n11514 ;
  assign n11935 = n11934 ^ n11520 ;
  assign n11936 = ~n11521 & n11935 ;
  assign n11937 = n11936 ^ n11520 ;
  assign n11938 = ~n11515 & n11937 ;
  assign n11939 = n11938 ^ x116 ;
  assign n11943 = n11942 ^ n11939 ;
  assign n12382 = n11939 ^ x117 ;
  assign n11947 = n11943 & n12382 ;
  assign n11944 = x118 ^ x117 ;
  assign n11948 = n11947 ^ n11944 ;
  assign n11949 = n11511 & n11948 ;
  assign n11950 = n11949 ^ n11510 ;
  assign n11951 = n11950 ^ n11068 ;
  assign n11952 = ~x119 & ~n11951 ;
  assign n11953 = n11952 ^ n11068 ;
  assign n11956 = x118 & ~n11510 ;
  assign n11957 = n137 & ~n11956 ;
  assign n11958 = n11510 ^ x118 ;
  assign n11959 = n11958 ^ n11956 ;
  assign n11960 = ~n11942 & ~n11959 ;
  assign n11961 = x117 & n11960 ;
  assign n11962 = n11957 & ~n11961 ;
  assign n11967 = x117 & x118 ;
  assign n11968 = n11967 ^ n11960 ;
  assign n11969 = n11939 & n11968 ;
  assign n11970 = n11962 & ~n11969 ;
  assign n12383 = n11970 & n12382 ;
  assign n12384 = n12383 ^ n11942 ;
  assign n12386 = n12384 ^ x117 ;
  assign n11955 = x117 & ~n11510 ;
  assign n11971 = n11939 & n11970 ;
  assign n11972 = n11955 & n11971 ;
  assign n11973 = n11972 ^ n11970 ;
  assign n12375 = n11933 ^ x115 ;
  assign n12376 = n11973 & n12375 ;
  assign n12377 = n12376 ^ n11518 ;
  assign n12360 = n11536 ^ x114 ;
  assign n12361 = n12360 ^ x113 ;
  assign n12362 = n12361 ^ n11927 ;
  assign n12363 = n12362 ^ n12360 ;
  assign n12366 = n12360 ^ n10259 ;
  assign n12367 = ~n12363 & ~n12366 ;
  assign n12368 = n12367 ^ n12360 ;
  assign n12369 = n11973 & ~n12368 ;
  assign n12370 = n12369 ^ n11532 ;
  assign n12353 = n11927 ^ x113 ;
  assign n12354 = n11973 & n12353 ;
  assign n12355 = n12354 ^ n11536 ;
  assign n12346 = n11920 ^ x112 ;
  assign n12347 = n11973 & n12346 ;
  assign n12348 = n12347 ^ n11923 ;
  assign n12339 = n11913 ^ x111 ;
  assign n12340 = n11973 & n12339 ;
  assign n12341 = n12340 ^ n11916 ;
  assign n12332 = n11906 ^ x110 ;
  assign n12333 = n11973 & n12332 ;
  assign n12334 = n12333 ^ n11909 ;
  assign n12325 = n11899 ^ x109 ;
  assign n12326 = n11973 & n12325 ;
  assign n12327 = n12326 ^ n11902 ;
  assign n12310 = n11546 ^ x108 ;
  assign n12311 = n12310 ^ x107 ;
  assign n12312 = n12311 ^ n11893 ;
  assign n12313 = n12312 ^ n12310 ;
  assign n12315 = x108 ^ x107 ;
  assign n12316 = n12315 ^ n12310 ;
  assign n12317 = ~n12313 & ~n12316 ;
  assign n12318 = n12317 ^ n12310 ;
  assign n12319 = n11973 & ~n12318 ;
  assign n12320 = n12319 ^ n11542 ;
  assign n12303 = n11893 ^ x107 ;
  assign n12304 = n11973 & n12303 ;
  assign n12305 = n12304 ^ n11546 ;
  assign n12296 = n11886 ^ x106 ;
  assign n12297 = n11973 & n12296 ;
  assign n12298 = n12297 ^ n11889 ;
  assign n12289 = n11879 ^ x105 ;
  assign n12290 = n11973 & n12289 ;
  assign n12291 = n12290 ^ n11882 ;
  assign n12282 = n11872 ^ x104 ;
  assign n12283 = n11973 & n12282 ;
  assign n12284 = n12283 ^ n11875 ;
  assign n12275 = n11865 ^ x103 ;
  assign n12276 = n11973 & n12275 ;
  assign n12277 = n12276 ^ n11868 ;
  assign n12268 = n11858 ^ x102 ;
  assign n12269 = n11973 & n12268 ;
  assign n12270 = n12269 ^ n11861 ;
  assign n12261 = n11851 ^ x101 ;
  assign n12262 = n11973 & n12261 ;
  assign n12263 = n12262 ^ n11854 ;
  assign n12254 = n11844 ^ x100 ;
  assign n12255 = n11973 & n12254 ;
  assign n12256 = n12255 ^ n11847 ;
  assign n12247 = n11837 ^ x99 ;
  assign n12248 = n11973 & n12247 ;
  assign n12249 = n12248 ^ n11840 ;
  assign n12240 = n11830 ^ x98 ;
  assign n12241 = n11973 & n12240 ;
  assign n12242 = n12241 ^ n11833 ;
  assign n12233 = n11823 ^ x97 ;
  assign n12234 = n11973 & n12233 ;
  assign n12235 = n12234 ^ n11826 ;
  assign n12226 = n11816 ^ x96 ;
  assign n12227 = n11973 & n12226 ;
  assign n12228 = n12227 ^ n11819 ;
  assign n12219 = n11809 ^ x95 ;
  assign n12220 = n11973 & n12219 ;
  assign n12221 = n12220 ^ n11812 ;
  assign n12212 = n11802 ^ x94 ;
  assign n12213 = n11973 & n12212 ;
  assign n12214 = n12213 ^ n11805 ;
  assign n11954 = n11795 ^ x93 ;
  assign n11974 = n11954 & n11973 ;
  assign n11975 = n11974 ^ n11798 ;
  assign n11976 = n11975 ^ x94 ;
  assign n11981 = n11975 ^ x93 ;
  assign n11977 = n11788 ^ x92 ;
  assign n11978 = n11973 & n11977 ;
  assign n11979 = n11978 ^ n11791 ;
  assign n11980 = n11979 ^ n11975 ;
  assign n11982 = n11981 ^ n11980 ;
  assign n12199 = n11781 ^ x91 ;
  assign n12200 = n11973 & n12199 ;
  assign n12201 = n12200 ^ n11784 ;
  assign n12192 = n11774 ^ x90 ;
  assign n12193 = n11973 & n12192 ;
  assign n12194 = n12193 ^ n11777 ;
  assign n12185 = n11767 ^ x89 ;
  assign n12186 = n11973 & n12185 ;
  assign n12187 = n12186 ^ n11770 ;
  assign n12178 = n11760 ^ x88 ;
  assign n12179 = n11973 & n12178 ;
  assign n12180 = n12179 ^ n11763 ;
  assign n12171 = n11753 ^ x87 ;
  assign n12172 = n11973 & n12171 ;
  assign n12173 = n12172 ^ n11756 ;
  assign n12164 = n11746 ^ x86 ;
  assign n12165 = n11973 & n12164 ;
  assign n12166 = n12165 ^ n11749 ;
  assign n12157 = n11739 ^ x85 ;
  assign n12158 = n11973 & n12157 ;
  assign n12159 = n12158 ^ n11742 ;
  assign n12150 = n11732 ^ x84 ;
  assign n12151 = n11973 & n12150 ;
  assign n12152 = n12151 ^ n11735 ;
  assign n12143 = n11725 ^ x83 ;
  assign n12144 = n11973 & n12143 ;
  assign n12145 = n12144 ^ n11728 ;
  assign n12136 = n11718 ^ x82 ;
  assign n12137 = n11973 & n12136 ;
  assign n12138 = n12137 ^ n11721 ;
  assign n12129 = n11711 ^ x81 ;
  assign n12130 = n11973 & n12129 ;
  assign n12131 = n12130 ^ n11714 ;
  assign n12122 = n11704 ^ x80 ;
  assign n12123 = n11973 & n12122 ;
  assign n12124 = n12123 ^ n11707 ;
  assign n12115 = n11697 ^ x79 ;
  assign n12116 = n11973 & n12115 ;
  assign n12117 = n12116 ^ n11700 ;
  assign n12108 = n11682 ^ x78 ;
  assign n12109 = n11973 & n12108 ;
  assign n12110 = n12109 ^ n11693 ;
  assign n12101 = n11675 ^ x77 ;
  assign n12102 = n11973 & n12101 ;
  assign n12103 = n12102 ^ n11678 ;
  assign n12094 = n11668 ^ x76 ;
  assign n12095 = n11973 & n12094 ;
  assign n12096 = n12095 ^ n11671 ;
  assign n12087 = n11661 ^ x75 ;
  assign n12088 = n11973 & n12087 ;
  assign n12089 = n12088 ^ n11664 ;
  assign n12080 = n11654 ^ x74 ;
  assign n12081 = n11973 & n12080 ;
  assign n12082 = n12081 ^ n11657 ;
  assign n12073 = n11647 ^ x73 ;
  assign n12074 = n11973 & n12073 ;
  assign n12075 = n12074 ^ n11650 ;
  assign n12066 = n11640 ^ x72 ;
  assign n12067 = n11973 & n12066 ;
  assign n12068 = n12067 ^ n11643 ;
  assign n12051 = n11555 ^ x71 ;
  assign n12052 = n12051 ^ x70 ;
  assign n12053 = n12052 ^ n11634 ;
  assign n12054 = n12053 ^ n12051 ;
  assign n12057 = n12051 ^ n711 ;
  assign n12058 = ~n12054 & ~n12057 ;
  assign n12059 = n12058 ^ n12051 ;
  assign n12060 = n11973 & ~n12059 ;
  assign n12061 = n12060 ^ n11551 ;
  assign n12044 = n11634 ^ x70 ;
  assign n12045 = n11973 & n12044 ;
  assign n12046 = n12045 ^ n11555 ;
  assign n12037 = n11627 ^ x69 ;
  assign n12038 = n11973 & n12037 ;
  assign n12039 = n12038 ^ n11630 ;
  assign n12030 = n11620 ^ x68 ;
  assign n12031 = n11973 & n12030 ;
  assign n12032 = n12031 ^ n11623 ;
  assign n12023 = n11613 ^ x67 ;
  assign n12024 = n11973 & n12023 ;
  assign n12025 = n12024 ^ n11616 ;
  assign n11984 = n11561 ^ x65 ;
  assign n11985 = n11973 & n11984 ;
  assign n11983 = n11595 ^ x10 ;
  assign n11986 = n11985 ^ n11983 ;
  assign n11987 = n11986 ^ x66 ;
  assign n11995 = x9 & x65 ;
  assign n11992 = x65 ^ x8 ;
  assign n11988 = x64 ^ x9 ;
  assign n11989 = n11988 ^ x65 ;
  assign n11993 = n11989 ^ n11973 ;
  assign n11994 = ~n11992 & n11993 ;
  assign n11996 = n11995 ^ n11994 ;
  assign n11997 = x64 & n11996 ;
  assign n11998 = n11997 ^ n11995 ;
  assign n11999 = n11998 ^ x65 ;
  assign n12000 = n11999 ^ n11986 ;
  assign n12001 = ~n11987 & n12000 ;
  assign n12002 = n12001 ^ x66 ;
  assign n12003 = n12002 ^ x67 ;
  assign n12018 = n11148 & n11508 ;
  assign n12013 = n11595 ^ n11565 ;
  assign n12014 = n11568 & n12013 ;
  assign n12005 = n11141 ^ x65 ;
  assign n12006 = n12005 ^ x10 ;
  assign n12009 = x9 & n12006 ;
  assign n12010 = n12009 ^ x10 ;
  assign n12011 = n11595 & ~n12010 ;
  assign n12012 = n12011 ^ x66 ;
  assign n12015 = n12014 ^ n12012 ;
  assign n12016 = n11973 & ~n12015 ;
  assign n12017 = n12016 ^ n11146 ;
  assign n12019 = n12018 ^ n12017 ;
  assign n12020 = n12019 ^ n12002 ;
  assign n12021 = n12003 & n12020 ;
  assign n12022 = n12021 ^ x67 ;
  assign n12026 = n12025 ^ n12022 ;
  assign n12027 = n12025 ^ x68 ;
  assign n12028 = n12026 & ~n12027 ;
  assign n12029 = n12028 ^ x68 ;
  assign n12033 = n12032 ^ n12029 ;
  assign n12034 = n12032 ^ x69 ;
  assign n12035 = n12033 & ~n12034 ;
  assign n12036 = n12035 ^ x69 ;
  assign n12040 = n12039 ^ n12036 ;
  assign n12041 = n12039 ^ x70 ;
  assign n12042 = n12040 & ~n12041 ;
  assign n12043 = n12042 ^ x70 ;
  assign n12047 = n12046 ^ n12043 ;
  assign n12048 = n12046 ^ x71 ;
  assign n12049 = n12047 & ~n12048 ;
  assign n12050 = n12049 ^ x71 ;
  assign n12062 = n12061 ^ n12050 ;
  assign n12063 = n12061 ^ x72 ;
  assign n12064 = n12062 & ~n12063 ;
  assign n12065 = n12064 ^ x72 ;
  assign n12069 = n12068 ^ n12065 ;
  assign n12070 = n12068 ^ x73 ;
  assign n12071 = n12069 & ~n12070 ;
  assign n12072 = n12071 ^ x73 ;
  assign n12076 = n12075 ^ n12072 ;
  assign n12077 = n12075 ^ x74 ;
  assign n12078 = n12076 & ~n12077 ;
  assign n12079 = n12078 ^ x74 ;
  assign n12083 = n12082 ^ n12079 ;
  assign n12084 = n12082 ^ x75 ;
  assign n12085 = n12083 & ~n12084 ;
  assign n12086 = n12085 ^ x75 ;
  assign n12090 = n12089 ^ n12086 ;
  assign n12091 = n12089 ^ x76 ;
  assign n12092 = n12090 & ~n12091 ;
  assign n12093 = n12092 ^ x76 ;
  assign n12097 = n12096 ^ n12093 ;
  assign n12098 = n12096 ^ x77 ;
  assign n12099 = n12097 & ~n12098 ;
  assign n12100 = n12099 ^ x77 ;
  assign n12104 = n12103 ^ n12100 ;
  assign n12105 = n12103 ^ x78 ;
  assign n12106 = n12104 & ~n12105 ;
  assign n12107 = n12106 ^ x78 ;
  assign n12111 = n12110 ^ n12107 ;
  assign n12112 = n12110 ^ x79 ;
  assign n12113 = n12111 & ~n12112 ;
  assign n12114 = n12113 ^ x79 ;
  assign n12118 = n12117 ^ n12114 ;
  assign n12119 = n12117 ^ x80 ;
  assign n12120 = n12118 & ~n12119 ;
  assign n12121 = n12120 ^ x80 ;
  assign n12125 = n12124 ^ n12121 ;
  assign n12126 = n12124 ^ x81 ;
  assign n12127 = n12125 & ~n12126 ;
  assign n12128 = n12127 ^ x81 ;
  assign n12132 = n12131 ^ n12128 ;
  assign n12133 = n12131 ^ x82 ;
  assign n12134 = n12132 & ~n12133 ;
  assign n12135 = n12134 ^ x82 ;
  assign n12139 = n12138 ^ n12135 ;
  assign n12140 = n12138 ^ x83 ;
  assign n12141 = n12139 & ~n12140 ;
  assign n12142 = n12141 ^ x83 ;
  assign n12146 = n12145 ^ n12142 ;
  assign n12147 = n12145 ^ x84 ;
  assign n12148 = n12146 & ~n12147 ;
  assign n12149 = n12148 ^ x84 ;
  assign n12153 = n12152 ^ n12149 ;
  assign n12154 = n12152 ^ x85 ;
  assign n12155 = n12153 & ~n12154 ;
  assign n12156 = n12155 ^ x85 ;
  assign n12160 = n12159 ^ n12156 ;
  assign n12161 = n12159 ^ x86 ;
  assign n12162 = n12160 & ~n12161 ;
  assign n12163 = n12162 ^ x86 ;
  assign n12167 = n12166 ^ n12163 ;
  assign n12168 = n12166 ^ x87 ;
  assign n12169 = n12167 & ~n12168 ;
  assign n12170 = n12169 ^ x87 ;
  assign n12174 = n12173 ^ n12170 ;
  assign n12175 = n12173 ^ x88 ;
  assign n12176 = n12174 & ~n12175 ;
  assign n12177 = n12176 ^ x88 ;
  assign n12181 = n12180 ^ n12177 ;
  assign n12182 = n12180 ^ x89 ;
  assign n12183 = n12181 & ~n12182 ;
  assign n12184 = n12183 ^ x89 ;
  assign n12188 = n12187 ^ n12184 ;
  assign n12189 = n12187 ^ x90 ;
  assign n12190 = n12188 & ~n12189 ;
  assign n12191 = n12190 ^ x90 ;
  assign n12195 = n12194 ^ n12191 ;
  assign n12196 = n12194 ^ x91 ;
  assign n12197 = n12195 & ~n12196 ;
  assign n12198 = n12197 ^ x91 ;
  assign n12202 = n12201 ^ n12198 ;
  assign n12203 = n12201 ^ x92 ;
  assign n12204 = n12202 & ~n12203 ;
  assign n12205 = n12204 ^ x92 ;
  assign n12206 = n12205 ^ n11975 ;
  assign n12207 = n12206 ^ n11981 ;
  assign n12208 = ~n11982 & n12207 ;
  assign n12209 = n12208 ^ n11981 ;
  assign n12210 = ~n11976 & n12209 ;
  assign n12211 = n12210 ^ x94 ;
  assign n12215 = n12214 ^ n12211 ;
  assign n12216 = n12214 ^ x95 ;
  assign n12217 = n12215 & ~n12216 ;
  assign n12218 = n12217 ^ x95 ;
  assign n12222 = n12221 ^ n12218 ;
  assign n12223 = n12221 ^ x96 ;
  assign n12224 = n12222 & ~n12223 ;
  assign n12225 = n12224 ^ x96 ;
  assign n12229 = n12228 ^ n12225 ;
  assign n12230 = n12228 ^ x97 ;
  assign n12231 = n12229 & ~n12230 ;
  assign n12232 = n12231 ^ x97 ;
  assign n12236 = n12235 ^ n12232 ;
  assign n12237 = n12235 ^ x98 ;
  assign n12238 = n12236 & ~n12237 ;
  assign n12239 = n12238 ^ x98 ;
  assign n12243 = n12242 ^ n12239 ;
  assign n12244 = n12242 ^ x99 ;
  assign n12245 = n12243 & ~n12244 ;
  assign n12246 = n12245 ^ x99 ;
  assign n12250 = n12249 ^ n12246 ;
  assign n12251 = n12249 ^ x100 ;
  assign n12252 = n12250 & ~n12251 ;
  assign n12253 = n12252 ^ x100 ;
  assign n12257 = n12256 ^ n12253 ;
  assign n12258 = n12256 ^ x101 ;
  assign n12259 = n12257 & ~n12258 ;
  assign n12260 = n12259 ^ x101 ;
  assign n12264 = n12263 ^ n12260 ;
  assign n12265 = n12263 ^ x102 ;
  assign n12266 = n12264 & ~n12265 ;
  assign n12267 = n12266 ^ x102 ;
  assign n12271 = n12270 ^ n12267 ;
  assign n12272 = n12270 ^ x103 ;
  assign n12273 = n12271 & ~n12272 ;
  assign n12274 = n12273 ^ x103 ;
  assign n12278 = n12277 ^ n12274 ;
  assign n12279 = n12277 ^ x104 ;
  assign n12280 = n12278 & ~n12279 ;
  assign n12281 = n12280 ^ x104 ;
  assign n12285 = n12284 ^ n12281 ;
  assign n12286 = n12284 ^ x105 ;
  assign n12287 = n12285 & ~n12286 ;
  assign n12288 = n12287 ^ x105 ;
  assign n12292 = n12291 ^ n12288 ;
  assign n12293 = n12291 ^ x106 ;
  assign n12294 = n12292 & ~n12293 ;
  assign n12295 = n12294 ^ x106 ;
  assign n12299 = n12298 ^ n12295 ;
  assign n12300 = n12298 ^ x107 ;
  assign n12301 = n12299 & ~n12300 ;
  assign n12302 = n12301 ^ x107 ;
  assign n12306 = n12305 ^ n12302 ;
  assign n12307 = n12305 ^ x108 ;
  assign n12308 = n12306 & ~n12307 ;
  assign n12309 = n12308 ^ x108 ;
  assign n12321 = n12320 ^ n12309 ;
  assign n12322 = n12320 ^ x109 ;
  assign n12323 = n12321 & ~n12322 ;
  assign n12324 = n12323 ^ x109 ;
  assign n12328 = n12327 ^ n12324 ;
  assign n12329 = n12327 ^ x110 ;
  assign n12330 = n12328 & ~n12329 ;
  assign n12331 = n12330 ^ x110 ;
  assign n12335 = n12334 ^ n12331 ;
  assign n12336 = n12334 ^ x111 ;
  assign n12337 = n12335 & ~n12336 ;
  assign n12338 = n12337 ^ x111 ;
  assign n12342 = n12341 ^ n12338 ;
  assign n12343 = n12341 ^ x112 ;
  assign n12344 = n12342 & ~n12343 ;
  assign n12345 = n12344 ^ x112 ;
  assign n12349 = n12348 ^ n12345 ;
  assign n12350 = n12348 ^ x113 ;
  assign n12351 = n12349 & ~n12350 ;
  assign n12352 = n12351 ^ x113 ;
  assign n12356 = n12355 ^ n12352 ;
  assign n12357 = n12355 ^ x114 ;
  assign n12358 = n12356 & ~n12357 ;
  assign n12359 = n12358 ^ x114 ;
  assign n12371 = n12370 ^ n12359 ;
  assign n12372 = n12370 ^ x115 ;
  assign n12373 = n12371 & ~n12372 ;
  assign n12374 = n12373 ^ x115 ;
  assign n12378 = n12377 ^ n12374 ;
  assign n12379 = n12377 ^ x116 ;
  assign n12380 = n12378 & ~n12379 ;
  assign n12381 = n12380 ^ x116 ;
  assign n12385 = n12384 ^ n12381 ;
  assign n12387 = n12386 ^ n12385 ;
  assign n12388 = n11518 ^ x116 ;
  assign n12389 = n12388 ^ x115 ;
  assign n12390 = n12389 ^ n11933 ;
  assign n12391 = n12390 ^ n12388 ;
  assign n12393 = x116 ^ x115 ;
  assign n12394 = n12393 ^ n12388 ;
  assign n12395 = ~n12391 & ~n12394 ;
  assign n12396 = n12395 ^ n12388 ;
  assign n12397 = n11973 & ~n12396 ;
  assign n12398 = n12397 ^ n11514 ;
  assign n12399 = n12398 ^ n12384 ;
  assign n12400 = n12399 ^ n12386 ;
  assign n12401 = n12387 & ~n12400 ;
  assign n12402 = n12401 ^ n12386 ;
  assign n12404 = x119 ^ x118 ;
  assign n12403 = n12384 ^ x119 ;
  assign n12405 = n12404 ^ n12403 ;
  assign n12406 = n12402 & ~n12405 ;
  assign n12407 = n12406 ^ n12404 ;
  assign n12410 = n12407 ^ n136 ;
  assign n12411 = n11953 & ~n12410 ;
  assign n12412 = n12411 ^ x119 ;
  assign n12413 = n136 & ~n12412 ;
  assign n12414 = n12398 ^ x118 ;
  assign n12415 = n12414 ^ n12381 ;
  assign n12416 = n12415 ^ x117 ;
  assign n12417 = n12416 ^ n12414 ;
  assign n12419 = n12381 ^ x118 ;
  assign n12420 = n12419 ^ n12414 ;
  assign n12421 = ~n12417 & ~n12420 ;
  assign n12422 = n12421 ^ n12414 ;
  assign n12423 = n12413 & ~n12422 ;
  assign n12424 = n12423 ^ n12384 ;
  assign n12425 = n12424 ^ x119 ;
  assign n12430 = n12424 ^ x118 ;
  assign n12426 = n12381 ^ x117 ;
  assign n12427 = n12413 & n12426 ;
  assign n12428 = n12427 ^ n12398 ;
  assign n12429 = n12428 ^ n12424 ;
  assign n12431 = n12430 ^ n12429 ;
  assign n12816 = n12374 ^ x116 ;
  assign n12817 = n12413 & n12816 ;
  assign n12818 = n12817 ^ n12377 ;
  assign n12809 = n12359 ^ x115 ;
  assign n12810 = n12413 & n12809 ;
  assign n12811 = n12810 ^ n12370 ;
  assign n12802 = n12352 ^ x114 ;
  assign n12803 = n12413 & n12802 ;
  assign n12804 = n12803 ^ n12355 ;
  assign n12795 = n12345 ^ x113 ;
  assign n12796 = n12413 & n12795 ;
  assign n12797 = n12796 ^ n12348 ;
  assign n12788 = n12338 ^ x112 ;
  assign n12789 = n12413 & n12788 ;
  assign n12790 = n12789 ^ n12341 ;
  assign n12781 = n12331 ^ x111 ;
  assign n12782 = n12413 & n12781 ;
  assign n12783 = n12782 ^ n12334 ;
  assign n12774 = n12324 ^ x110 ;
  assign n12775 = n12413 & n12774 ;
  assign n12776 = n12775 ^ n12327 ;
  assign n12767 = n12309 ^ x109 ;
  assign n12768 = n12413 & n12767 ;
  assign n12769 = n12768 ^ n12320 ;
  assign n12760 = n12302 ^ x108 ;
  assign n12761 = n12413 & n12760 ;
  assign n12762 = n12761 ^ n12305 ;
  assign n12432 = n12295 ^ x107 ;
  assign n12433 = n12413 & n12432 ;
  assign n12434 = n12433 ^ n12298 ;
  assign n12435 = n12434 ^ x108 ;
  assign n12440 = n12434 ^ x107 ;
  assign n12436 = n12288 ^ x106 ;
  assign n12437 = n12413 & n12436 ;
  assign n12438 = n12437 ^ n12291 ;
  assign n12439 = n12438 ^ n12434 ;
  assign n12441 = n12440 ^ n12439 ;
  assign n12747 = n12281 ^ x105 ;
  assign n12748 = n12413 & n12747 ;
  assign n12749 = n12748 ^ n12284 ;
  assign n12740 = n12274 ^ x104 ;
  assign n12741 = n12413 & n12740 ;
  assign n12742 = n12741 ^ n12277 ;
  assign n12733 = n12267 ^ x103 ;
  assign n12734 = n12413 & n12733 ;
  assign n12735 = n12734 ^ n12270 ;
  assign n12726 = n12260 ^ x102 ;
  assign n12727 = n12413 & n12726 ;
  assign n12728 = n12727 ^ n12263 ;
  assign n12719 = n12253 ^ x101 ;
  assign n12720 = n12413 & n12719 ;
  assign n12721 = n12720 ^ n12256 ;
  assign n12712 = n12246 ^ x100 ;
  assign n12713 = n12413 & n12712 ;
  assign n12714 = n12713 ^ n12249 ;
  assign n12705 = n12239 ^ x99 ;
  assign n12706 = n12413 & n12705 ;
  assign n12707 = n12706 ^ n12242 ;
  assign n12698 = n12232 ^ x98 ;
  assign n12699 = n12413 & n12698 ;
  assign n12700 = n12699 ^ n12235 ;
  assign n12442 = n12225 ^ x97 ;
  assign n12443 = n12413 & n12442 ;
  assign n12444 = n12443 ^ n12228 ;
  assign n12445 = n12444 ^ x98 ;
  assign n12446 = n12218 ^ x96 ;
  assign n12447 = n12413 & n12446 ;
  assign n12448 = n12447 ^ n12221 ;
  assign n12449 = n12448 ^ x97 ;
  assign n12685 = n12211 ^ x95 ;
  assign n12686 = n12413 & n12685 ;
  assign n12687 = n12686 ^ n12214 ;
  assign n12670 = n11979 ^ x94 ;
  assign n12671 = n12670 ^ n12205 ;
  assign n12672 = n12671 ^ x93 ;
  assign n12673 = n12672 ^ n12670 ;
  assign n12675 = n12205 ^ x94 ;
  assign n12676 = n12675 ^ n12670 ;
  assign n12677 = ~n12673 & ~n12676 ;
  assign n12678 = n12677 ^ n12670 ;
  assign n12679 = n12413 & ~n12678 ;
  assign n12680 = n12679 ^ n11975 ;
  assign n12663 = n12205 ^ x93 ;
  assign n12664 = n12413 & n12663 ;
  assign n12665 = n12664 ^ n11979 ;
  assign n12656 = n12198 ^ x92 ;
  assign n12657 = n12413 & n12656 ;
  assign n12658 = n12657 ^ n12201 ;
  assign n12649 = n12191 ^ x91 ;
  assign n12650 = n12413 & n12649 ;
  assign n12651 = n12650 ^ n12194 ;
  assign n12642 = n12184 ^ x90 ;
  assign n12643 = n12413 & n12642 ;
  assign n12644 = n12643 ^ n12187 ;
  assign n12635 = n12177 ^ x89 ;
  assign n12636 = n12413 & n12635 ;
  assign n12637 = n12636 ^ n12180 ;
  assign n12628 = n12170 ^ x88 ;
  assign n12629 = n12413 & n12628 ;
  assign n12630 = n12629 ^ n12173 ;
  assign n12621 = n12163 ^ x87 ;
  assign n12622 = n12413 & n12621 ;
  assign n12623 = n12622 ^ n12166 ;
  assign n12614 = n12156 ^ x86 ;
  assign n12615 = n12413 & n12614 ;
  assign n12616 = n12615 ^ n12159 ;
  assign n12607 = n12149 ^ x85 ;
  assign n12608 = n12413 & n12607 ;
  assign n12609 = n12608 ^ n12152 ;
  assign n12600 = n12142 ^ x84 ;
  assign n12601 = n12413 & n12600 ;
  assign n12602 = n12601 ^ n12145 ;
  assign n12593 = n12135 ^ x83 ;
  assign n12594 = n12413 & n12593 ;
  assign n12595 = n12594 ^ n12138 ;
  assign n12586 = n12128 ^ x82 ;
  assign n12587 = n12413 & n12586 ;
  assign n12588 = n12587 ^ n12131 ;
  assign n12579 = n12121 ^ x81 ;
  assign n12580 = n12413 & n12579 ;
  assign n12581 = n12580 ^ n12124 ;
  assign n12572 = n12114 ^ x80 ;
  assign n12573 = n12413 & n12572 ;
  assign n12574 = n12573 ^ n12117 ;
  assign n12450 = n12107 ^ x79 ;
  assign n12451 = n12413 & n12450 ;
  assign n12452 = n12451 ^ n12110 ;
  assign n12453 = n12452 ^ x80 ;
  assign n12458 = n12452 ^ x79 ;
  assign n12454 = n12100 ^ x78 ;
  assign n12455 = n12413 & n12454 ;
  assign n12456 = n12455 ^ n12103 ;
  assign n12457 = n12456 ^ n12452 ;
  assign n12459 = n12458 ^ n12457 ;
  assign n12559 = n12093 ^ x77 ;
  assign n12560 = n12413 & n12559 ;
  assign n12561 = n12560 ^ n12096 ;
  assign n12552 = n12086 ^ x76 ;
  assign n12553 = n12413 & n12552 ;
  assign n12554 = n12553 ^ n12089 ;
  assign n12545 = n12079 ^ x75 ;
  assign n12546 = n12413 & n12545 ;
  assign n12547 = n12546 ^ n12082 ;
  assign n12538 = n12072 ^ x74 ;
  assign n12539 = n12413 & n12538 ;
  assign n12540 = n12539 ^ n12075 ;
  assign n12531 = n12065 ^ x73 ;
  assign n12532 = n12413 & n12531 ;
  assign n12533 = n12532 ^ n12068 ;
  assign n12460 = n12050 ^ x72 ;
  assign n12461 = n12413 & n12460 ;
  assign n12462 = n12461 ^ n12061 ;
  assign n12463 = n12462 ^ x73 ;
  assign n12464 = n12043 ^ x71 ;
  assign n12465 = n12413 & n12464 ;
  assign n12466 = n12465 ^ n12046 ;
  assign n12467 = n12466 ^ x72 ;
  assign n12518 = n12036 ^ x70 ;
  assign n12519 = n12413 & n12518 ;
  assign n12520 = n12519 ^ n12039 ;
  assign n12511 = n12029 ^ x69 ;
  assign n12512 = n12413 & n12511 ;
  assign n12513 = n12512 ^ n12032 ;
  assign n12504 = n12022 ^ x68 ;
  assign n12505 = n12413 & n12504 ;
  assign n12506 = n12505 ^ n12025 ;
  assign n12481 = x65 ^ x7 ;
  assign n12482 = x64 ^ x8 ;
  assign n12483 = n12482 ^ x65 ;
  assign n12484 = n12483 ^ n12413 ;
  assign n12485 = ~n12481 & n12484 ;
  assign n12480 = x8 & x65 ;
  assign n12486 = n12485 ^ n12480 ;
  assign n12489 = x64 & n12486 ;
  assign n12490 = n12489 ^ n12480 ;
  assign n12491 = n12490 ^ x65 ;
  assign n12478 = x64 & n11973 ;
  assign n12474 = ~x8 & x64 ;
  assign n12475 = n12474 ^ x65 ;
  assign n12476 = n12413 & n12475 ;
  assign n12477 = n12476 ^ x9 ;
  assign n12479 = n12478 ^ n12477 ;
  assign n12492 = n12491 ^ n12479 ;
  assign n12493 = n12491 ^ x66 ;
  assign n12494 = n12492 & n12493 ;
  assign n12495 = n12494 ^ x66 ;
  assign n12470 = n11999 ^ x66 ;
  assign n12471 = n12413 & n12470 ;
  assign n12472 = n12471 ^ n11986 ;
  assign n12496 = n12495 ^ n12472 ;
  assign n12497 = n12495 ^ x67 ;
  assign n12498 = n12496 & n12497 ;
  assign n12499 = n12498 ^ x67 ;
  assign n12468 = n12003 & n12413 ;
  assign n12469 = n12468 ^ n12019 ;
  assign n12500 = n12499 ^ n12469 ;
  assign n12501 = n12499 ^ x68 ;
  assign n12502 = n12500 & n12501 ;
  assign n12503 = n12502 ^ x68 ;
  assign n12507 = n12506 ^ n12503 ;
  assign n12508 = n12506 ^ x69 ;
  assign n12509 = n12507 & ~n12508 ;
  assign n12510 = n12509 ^ x69 ;
  assign n12514 = n12513 ^ n12510 ;
  assign n12515 = n12513 ^ x70 ;
  assign n12516 = n12514 & ~n12515 ;
  assign n12517 = n12516 ^ x70 ;
  assign n12521 = n12520 ^ n12517 ;
  assign n12522 = n12520 ^ x71 ;
  assign n12523 = n12521 & ~n12522 ;
  assign n12524 = n12523 ^ x71 ;
  assign n12525 = n12524 ^ n12466 ;
  assign n12526 = ~n12467 & n12525 ;
  assign n12527 = n12526 ^ x72 ;
  assign n12528 = n12527 ^ n12462 ;
  assign n12529 = ~n12463 & n12528 ;
  assign n12530 = n12529 ^ x73 ;
  assign n12534 = n12533 ^ n12530 ;
  assign n12535 = n12533 ^ x74 ;
  assign n12536 = n12534 & ~n12535 ;
  assign n12537 = n12536 ^ x74 ;
  assign n12541 = n12540 ^ n12537 ;
  assign n12542 = n12540 ^ x75 ;
  assign n12543 = n12541 & ~n12542 ;
  assign n12544 = n12543 ^ x75 ;
  assign n12548 = n12547 ^ n12544 ;
  assign n12549 = n12547 ^ x76 ;
  assign n12550 = n12548 & ~n12549 ;
  assign n12551 = n12550 ^ x76 ;
  assign n12555 = n12554 ^ n12551 ;
  assign n12556 = n12554 ^ x77 ;
  assign n12557 = n12555 & ~n12556 ;
  assign n12558 = n12557 ^ x77 ;
  assign n12562 = n12561 ^ n12558 ;
  assign n12563 = n12561 ^ x78 ;
  assign n12564 = n12562 & ~n12563 ;
  assign n12565 = n12564 ^ x78 ;
  assign n12566 = n12565 ^ n12452 ;
  assign n12567 = n12566 ^ n12458 ;
  assign n12568 = ~n12459 & n12567 ;
  assign n12569 = n12568 ^ n12458 ;
  assign n12570 = ~n12453 & n12569 ;
  assign n12571 = n12570 ^ x80 ;
  assign n12575 = n12574 ^ n12571 ;
  assign n12576 = n12574 ^ x81 ;
  assign n12577 = n12575 & ~n12576 ;
  assign n12578 = n12577 ^ x81 ;
  assign n12582 = n12581 ^ n12578 ;
  assign n12583 = n12581 ^ x82 ;
  assign n12584 = n12582 & ~n12583 ;
  assign n12585 = n12584 ^ x82 ;
  assign n12589 = n12588 ^ n12585 ;
  assign n12590 = n12588 ^ x83 ;
  assign n12591 = n12589 & ~n12590 ;
  assign n12592 = n12591 ^ x83 ;
  assign n12596 = n12595 ^ n12592 ;
  assign n12597 = n12595 ^ x84 ;
  assign n12598 = n12596 & ~n12597 ;
  assign n12599 = n12598 ^ x84 ;
  assign n12603 = n12602 ^ n12599 ;
  assign n12604 = n12602 ^ x85 ;
  assign n12605 = n12603 & ~n12604 ;
  assign n12606 = n12605 ^ x85 ;
  assign n12610 = n12609 ^ n12606 ;
  assign n12611 = n12609 ^ x86 ;
  assign n12612 = n12610 & ~n12611 ;
  assign n12613 = n12612 ^ x86 ;
  assign n12617 = n12616 ^ n12613 ;
  assign n12618 = n12616 ^ x87 ;
  assign n12619 = n12617 & ~n12618 ;
  assign n12620 = n12619 ^ x87 ;
  assign n12624 = n12623 ^ n12620 ;
  assign n12625 = n12623 ^ x88 ;
  assign n12626 = n12624 & ~n12625 ;
  assign n12627 = n12626 ^ x88 ;
  assign n12631 = n12630 ^ n12627 ;
  assign n12632 = n12630 ^ x89 ;
  assign n12633 = n12631 & ~n12632 ;
  assign n12634 = n12633 ^ x89 ;
  assign n12638 = n12637 ^ n12634 ;
  assign n12639 = n12637 ^ x90 ;
  assign n12640 = n12638 & ~n12639 ;
  assign n12641 = n12640 ^ x90 ;
  assign n12645 = n12644 ^ n12641 ;
  assign n12646 = n12644 ^ x91 ;
  assign n12647 = n12645 & ~n12646 ;
  assign n12648 = n12647 ^ x91 ;
  assign n12652 = n12651 ^ n12648 ;
  assign n12653 = n12651 ^ x92 ;
  assign n12654 = n12652 & ~n12653 ;
  assign n12655 = n12654 ^ x92 ;
  assign n12659 = n12658 ^ n12655 ;
  assign n12660 = n12658 ^ x93 ;
  assign n12661 = n12659 & ~n12660 ;
  assign n12662 = n12661 ^ x93 ;
  assign n12666 = n12665 ^ n12662 ;
  assign n12667 = n12665 ^ x94 ;
  assign n12668 = n12666 & ~n12667 ;
  assign n12669 = n12668 ^ x94 ;
  assign n12681 = n12680 ^ n12669 ;
  assign n12682 = n12680 ^ x95 ;
  assign n12683 = n12681 & ~n12682 ;
  assign n12684 = n12683 ^ x95 ;
  assign n12688 = n12687 ^ n12684 ;
  assign n12689 = n12687 ^ x96 ;
  assign n12690 = n12688 & ~n12689 ;
  assign n12691 = n12690 ^ x96 ;
  assign n12692 = n12691 ^ n12448 ;
  assign n12693 = ~n12449 & n12692 ;
  assign n12694 = n12693 ^ x97 ;
  assign n12695 = n12694 ^ n12444 ;
  assign n12696 = ~n12445 & n12695 ;
  assign n12697 = n12696 ^ x98 ;
  assign n12701 = n12700 ^ n12697 ;
  assign n12702 = n12700 ^ x99 ;
  assign n12703 = n12701 & ~n12702 ;
  assign n12704 = n12703 ^ x99 ;
  assign n12708 = n12707 ^ n12704 ;
  assign n12709 = n12707 ^ x100 ;
  assign n12710 = n12708 & ~n12709 ;
  assign n12711 = n12710 ^ x100 ;
  assign n12715 = n12714 ^ n12711 ;
  assign n12716 = n12714 ^ x101 ;
  assign n12717 = n12715 & ~n12716 ;
  assign n12718 = n12717 ^ x101 ;
  assign n12722 = n12721 ^ n12718 ;
  assign n12723 = n12721 ^ x102 ;
  assign n12724 = n12722 & ~n12723 ;
  assign n12725 = n12724 ^ x102 ;
  assign n12729 = n12728 ^ n12725 ;
  assign n12730 = n12728 ^ x103 ;
  assign n12731 = n12729 & ~n12730 ;
  assign n12732 = n12731 ^ x103 ;
  assign n12736 = n12735 ^ n12732 ;
  assign n12737 = n12735 ^ x104 ;
  assign n12738 = n12736 & ~n12737 ;
  assign n12739 = n12738 ^ x104 ;
  assign n12743 = n12742 ^ n12739 ;
  assign n12744 = n12742 ^ x105 ;
  assign n12745 = n12743 & ~n12744 ;
  assign n12746 = n12745 ^ x105 ;
  assign n12750 = n12749 ^ n12746 ;
  assign n12751 = n12749 ^ x106 ;
  assign n12752 = n12750 & ~n12751 ;
  assign n12753 = n12752 ^ x106 ;
  assign n12754 = n12753 ^ n12434 ;
  assign n12755 = n12754 ^ n12440 ;
  assign n12756 = ~n12441 & n12755 ;
  assign n12757 = n12756 ^ n12440 ;
  assign n12758 = ~n12435 & n12757 ;
  assign n12759 = n12758 ^ x108 ;
  assign n12763 = n12762 ^ n12759 ;
  assign n12764 = n12762 ^ x109 ;
  assign n12765 = n12763 & ~n12764 ;
  assign n12766 = n12765 ^ x109 ;
  assign n12770 = n12769 ^ n12766 ;
  assign n12771 = n12769 ^ x110 ;
  assign n12772 = n12770 & ~n12771 ;
  assign n12773 = n12772 ^ x110 ;
  assign n12777 = n12776 ^ n12773 ;
  assign n12778 = n12776 ^ x111 ;
  assign n12779 = n12777 & ~n12778 ;
  assign n12780 = n12779 ^ x111 ;
  assign n12784 = n12783 ^ n12780 ;
  assign n12785 = n12783 ^ x112 ;
  assign n12786 = n12784 & ~n12785 ;
  assign n12787 = n12786 ^ x112 ;
  assign n12791 = n12790 ^ n12787 ;
  assign n12792 = n12790 ^ x113 ;
  assign n12793 = n12791 & ~n12792 ;
  assign n12794 = n12793 ^ x113 ;
  assign n12798 = n12797 ^ n12794 ;
  assign n12799 = n12797 ^ x114 ;
  assign n12800 = n12798 & ~n12799 ;
  assign n12801 = n12800 ^ x114 ;
  assign n12805 = n12804 ^ n12801 ;
  assign n12806 = n12804 ^ x115 ;
  assign n12807 = n12805 & ~n12806 ;
  assign n12808 = n12807 ^ x115 ;
  assign n12812 = n12811 ^ n12808 ;
  assign n12813 = n12811 ^ x116 ;
  assign n12814 = n12812 & ~n12813 ;
  assign n12815 = n12814 ^ x116 ;
  assign n12819 = n12818 ^ n12815 ;
  assign n12820 = n12818 ^ x117 ;
  assign n12821 = n12819 & ~n12820 ;
  assign n12822 = n12821 ^ x117 ;
  assign n12823 = n12822 ^ n12424 ;
  assign n12824 = n12823 ^ n12430 ;
  assign n12825 = ~n12431 & n12824 ;
  assign n12826 = n12825 ^ n12430 ;
  assign n12827 = ~n12425 & n12826 ;
  assign n12828 = n12827 ^ x119 ;
  assign n12829 = n12828 ^ x120 ;
  assign n12830 = n136 & n11950 ;
  assign n12831 = n12407 & n12830 ;
  assign n12832 = n12831 ^ n11950 ;
  assign n12833 = n135 & n12832 ;
  assign n12834 = n12829 & n12833 ;
  assign n12835 = n12834 ^ n12832 ;
  assign n12836 = x124 & n131 ;
  assign n12837 = ~n12835 & n12836 ;
  assign n12838 = n12837 ^ n131 ;
  assign n12840 = x120 & n135 ;
  assign n12841 = ~n11510 & n12840 ;
  assign n12842 = n12841 ^ n135 ;
  assign n12843 = n12828 & n12842 ;
  assign n12844 = n12832 ^ x120 ;
  assign n12845 = n12844 ^ n12841 ;
  assign n12846 = n12843 & ~n12845 ;
  assign n12847 = n12846 ^ n12842 ;
  assign n13258 = n12428 ^ x119 ;
  assign n13259 = n13258 ^ n12822 ;
  assign n13260 = n13259 ^ x118 ;
  assign n13261 = n13260 ^ n13258 ;
  assign n13263 = n12822 ^ x119 ;
  assign n13264 = n13263 ^ n13258 ;
  assign n13265 = ~n13261 & ~n13264 ;
  assign n13266 = n13265 ^ n13258 ;
  assign n13267 = n12847 & ~n13266 ;
  assign n13268 = n13267 ^ n12424 ;
  assign n13251 = n12822 ^ x118 ;
  assign n13252 = n12847 & n13251 ;
  assign n13253 = n13252 ^ n12428 ;
  assign n13244 = n12815 ^ x117 ;
  assign n13245 = n12847 & n13244 ;
  assign n13246 = n13245 ^ n12818 ;
  assign n13237 = n12808 ^ x116 ;
  assign n13238 = n12847 & n13237 ;
  assign n13239 = n13238 ^ n12811 ;
  assign n13230 = n12801 ^ x115 ;
  assign n13231 = n12847 & n13230 ;
  assign n13232 = n13231 ^ n12804 ;
  assign n13223 = n12794 ^ x114 ;
  assign n13224 = n12847 & n13223 ;
  assign n13225 = n13224 ^ n12797 ;
  assign n13216 = n12787 ^ x113 ;
  assign n13217 = n12847 & n13216 ;
  assign n13218 = n13217 ^ n12790 ;
  assign n13155 = n12780 ^ x112 ;
  assign n13156 = n12847 & n13155 ;
  assign n13157 = n13156 ^ n12783 ;
  assign n13158 = n13157 ^ x113 ;
  assign n13163 = n13157 ^ x112 ;
  assign n13159 = n12773 ^ x111 ;
  assign n13160 = n12847 & n13159 ;
  assign n13161 = n13160 ^ n12776 ;
  assign n13162 = n13161 ^ n13157 ;
  assign n13164 = n13163 ^ n13162 ;
  assign n13199 = n12759 ^ x109 ;
  assign n13200 = n12847 & n13199 ;
  assign n13201 = n13200 ^ n12762 ;
  assign n13168 = n12438 ^ x108 ;
  assign n13169 = n13168 ^ n12753 ;
  assign n13170 = n13169 ^ x107 ;
  assign n13171 = n13170 ^ n13168 ;
  assign n13173 = n12753 ^ x108 ;
  assign n13174 = n13173 ^ n13168 ;
  assign n13175 = ~n13171 & ~n13174 ;
  assign n13176 = n13175 ^ n13168 ;
  assign n13177 = n12847 & ~n13176 ;
  assign n13178 = n13177 ^ n12434 ;
  assign n13179 = n13178 ^ x109 ;
  assign n13184 = n13178 ^ x108 ;
  assign n13180 = n12753 ^ x107 ;
  assign n13181 = n12847 & n13180 ;
  assign n13182 = n13181 ^ n12438 ;
  assign n13183 = n13182 ^ n13178 ;
  assign n13185 = n13184 ^ n13183 ;
  assign n13186 = n12746 ^ x106 ;
  assign n13187 = n12847 & n13186 ;
  assign n13188 = n13187 ^ n12749 ;
  assign n13144 = n12739 ^ x105 ;
  assign n13145 = n12847 & n13144 ;
  assign n13146 = n13145 ^ n12742 ;
  assign n13137 = n12732 ^ x104 ;
  assign n13138 = n12847 & n13137 ;
  assign n13139 = n13138 ^ n12735 ;
  assign n13130 = n12725 ^ x103 ;
  assign n13131 = n12847 & n13130 ;
  assign n13132 = n13131 ^ n12728 ;
  assign n13123 = n12718 ^ x102 ;
  assign n13124 = n12847 & n13123 ;
  assign n13125 = n13124 ^ n12721 ;
  assign n13116 = n12711 ^ x101 ;
  assign n13117 = n12847 & n13116 ;
  assign n13118 = n13117 ^ n12714 ;
  assign n13109 = n12704 ^ x100 ;
  assign n13110 = n12847 & n13109 ;
  assign n13111 = n13110 ^ n12707 ;
  assign n12839 = n12697 ^ x99 ;
  assign n12848 = n12839 & n12847 ;
  assign n12849 = n12848 ^ n12700 ;
  assign n12850 = n12849 ^ x100 ;
  assign n12851 = n12694 ^ x98 ;
  assign n12852 = n12847 & n12851 ;
  assign n12853 = n12852 ^ n12444 ;
  assign n12854 = n12853 ^ x99 ;
  assign n13096 = n12691 ^ x97 ;
  assign n13097 = n12847 & n13096 ;
  assign n13098 = n13097 ^ n12448 ;
  assign n13089 = n12684 ^ x96 ;
  assign n13090 = n12847 & n13089 ;
  assign n13091 = n13090 ^ n12687 ;
  assign n12855 = n12669 ^ x95 ;
  assign n12856 = n12847 & n12855 ;
  assign n12857 = n12856 ^ n12680 ;
  assign n12858 = n12857 ^ x96 ;
  assign n12859 = n12662 ^ x94 ;
  assign n12860 = n12847 & n12859 ;
  assign n12861 = n12860 ^ n12665 ;
  assign n12862 = n12861 ^ x95 ;
  assign n13076 = n12655 ^ x93 ;
  assign n13077 = n12847 & n13076 ;
  assign n13078 = n13077 ^ n12658 ;
  assign n13069 = n12648 ^ x92 ;
  assign n13070 = n12847 & n13069 ;
  assign n13071 = n13070 ^ n12651 ;
  assign n13062 = n12641 ^ x91 ;
  assign n13063 = n12847 & n13062 ;
  assign n13064 = n13063 ^ n12644 ;
  assign n13055 = n12634 ^ x90 ;
  assign n13056 = n12847 & n13055 ;
  assign n13057 = n13056 ^ n12637 ;
  assign n12863 = n12620 ^ x88 ;
  assign n12864 = n12847 & n12863 ;
  assign n12865 = n12864 ^ n12623 ;
  assign n12866 = n12865 ^ x89 ;
  assign n13038 = n12613 ^ x87 ;
  assign n13039 = n12847 & n13038 ;
  assign n13040 = n13039 ^ n12616 ;
  assign n13031 = n12606 ^ x86 ;
  assign n13032 = n12847 & n13031 ;
  assign n13033 = n13032 ^ n12609 ;
  assign n13024 = n12599 ^ x85 ;
  assign n13025 = n12847 & n13024 ;
  assign n13026 = n13025 ^ n12602 ;
  assign n13017 = n12592 ^ x84 ;
  assign n13018 = n12847 & n13017 ;
  assign n13019 = n13018 ^ n12595 ;
  assign n13010 = n12585 ^ x83 ;
  assign n13011 = n12847 & n13010 ;
  assign n13012 = n13011 ^ n12588 ;
  assign n13003 = n12578 ^ x82 ;
  assign n13004 = n12847 & n13003 ;
  assign n13005 = n13004 ^ n12581 ;
  assign n12996 = n12571 ^ x81 ;
  assign n12997 = n12847 & n12996 ;
  assign n12998 = n12997 ^ n12574 ;
  assign n12981 = n12456 ^ x80 ;
  assign n12982 = n12981 ^ n12565 ;
  assign n12983 = n12982 ^ x79 ;
  assign n12984 = n12983 ^ n12981 ;
  assign n12986 = n12565 ^ x80 ;
  assign n12987 = n12986 ^ n12981 ;
  assign n12988 = ~n12984 & ~n12987 ;
  assign n12989 = n12988 ^ n12981 ;
  assign n12990 = n12847 & ~n12989 ;
  assign n12991 = n12990 ^ n12452 ;
  assign n12974 = n12565 ^ x79 ;
  assign n12975 = n12847 & n12974 ;
  assign n12976 = n12975 ^ n12456 ;
  assign n12967 = n12558 ^ x78 ;
  assign n12968 = n12847 & n12967 ;
  assign n12969 = n12968 ^ n12561 ;
  assign n12960 = n12551 ^ x77 ;
  assign n12961 = n12847 & n12960 ;
  assign n12962 = n12961 ^ n12554 ;
  assign n12867 = n12544 ^ x76 ;
  assign n12868 = n12847 & n12867 ;
  assign n12869 = n12868 ^ n12547 ;
  assign n12870 = n12869 ^ x77 ;
  assign n12875 = n12869 ^ x76 ;
  assign n12871 = n12537 ^ x75 ;
  assign n12872 = n12847 & n12871 ;
  assign n12873 = n12872 ^ n12540 ;
  assign n12874 = n12873 ^ n12869 ;
  assign n12876 = n12875 ^ n12874 ;
  assign n12947 = n12530 ^ x74 ;
  assign n12948 = n12847 & n12947 ;
  assign n12949 = n12948 ^ n12533 ;
  assign n12940 = n12527 ^ x73 ;
  assign n12941 = n12847 & n12940 ;
  assign n12942 = n12941 ^ n12462 ;
  assign n12933 = n12524 ^ x72 ;
  assign n12934 = n12847 & n12933 ;
  assign n12935 = n12934 ^ n12466 ;
  assign n12926 = n12517 ^ x71 ;
  assign n12927 = n12847 & n12926 ;
  assign n12928 = n12927 ^ n12520 ;
  assign n12919 = n12510 ^ x70 ;
  assign n12920 = n12847 & n12919 ;
  assign n12921 = n12920 ^ n12513 ;
  assign n12912 = n12503 ^ x69 ;
  assign n12913 = n12847 & n12912 ;
  assign n12914 = n12913 ^ n12506 ;
  assign n12906 = n12501 & n12847 ;
  assign n12907 = n12906 ^ n12469 ;
  assign n12900 = n12497 & n12847 ;
  assign n12901 = n12900 ^ n12472 ;
  assign n12894 = n12493 & n12847 ;
  assign n12895 = n12894 ^ n12479 ;
  assign n12881 = x64 & n12847 ;
  assign n12882 = ~x7 & n12881 ;
  assign n12878 = x64 & n12413 ;
  assign n12877 = x65 & n12847 ;
  assign n12879 = n12878 ^ n12877 ;
  assign n12880 = n12879 ^ x8 ;
  assign n12883 = n12882 ^ n12880 ;
  assign n12884 = n12883 ^ x66 ;
  assign n12885 = ~x6 & x64 ;
  assign n12886 = n12885 ^ x65 ;
  assign n12887 = n12881 ^ x65 ;
  assign n12888 = n12887 ^ x7 ;
  assign n12889 = n12886 & ~n12888 ;
  assign n12890 = n12889 ^ x65 ;
  assign n12891 = n12890 ^ n12883 ;
  assign n12892 = ~n12884 & n12891 ;
  assign n12893 = n12892 ^ x66 ;
  assign n12896 = n12895 ^ n12893 ;
  assign n12897 = n12895 ^ x67 ;
  assign n12898 = n12896 & ~n12897 ;
  assign n12899 = n12898 ^ x67 ;
  assign n12902 = n12901 ^ n12899 ;
  assign n12903 = n12901 ^ x68 ;
  assign n12904 = n12902 & ~n12903 ;
  assign n12905 = n12904 ^ x68 ;
  assign n12908 = n12907 ^ n12905 ;
  assign n12909 = n12907 ^ x69 ;
  assign n12910 = n12908 & ~n12909 ;
  assign n12911 = n12910 ^ x69 ;
  assign n12915 = n12914 ^ n12911 ;
  assign n12916 = n12914 ^ x70 ;
  assign n12917 = n12915 & ~n12916 ;
  assign n12918 = n12917 ^ x70 ;
  assign n12922 = n12921 ^ n12918 ;
  assign n12923 = n12921 ^ x71 ;
  assign n12924 = n12922 & ~n12923 ;
  assign n12925 = n12924 ^ x71 ;
  assign n12929 = n12928 ^ n12925 ;
  assign n12930 = n12928 ^ x72 ;
  assign n12931 = n12929 & ~n12930 ;
  assign n12932 = n12931 ^ x72 ;
  assign n12936 = n12935 ^ n12932 ;
  assign n12937 = n12935 ^ x73 ;
  assign n12938 = n12936 & ~n12937 ;
  assign n12939 = n12938 ^ x73 ;
  assign n12943 = n12942 ^ n12939 ;
  assign n12944 = n12942 ^ x74 ;
  assign n12945 = n12943 & ~n12944 ;
  assign n12946 = n12945 ^ x74 ;
  assign n12950 = n12949 ^ n12946 ;
  assign n12951 = n12949 ^ x75 ;
  assign n12952 = n12950 & ~n12951 ;
  assign n12953 = n12952 ^ x75 ;
  assign n12954 = n12953 ^ n12869 ;
  assign n12955 = n12954 ^ n12875 ;
  assign n12956 = ~n12876 & n12955 ;
  assign n12957 = n12956 ^ n12875 ;
  assign n12958 = ~n12870 & n12957 ;
  assign n12959 = n12958 ^ x77 ;
  assign n12963 = n12962 ^ n12959 ;
  assign n12964 = n12962 ^ x78 ;
  assign n12965 = n12963 & ~n12964 ;
  assign n12966 = n12965 ^ x78 ;
  assign n12970 = n12969 ^ n12966 ;
  assign n12971 = n12969 ^ x79 ;
  assign n12972 = n12970 & ~n12971 ;
  assign n12973 = n12972 ^ x79 ;
  assign n12977 = n12976 ^ n12973 ;
  assign n12978 = n12976 ^ x80 ;
  assign n12979 = n12977 & ~n12978 ;
  assign n12980 = n12979 ^ x80 ;
  assign n12992 = n12991 ^ n12980 ;
  assign n12993 = n12991 ^ x81 ;
  assign n12994 = n12992 & ~n12993 ;
  assign n12995 = n12994 ^ x81 ;
  assign n12999 = n12998 ^ n12995 ;
  assign n13000 = n12998 ^ x82 ;
  assign n13001 = n12999 & ~n13000 ;
  assign n13002 = n13001 ^ x82 ;
  assign n13006 = n13005 ^ n13002 ;
  assign n13007 = n13005 ^ x83 ;
  assign n13008 = n13006 & ~n13007 ;
  assign n13009 = n13008 ^ x83 ;
  assign n13013 = n13012 ^ n13009 ;
  assign n13014 = n13012 ^ x84 ;
  assign n13015 = n13013 & ~n13014 ;
  assign n13016 = n13015 ^ x84 ;
  assign n13020 = n13019 ^ n13016 ;
  assign n13021 = n13019 ^ x85 ;
  assign n13022 = n13020 & ~n13021 ;
  assign n13023 = n13022 ^ x85 ;
  assign n13027 = n13026 ^ n13023 ;
  assign n13028 = n13026 ^ x86 ;
  assign n13029 = n13027 & ~n13028 ;
  assign n13030 = n13029 ^ x86 ;
  assign n13034 = n13033 ^ n13030 ;
  assign n13035 = n13033 ^ x87 ;
  assign n13036 = n13034 & ~n13035 ;
  assign n13037 = n13036 ^ x87 ;
  assign n13041 = n13040 ^ n13037 ;
  assign n13042 = n13040 ^ x88 ;
  assign n13043 = n13041 & ~n13042 ;
  assign n13044 = n13043 ^ x88 ;
  assign n13045 = n13044 ^ n12865 ;
  assign n13046 = ~n12866 & n13045 ;
  assign n13047 = n13046 ^ x89 ;
  assign n13048 = n13047 ^ x90 ;
  assign n13049 = n12627 ^ x89 ;
  assign n13050 = n12847 & n13049 ;
  assign n13051 = n13050 ^ n12630 ;
  assign n13052 = n13051 ^ n13047 ;
  assign n13053 = n13048 & n13052 ;
  assign n13054 = n13053 ^ x90 ;
  assign n13058 = n13057 ^ n13054 ;
  assign n13059 = n13057 ^ x91 ;
  assign n13060 = n13058 & ~n13059 ;
  assign n13061 = n13060 ^ x91 ;
  assign n13065 = n13064 ^ n13061 ;
  assign n13066 = n13064 ^ x92 ;
  assign n13067 = n13065 & ~n13066 ;
  assign n13068 = n13067 ^ x92 ;
  assign n13072 = n13071 ^ n13068 ;
  assign n13073 = n13071 ^ x93 ;
  assign n13074 = n13072 & ~n13073 ;
  assign n13075 = n13074 ^ x93 ;
  assign n13079 = n13078 ^ n13075 ;
  assign n13080 = n13078 ^ x94 ;
  assign n13081 = n13079 & ~n13080 ;
  assign n13082 = n13081 ^ x94 ;
  assign n13083 = n13082 ^ n12861 ;
  assign n13084 = ~n12862 & n13083 ;
  assign n13085 = n13084 ^ x95 ;
  assign n13086 = n13085 ^ n12857 ;
  assign n13087 = ~n12858 & n13086 ;
  assign n13088 = n13087 ^ x96 ;
  assign n13092 = n13091 ^ n13088 ;
  assign n13093 = n13091 ^ x97 ;
  assign n13094 = n13092 & ~n13093 ;
  assign n13095 = n13094 ^ x97 ;
  assign n13099 = n13098 ^ n13095 ;
  assign n13100 = n13098 ^ x98 ;
  assign n13101 = n13099 & ~n13100 ;
  assign n13102 = n13101 ^ x98 ;
  assign n13103 = n13102 ^ n12853 ;
  assign n13104 = ~n12854 & n13103 ;
  assign n13105 = n13104 ^ x99 ;
  assign n13106 = n13105 ^ n12849 ;
  assign n13107 = ~n12850 & n13106 ;
  assign n13108 = n13107 ^ x100 ;
  assign n13112 = n13111 ^ n13108 ;
  assign n13113 = n13111 ^ x101 ;
  assign n13114 = n13112 & ~n13113 ;
  assign n13115 = n13114 ^ x101 ;
  assign n13119 = n13118 ^ n13115 ;
  assign n13120 = n13118 ^ x102 ;
  assign n13121 = n13119 & ~n13120 ;
  assign n13122 = n13121 ^ x102 ;
  assign n13126 = n13125 ^ n13122 ;
  assign n13127 = n13125 ^ x103 ;
  assign n13128 = n13126 & ~n13127 ;
  assign n13129 = n13128 ^ x103 ;
  assign n13133 = n13132 ^ n13129 ;
  assign n13134 = n13132 ^ x104 ;
  assign n13135 = n13133 & ~n13134 ;
  assign n13136 = n13135 ^ x104 ;
  assign n13140 = n13139 ^ n13136 ;
  assign n13141 = n13139 ^ x105 ;
  assign n13142 = n13140 & ~n13141 ;
  assign n13143 = n13142 ^ x105 ;
  assign n13147 = n13146 ^ n13143 ;
  assign n13148 = n13146 ^ x106 ;
  assign n13149 = n13147 & ~n13148 ;
  assign n13150 = n13149 ^ x106 ;
  assign n13189 = n13188 ^ n13150 ;
  assign n13190 = n13188 ^ x107 ;
  assign n13191 = n13189 & ~n13190 ;
  assign n13192 = n13191 ^ x107 ;
  assign n13193 = n13192 ^ n13178 ;
  assign n13194 = n13193 ^ n13184 ;
  assign n13195 = ~n13185 & n13194 ;
  assign n13196 = n13195 ^ n13184 ;
  assign n13197 = ~n13179 & n13196 ;
  assign n13198 = n13197 ^ x109 ;
  assign n13202 = n13201 ^ n13198 ;
  assign n13203 = n13201 ^ x110 ;
  assign n13204 = n13202 & ~n13203 ;
  assign n13205 = n13204 ^ x110 ;
  assign n13165 = n12766 ^ x110 ;
  assign n13166 = n12847 & n13165 ;
  assign n13167 = n13166 ^ n12769 ;
  assign n13206 = n13205 ^ n13167 ;
  assign n13207 = n13205 ^ x111 ;
  assign n13208 = n13206 & n13207 ;
  assign n13209 = n13208 ^ x111 ;
  assign n13210 = n13209 ^ n13157 ;
  assign n13211 = n13210 ^ n13163 ;
  assign n13212 = ~n13164 & n13211 ;
  assign n13213 = n13212 ^ n13163 ;
  assign n13214 = ~n13158 & n13213 ;
  assign n13215 = n13214 ^ x113 ;
  assign n13219 = n13218 ^ n13215 ;
  assign n13220 = n13218 ^ x114 ;
  assign n13221 = n13219 & ~n13220 ;
  assign n13222 = n13221 ^ x114 ;
  assign n13226 = n13225 ^ n13222 ;
  assign n13227 = n13225 ^ x115 ;
  assign n13228 = n13226 & ~n13227 ;
  assign n13229 = n13228 ^ x115 ;
  assign n13233 = n13232 ^ n13229 ;
  assign n13234 = n13232 ^ x116 ;
  assign n13235 = n13233 & ~n13234 ;
  assign n13236 = n13235 ^ x116 ;
  assign n13240 = n13239 ^ n13236 ;
  assign n13241 = n13239 ^ x117 ;
  assign n13242 = n13240 & ~n13241 ;
  assign n13243 = n13242 ^ x117 ;
  assign n13247 = n13246 ^ n13243 ;
  assign n13248 = n13246 ^ x118 ;
  assign n13249 = n13247 & ~n13248 ;
  assign n13250 = n13249 ^ x118 ;
  assign n13254 = n13253 ^ n13250 ;
  assign n13255 = n13253 ^ x119 ;
  assign n13256 = n13254 & ~n13255 ;
  assign n13257 = n13256 ^ x119 ;
  assign n13269 = n13268 ^ n13257 ;
  assign n13270 = n13268 ^ x120 ;
  assign n13271 = n13269 & ~n13270 ;
  assign n13272 = n13271 ^ x120 ;
  assign n14064 = ~x121 & n12835 ;
  assign n14065 = ~n13272 & n14064 ;
  assign n13152 = n12835 ^ n11950 ;
  assign n13153 = ~x121 & ~n13152 ;
  assign n13154 = n13153 ^ n11950 ;
  assign n13273 = n13272 ^ x121 ;
  assign n13274 = n13273 ^ n134 ;
  assign n13275 = n13154 & ~n13274 ;
  assign n13276 = n13275 ^ x121 ;
  assign n13277 = n134 & ~n13276 ;
  assign n13697 = n13257 ^ x120 ;
  assign n13698 = n13277 & n13697 ;
  assign n13699 = n13698 ^ n13268 ;
  assign n13605 = n13250 ^ x119 ;
  assign n13606 = n13277 & n13605 ;
  assign n13607 = n13606 ^ n13253 ;
  assign n13608 = n13607 ^ x120 ;
  assign n13609 = n13243 ^ x118 ;
  assign n13610 = n13277 & n13609 ;
  assign n13611 = n13610 ^ n13246 ;
  assign n13612 = n13611 ^ x119 ;
  assign n13613 = n13236 ^ x117 ;
  assign n13614 = n13277 & n13613 ;
  assign n13615 = n13614 ^ n13239 ;
  assign n13616 = n13615 ^ x118 ;
  assign n13681 = n13229 ^ x116 ;
  assign n13682 = n13277 & n13681 ;
  assign n13683 = n13682 ^ n13232 ;
  assign n13674 = n13222 ^ x115 ;
  assign n13675 = n13277 & n13674 ;
  assign n13676 = n13675 ^ n13225 ;
  assign n13617 = n13215 ^ x114 ;
  assign n13618 = n13277 & n13617 ;
  assign n13619 = n13618 ^ n13218 ;
  assign n13620 = n13619 ^ x115 ;
  assign n13656 = n13161 ^ x113 ;
  assign n13657 = n13656 ^ n13209 ;
  assign n13658 = n13657 ^ x112 ;
  assign n13659 = n13658 ^ n13656 ;
  assign n13661 = n13209 ^ x113 ;
  assign n13662 = n13661 ^ n13656 ;
  assign n13663 = ~n13659 & ~n13662 ;
  assign n13664 = n13663 ^ n13656 ;
  assign n13665 = n13277 & ~n13664 ;
  assign n13666 = n13665 ^ n13157 ;
  assign n13649 = n13209 ^ x112 ;
  assign n13650 = n13277 & n13649 ;
  assign n13651 = n13650 ^ n13161 ;
  assign n13643 = n13207 & n13277 ;
  assign n13644 = n13643 ^ n13167 ;
  assign n13636 = n13198 ^ x110 ;
  assign n13637 = n13277 & n13636 ;
  assign n13638 = n13637 ^ n13201 ;
  assign n13621 = n13182 ^ x109 ;
  assign n13622 = n13621 ^ n13192 ;
  assign n13623 = n13622 ^ x108 ;
  assign n13624 = n13623 ^ n13621 ;
  assign n13626 = n13192 ^ x109 ;
  assign n13627 = n13626 ^ n13621 ;
  assign n13628 = ~n13624 & ~n13627 ;
  assign n13629 = n13628 ^ n13621 ;
  assign n13630 = n13277 & ~n13629 ;
  assign n13631 = n13630 ^ n13178 ;
  assign n13596 = n13192 ^ x108 ;
  assign n13597 = n13277 & n13596 ;
  assign n13598 = n13597 ^ n13182 ;
  assign n13151 = n13150 ^ x107 ;
  assign n13278 = n13151 & n13277 ;
  assign n13279 = n13278 ^ n13188 ;
  assign n13280 = n13279 ^ x108 ;
  assign n13285 = n13279 ^ x107 ;
  assign n13281 = n13143 ^ x106 ;
  assign n13282 = n13277 & n13281 ;
  assign n13283 = n13282 ^ n13146 ;
  assign n13284 = n13283 ^ n13279 ;
  assign n13286 = n13285 ^ n13284 ;
  assign n13583 = n13136 ^ x105 ;
  assign n13584 = n13277 & n13583 ;
  assign n13585 = n13584 ^ n13139 ;
  assign n13576 = n13129 ^ x104 ;
  assign n13577 = n13277 & n13576 ;
  assign n13578 = n13577 ^ n13132 ;
  assign n13569 = n13122 ^ x103 ;
  assign n13570 = n13277 & n13569 ;
  assign n13571 = n13570 ^ n13125 ;
  assign n13562 = n13115 ^ x102 ;
  assign n13563 = n13277 & n13562 ;
  assign n13564 = n13563 ^ n13118 ;
  assign n13555 = n13108 ^ x101 ;
  assign n13556 = n13277 & n13555 ;
  assign n13557 = n13556 ^ n13111 ;
  assign n13548 = n13105 ^ x100 ;
  assign n13549 = n13277 & n13548 ;
  assign n13550 = n13549 ^ n12849 ;
  assign n13541 = n13102 ^ x99 ;
  assign n13542 = n13277 & n13541 ;
  assign n13543 = n13542 ^ n12853 ;
  assign n13534 = n13095 ^ x98 ;
  assign n13535 = n13277 & n13534 ;
  assign n13536 = n13535 ^ n13098 ;
  assign n13527 = n13088 ^ x97 ;
  assign n13528 = n13277 & n13527 ;
  assign n13529 = n13528 ^ n13091 ;
  assign n13520 = n13085 ^ x96 ;
  assign n13521 = n13277 & n13520 ;
  assign n13522 = n13521 ^ n12857 ;
  assign n13513 = n13082 ^ x95 ;
  assign n13514 = n13277 & n13513 ;
  assign n13515 = n13514 ^ n12861 ;
  assign n13506 = n13075 ^ x94 ;
  assign n13507 = n13277 & n13506 ;
  assign n13508 = n13507 ^ n13078 ;
  assign n13287 = n13068 ^ x93 ;
  assign n13288 = n13277 & n13287 ;
  assign n13289 = n13288 ^ n13071 ;
  assign n13290 = n13289 ^ x94 ;
  assign n13291 = n13061 ^ x92 ;
  assign n13292 = n13277 & n13291 ;
  assign n13293 = n13292 ^ n13064 ;
  assign n13294 = n13293 ^ x93 ;
  assign n13493 = n13054 ^ x91 ;
  assign n13494 = n13277 & n13493 ;
  assign n13495 = n13494 ^ n13057 ;
  assign n13487 = n13048 & n13277 ;
  assign n13488 = n13487 ^ n13051 ;
  assign n13480 = n13044 ^ x89 ;
  assign n13481 = n13277 & n13480 ;
  assign n13482 = n13481 ^ n12865 ;
  assign n13473 = n13037 ^ x88 ;
  assign n13474 = n13277 & n13473 ;
  assign n13475 = n13474 ^ n13040 ;
  assign n13295 = n13030 ^ x87 ;
  assign n13296 = n13277 & n13295 ;
  assign n13297 = n13296 ^ n13033 ;
  assign n13298 = n13297 ^ x88 ;
  assign n13299 = n13023 ^ x86 ;
  assign n13300 = n13277 & n13299 ;
  assign n13301 = n13300 ^ n13026 ;
  assign n13302 = n13301 ^ x87 ;
  assign n13460 = n13016 ^ x85 ;
  assign n13461 = n13277 & n13460 ;
  assign n13462 = n13461 ^ n13019 ;
  assign n13453 = n13009 ^ x84 ;
  assign n13454 = n13277 & n13453 ;
  assign n13455 = n13454 ^ n13012 ;
  assign n13446 = n13002 ^ x83 ;
  assign n13447 = n13277 & n13446 ;
  assign n13448 = n13447 ^ n13005 ;
  assign n13439 = n12995 ^ x82 ;
  assign n13440 = n13277 & n13439 ;
  assign n13441 = n13440 ^ n12998 ;
  assign n13432 = n12980 ^ x81 ;
  assign n13433 = n13277 & n13432 ;
  assign n13434 = n13433 ^ n12991 ;
  assign n13425 = n12973 ^ x80 ;
  assign n13426 = n13277 & n13425 ;
  assign n13427 = n13426 ^ n12976 ;
  assign n13418 = n12966 ^ x79 ;
  assign n13419 = n13277 & n13418 ;
  assign n13420 = n13419 ^ n12969 ;
  assign n13411 = n12959 ^ x78 ;
  assign n13412 = n13277 & n13411 ;
  assign n13413 = n13412 ^ n12962 ;
  assign n13396 = n12873 ^ x77 ;
  assign n13397 = n13396 ^ n12953 ;
  assign n13398 = n13397 ^ x76 ;
  assign n13399 = n13398 ^ n13396 ;
  assign n13401 = n12953 ^ x77 ;
  assign n13402 = n13401 ^ n13396 ;
  assign n13403 = ~n13399 & ~n13402 ;
  assign n13404 = n13403 ^ n13396 ;
  assign n13405 = n13277 & ~n13404 ;
  assign n13406 = n13405 ^ n12869 ;
  assign n13303 = n12953 ^ x76 ;
  assign n13304 = n13277 & n13303 ;
  assign n13305 = n13304 ^ n12873 ;
  assign n13306 = n13305 ^ x77 ;
  assign n13307 = n12946 ^ x75 ;
  assign n13308 = n13277 & n13307 ;
  assign n13309 = n13308 ^ n12949 ;
  assign n13310 = n13309 ^ x76 ;
  assign n13383 = n12939 ^ x74 ;
  assign n13384 = n13277 & n13383 ;
  assign n13385 = n13384 ^ n12942 ;
  assign n13376 = n12932 ^ x73 ;
  assign n13377 = n13277 & n13376 ;
  assign n13378 = n13377 ^ n12935 ;
  assign n13369 = n12925 ^ x72 ;
  assign n13370 = n13277 & n13369 ;
  assign n13371 = n13370 ^ n12928 ;
  assign n13362 = n12918 ^ x71 ;
  assign n13363 = n13277 & n13362 ;
  assign n13364 = n13363 ^ n12921 ;
  assign n13355 = n12911 ^ x70 ;
  assign n13356 = n13277 & n13355 ;
  assign n13357 = n13356 ^ n12914 ;
  assign n13348 = n12905 ^ x69 ;
  assign n13349 = n13277 & n13348 ;
  assign n13350 = n13349 ^ n12907 ;
  assign n13341 = n12899 ^ x68 ;
  assign n13342 = n13277 & n13341 ;
  assign n13343 = n13342 ^ n12901 ;
  assign n13334 = n12893 ^ x67 ;
  assign n13335 = n13277 & n13334 ;
  assign n13336 = n13335 ^ n12895 ;
  assign n13327 = n12890 ^ x66 ;
  assign n13328 = n13277 & n13327 ;
  assign n13329 = n13328 ^ n12883 ;
  assign n13312 = n12886 & n13277 ;
  assign n13311 = n12881 ^ x7 ;
  assign n13313 = n13312 ^ n13311 ;
  assign n13314 = n13313 ^ x66 ;
  assign n13317 = ~x5 & x64 ;
  assign n13315 = x64 & n13277 ;
  assign n13320 = n13317 ^ n13315 ;
  assign n13321 = ~x65 & ~n13320 ;
  assign n13318 = n13317 ^ x65 ;
  assign n13319 = x6 & n13318 ;
  assign n13322 = n13321 ^ n13319 ;
  assign n13316 = x5 & n13315 ;
  assign n13323 = n13322 ^ n13316 ;
  assign n13324 = n13323 ^ n13313 ;
  assign n13325 = ~n13314 & ~n13324 ;
  assign n13326 = n13325 ^ x66 ;
  assign n13330 = n13329 ^ n13326 ;
  assign n13331 = n13329 ^ x67 ;
  assign n13332 = n13330 & ~n13331 ;
  assign n13333 = n13332 ^ x67 ;
  assign n13337 = n13336 ^ n13333 ;
  assign n13338 = n13336 ^ x68 ;
  assign n13339 = n13337 & ~n13338 ;
  assign n13340 = n13339 ^ x68 ;
  assign n13344 = n13343 ^ n13340 ;
  assign n13345 = n13343 ^ x69 ;
  assign n13346 = n13344 & ~n13345 ;
  assign n13347 = n13346 ^ x69 ;
  assign n13351 = n13350 ^ n13347 ;
  assign n13352 = n13350 ^ x70 ;
  assign n13353 = n13351 & ~n13352 ;
  assign n13354 = n13353 ^ x70 ;
  assign n13358 = n13357 ^ n13354 ;
  assign n13359 = n13357 ^ x71 ;
  assign n13360 = n13358 & ~n13359 ;
  assign n13361 = n13360 ^ x71 ;
  assign n13365 = n13364 ^ n13361 ;
  assign n13366 = n13364 ^ x72 ;
  assign n13367 = n13365 & ~n13366 ;
  assign n13368 = n13367 ^ x72 ;
  assign n13372 = n13371 ^ n13368 ;
  assign n13373 = n13371 ^ x73 ;
  assign n13374 = n13372 & ~n13373 ;
  assign n13375 = n13374 ^ x73 ;
  assign n13379 = n13378 ^ n13375 ;
  assign n13380 = n13378 ^ x74 ;
  assign n13381 = n13379 & ~n13380 ;
  assign n13382 = n13381 ^ x74 ;
  assign n13386 = n13385 ^ n13382 ;
  assign n13387 = n13385 ^ x75 ;
  assign n13388 = n13386 & ~n13387 ;
  assign n13389 = n13388 ^ x75 ;
  assign n13390 = n13389 ^ n13309 ;
  assign n13391 = ~n13310 & n13390 ;
  assign n13392 = n13391 ^ x76 ;
  assign n13393 = n13392 ^ n13305 ;
  assign n13394 = ~n13306 & n13393 ;
  assign n13395 = n13394 ^ x77 ;
  assign n13407 = n13406 ^ n13395 ;
  assign n13408 = n13406 ^ x78 ;
  assign n13409 = n13407 & ~n13408 ;
  assign n13410 = n13409 ^ x78 ;
  assign n13414 = n13413 ^ n13410 ;
  assign n13415 = n13413 ^ x79 ;
  assign n13416 = n13414 & ~n13415 ;
  assign n13417 = n13416 ^ x79 ;
  assign n13421 = n13420 ^ n13417 ;
  assign n13422 = n13420 ^ x80 ;
  assign n13423 = n13421 & ~n13422 ;
  assign n13424 = n13423 ^ x80 ;
  assign n13428 = n13427 ^ n13424 ;
  assign n13429 = n13427 ^ x81 ;
  assign n13430 = n13428 & ~n13429 ;
  assign n13431 = n13430 ^ x81 ;
  assign n13435 = n13434 ^ n13431 ;
  assign n13436 = n13434 ^ x82 ;
  assign n13437 = n13435 & ~n13436 ;
  assign n13438 = n13437 ^ x82 ;
  assign n13442 = n13441 ^ n13438 ;
  assign n13443 = n13441 ^ x83 ;
  assign n13444 = n13442 & ~n13443 ;
  assign n13445 = n13444 ^ x83 ;
  assign n13449 = n13448 ^ n13445 ;
  assign n13450 = n13448 ^ x84 ;
  assign n13451 = n13449 & ~n13450 ;
  assign n13452 = n13451 ^ x84 ;
  assign n13456 = n13455 ^ n13452 ;
  assign n13457 = n13455 ^ x85 ;
  assign n13458 = n13456 & ~n13457 ;
  assign n13459 = n13458 ^ x85 ;
  assign n13463 = n13462 ^ n13459 ;
  assign n13464 = n13462 ^ x86 ;
  assign n13465 = n13463 & ~n13464 ;
  assign n13466 = n13465 ^ x86 ;
  assign n13467 = n13466 ^ n13301 ;
  assign n13468 = ~n13302 & n13467 ;
  assign n13469 = n13468 ^ x87 ;
  assign n13470 = n13469 ^ n13297 ;
  assign n13471 = ~n13298 & n13470 ;
  assign n13472 = n13471 ^ x88 ;
  assign n13476 = n13475 ^ n13472 ;
  assign n13477 = n13475 ^ x89 ;
  assign n13478 = n13476 & ~n13477 ;
  assign n13479 = n13478 ^ x89 ;
  assign n13483 = n13482 ^ n13479 ;
  assign n13484 = n13482 ^ x90 ;
  assign n13485 = n13483 & ~n13484 ;
  assign n13486 = n13485 ^ x90 ;
  assign n13489 = n13488 ^ n13486 ;
  assign n13490 = n13488 ^ x91 ;
  assign n13491 = n13489 & ~n13490 ;
  assign n13492 = n13491 ^ x91 ;
  assign n13496 = n13495 ^ n13492 ;
  assign n13497 = n13495 ^ x92 ;
  assign n13498 = n13496 & ~n13497 ;
  assign n13499 = n13498 ^ x92 ;
  assign n13500 = n13499 ^ n13293 ;
  assign n13501 = ~n13294 & n13500 ;
  assign n13502 = n13501 ^ x93 ;
  assign n13503 = n13502 ^ n13289 ;
  assign n13504 = ~n13290 & n13503 ;
  assign n13505 = n13504 ^ x94 ;
  assign n13509 = n13508 ^ n13505 ;
  assign n13510 = n13508 ^ x95 ;
  assign n13511 = n13509 & ~n13510 ;
  assign n13512 = n13511 ^ x95 ;
  assign n13516 = n13515 ^ n13512 ;
  assign n13517 = n13515 ^ x96 ;
  assign n13518 = n13516 & ~n13517 ;
  assign n13519 = n13518 ^ x96 ;
  assign n13523 = n13522 ^ n13519 ;
  assign n13524 = n13522 ^ x97 ;
  assign n13525 = n13523 & ~n13524 ;
  assign n13526 = n13525 ^ x97 ;
  assign n13530 = n13529 ^ n13526 ;
  assign n13531 = n13529 ^ x98 ;
  assign n13532 = n13530 & ~n13531 ;
  assign n13533 = n13532 ^ x98 ;
  assign n13537 = n13536 ^ n13533 ;
  assign n13538 = n13536 ^ x99 ;
  assign n13539 = n13537 & ~n13538 ;
  assign n13540 = n13539 ^ x99 ;
  assign n13544 = n13543 ^ n13540 ;
  assign n13545 = n13543 ^ x100 ;
  assign n13546 = n13544 & ~n13545 ;
  assign n13547 = n13546 ^ x100 ;
  assign n13551 = n13550 ^ n13547 ;
  assign n13552 = n13550 ^ x101 ;
  assign n13553 = n13551 & ~n13552 ;
  assign n13554 = n13553 ^ x101 ;
  assign n13558 = n13557 ^ n13554 ;
  assign n13559 = n13557 ^ x102 ;
  assign n13560 = n13558 & ~n13559 ;
  assign n13561 = n13560 ^ x102 ;
  assign n13565 = n13564 ^ n13561 ;
  assign n13566 = n13564 ^ x103 ;
  assign n13567 = n13565 & ~n13566 ;
  assign n13568 = n13567 ^ x103 ;
  assign n13572 = n13571 ^ n13568 ;
  assign n13573 = n13571 ^ x104 ;
  assign n13574 = n13572 & ~n13573 ;
  assign n13575 = n13574 ^ x104 ;
  assign n13579 = n13578 ^ n13575 ;
  assign n13580 = n13578 ^ x105 ;
  assign n13581 = n13579 & ~n13580 ;
  assign n13582 = n13581 ^ x105 ;
  assign n13586 = n13585 ^ n13582 ;
  assign n13587 = n13585 ^ x106 ;
  assign n13588 = n13586 & ~n13587 ;
  assign n13589 = n13588 ^ x106 ;
  assign n13590 = n13589 ^ n13279 ;
  assign n13591 = n13590 ^ n13285 ;
  assign n13592 = ~n13286 & n13591 ;
  assign n13593 = n13592 ^ n13285 ;
  assign n13594 = ~n13280 & n13593 ;
  assign n13595 = n13594 ^ x108 ;
  assign n13599 = n13598 ^ n13595 ;
  assign n13600 = n13598 ^ x109 ;
  assign n13601 = n13599 & ~n13600 ;
  assign n13602 = n13601 ^ x109 ;
  assign n13632 = n13631 ^ n13602 ;
  assign n13633 = n13631 ^ x110 ;
  assign n13634 = n13632 & ~n13633 ;
  assign n13635 = n13634 ^ x110 ;
  assign n13639 = n13638 ^ n13635 ;
  assign n13640 = n13638 ^ x111 ;
  assign n13641 = n13639 & ~n13640 ;
  assign n13642 = n13641 ^ x111 ;
  assign n13645 = n13644 ^ n13642 ;
  assign n13646 = n13644 ^ x112 ;
  assign n13647 = n13645 & ~n13646 ;
  assign n13648 = n13647 ^ x112 ;
  assign n13652 = n13651 ^ n13648 ;
  assign n13653 = n13651 ^ x113 ;
  assign n13654 = n13652 & ~n13653 ;
  assign n13655 = n13654 ^ x113 ;
  assign n13667 = n13666 ^ n13655 ;
  assign n13668 = n13666 ^ x114 ;
  assign n13669 = n13667 & ~n13668 ;
  assign n13670 = n13669 ^ x114 ;
  assign n13671 = n13670 ^ n13619 ;
  assign n13672 = ~n13620 & n13671 ;
  assign n13673 = n13672 ^ x115 ;
  assign n13677 = n13676 ^ n13673 ;
  assign n13678 = n13676 ^ x116 ;
  assign n13679 = n13677 & ~n13678 ;
  assign n13680 = n13679 ^ x116 ;
  assign n13684 = n13683 ^ n13680 ;
  assign n13685 = n13683 ^ x117 ;
  assign n13686 = n13684 & ~n13685 ;
  assign n13687 = n13686 ^ x117 ;
  assign n13688 = n13687 ^ n13615 ;
  assign n13689 = ~n13616 & n13688 ;
  assign n13690 = n13689 ^ x118 ;
  assign n13691 = n13690 ^ n13611 ;
  assign n13692 = ~n13612 & n13691 ;
  assign n13693 = n13692 ^ x119 ;
  assign n13694 = n13693 ^ n13607 ;
  assign n13695 = ~n13608 & n13694 ;
  assign n13696 = n13695 ^ x120 ;
  assign n13700 = n13699 ^ n13696 ;
  assign n13701 = n13699 ^ x121 ;
  assign n13702 = n13700 & ~n13701 ;
  assign n13703 = n13702 ^ x121 ;
  assign n14066 = n14065 ^ n13703 ;
  assign n14073 = ~n134 & n11950 ;
  assign n14067 = n14066 ^ n134 ;
  assign n14068 = n14067 ^ n133 ;
  assign n14074 = n14073 ^ n14068 ;
  assign n14075 = ~n14065 & n14074 ;
  assign n14076 = n14075 ^ n14068 ;
  assign n14077 = n14076 ^ n13703 ;
  assign n14078 = ~n14075 & n14077 ;
  assign n14079 = ~n14066 & n14078 ;
  assign n14080 = n14079 ^ n14076 ;
  assign n14081 = n14080 ^ x123 ;
  assign n13604 = n134 & n12835 ;
  assign n13704 = n133 & ~n13703 ;
  assign n13705 = x122 & ~n12832 ;
  assign n13706 = n13704 & n13705 ;
  assign n13707 = n13706 ^ n13704 ;
  assign n13708 = ~n13273 & ~n13707 ;
  assign n13709 = n13604 & n13708 ;
  assign n13710 = n13709 ^ n13707 ;
  assign n14152 = n13696 ^ x121 ;
  assign n14153 = n13710 & n14152 ;
  assign n14154 = n14153 ^ n13699 ;
  assign n14145 = n13693 ^ x120 ;
  assign n14146 = n13710 & n14145 ;
  assign n14147 = n14146 ^ n13607 ;
  assign n14138 = n13690 ^ x119 ;
  assign n14139 = n13710 & n14138 ;
  assign n14140 = n14139 ^ n13611 ;
  assign n14131 = n13687 ^ x118 ;
  assign n14132 = n13710 & n14131 ;
  assign n14133 = n14132 ^ n13615 ;
  assign n14124 = n13680 ^ x117 ;
  assign n14125 = n13710 & n14124 ;
  assign n14126 = n14125 ^ n13683 ;
  assign n14117 = n13673 ^ x116 ;
  assign n14118 = n13710 & n14117 ;
  assign n14119 = n14118 ^ n13676 ;
  assign n14110 = n13670 ^ x115 ;
  assign n14111 = n13710 & n14110 ;
  assign n14112 = n14111 ^ n13619 ;
  assign n14082 = n13655 ^ x114 ;
  assign n14083 = n13710 & n14082 ;
  assign n14084 = n14083 ^ n13666 ;
  assign n14085 = n14084 ^ x115 ;
  assign n14086 = n13648 ^ x113 ;
  assign n14087 = n13710 & n14086 ;
  assign n14088 = n14087 ^ n13651 ;
  assign n14089 = n14088 ^ x114 ;
  assign n14097 = n13642 ^ x112 ;
  assign n14098 = n13710 & n14097 ;
  assign n14099 = n14098 ^ n13644 ;
  assign n14090 = n13635 ^ x111 ;
  assign n14091 = n13710 & n14090 ;
  assign n14092 = n14091 ^ n13638 ;
  assign n14052 = n13595 ^ x109 ;
  assign n14053 = n13710 & n14052 ;
  assign n14054 = n14053 ^ n13598 ;
  assign n13713 = n13283 ^ x108 ;
  assign n13714 = n13713 ^ x107 ;
  assign n13715 = n13714 ^ n13589 ;
  assign n13716 = n13715 ^ n13713 ;
  assign n13719 = n13713 ^ n12315 ;
  assign n13720 = ~n13716 & ~n13719 ;
  assign n13721 = n13720 ^ n13713 ;
  assign n13722 = n13710 & ~n13721 ;
  assign n13723 = n13722 ^ n13279 ;
  assign n13724 = n13723 ^ x109 ;
  assign n13729 = n13723 ^ x108 ;
  assign n13725 = n13589 ^ x107 ;
  assign n13726 = n13710 & n13725 ;
  assign n13727 = n13726 ^ n13283 ;
  assign n13728 = n13727 ^ n13723 ;
  assign n13730 = n13729 ^ n13728 ;
  assign n14039 = n13582 ^ x106 ;
  assign n14040 = n13710 & n14039 ;
  assign n14041 = n14040 ^ n13585 ;
  assign n14032 = n13575 ^ x105 ;
  assign n14033 = n13710 & n14032 ;
  assign n14034 = n14033 ^ n13578 ;
  assign n14025 = n13568 ^ x104 ;
  assign n14026 = n13710 & n14025 ;
  assign n14027 = n14026 ^ n13571 ;
  assign n14018 = n13561 ^ x103 ;
  assign n14019 = n13710 & n14018 ;
  assign n14020 = n14019 ^ n13564 ;
  assign n14011 = n13554 ^ x102 ;
  assign n14012 = n13710 & n14011 ;
  assign n14013 = n14012 ^ n13557 ;
  assign n14004 = n13547 ^ x101 ;
  assign n14005 = n13710 & n14004 ;
  assign n14006 = n14005 ^ n13550 ;
  assign n13731 = n13540 ^ x100 ;
  assign n13732 = n13710 & n13731 ;
  assign n13733 = n13732 ^ n13543 ;
  assign n13734 = n13733 ^ x101 ;
  assign n13735 = n13533 ^ x99 ;
  assign n13736 = n13710 & n13735 ;
  assign n13737 = n13736 ^ n13536 ;
  assign n13738 = n13737 ^ x100 ;
  assign n13991 = n13526 ^ x98 ;
  assign n13992 = n13710 & n13991 ;
  assign n13993 = n13992 ^ n13529 ;
  assign n13984 = n13519 ^ x97 ;
  assign n13985 = n13710 & n13984 ;
  assign n13986 = n13985 ^ n13522 ;
  assign n13977 = n13512 ^ x96 ;
  assign n13978 = n13710 & n13977 ;
  assign n13979 = n13978 ^ n13515 ;
  assign n13970 = n13505 ^ x95 ;
  assign n13971 = n13710 & n13970 ;
  assign n13972 = n13971 ^ n13508 ;
  assign n13963 = n13502 ^ x94 ;
  assign n13964 = n13710 & n13963 ;
  assign n13965 = n13964 ^ n13289 ;
  assign n13952 = n13492 ^ x92 ;
  assign n13953 = n13710 & n13952 ;
  assign n13954 = n13953 ^ n13495 ;
  assign n13742 = n13486 ^ x91 ;
  assign n13743 = n13710 & n13742 ;
  assign n13744 = n13743 ^ n13488 ;
  assign n13745 = n13744 ^ x92 ;
  assign n13750 = n13744 ^ x91 ;
  assign n13746 = n13479 ^ x90 ;
  assign n13747 = n13710 & n13746 ;
  assign n13748 = n13747 ^ n13482 ;
  assign n13749 = n13748 ^ n13744 ;
  assign n13751 = n13750 ^ n13749 ;
  assign n13939 = n13472 ^ x89 ;
  assign n13940 = n13710 & n13939 ;
  assign n13941 = n13940 ^ n13475 ;
  assign n13932 = n13469 ^ x88 ;
  assign n13933 = n13710 & n13932 ;
  assign n13934 = n13933 ^ n13297 ;
  assign n13925 = n13466 ^ x87 ;
  assign n13926 = n13710 & n13925 ;
  assign n13927 = n13926 ^ n13301 ;
  assign n13918 = n13459 ^ x86 ;
  assign n13919 = n13710 & n13918 ;
  assign n13920 = n13919 ^ n13462 ;
  assign n13911 = n13452 ^ x85 ;
  assign n13912 = n13710 & n13911 ;
  assign n13913 = n13912 ^ n13455 ;
  assign n13752 = n13445 ^ x84 ;
  assign n13753 = n13710 & n13752 ;
  assign n13754 = n13753 ^ n13448 ;
  assign n13755 = n13754 ^ x85 ;
  assign n13760 = n13754 ^ x84 ;
  assign n13756 = n13438 ^ x83 ;
  assign n13757 = n13710 & n13756 ;
  assign n13758 = n13757 ^ n13441 ;
  assign n13759 = n13758 ^ n13754 ;
  assign n13761 = n13760 ^ n13759 ;
  assign n13762 = n13431 ^ x82 ;
  assign n13763 = n13710 & n13762 ;
  assign n13764 = n13763 ^ n13434 ;
  assign n13765 = n13764 ^ x83 ;
  assign n13770 = n13764 ^ x82 ;
  assign n13766 = n13424 ^ x81 ;
  assign n13767 = n13710 & n13766 ;
  assign n13768 = n13767 ^ n13427 ;
  assign n13769 = n13768 ^ n13764 ;
  assign n13771 = n13770 ^ n13769 ;
  assign n13772 = n13417 ^ x80 ;
  assign n13773 = n13710 & n13772 ;
  assign n13774 = n13773 ^ n13420 ;
  assign n13775 = n13774 ^ x81 ;
  assign n13776 = n13410 ^ x79 ;
  assign n13777 = n13710 & n13776 ;
  assign n13778 = n13777 ^ n13413 ;
  assign n13779 = n13778 ^ x80 ;
  assign n13886 = n13395 ^ x78 ;
  assign n13887 = n13710 & n13886 ;
  assign n13888 = n13887 ^ n13406 ;
  assign n13879 = n13392 ^ x77 ;
  assign n13880 = n13710 & n13879 ;
  assign n13881 = n13880 ^ n13305 ;
  assign n13872 = n13389 ^ x76 ;
  assign n13873 = n13710 & n13872 ;
  assign n13874 = n13873 ^ n13309 ;
  assign n13865 = n13382 ^ x75 ;
  assign n13866 = n13710 & n13865 ;
  assign n13867 = n13866 ^ n13385 ;
  assign n13858 = n13375 ^ x74 ;
  assign n13859 = n13710 & n13858 ;
  assign n13860 = n13859 ^ n13378 ;
  assign n13780 = n13368 ^ x73 ;
  assign n13781 = n13710 & n13780 ;
  assign n13782 = n13781 ^ n13371 ;
  assign n13783 = n13782 ^ x74 ;
  assign n13784 = n13361 ^ x72 ;
  assign n13785 = n13710 & n13784 ;
  assign n13786 = n13785 ^ n13364 ;
  assign n13787 = n13786 ^ x73 ;
  assign n13845 = n13354 ^ x71 ;
  assign n13846 = n13710 & n13845 ;
  assign n13847 = n13846 ^ n13357 ;
  assign n13838 = n13347 ^ x70 ;
  assign n13839 = n13710 & n13838 ;
  assign n13840 = n13839 ^ n13350 ;
  assign n13831 = n13340 ^ x69 ;
  assign n13832 = n13710 & n13831 ;
  assign n13833 = n13832 ^ n13343 ;
  assign n13824 = n13333 ^ x68 ;
  assign n13825 = n13710 & n13824 ;
  assign n13826 = n13825 ^ n13336 ;
  assign n13817 = n13326 ^ x67 ;
  assign n13818 = n13710 & n13817 ;
  assign n13819 = n13818 ^ n13329 ;
  assign n13810 = n13323 ^ x66 ;
  assign n13811 = n13710 & ~n13810 ;
  assign n13812 = n13811 ^ n13313 ;
  assign n13790 = n13710 ^ n13277 ;
  assign n13791 = n13317 & n13790 ;
  assign n13789 = n13316 ^ x6 ;
  assign n13792 = n13791 ^ n13789 ;
  assign n13788 = x65 & n13710 ;
  assign n13793 = n13792 ^ n13788 ;
  assign n13794 = n13793 ^ x66 ;
  assign n13796 = x65 ^ x4 ;
  assign n13797 = x64 ^ x5 ;
  assign n13798 = n13797 ^ x65 ;
  assign n13799 = n13798 ^ n13710 ;
  assign n13800 = ~n13796 & n13799 ;
  assign n13795 = x5 & x65 ;
  assign n13801 = n13800 ^ n13795 ;
  assign n13804 = x64 & n13801 ;
  assign n13805 = n13804 ^ n13795 ;
  assign n13806 = n13805 ^ x65 ;
  assign n13807 = n13806 ^ n13793 ;
  assign n13808 = ~n13794 & n13807 ;
  assign n13809 = n13808 ^ x66 ;
  assign n13813 = n13812 ^ n13809 ;
  assign n13814 = n13812 ^ x67 ;
  assign n13815 = n13813 & ~n13814 ;
  assign n13816 = n13815 ^ x67 ;
  assign n13820 = n13819 ^ n13816 ;
  assign n13821 = n13819 ^ x68 ;
  assign n13822 = n13820 & ~n13821 ;
  assign n13823 = n13822 ^ x68 ;
  assign n13827 = n13826 ^ n13823 ;
  assign n13828 = n13826 ^ x69 ;
  assign n13829 = n13827 & ~n13828 ;
  assign n13830 = n13829 ^ x69 ;
  assign n13834 = n13833 ^ n13830 ;
  assign n13835 = n13833 ^ x70 ;
  assign n13836 = n13834 & ~n13835 ;
  assign n13837 = n13836 ^ x70 ;
  assign n13841 = n13840 ^ n13837 ;
  assign n13842 = n13840 ^ x71 ;
  assign n13843 = n13841 & ~n13842 ;
  assign n13844 = n13843 ^ x71 ;
  assign n13848 = n13847 ^ n13844 ;
  assign n13849 = n13847 ^ x72 ;
  assign n13850 = n13848 & ~n13849 ;
  assign n13851 = n13850 ^ x72 ;
  assign n13852 = n13851 ^ n13786 ;
  assign n13853 = ~n13787 & n13852 ;
  assign n13854 = n13853 ^ x73 ;
  assign n13855 = n13854 ^ n13782 ;
  assign n13856 = ~n13783 & n13855 ;
  assign n13857 = n13856 ^ x74 ;
  assign n13861 = n13860 ^ n13857 ;
  assign n13862 = n13860 ^ x75 ;
  assign n13863 = n13861 & ~n13862 ;
  assign n13864 = n13863 ^ x75 ;
  assign n13868 = n13867 ^ n13864 ;
  assign n13869 = n13867 ^ x76 ;
  assign n13870 = n13868 & ~n13869 ;
  assign n13871 = n13870 ^ x76 ;
  assign n13875 = n13874 ^ n13871 ;
  assign n13876 = n13874 ^ x77 ;
  assign n13877 = n13875 & ~n13876 ;
  assign n13878 = n13877 ^ x77 ;
  assign n13882 = n13881 ^ n13878 ;
  assign n13883 = n13881 ^ x78 ;
  assign n13884 = n13882 & ~n13883 ;
  assign n13885 = n13884 ^ x78 ;
  assign n13889 = n13888 ^ n13885 ;
  assign n13890 = n13888 ^ x79 ;
  assign n13891 = n13889 & ~n13890 ;
  assign n13892 = n13891 ^ x79 ;
  assign n13893 = n13892 ^ n13778 ;
  assign n13894 = ~n13779 & n13893 ;
  assign n13895 = n13894 ^ x80 ;
  assign n13896 = n13895 ^ n13774 ;
  assign n13897 = ~n13775 & n13896 ;
  assign n13898 = n13897 ^ x81 ;
  assign n13899 = n13898 ^ n13764 ;
  assign n13900 = n13899 ^ n13770 ;
  assign n13901 = ~n13771 & n13900 ;
  assign n13902 = n13901 ^ n13770 ;
  assign n13903 = ~n13765 & n13902 ;
  assign n13904 = n13903 ^ x83 ;
  assign n13905 = n13904 ^ n13754 ;
  assign n13906 = n13905 ^ n13760 ;
  assign n13907 = ~n13761 & n13906 ;
  assign n13908 = n13907 ^ n13760 ;
  assign n13909 = ~n13755 & n13908 ;
  assign n13910 = n13909 ^ x85 ;
  assign n13914 = n13913 ^ n13910 ;
  assign n13915 = n13913 ^ x86 ;
  assign n13916 = n13914 & ~n13915 ;
  assign n13917 = n13916 ^ x86 ;
  assign n13921 = n13920 ^ n13917 ;
  assign n13922 = n13920 ^ x87 ;
  assign n13923 = n13921 & ~n13922 ;
  assign n13924 = n13923 ^ x87 ;
  assign n13928 = n13927 ^ n13924 ;
  assign n13929 = n13927 ^ x88 ;
  assign n13930 = n13928 & ~n13929 ;
  assign n13931 = n13930 ^ x88 ;
  assign n13935 = n13934 ^ n13931 ;
  assign n13936 = n13934 ^ x89 ;
  assign n13937 = n13935 & ~n13936 ;
  assign n13938 = n13937 ^ x89 ;
  assign n13942 = n13941 ^ n13938 ;
  assign n13943 = n13941 ^ x90 ;
  assign n13944 = n13942 & ~n13943 ;
  assign n13945 = n13944 ^ x90 ;
  assign n13946 = n13945 ^ n13744 ;
  assign n13947 = n13946 ^ n13750 ;
  assign n13948 = ~n13751 & n13947 ;
  assign n13949 = n13948 ^ n13750 ;
  assign n13950 = ~n13745 & n13949 ;
  assign n13951 = n13950 ^ x92 ;
  assign n13955 = n13954 ^ n13951 ;
  assign n13956 = n13954 ^ x93 ;
  assign n13957 = n13955 & ~n13956 ;
  assign n13958 = n13957 ^ x93 ;
  assign n13739 = n13499 ^ x93 ;
  assign n13740 = n13710 & n13739 ;
  assign n13741 = n13740 ^ n13293 ;
  assign n13959 = n13958 ^ n13741 ;
  assign n13960 = n13958 ^ x94 ;
  assign n13961 = n13959 & n13960 ;
  assign n13962 = n13961 ^ x94 ;
  assign n13966 = n13965 ^ n13962 ;
  assign n13967 = n13965 ^ x95 ;
  assign n13968 = n13966 & ~n13967 ;
  assign n13969 = n13968 ^ x95 ;
  assign n13973 = n13972 ^ n13969 ;
  assign n13974 = n13972 ^ x96 ;
  assign n13975 = n13973 & ~n13974 ;
  assign n13976 = n13975 ^ x96 ;
  assign n13980 = n13979 ^ n13976 ;
  assign n13981 = n13979 ^ x97 ;
  assign n13982 = n13980 & ~n13981 ;
  assign n13983 = n13982 ^ x97 ;
  assign n13987 = n13986 ^ n13983 ;
  assign n13988 = n13986 ^ x98 ;
  assign n13989 = n13987 & ~n13988 ;
  assign n13990 = n13989 ^ x98 ;
  assign n13994 = n13993 ^ n13990 ;
  assign n13995 = n13993 ^ x99 ;
  assign n13996 = n13994 & ~n13995 ;
  assign n13997 = n13996 ^ x99 ;
  assign n13998 = n13997 ^ n13737 ;
  assign n13999 = ~n13738 & n13998 ;
  assign n14000 = n13999 ^ x100 ;
  assign n14001 = n14000 ^ n13733 ;
  assign n14002 = ~n13734 & n14001 ;
  assign n14003 = n14002 ^ x101 ;
  assign n14007 = n14006 ^ n14003 ;
  assign n14008 = n14006 ^ x102 ;
  assign n14009 = n14007 & ~n14008 ;
  assign n14010 = n14009 ^ x102 ;
  assign n14014 = n14013 ^ n14010 ;
  assign n14015 = n14013 ^ x103 ;
  assign n14016 = n14014 & ~n14015 ;
  assign n14017 = n14016 ^ x103 ;
  assign n14021 = n14020 ^ n14017 ;
  assign n14022 = n14020 ^ x104 ;
  assign n14023 = n14021 & ~n14022 ;
  assign n14024 = n14023 ^ x104 ;
  assign n14028 = n14027 ^ n14024 ;
  assign n14029 = n14027 ^ x105 ;
  assign n14030 = n14028 & ~n14029 ;
  assign n14031 = n14030 ^ x105 ;
  assign n14035 = n14034 ^ n14031 ;
  assign n14036 = n14034 ^ x106 ;
  assign n14037 = n14035 & ~n14036 ;
  assign n14038 = n14037 ^ x106 ;
  assign n14042 = n14041 ^ n14038 ;
  assign n14043 = n14041 ^ x107 ;
  assign n14044 = n14042 & ~n14043 ;
  assign n14045 = n14044 ^ x107 ;
  assign n14046 = n14045 ^ n13723 ;
  assign n14047 = n14046 ^ n13729 ;
  assign n14048 = ~n13730 & n14047 ;
  assign n14049 = n14048 ^ n13729 ;
  assign n14050 = ~n13724 & n14049 ;
  assign n14051 = n14050 ^ x109 ;
  assign n14055 = n14054 ^ n14051 ;
  assign n14056 = n14054 ^ x110 ;
  assign n14057 = n14055 & ~n14056 ;
  assign n14058 = n14057 ^ x110 ;
  assign n13603 = n13602 ^ x110 ;
  assign n13711 = n13603 & n13710 ;
  assign n13712 = n13711 ^ n13631 ;
  assign n14059 = n14058 ^ n13712 ;
  assign n14060 = n14058 ^ x111 ;
  assign n14061 = n14059 & n14060 ;
  assign n14062 = n14061 ^ x111 ;
  assign n14093 = n14092 ^ n14062 ;
  assign n14094 = n14092 ^ x112 ;
  assign n14095 = n14093 & ~n14094 ;
  assign n14096 = n14095 ^ x112 ;
  assign n14100 = n14099 ^ n14096 ;
  assign n14101 = n14099 ^ x113 ;
  assign n14102 = n14100 & ~n14101 ;
  assign n14103 = n14102 ^ x113 ;
  assign n14104 = n14103 ^ n14088 ;
  assign n14105 = ~n14089 & n14104 ;
  assign n14106 = n14105 ^ x114 ;
  assign n14107 = n14106 ^ n14084 ;
  assign n14108 = ~n14085 & n14107 ;
  assign n14109 = n14108 ^ x115 ;
  assign n14113 = n14112 ^ n14109 ;
  assign n14114 = n14112 ^ x116 ;
  assign n14115 = n14113 & ~n14114 ;
  assign n14116 = n14115 ^ x116 ;
  assign n14120 = n14119 ^ n14116 ;
  assign n14121 = n14119 ^ x117 ;
  assign n14122 = n14120 & ~n14121 ;
  assign n14123 = n14122 ^ x117 ;
  assign n14127 = n14126 ^ n14123 ;
  assign n14128 = n14126 ^ x118 ;
  assign n14129 = n14127 & ~n14128 ;
  assign n14130 = n14129 ^ x118 ;
  assign n14134 = n14133 ^ n14130 ;
  assign n14135 = n14133 ^ x119 ;
  assign n14136 = n14134 & ~n14135 ;
  assign n14137 = n14136 ^ x119 ;
  assign n14141 = n14140 ^ n14137 ;
  assign n14142 = n14140 ^ x120 ;
  assign n14143 = n14141 & ~n14142 ;
  assign n14144 = n14143 ^ x120 ;
  assign n14148 = n14147 ^ n14144 ;
  assign n14149 = n14147 ^ x121 ;
  assign n14150 = n14148 & ~n14149 ;
  assign n14151 = n14150 ^ x121 ;
  assign n14155 = n14154 ^ n14151 ;
  assign n14618 = n14151 ^ x122 ;
  assign n14159 = n14155 & n14618 ;
  assign n14156 = x123 ^ x122 ;
  assign n14160 = n14159 ^ n14156 ;
  assign n14163 = ~n14081 & n14160 ;
  assign n14164 = n14163 ^ x123 ;
  assign n14165 = n132 & ~n14164 ;
  assign n14619 = n14165 & n14618 ;
  assign n14620 = n14619 ^ n14154 ;
  assign n14611 = n14144 ^ x121 ;
  assign n14612 = n14165 & n14611 ;
  assign n14613 = n14612 ^ n14147 ;
  assign n14604 = n14137 ^ x120 ;
  assign n14605 = n14165 & n14604 ;
  assign n14606 = n14605 ^ n14140 ;
  assign n14597 = n14130 ^ x119 ;
  assign n14598 = n14165 & n14597 ;
  assign n14599 = n14598 ^ n14133 ;
  assign n14590 = n14123 ^ x118 ;
  assign n14591 = n14165 & n14590 ;
  assign n14592 = n14591 ^ n14126 ;
  assign n14583 = n14116 ^ x117 ;
  assign n14584 = n14165 & n14583 ;
  assign n14585 = n14584 ^ n14119 ;
  assign n14576 = n14109 ^ x116 ;
  assign n14577 = n14165 & n14576 ;
  assign n14578 = n14577 ^ n14112 ;
  assign n14569 = n14106 ^ x115 ;
  assign n14570 = n14165 & n14569 ;
  assign n14571 = n14570 ^ n14084 ;
  assign n14562 = n14103 ^ x114 ;
  assign n14563 = n14165 & n14562 ;
  assign n14564 = n14563 ^ n14088 ;
  assign n14555 = n14096 ^ x113 ;
  assign n14556 = n14165 & n14555 ;
  assign n14557 = n14556 ^ n14099 ;
  assign n14063 = n14062 ^ x112 ;
  assign n14166 = n14063 & n14165 ;
  assign n14167 = n14166 ^ n14092 ;
  assign n14168 = n14167 ^ x113 ;
  assign n14169 = n14060 & n14165 ;
  assign n14170 = n14169 ^ n13712 ;
  assign n14171 = n14170 ^ x112 ;
  assign n14542 = n14051 ^ x110 ;
  assign n14543 = n14165 & n14542 ;
  assign n14544 = n14543 ^ n14054 ;
  assign n14527 = n13727 ^ x109 ;
  assign n14528 = n14527 ^ n14045 ;
  assign n14529 = n14528 ^ x108 ;
  assign n14530 = n14529 ^ n14527 ;
  assign n14532 = n14045 ^ x109 ;
  assign n14533 = n14532 ^ n14527 ;
  assign n14534 = ~n14530 & ~n14533 ;
  assign n14535 = n14534 ^ n14527 ;
  assign n14536 = n14165 & ~n14535 ;
  assign n14537 = n14536 ^ n13723 ;
  assign n14520 = n14045 ^ x108 ;
  assign n14521 = n14165 & n14520 ;
  assign n14522 = n14521 ^ n13727 ;
  assign n14513 = n14038 ^ x107 ;
  assign n14514 = n14165 & n14513 ;
  assign n14515 = n14514 ^ n14041 ;
  assign n14506 = n14031 ^ x106 ;
  assign n14507 = n14165 & n14506 ;
  assign n14508 = n14507 ^ n14034 ;
  assign n14499 = n14024 ^ x105 ;
  assign n14500 = n14165 & n14499 ;
  assign n14501 = n14500 ^ n14027 ;
  assign n14492 = n14017 ^ x104 ;
  assign n14493 = n14165 & n14492 ;
  assign n14494 = n14493 ^ n14020 ;
  assign n14485 = n14010 ^ x103 ;
  assign n14486 = n14165 & n14485 ;
  assign n14487 = n14486 ^ n14013 ;
  assign n14478 = n14003 ^ x102 ;
  assign n14479 = n14165 & n14478 ;
  assign n14480 = n14479 ^ n14006 ;
  assign n14471 = n14000 ^ x101 ;
  assign n14472 = n14165 & n14471 ;
  assign n14473 = n14472 ^ n13733 ;
  assign n14464 = n13997 ^ x100 ;
  assign n14465 = n14165 & n14464 ;
  assign n14466 = n14465 ^ n13737 ;
  assign n14457 = n13990 ^ x99 ;
  assign n14458 = n14165 & n14457 ;
  assign n14459 = n14458 ^ n13993 ;
  assign n14450 = n13983 ^ x98 ;
  assign n14451 = n14165 & n14450 ;
  assign n14452 = n14451 ^ n13986 ;
  assign n14443 = n13976 ^ x97 ;
  assign n14444 = n14165 & n14443 ;
  assign n14445 = n14444 ^ n13979 ;
  assign n14436 = n13969 ^ x96 ;
  assign n14437 = n14165 & n14436 ;
  assign n14438 = n14437 ^ n13972 ;
  assign n14172 = n13962 ^ x95 ;
  assign n14173 = n14165 & n14172 ;
  assign n14174 = n14173 ^ n13965 ;
  assign n14175 = n14174 ^ x96 ;
  assign n14179 = n14174 ^ x95 ;
  assign n14176 = n13960 & n14165 ;
  assign n14177 = n14176 ^ n13741 ;
  assign n14178 = n14177 ^ n14174 ;
  assign n14180 = n14179 ^ n14178 ;
  assign n14423 = n13951 ^ x93 ;
  assign n14424 = n14165 & n14423 ;
  assign n14425 = n14424 ^ n13954 ;
  assign n14408 = n13748 ^ x92 ;
  assign n14409 = n14408 ^ n13945 ;
  assign n14410 = n14409 ^ x91 ;
  assign n14411 = n14410 ^ n14408 ;
  assign n14413 = n13945 ^ x92 ;
  assign n14414 = n14413 ^ n14408 ;
  assign n14415 = ~n14411 & ~n14414 ;
  assign n14416 = n14415 ^ n14408 ;
  assign n14417 = n14165 & ~n14416 ;
  assign n14418 = n14417 ^ n13744 ;
  assign n14401 = n13945 ^ x91 ;
  assign n14402 = n14165 & n14401 ;
  assign n14403 = n14402 ^ n13748 ;
  assign n14394 = n13938 ^ x90 ;
  assign n14395 = n14165 & n14394 ;
  assign n14396 = n14395 ^ n13941 ;
  assign n14387 = n13931 ^ x89 ;
  assign n14388 = n14165 & n14387 ;
  assign n14389 = n14388 ^ n13934 ;
  assign n14181 = n13924 ^ x88 ;
  assign n14182 = n14165 & n14181 ;
  assign n14183 = n14182 ^ n13927 ;
  assign n14184 = n14183 ^ x89 ;
  assign n14189 = n14183 ^ x88 ;
  assign n14185 = n13917 ^ x87 ;
  assign n14186 = n14165 & n14185 ;
  assign n14187 = n14186 ^ n13920 ;
  assign n14188 = n14187 ^ n14183 ;
  assign n14190 = n14189 ^ n14188 ;
  assign n14374 = n13910 ^ x86 ;
  assign n14375 = n14165 & n14374 ;
  assign n14376 = n14375 ^ n13913 ;
  assign n14359 = n13758 ^ x85 ;
  assign n14360 = n14359 ^ n13904 ;
  assign n14361 = n14360 ^ x84 ;
  assign n14362 = n14361 ^ n14359 ;
  assign n14364 = n13904 ^ x85 ;
  assign n14365 = n14364 ^ n14359 ;
  assign n14366 = ~n14362 & ~n14365 ;
  assign n14367 = n14366 ^ n14359 ;
  assign n14368 = n14165 & ~n14367 ;
  assign n14369 = n14368 ^ n13754 ;
  assign n14352 = n13904 ^ x84 ;
  assign n14353 = n14165 & n14352 ;
  assign n14354 = n14353 ^ n13758 ;
  assign n14337 = n13768 ^ x83 ;
  assign n14338 = n14337 ^ n13898 ;
  assign n14339 = n14338 ^ x82 ;
  assign n14340 = n14339 ^ n14337 ;
  assign n14342 = n13898 ^ x83 ;
  assign n14343 = n14342 ^ n14337 ;
  assign n14344 = ~n14340 & ~n14343 ;
  assign n14345 = n14344 ^ n14337 ;
  assign n14346 = n14165 & ~n14345 ;
  assign n14347 = n14346 ^ n13764 ;
  assign n14330 = n13898 ^ x82 ;
  assign n14331 = n14165 & n14330 ;
  assign n14332 = n14331 ^ n13768 ;
  assign n14323 = n13895 ^ x81 ;
  assign n14324 = n14165 & n14323 ;
  assign n14325 = n14324 ^ n13774 ;
  assign n14316 = n13892 ^ x80 ;
  assign n14317 = n14165 & n14316 ;
  assign n14318 = n14317 ^ n13778 ;
  assign n14309 = n13885 ^ x79 ;
  assign n14310 = n14165 & n14309 ;
  assign n14311 = n14310 ^ n13888 ;
  assign n14302 = n13878 ^ x78 ;
  assign n14303 = n14165 & n14302 ;
  assign n14304 = n14303 ^ n13881 ;
  assign n14295 = n13871 ^ x77 ;
  assign n14296 = n14165 & n14295 ;
  assign n14297 = n14296 ^ n13874 ;
  assign n14288 = n13864 ^ x76 ;
  assign n14289 = n14165 & n14288 ;
  assign n14290 = n14289 ^ n13867 ;
  assign n14281 = n13857 ^ x75 ;
  assign n14282 = n14165 & n14281 ;
  assign n14283 = n14282 ^ n13860 ;
  assign n14191 = n13854 ^ x74 ;
  assign n14192 = n14165 & n14191 ;
  assign n14193 = n14192 ^ n13782 ;
  assign n14194 = n14193 ^ x75 ;
  assign n14199 = n14193 ^ x74 ;
  assign n14195 = n13851 ^ x73 ;
  assign n14196 = n14165 & n14195 ;
  assign n14197 = n14196 ^ n13786 ;
  assign n14198 = n14197 ^ n14193 ;
  assign n14200 = n14199 ^ n14198 ;
  assign n14268 = n13844 ^ x72 ;
  assign n14269 = n14165 & n14268 ;
  assign n14270 = n14269 ^ n13847 ;
  assign n14261 = n13837 ^ x71 ;
  assign n14262 = n14165 & n14261 ;
  assign n14263 = n14262 ^ n13840 ;
  assign n14254 = n13830 ^ x70 ;
  assign n14255 = n14165 & n14254 ;
  assign n14256 = n14255 ^ n13833 ;
  assign n14247 = n13823 ^ x69 ;
  assign n14248 = n14165 & n14247 ;
  assign n14249 = n14248 ^ n13826 ;
  assign n14240 = n13816 ^ x68 ;
  assign n14241 = n14165 & n14240 ;
  assign n14242 = n14241 ^ n13819 ;
  assign n14233 = n13809 ^ x67 ;
  assign n14234 = n14165 & n14233 ;
  assign n14235 = n14234 ^ n13812 ;
  assign n14226 = n13806 ^ x66 ;
  assign n14227 = n14165 & n14226 ;
  assign n14228 = n14227 ^ n13793 ;
  assign n14201 = ~x3 & x64 ;
  assign n14202 = n14201 ^ x65 ;
  assign n14203 = x64 & n14165 ;
  assign n14204 = n14203 ^ x4 ;
  assign n14205 = n14204 ^ n14201 ;
  assign n14206 = n14202 & n14205 ;
  assign n14207 = n14206 ^ x65 ;
  assign n14208 = n14207 ^ x66 ;
  assign n14211 = x65 & n14165 ;
  assign n14220 = n14211 ^ x5 ;
  assign n14212 = n14165 ^ n13710 ;
  assign n14213 = n14212 ^ n14211 ;
  assign n14214 = n14213 ^ n14212 ;
  assign n14215 = n14212 ^ x4 ;
  assign n14216 = n14215 ^ n14212 ;
  assign n14217 = n14214 & n14216 ;
  assign n14218 = n14217 ^ n14212 ;
  assign n14219 = x64 & n14218 ;
  assign n14221 = n14220 ^ n14219 ;
  assign n14209 = x4 & n3862 ;
  assign n14210 = n14165 & n14209 ;
  assign n14222 = n14221 ^ n14210 ;
  assign n14223 = n14222 ^ n14207 ;
  assign n14224 = n14208 & n14223 ;
  assign n14225 = n14224 ^ x66 ;
  assign n14229 = n14228 ^ n14225 ;
  assign n14230 = n14228 ^ x67 ;
  assign n14231 = n14229 & ~n14230 ;
  assign n14232 = n14231 ^ x67 ;
  assign n14236 = n14235 ^ n14232 ;
  assign n14237 = n14235 ^ x68 ;
  assign n14238 = n14236 & ~n14237 ;
  assign n14239 = n14238 ^ x68 ;
  assign n14243 = n14242 ^ n14239 ;
  assign n14244 = n14242 ^ x69 ;
  assign n14245 = n14243 & ~n14244 ;
  assign n14246 = n14245 ^ x69 ;
  assign n14250 = n14249 ^ n14246 ;
  assign n14251 = n14249 ^ x70 ;
  assign n14252 = n14250 & ~n14251 ;
  assign n14253 = n14252 ^ x70 ;
  assign n14257 = n14256 ^ n14253 ;
  assign n14258 = n14256 ^ x71 ;
  assign n14259 = n14257 & ~n14258 ;
  assign n14260 = n14259 ^ x71 ;
  assign n14264 = n14263 ^ n14260 ;
  assign n14265 = n14263 ^ x72 ;
  assign n14266 = n14264 & ~n14265 ;
  assign n14267 = n14266 ^ x72 ;
  assign n14271 = n14270 ^ n14267 ;
  assign n14272 = n14270 ^ x73 ;
  assign n14273 = n14271 & ~n14272 ;
  assign n14274 = n14273 ^ x73 ;
  assign n14275 = n14274 ^ n14193 ;
  assign n14276 = n14275 ^ n14199 ;
  assign n14277 = ~n14200 & n14276 ;
  assign n14278 = n14277 ^ n14199 ;
  assign n14279 = ~n14194 & n14278 ;
  assign n14280 = n14279 ^ x75 ;
  assign n14284 = n14283 ^ n14280 ;
  assign n14285 = n14283 ^ x76 ;
  assign n14286 = n14284 & ~n14285 ;
  assign n14287 = n14286 ^ x76 ;
  assign n14291 = n14290 ^ n14287 ;
  assign n14292 = n14290 ^ x77 ;
  assign n14293 = n14291 & ~n14292 ;
  assign n14294 = n14293 ^ x77 ;
  assign n14298 = n14297 ^ n14294 ;
  assign n14299 = n14297 ^ x78 ;
  assign n14300 = n14298 & ~n14299 ;
  assign n14301 = n14300 ^ x78 ;
  assign n14305 = n14304 ^ n14301 ;
  assign n14306 = n14304 ^ x79 ;
  assign n14307 = n14305 & ~n14306 ;
  assign n14308 = n14307 ^ x79 ;
  assign n14312 = n14311 ^ n14308 ;
  assign n14313 = n14311 ^ x80 ;
  assign n14314 = n14312 & ~n14313 ;
  assign n14315 = n14314 ^ x80 ;
  assign n14319 = n14318 ^ n14315 ;
  assign n14320 = n14318 ^ x81 ;
  assign n14321 = n14319 & ~n14320 ;
  assign n14322 = n14321 ^ x81 ;
  assign n14326 = n14325 ^ n14322 ;
  assign n14327 = n14325 ^ x82 ;
  assign n14328 = n14326 & ~n14327 ;
  assign n14329 = n14328 ^ x82 ;
  assign n14333 = n14332 ^ n14329 ;
  assign n14334 = n14332 ^ x83 ;
  assign n14335 = n14333 & ~n14334 ;
  assign n14336 = n14335 ^ x83 ;
  assign n14348 = n14347 ^ n14336 ;
  assign n14349 = n14347 ^ x84 ;
  assign n14350 = n14348 & ~n14349 ;
  assign n14351 = n14350 ^ x84 ;
  assign n14355 = n14354 ^ n14351 ;
  assign n14356 = n14354 ^ x85 ;
  assign n14357 = n14355 & ~n14356 ;
  assign n14358 = n14357 ^ x85 ;
  assign n14370 = n14369 ^ n14358 ;
  assign n14371 = n14369 ^ x86 ;
  assign n14372 = n14370 & ~n14371 ;
  assign n14373 = n14372 ^ x86 ;
  assign n14377 = n14376 ^ n14373 ;
  assign n14378 = n14376 ^ x87 ;
  assign n14379 = n14377 & ~n14378 ;
  assign n14380 = n14379 ^ x87 ;
  assign n14381 = n14380 ^ n14183 ;
  assign n14382 = n14381 ^ n14189 ;
  assign n14383 = ~n14190 & n14382 ;
  assign n14384 = n14383 ^ n14189 ;
  assign n14385 = ~n14184 & n14384 ;
  assign n14386 = n14385 ^ x89 ;
  assign n14390 = n14389 ^ n14386 ;
  assign n14391 = n14389 ^ x90 ;
  assign n14392 = n14390 & ~n14391 ;
  assign n14393 = n14392 ^ x90 ;
  assign n14397 = n14396 ^ n14393 ;
  assign n14398 = n14396 ^ x91 ;
  assign n14399 = n14397 & ~n14398 ;
  assign n14400 = n14399 ^ x91 ;
  assign n14404 = n14403 ^ n14400 ;
  assign n14405 = n14403 ^ x92 ;
  assign n14406 = n14404 & ~n14405 ;
  assign n14407 = n14406 ^ x92 ;
  assign n14419 = n14418 ^ n14407 ;
  assign n14420 = n14418 ^ x93 ;
  assign n14421 = n14419 & ~n14420 ;
  assign n14422 = n14421 ^ x93 ;
  assign n14426 = n14425 ^ n14422 ;
  assign n14427 = n14425 ^ x94 ;
  assign n14428 = n14426 & ~n14427 ;
  assign n14429 = n14428 ^ x94 ;
  assign n14430 = n14429 ^ n14174 ;
  assign n14431 = n14430 ^ n14179 ;
  assign n14432 = ~n14180 & n14431 ;
  assign n14433 = n14432 ^ n14179 ;
  assign n14434 = ~n14175 & n14433 ;
  assign n14435 = n14434 ^ x96 ;
  assign n14439 = n14438 ^ n14435 ;
  assign n14440 = n14438 ^ x97 ;
  assign n14441 = n14439 & ~n14440 ;
  assign n14442 = n14441 ^ x97 ;
  assign n14446 = n14445 ^ n14442 ;
  assign n14447 = n14445 ^ x98 ;
  assign n14448 = n14446 & ~n14447 ;
  assign n14449 = n14448 ^ x98 ;
  assign n14453 = n14452 ^ n14449 ;
  assign n14454 = n14452 ^ x99 ;
  assign n14455 = n14453 & ~n14454 ;
  assign n14456 = n14455 ^ x99 ;
  assign n14460 = n14459 ^ n14456 ;
  assign n14461 = n14459 ^ x100 ;
  assign n14462 = n14460 & ~n14461 ;
  assign n14463 = n14462 ^ x100 ;
  assign n14467 = n14466 ^ n14463 ;
  assign n14468 = n14466 ^ x101 ;
  assign n14469 = n14467 & ~n14468 ;
  assign n14470 = n14469 ^ x101 ;
  assign n14474 = n14473 ^ n14470 ;
  assign n14475 = n14473 ^ x102 ;
  assign n14476 = n14474 & ~n14475 ;
  assign n14477 = n14476 ^ x102 ;
  assign n14481 = n14480 ^ n14477 ;
  assign n14482 = n14480 ^ x103 ;
  assign n14483 = n14481 & ~n14482 ;
  assign n14484 = n14483 ^ x103 ;
  assign n14488 = n14487 ^ n14484 ;
  assign n14489 = n14487 ^ x104 ;
  assign n14490 = n14488 & ~n14489 ;
  assign n14491 = n14490 ^ x104 ;
  assign n14495 = n14494 ^ n14491 ;
  assign n14496 = n14494 ^ x105 ;
  assign n14497 = n14495 & ~n14496 ;
  assign n14498 = n14497 ^ x105 ;
  assign n14502 = n14501 ^ n14498 ;
  assign n14503 = n14501 ^ x106 ;
  assign n14504 = n14502 & ~n14503 ;
  assign n14505 = n14504 ^ x106 ;
  assign n14509 = n14508 ^ n14505 ;
  assign n14510 = n14508 ^ x107 ;
  assign n14511 = n14509 & ~n14510 ;
  assign n14512 = n14511 ^ x107 ;
  assign n14516 = n14515 ^ n14512 ;
  assign n14517 = n14515 ^ x108 ;
  assign n14518 = n14516 & ~n14517 ;
  assign n14519 = n14518 ^ x108 ;
  assign n14523 = n14522 ^ n14519 ;
  assign n14524 = n14522 ^ x109 ;
  assign n14525 = n14523 & ~n14524 ;
  assign n14526 = n14525 ^ x109 ;
  assign n14538 = n14537 ^ n14526 ;
  assign n14539 = n14537 ^ x110 ;
  assign n14540 = n14538 & ~n14539 ;
  assign n14541 = n14540 ^ x110 ;
  assign n14545 = n14544 ^ n14541 ;
  assign n14546 = n14544 ^ x111 ;
  assign n14547 = n14545 & ~n14546 ;
  assign n14548 = n14547 ^ x111 ;
  assign n14549 = n14548 ^ n14170 ;
  assign n14550 = ~n14171 & n14549 ;
  assign n14551 = n14550 ^ x112 ;
  assign n14552 = n14551 ^ n14167 ;
  assign n14553 = ~n14168 & n14552 ;
  assign n14554 = n14553 ^ x113 ;
  assign n14558 = n14557 ^ n14554 ;
  assign n14559 = n14557 ^ x114 ;
  assign n14560 = n14558 & ~n14559 ;
  assign n14561 = n14560 ^ x114 ;
  assign n14565 = n14564 ^ n14561 ;
  assign n14566 = n14564 ^ x115 ;
  assign n14567 = n14565 & ~n14566 ;
  assign n14568 = n14567 ^ x115 ;
  assign n14572 = n14571 ^ n14568 ;
  assign n14573 = n14571 ^ x116 ;
  assign n14574 = n14572 & ~n14573 ;
  assign n14575 = n14574 ^ x116 ;
  assign n14579 = n14578 ^ n14575 ;
  assign n14580 = n14578 ^ x117 ;
  assign n14581 = n14579 & ~n14580 ;
  assign n14582 = n14581 ^ x117 ;
  assign n14586 = n14585 ^ n14582 ;
  assign n14587 = n14585 ^ x118 ;
  assign n14588 = n14586 & ~n14587 ;
  assign n14589 = n14588 ^ x118 ;
  assign n14593 = n14592 ^ n14589 ;
  assign n14594 = n14592 ^ x119 ;
  assign n14595 = n14593 & ~n14594 ;
  assign n14596 = n14595 ^ x119 ;
  assign n14600 = n14599 ^ n14596 ;
  assign n14601 = n14599 ^ x120 ;
  assign n14602 = n14600 & ~n14601 ;
  assign n14603 = n14602 ^ x120 ;
  assign n14607 = n14606 ^ n14603 ;
  assign n14608 = n14606 ^ x121 ;
  assign n14609 = n14607 & ~n14608 ;
  assign n14610 = n14609 ^ x121 ;
  assign n14614 = n14613 ^ n14610 ;
  assign n14615 = n14613 ^ x122 ;
  assign n14616 = n14614 & ~n14615 ;
  assign n14617 = n14616 ^ x122 ;
  assign n14621 = n14620 ^ n14617 ;
  assign n14622 = n14620 ^ x123 ;
  assign n14623 = n14621 & ~n14622 ;
  assign n14624 = n14623 ^ x123 ;
  assign n14625 = n12838 & n14624 ;
  assign n14626 = n132 & n14080 ;
  assign n14627 = n14160 & n14626 ;
  assign n14628 = n14627 ^ n14080 ;
  assign n14629 = n14628 ^ x124 ;
  assign n14630 = n14629 ^ n12837 ;
  assign n14631 = n14625 & ~n14630 ;
  assign n14632 = n14631 ^ n12838 ;
  assign n15110 = n14617 ^ x123 ;
  assign n15111 = n14632 & n15110 ;
  assign n15112 = n15111 ^ n14620 ;
  assign n15103 = n14610 ^ x122 ;
  assign n15104 = n14632 & n15103 ;
  assign n15105 = n15104 ^ n14613 ;
  assign n15096 = n14603 ^ x121 ;
  assign n15097 = n14632 & n15096 ;
  assign n15098 = n15097 ^ n14606 ;
  assign n15089 = n14596 ^ x120 ;
  assign n15090 = n14632 & n15089 ;
  assign n15091 = n15090 ^ n14599 ;
  assign n15082 = n14589 ^ x119 ;
  assign n15083 = n14632 & n15082 ;
  assign n15084 = n15083 ^ n14592 ;
  assign n15075 = n14582 ^ x118 ;
  assign n15076 = n14632 & n15075 ;
  assign n15077 = n15076 ^ n14585 ;
  assign n15068 = n14575 ^ x117 ;
  assign n15069 = n14632 & n15068 ;
  assign n15070 = n15069 ^ n14578 ;
  assign n15061 = n14568 ^ x116 ;
  assign n15062 = n14632 & n15061 ;
  assign n15063 = n15062 ^ n14571 ;
  assign n14687 = n14561 ^ x115 ;
  assign n14688 = n14632 & n14687 ;
  assign n14689 = n14688 ^ n14564 ;
  assign n14690 = n14689 ^ x116 ;
  assign n14695 = n14689 ^ x115 ;
  assign n14691 = n14554 ^ x114 ;
  assign n14692 = n14632 & n14691 ;
  assign n14693 = n14692 ^ n14557 ;
  assign n14694 = n14693 ^ n14689 ;
  assign n14696 = n14695 ^ n14694 ;
  assign n15048 = n14551 ^ x113 ;
  assign n15049 = n14632 & n15048 ;
  assign n15050 = n15049 ^ n14167 ;
  assign n15041 = n14548 ^ x112 ;
  assign n15042 = n14632 & n15041 ;
  assign n15043 = n15042 ^ n14170 ;
  assign n15034 = n14541 ^ x111 ;
  assign n15035 = n14632 & n15034 ;
  assign n15036 = n15035 ^ n14544 ;
  assign n15027 = n14526 ^ x110 ;
  assign n15028 = n14632 & n15027 ;
  assign n15029 = n15028 ^ n14537 ;
  assign n15020 = n14519 ^ x109 ;
  assign n15021 = n14632 & n15020 ;
  assign n15022 = n15021 ^ n14522 ;
  assign n15013 = n14512 ^ x108 ;
  assign n15014 = n14632 & n15013 ;
  assign n15015 = n15014 ^ n14515 ;
  assign n15006 = n14505 ^ x107 ;
  assign n15007 = n14632 & n15006 ;
  assign n15008 = n15007 ^ n14508 ;
  assign n14999 = n14498 ^ x106 ;
  assign n15000 = n14632 & n14999 ;
  assign n15001 = n15000 ^ n14501 ;
  assign n14992 = n14491 ^ x105 ;
  assign n14993 = n14632 & n14992 ;
  assign n14994 = n14993 ^ n14494 ;
  assign n14985 = n14484 ^ x104 ;
  assign n14986 = n14632 & n14985 ;
  assign n14987 = n14986 ^ n14487 ;
  assign n14978 = n14477 ^ x103 ;
  assign n14979 = n14632 & n14978 ;
  assign n14980 = n14979 ^ n14480 ;
  assign n14697 = n14470 ^ x102 ;
  assign n14698 = n14632 & n14697 ;
  assign n14699 = n14698 ^ n14473 ;
  assign n14700 = n14699 ^ x103 ;
  assign n14705 = n14699 ^ x102 ;
  assign n14701 = n14463 ^ x101 ;
  assign n14702 = n14632 & n14701 ;
  assign n14703 = n14702 ^ n14466 ;
  assign n14704 = n14703 ^ n14699 ;
  assign n14706 = n14705 ^ n14704 ;
  assign n14965 = n14456 ^ x100 ;
  assign n14966 = n14632 & n14965 ;
  assign n14967 = n14966 ^ n14459 ;
  assign n14707 = n14449 ^ x99 ;
  assign n14708 = n14632 & n14707 ;
  assign n14709 = n14708 ^ n14452 ;
  assign n14710 = n14709 ^ x100 ;
  assign n14715 = n14709 ^ x99 ;
  assign n14711 = n14442 ^ x98 ;
  assign n14712 = n14632 & n14711 ;
  assign n14713 = n14712 ^ n14445 ;
  assign n14714 = n14713 ^ n14709 ;
  assign n14716 = n14715 ^ n14714 ;
  assign n14952 = n14435 ^ x97 ;
  assign n14953 = n14632 & n14952 ;
  assign n14954 = n14953 ^ n14438 ;
  assign n14937 = n14177 ^ x96 ;
  assign n14938 = n14937 ^ n14429 ;
  assign n14939 = n14938 ^ x95 ;
  assign n14940 = n14939 ^ n14937 ;
  assign n14942 = n14429 ^ x96 ;
  assign n14943 = n14942 ^ n14937 ;
  assign n14944 = ~n14940 & ~n14943 ;
  assign n14945 = n14944 ^ n14937 ;
  assign n14946 = n14632 & ~n14945 ;
  assign n14947 = n14946 ^ n14174 ;
  assign n14930 = n14429 ^ x95 ;
  assign n14931 = n14632 & n14930 ;
  assign n14932 = n14931 ^ n14177 ;
  assign n14923 = n14422 ^ x94 ;
  assign n14924 = n14632 & n14923 ;
  assign n14925 = n14924 ^ n14425 ;
  assign n14717 = n14400 ^ x92 ;
  assign n14718 = n14632 & n14717 ;
  assign n14719 = n14718 ^ n14403 ;
  assign n14720 = n14719 ^ x93 ;
  assign n14906 = n14393 ^ x91 ;
  assign n14907 = n14632 & n14906 ;
  assign n14908 = n14907 ^ n14396 ;
  assign n14899 = n14386 ^ x90 ;
  assign n14900 = n14632 & n14899 ;
  assign n14901 = n14900 ^ n14389 ;
  assign n14884 = n14187 ^ x89 ;
  assign n14885 = n14884 ^ n14380 ;
  assign n14886 = n14885 ^ x88 ;
  assign n14887 = n14886 ^ n14884 ;
  assign n14889 = n14380 ^ x89 ;
  assign n14890 = n14889 ^ n14884 ;
  assign n14891 = ~n14887 & ~n14890 ;
  assign n14892 = n14891 ^ n14884 ;
  assign n14893 = n14632 & ~n14892 ;
  assign n14894 = n14893 ^ n14183 ;
  assign n14877 = n14380 ^ x88 ;
  assign n14878 = n14632 & n14877 ;
  assign n14879 = n14878 ^ n14187 ;
  assign n14870 = n14373 ^ x87 ;
  assign n14871 = n14632 & n14870 ;
  assign n14872 = n14871 ^ n14376 ;
  assign n14863 = n14358 ^ x86 ;
  assign n14864 = n14632 & n14863 ;
  assign n14865 = n14864 ^ n14369 ;
  assign n14856 = n14351 ^ x85 ;
  assign n14857 = n14632 & n14856 ;
  assign n14858 = n14857 ^ n14354 ;
  assign n14849 = n14336 ^ x84 ;
  assign n14850 = n14632 & n14849 ;
  assign n14851 = n14850 ^ n14347 ;
  assign n14842 = n14329 ^ x83 ;
  assign n14843 = n14632 & n14842 ;
  assign n14844 = n14843 ^ n14332 ;
  assign n14835 = n14322 ^ x82 ;
  assign n14836 = n14632 & n14835 ;
  assign n14837 = n14836 ^ n14325 ;
  assign n14828 = n14315 ^ x81 ;
  assign n14829 = n14632 & n14828 ;
  assign n14830 = n14829 ^ n14318 ;
  assign n14821 = n14308 ^ x80 ;
  assign n14822 = n14632 & n14821 ;
  assign n14823 = n14822 ^ n14311 ;
  assign n14814 = n14301 ^ x79 ;
  assign n14815 = n14632 & n14814 ;
  assign n14816 = n14815 ^ n14304 ;
  assign n14807 = n14294 ^ x78 ;
  assign n14808 = n14632 & n14807 ;
  assign n14809 = n14808 ^ n14297 ;
  assign n14800 = n14287 ^ x77 ;
  assign n14801 = n14632 & n14800 ;
  assign n14802 = n14801 ^ n14290 ;
  assign n14793 = n14280 ^ x76 ;
  assign n14794 = n14632 & n14793 ;
  assign n14795 = n14794 ^ n14283 ;
  assign n14778 = n14197 ^ x75 ;
  assign n14779 = n14778 ^ n14274 ;
  assign n14780 = n14779 ^ x74 ;
  assign n14781 = n14780 ^ n14778 ;
  assign n14783 = n14274 ^ x75 ;
  assign n14784 = n14783 ^ n14778 ;
  assign n14785 = ~n14781 & ~n14784 ;
  assign n14786 = n14785 ^ n14778 ;
  assign n14787 = n14632 & ~n14786 ;
  assign n14788 = n14787 ^ n14193 ;
  assign n14771 = n14274 ^ x74 ;
  assign n14772 = n14632 & n14771 ;
  assign n14773 = n14772 ^ n14197 ;
  assign n14764 = n14267 ^ x73 ;
  assign n14765 = n14632 & n14764 ;
  assign n14766 = n14765 ^ n14270 ;
  assign n14753 = n14253 ^ x71 ;
  assign n14754 = n14632 & n14753 ;
  assign n14755 = n14754 ^ n14256 ;
  assign n14724 = n14246 ^ x70 ;
  assign n14725 = n14632 & n14724 ;
  assign n14726 = n14725 ^ n14249 ;
  assign n14727 = n14726 ^ x71 ;
  assign n14732 = n14726 ^ x70 ;
  assign n14728 = n14239 ^ x69 ;
  assign n14729 = n14632 & n14728 ;
  assign n14730 = n14729 ^ n14242 ;
  assign n14731 = n14730 ^ n14726 ;
  assign n14733 = n14732 ^ n14731 ;
  assign n14740 = n14232 ^ x68 ;
  assign n14741 = n14632 & n14740 ;
  assign n14742 = n14741 ^ n14235 ;
  assign n14647 = x3 & ~x4 ;
  assign n14648 = n926 & n14647 ;
  assign n14642 = n14204 ^ x65 ;
  assign n14643 = n14201 & ~n14642 ;
  assign n14644 = ~x2 & n14204 ;
  assign n14645 = n14643 & n14644 ;
  assign n14646 = n14645 ^ n14643 ;
  assign n14649 = n14648 ^ n14646 ;
  assign n14650 = n14632 & n14649 ;
  assign n129 = ~x2 & x64 ;
  assign n14633 = x3 & ~x65 ;
  assign n14634 = n14633 ^ n14632 ;
  assign n14635 = n129 & ~n14634 ;
  assign n14636 = x65 ^ x3 ;
  assign n14637 = n14636 ^ n14633 ;
  assign n14638 = n14204 & ~n14637 ;
  assign n14639 = n14202 & n14632 ;
  assign n14640 = n14638 & ~n14639 ;
  assign n14641 = ~n14635 & n14640 ;
  assign n14651 = n14650 ^ n14641 ;
  assign n14652 = ~x66 & n14637 ;
  assign n14653 = x64 & n14632 ;
  assign n14654 = n14632 ^ n14204 ;
  assign n14655 = ~n14653 & ~n14654 ;
  assign n14656 = n14652 & n14655 ;
  assign n14657 = n14656 ^ x66 ;
  assign n14658 = x64 & ~n14657 ;
  assign n14659 = n14204 ^ x2 ;
  assign n14660 = n14659 ^ x65 ;
  assign n14661 = n14660 ^ x3 ;
  assign n14662 = n14661 ^ n14632 ;
  assign n14663 = ~x2 & ~n14662 ;
  assign n14664 = n14663 ^ n14659 ;
  assign n14665 = n14632 ^ x3 ;
  assign n14666 = n14659 ^ n14632 ;
  assign n14667 = n14666 ^ x2 ;
  assign n14668 = ~n14665 & ~n14667 ;
  assign n14669 = n14668 ^ n14659 ;
  assign n14670 = ~n14664 & ~n14669 ;
  assign n14671 = n14670 ^ n14659 ;
  assign n14672 = n14658 & ~n14671 ;
  assign n14673 = n14672 ^ n14657 ;
  assign n14674 = ~n14651 & n14673 ;
  assign n14675 = n14674 ^ x67 ;
  assign n14676 = n14208 & n14632 ;
  assign n14677 = n14676 ^ n14222 ;
  assign n14678 = n14677 ^ n14674 ;
  assign n14679 = n14675 & n14678 ;
  assign n14680 = n14679 ^ x67 ;
  assign n14681 = n14680 ^ x68 ;
  assign n14734 = n14225 ^ x67 ;
  assign n14735 = n14632 & n14734 ;
  assign n14736 = n14735 ^ n14228 ;
  assign n14737 = n14736 ^ n14680 ;
  assign n14738 = n14681 & n14737 ;
  assign n14739 = n14738 ^ x68 ;
  assign n14743 = n14742 ^ n14739 ;
  assign n14744 = n14742 ^ x69 ;
  assign n14745 = n14743 & ~n14744 ;
  assign n14746 = n14745 ^ x69 ;
  assign n14747 = n14746 ^ n14726 ;
  assign n14748 = n14747 ^ n14732 ;
  assign n14749 = ~n14733 & n14748 ;
  assign n14750 = n14749 ^ n14732 ;
  assign n14751 = ~n14727 & n14750 ;
  assign n14752 = n14751 ^ x71 ;
  assign n14756 = n14755 ^ n14752 ;
  assign n14757 = n14755 ^ x72 ;
  assign n14758 = n14756 & ~n14757 ;
  assign n14759 = n14758 ^ x72 ;
  assign n14721 = n14260 ^ x72 ;
  assign n14722 = n14632 & n14721 ;
  assign n14723 = n14722 ^ n14263 ;
  assign n14760 = n14759 ^ n14723 ;
  assign n14761 = n14759 ^ x73 ;
  assign n14762 = n14760 & n14761 ;
  assign n14763 = n14762 ^ x73 ;
  assign n14767 = n14766 ^ n14763 ;
  assign n14768 = n14766 ^ x74 ;
  assign n14769 = n14767 & ~n14768 ;
  assign n14770 = n14769 ^ x74 ;
  assign n14774 = n14773 ^ n14770 ;
  assign n14775 = n14773 ^ x75 ;
  assign n14776 = n14774 & ~n14775 ;
  assign n14777 = n14776 ^ x75 ;
  assign n14789 = n14788 ^ n14777 ;
  assign n14790 = n14788 ^ x76 ;
  assign n14791 = n14789 & ~n14790 ;
  assign n14792 = n14791 ^ x76 ;
  assign n14796 = n14795 ^ n14792 ;
  assign n14797 = n14795 ^ x77 ;
  assign n14798 = n14796 & ~n14797 ;
  assign n14799 = n14798 ^ x77 ;
  assign n14803 = n14802 ^ n14799 ;
  assign n14804 = n14802 ^ x78 ;
  assign n14805 = n14803 & ~n14804 ;
  assign n14806 = n14805 ^ x78 ;
  assign n14810 = n14809 ^ n14806 ;
  assign n14811 = n14809 ^ x79 ;
  assign n14812 = n14810 & ~n14811 ;
  assign n14813 = n14812 ^ x79 ;
  assign n14817 = n14816 ^ n14813 ;
  assign n14818 = n14816 ^ x80 ;
  assign n14819 = n14817 & ~n14818 ;
  assign n14820 = n14819 ^ x80 ;
  assign n14824 = n14823 ^ n14820 ;
  assign n14825 = n14823 ^ x81 ;
  assign n14826 = n14824 & ~n14825 ;
  assign n14827 = n14826 ^ x81 ;
  assign n14831 = n14830 ^ n14827 ;
  assign n14832 = n14830 ^ x82 ;
  assign n14833 = n14831 & ~n14832 ;
  assign n14834 = n14833 ^ x82 ;
  assign n14838 = n14837 ^ n14834 ;
  assign n14839 = n14837 ^ x83 ;
  assign n14840 = n14838 & ~n14839 ;
  assign n14841 = n14840 ^ x83 ;
  assign n14845 = n14844 ^ n14841 ;
  assign n14846 = n14844 ^ x84 ;
  assign n14847 = n14845 & ~n14846 ;
  assign n14848 = n14847 ^ x84 ;
  assign n14852 = n14851 ^ n14848 ;
  assign n14853 = n14851 ^ x85 ;
  assign n14854 = n14852 & ~n14853 ;
  assign n14855 = n14854 ^ x85 ;
  assign n14859 = n14858 ^ n14855 ;
  assign n14860 = n14858 ^ x86 ;
  assign n14861 = n14859 & ~n14860 ;
  assign n14862 = n14861 ^ x86 ;
  assign n14866 = n14865 ^ n14862 ;
  assign n14867 = n14865 ^ x87 ;
  assign n14868 = n14866 & ~n14867 ;
  assign n14869 = n14868 ^ x87 ;
  assign n14873 = n14872 ^ n14869 ;
  assign n14874 = n14872 ^ x88 ;
  assign n14875 = n14873 & ~n14874 ;
  assign n14876 = n14875 ^ x88 ;
  assign n14880 = n14879 ^ n14876 ;
  assign n14881 = n14879 ^ x89 ;
  assign n14882 = n14880 & ~n14881 ;
  assign n14883 = n14882 ^ x89 ;
  assign n14895 = n14894 ^ n14883 ;
  assign n14896 = n14894 ^ x90 ;
  assign n14897 = n14895 & ~n14896 ;
  assign n14898 = n14897 ^ x90 ;
  assign n14902 = n14901 ^ n14898 ;
  assign n14903 = n14901 ^ x91 ;
  assign n14904 = n14902 & ~n14903 ;
  assign n14905 = n14904 ^ x91 ;
  assign n14909 = n14908 ^ n14905 ;
  assign n14910 = n14908 ^ x92 ;
  assign n14911 = n14909 & ~n14910 ;
  assign n14912 = n14911 ^ x92 ;
  assign n14913 = n14912 ^ n14719 ;
  assign n14914 = ~n14720 & n14913 ;
  assign n14915 = n14914 ^ x93 ;
  assign n14916 = n14915 ^ x94 ;
  assign n14917 = n14407 ^ x93 ;
  assign n14918 = n14632 & n14917 ;
  assign n14919 = n14918 ^ n14418 ;
  assign n14920 = n14919 ^ n14915 ;
  assign n14921 = n14916 & n14920 ;
  assign n14922 = n14921 ^ x94 ;
  assign n14926 = n14925 ^ n14922 ;
  assign n14927 = n14925 ^ x95 ;
  assign n14928 = n14926 & ~n14927 ;
  assign n14929 = n14928 ^ x95 ;
  assign n14933 = n14932 ^ n14929 ;
  assign n14934 = n14932 ^ x96 ;
  assign n14935 = n14933 & ~n14934 ;
  assign n14936 = n14935 ^ x96 ;
  assign n14948 = n14947 ^ n14936 ;
  assign n14949 = n14947 ^ x97 ;
  assign n14950 = n14948 & ~n14949 ;
  assign n14951 = n14950 ^ x97 ;
  assign n14955 = n14954 ^ n14951 ;
  assign n14956 = n14954 ^ x98 ;
  assign n14957 = n14955 & ~n14956 ;
  assign n14958 = n14957 ^ x98 ;
  assign n14959 = n14958 ^ n14709 ;
  assign n14960 = n14959 ^ n14715 ;
  assign n14961 = ~n14716 & n14960 ;
  assign n14962 = n14961 ^ n14715 ;
  assign n14963 = ~n14710 & n14962 ;
  assign n14964 = n14963 ^ x100 ;
  assign n14968 = n14967 ^ n14964 ;
  assign n14969 = n14967 ^ x101 ;
  assign n14970 = n14968 & ~n14969 ;
  assign n14971 = n14970 ^ x101 ;
  assign n14972 = n14971 ^ n14699 ;
  assign n14973 = n14972 ^ n14705 ;
  assign n14974 = ~n14706 & n14973 ;
  assign n14975 = n14974 ^ n14705 ;
  assign n14976 = ~n14700 & n14975 ;
  assign n14977 = n14976 ^ x103 ;
  assign n14981 = n14980 ^ n14977 ;
  assign n14982 = n14980 ^ x104 ;
  assign n14983 = n14981 & ~n14982 ;
  assign n14984 = n14983 ^ x104 ;
  assign n14988 = n14987 ^ n14984 ;
  assign n14989 = n14987 ^ x105 ;
  assign n14990 = n14988 & ~n14989 ;
  assign n14991 = n14990 ^ x105 ;
  assign n14995 = n14994 ^ n14991 ;
  assign n14996 = n14994 ^ x106 ;
  assign n14997 = n14995 & ~n14996 ;
  assign n14998 = n14997 ^ x106 ;
  assign n15002 = n15001 ^ n14998 ;
  assign n15003 = n15001 ^ x107 ;
  assign n15004 = n15002 & ~n15003 ;
  assign n15005 = n15004 ^ x107 ;
  assign n15009 = n15008 ^ n15005 ;
  assign n15010 = n15008 ^ x108 ;
  assign n15011 = n15009 & ~n15010 ;
  assign n15012 = n15011 ^ x108 ;
  assign n15016 = n15015 ^ n15012 ;
  assign n15017 = n15015 ^ x109 ;
  assign n15018 = n15016 & ~n15017 ;
  assign n15019 = n15018 ^ x109 ;
  assign n15023 = n15022 ^ n15019 ;
  assign n15024 = n15022 ^ x110 ;
  assign n15025 = n15023 & ~n15024 ;
  assign n15026 = n15025 ^ x110 ;
  assign n15030 = n15029 ^ n15026 ;
  assign n15031 = n15029 ^ x111 ;
  assign n15032 = n15030 & ~n15031 ;
  assign n15033 = n15032 ^ x111 ;
  assign n15037 = n15036 ^ n15033 ;
  assign n15038 = n15036 ^ x112 ;
  assign n15039 = n15037 & ~n15038 ;
  assign n15040 = n15039 ^ x112 ;
  assign n15044 = n15043 ^ n15040 ;
  assign n15045 = n15043 ^ x113 ;
  assign n15046 = n15044 & ~n15045 ;
  assign n15047 = n15046 ^ x113 ;
  assign n15051 = n15050 ^ n15047 ;
  assign n15052 = n15050 ^ x114 ;
  assign n15053 = n15051 & ~n15052 ;
  assign n15054 = n15053 ^ x114 ;
  assign n15055 = n15054 ^ n14689 ;
  assign n15056 = n15055 ^ n14695 ;
  assign n15057 = ~n14696 & n15056 ;
  assign n15058 = n15057 ^ n14695 ;
  assign n15059 = ~n14690 & n15058 ;
  assign n15060 = n15059 ^ x116 ;
  assign n15064 = n15063 ^ n15060 ;
  assign n15065 = n15063 ^ x117 ;
  assign n15066 = n15064 & ~n15065 ;
  assign n15067 = n15066 ^ x117 ;
  assign n15071 = n15070 ^ n15067 ;
  assign n15072 = n15070 ^ x118 ;
  assign n15073 = n15071 & ~n15072 ;
  assign n15074 = n15073 ^ x118 ;
  assign n15078 = n15077 ^ n15074 ;
  assign n15079 = n15077 ^ x119 ;
  assign n15080 = n15078 & ~n15079 ;
  assign n15081 = n15080 ^ x119 ;
  assign n15085 = n15084 ^ n15081 ;
  assign n15086 = n15084 ^ x120 ;
  assign n15087 = n15085 & ~n15086 ;
  assign n15088 = n15087 ^ x120 ;
  assign n15092 = n15091 ^ n15088 ;
  assign n15093 = n15091 ^ x121 ;
  assign n15094 = n15092 & ~n15093 ;
  assign n15095 = n15094 ^ x121 ;
  assign n15099 = n15098 ^ n15095 ;
  assign n15100 = n15098 ^ x122 ;
  assign n15101 = n15099 & ~n15100 ;
  assign n15102 = n15101 ^ x122 ;
  assign n15106 = n15105 ^ n15102 ;
  assign n15107 = n15105 ^ x123 ;
  assign n15108 = n15106 & ~n15107 ;
  assign n15109 = n15108 ^ x123 ;
  assign n15113 = n15112 ^ n15109 ;
  assign n15603 = n15109 ^ x124 ;
  assign n15117 = n15113 & n15603 ;
  assign n15114 = x125 ^ x124 ;
  assign n15118 = n15117 ^ n15114 ;
  assign n14682 = n14624 ^ x124 ;
  assign n14683 = n131 & n14628 ;
  assign n14684 = n14682 & n14683 ;
  assign n14685 = n14684 ^ n14628 ;
  assign n15299 = n130 & n14685 ;
  assign n15300 = n15118 & n15299 ;
  assign n15301 = n15300 ^ n14685 ;
  assign n15302 = n15301 ^ x126 ;
  assign n14686 = n14685 ^ x125 ;
  assign n15121 = ~n14686 & n15118 ;
  assign n15122 = n15121 ^ x125 ;
  assign n15123 = n130 & ~n15122 ;
  assign n15604 = n15123 & n15603 ;
  assign n15605 = n15604 ^ n15112 ;
  assign n15596 = n15102 ^ x123 ;
  assign n15597 = n15123 & n15596 ;
  assign n15598 = n15597 ^ n15105 ;
  assign n15589 = n15095 ^ x122 ;
  assign n15590 = n15123 & n15589 ;
  assign n15591 = n15590 ^ n15098 ;
  assign n15582 = n15088 ^ x121 ;
  assign n15583 = n15123 & n15582 ;
  assign n15584 = n15583 ^ n15091 ;
  assign n15575 = n15081 ^ x120 ;
  assign n15576 = n15123 & n15575 ;
  assign n15577 = n15576 ^ n15084 ;
  assign n15568 = n15074 ^ x119 ;
  assign n15569 = n15123 & n15568 ;
  assign n15570 = n15569 ^ n15077 ;
  assign n15303 = n15067 ^ x118 ;
  assign n15304 = n15123 & n15303 ;
  assign n15305 = n15304 ^ n15070 ;
  assign n15306 = n15305 ^ x119 ;
  assign n15311 = n15305 ^ x118 ;
  assign n15307 = n15060 ^ x117 ;
  assign n15308 = n15123 & n15307 ;
  assign n15309 = n15308 ^ n15063 ;
  assign n15310 = n15309 ^ n15305 ;
  assign n15312 = n15311 ^ n15310 ;
  assign n15547 = n14693 ^ x116 ;
  assign n15548 = n15547 ^ n15054 ;
  assign n15549 = n15548 ^ x115 ;
  assign n15550 = n15549 ^ n15547 ;
  assign n15552 = n15054 ^ x116 ;
  assign n15553 = n15552 ^ n15547 ;
  assign n15554 = ~n15550 & ~n15553 ;
  assign n15555 = n15554 ^ n15547 ;
  assign n15556 = n15123 & ~n15555 ;
  assign n15557 = n15556 ^ n14689 ;
  assign n15540 = n15054 ^ x115 ;
  assign n15541 = n15123 & n15540 ;
  assign n15542 = n15541 ^ n14693 ;
  assign n15533 = n15047 ^ x114 ;
  assign n15534 = n15123 & n15533 ;
  assign n15535 = n15534 ^ n15050 ;
  assign n15313 = n15040 ^ x113 ;
  assign n15314 = n15123 & n15313 ;
  assign n15315 = n15314 ^ n15043 ;
  assign n15316 = n15315 ^ x114 ;
  assign n15321 = n15315 ^ x113 ;
  assign n15317 = n15033 ^ x112 ;
  assign n15318 = n15123 & n15317 ;
  assign n15319 = n15318 ^ n15036 ;
  assign n15320 = n15319 ^ n15315 ;
  assign n15322 = n15321 ^ n15320 ;
  assign n15520 = n15026 ^ x111 ;
  assign n15521 = n15123 & n15520 ;
  assign n15522 = n15521 ^ n15029 ;
  assign n15513 = n15019 ^ x110 ;
  assign n15514 = n15123 & n15513 ;
  assign n15515 = n15514 ^ n15022 ;
  assign n15506 = n15012 ^ x109 ;
  assign n15507 = n15123 & n15506 ;
  assign n15508 = n15507 ^ n15015 ;
  assign n15499 = n15005 ^ x108 ;
  assign n15500 = n15123 & n15499 ;
  assign n15501 = n15500 ^ n15008 ;
  assign n15492 = n14998 ^ x107 ;
  assign n15493 = n15123 & n15492 ;
  assign n15494 = n15493 ^ n15001 ;
  assign n15485 = n14991 ^ x106 ;
  assign n15486 = n15123 & n15485 ;
  assign n15487 = n15486 ^ n14994 ;
  assign n15478 = n14984 ^ x105 ;
  assign n15479 = n15123 & n15478 ;
  assign n15480 = n15479 ^ n14987 ;
  assign n15471 = n14977 ^ x104 ;
  assign n15472 = n15123 & n15471 ;
  assign n15473 = n15472 ^ n14980 ;
  assign n15323 = n14703 ^ x103 ;
  assign n15324 = n15323 ^ n14971 ;
  assign n15325 = n15324 ^ x102 ;
  assign n15326 = n15325 ^ n15323 ;
  assign n15328 = n14971 ^ x103 ;
  assign n15329 = n15328 ^ n15323 ;
  assign n15330 = ~n15326 & ~n15329 ;
  assign n15331 = n15330 ^ n15323 ;
  assign n15332 = n15123 & ~n15331 ;
  assign n15333 = n15332 ^ n14699 ;
  assign n15334 = n15333 ^ x104 ;
  assign n15335 = n14971 ^ x102 ;
  assign n15336 = n15123 & n15335 ;
  assign n15337 = n15336 ^ n14703 ;
  assign n15338 = n15337 ^ x103 ;
  assign n15458 = n14964 ^ x101 ;
  assign n15459 = n15123 & n15458 ;
  assign n15460 = n15459 ^ n14967 ;
  assign n15443 = n14713 ^ x100 ;
  assign n15444 = n15443 ^ n14958 ;
  assign n15445 = n15444 ^ x99 ;
  assign n15446 = n15445 ^ n15443 ;
  assign n15448 = n14958 ^ x100 ;
  assign n15449 = n15448 ^ n15443 ;
  assign n15450 = ~n15446 & ~n15449 ;
  assign n15451 = n15450 ^ n15443 ;
  assign n15452 = n15123 & ~n15451 ;
  assign n15453 = n15452 ^ n14709 ;
  assign n15436 = n14958 ^ x99 ;
  assign n15437 = n15123 & n15436 ;
  assign n15438 = n15437 ^ n14713 ;
  assign n15429 = n14951 ^ x98 ;
  assign n15430 = n15123 & n15429 ;
  assign n15431 = n15430 ^ n14954 ;
  assign n15422 = n14936 ^ x97 ;
  assign n15423 = n15123 & n15422 ;
  assign n15424 = n15423 ^ n14947 ;
  assign n15415 = n14929 ^ x96 ;
  assign n15416 = n15123 & n15415 ;
  assign n15417 = n15416 ^ n14932 ;
  assign n15408 = n14922 ^ x95 ;
  assign n15409 = n15123 & n15408 ;
  assign n15410 = n15409 ^ n14925 ;
  assign n15402 = n14916 & n15123 ;
  assign n15403 = n15402 ^ n14919 ;
  assign n15395 = n14912 ^ x93 ;
  assign n15396 = n15123 & n15395 ;
  assign n15397 = n15396 ^ n14719 ;
  assign n15388 = n14905 ^ x92 ;
  assign n15389 = n15123 & n15388 ;
  assign n15390 = n15389 ^ n14908 ;
  assign n15381 = n14898 ^ x91 ;
  assign n15382 = n15123 & n15381 ;
  assign n15383 = n15382 ^ n14901 ;
  assign n15374 = n14883 ^ x90 ;
  assign n15375 = n15123 & n15374 ;
  assign n15376 = n15375 ^ n14894 ;
  assign n15367 = n14876 ^ x89 ;
  assign n15368 = n15123 & n15367 ;
  assign n15369 = n15368 ^ n14879 ;
  assign n15360 = n14869 ^ x88 ;
  assign n15361 = n15123 & n15360 ;
  assign n15362 = n15361 ^ n14872 ;
  assign n15353 = n14862 ^ x87 ;
  assign n15354 = n15123 & n15353 ;
  assign n15355 = n15354 ^ n14865 ;
  assign n15346 = n14855 ^ x86 ;
  assign n15347 = n15123 & n15346 ;
  assign n15348 = n15347 ^ n14858 ;
  assign n15339 = n14848 ^ x85 ;
  assign n15340 = n15123 & n15339 ;
  assign n15341 = n15340 ^ n14851 ;
  assign n15291 = n14841 ^ x84 ;
  assign n15292 = n15123 & n15291 ;
  assign n15293 = n15292 ^ n14844 ;
  assign n15284 = n14834 ^ x83 ;
  assign n15285 = n15123 & n15284 ;
  assign n15286 = n15285 ^ n14837 ;
  assign n15277 = n14827 ^ x82 ;
  assign n15278 = n15123 & n15277 ;
  assign n15279 = n15278 ^ n14830 ;
  assign n15270 = n14820 ^ x81 ;
  assign n15271 = n15123 & n15270 ;
  assign n15272 = n15271 ^ n14823 ;
  assign n15263 = n14813 ^ x80 ;
  assign n15264 = n15123 & n15263 ;
  assign n15265 = n15264 ^ n14816 ;
  assign n15256 = n14806 ^ x79 ;
  assign n15257 = n15123 & n15256 ;
  assign n15258 = n15257 ^ n14809 ;
  assign n15249 = n14799 ^ x78 ;
  assign n15250 = n15123 & n15249 ;
  assign n15251 = n15250 ^ n14802 ;
  assign n15242 = n14792 ^ x77 ;
  assign n15243 = n15123 & n15242 ;
  assign n15244 = n15243 ^ n14795 ;
  assign n15235 = n14777 ^ x76 ;
  assign n15236 = n15123 & n15235 ;
  assign n15237 = n15236 ^ n14788 ;
  assign n15228 = n14770 ^ x75 ;
  assign n15229 = n15123 & n15228 ;
  assign n15230 = n15229 ^ n14773 ;
  assign n15221 = n14763 ^ x74 ;
  assign n15222 = n15123 & n15221 ;
  assign n15223 = n15222 ^ n14766 ;
  assign n15215 = n14761 & n15123 ;
  assign n15216 = n15215 ^ n14723 ;
  assign n15208 = n14752 ^ x72 ;
  assign n15209 = n15123 & n15208 ;
  assign n15210 = n15209 ^ n14755 ;
  assign n15193 = n14730 ^ x71 ;
  assign n15194 = n15193 ^ n14746 ;
  assign n15195 = n15194 ^ x70 ;
  assign n15196 = n15195 ^ n15193 ;
  assign n15198 = n14746 ^ x71 ;
  assign n15199 = n15198 ^ n15193 ;
  assign n15200 = ~n15196 & ~n15199 ;
  assign n15201 = n15200 ^ n15193 ;
  assign n15202 = n15123 & ~n15201 ;
  assign n15203 = n15202 ^ n14726 ;
  assign n15186 = n14746 ^ x70 ;
  assign n15187 = n15123 & n15186 ;
  assign n15188 = n15187 ^ n14730 ;
  assign n15179 = n14739 ^ x69 ;
  assign n15180 = n15123 & n15179 ;
  assign n15181 = n15180 ^ n14742 ;
  assign n15124 = n14681 & n15123 ;
  assign n15125 = n15124 ^ n14736 ;
  assign n15126 = n15125 ^ x69 ;
  assign n15130 = n15125 ^ x68 ;
  assign n15127 = n14675 & n15123 ;
  assign n15128 = n15127 ^ n14677 ;
  assign n15129 = n15128 ^ n15125 ;
  assign n15131 = n15130 ^ n15129 ;
  assign n15167 = n14639 ^ n14204 ;
  assign n15162 = x3 & x65 ;
  assign n15152 = x65 ^ x2 ;
  assign n15153 = x64 ^ x3 ;
  assign n15154 = n15153 ^ x65 ;
  assign n15155 = n15154 ^ n14632 ;
  assign n15156 = ~n15152 & n15155 ;
  assign n15163 = n15162 ^ n15156 ;
  assign n15164 = ~x64 & n15163 ;
  assign n15159 = n15156 ^ n7358 ;
  assign n15165 = n15164 ^ n15159 ;
  assign n15166 = n15123 & n15165 ;
  assign n15168 = n15167 ^ n15166 ;
  assign n15145 = n129 ^ x65 ;
  assign n15146 = n15123 & n15145 ;
  assign n15144 = n14653 ^ x3 ;
  assign n15147 = n15146 ^ n15144 ;
  assign n15139 = x2 & x65 ;
  assign n15136 = x65 ^ x1 ;
  assign n15132 = x64 ^ x2 ;
  assign n15133 = n15132 ^ x65 ;
  assign n15137 = n15133 ^ n15123 ;
  assign n15138 = ~n15136 & n15137 ;
  assign n15140 = n15139 ^ n15138 ;
  assign n15141 = x64 & n15140 ;
  assign n15142 = n15141 ^ n15139 ;
  assign n15143 = n15142 ^ x65 ;
  assign n15148 = n15147 ^ n15143 ;
  assign n15149 = n15147 ^ x66 ;
  assign n15150 = n15148 & ~n15149 ;
  assign n15151 = n15150 ^ x66 ;
  assign n15169 = n15168 ^ n15151 ;
  assign n15170 = n15168 ^ x67 ;
  assign n15171 = n15169 & ~n15170 ;
  assign n15172 = n15171 ^ x67 ;
  assign n15173 = n15172 ^ n15125 ;
  assign n15174 = n15173 ^ n15130 ;
  assign n15175 = ~n15131 & n15174 ;
  assign n15176 = n15175 ^ n15130 ;
  assign n15177 = ~n15126 & n15176 ;
  assign n15178 = n15177 ^ x69 ;
  assign n15182 = n15181 ^ n15178 ;
  assign n15183 = n15181 ^ x70 ;
  assign n15184 = n15182 & ~n15183 ;
  assign n15185 = n15184 ^ x70 ;
  assign n15189 = n15188 ^ n15185 ;
  assign n15190 = n15188 ^ x71 ;
  assign n15191 = n15189 & ~n15190 ;
  assign n15192 = n15191 ^ x71 ;
  assign n15204 = n15203 ^ n15192 ;
  assign n15205 = n15203 ^ x72 ;
  assign n15206 = n15204 & ~n15205 ;
  assign n15207 = n15206 ^ x72 ;
  assign n15211 = n15210 ^ n15207 ;
  assign n15212 = n15210 ^ x73 ;
  assign n15213 = n15211 & ~n15212 ;
  assign n15214 = n15213 ^ x73 ;
  assign n15217 = n15216 ^ n15214 ;
  assign n15218 = n15216 ^ x74 ;
  assign n15219 = n15217 & ~n15218 ;
  assign n15220 = n15219 ^ x74 ;
  assign n15224 = n15223 ^ n15220 ;
  assign n15225 = n15223 ^ x75 ;
  assign n15226 = n15224 & ~n15225 ;
  assign n15227 = n15226 ^ x75 ;
  assign n15231 = n15230 ^ n15227 ;
  assign n15232 = n15230 ^ x76 ;
  assign n15233 = n15231 & ~n15232 ;
  assign n15234 = n15233 ^ x76 ;
  assign n15238 = n15237 ^ n15234 ;
  assign n15239 = n15237 ^ x77 ;
  assign n15240 = n15238 & ~n15239 ;
  assign n15241 = n15240 ^ x77 ;
  assign n15245 = n15244 ^ n15241 ;
  assign n15246 = n15244 ^ x78 ;
  assign n15247 = n15245 & ~n15246 ;
  assign n15248 = n15247 ^ x78 ;
  assign n15252 = n15251 ^ n15248 ;
  assign n15253 = n15251 ^ x79 ;
  assign n15254 = n15252 & ~n15253 ;
  assign n15255 = n15254 ^ x79 ;
  assign n15259 = n15258 ^ n15255 ;
  assign n15260 = n15258 ^ x80 ;
  assign n15261 = n15259 & ~n15260 ;
  assign n15262 = n15261 ^ x80 ;
  assign n15266 = n15265 ^ n15262 ;
  assign n15267 = n15265 ^ x81 ;
  assign n15268 = n15266 & ~n15267 ;
  assign n15269 = n15268 ^ x81 ;
  assign n15273 = n15272 ^ n15269 ;
  assign n15274 = n15272 ^ x82 ;
  assign n15275 = n15273 & ~n15274 ;
  assign n15276 = n15275 ^ x82 ;
  assign n15280 = n15279 ^ n15276 ;
  assign n15281 = n15279 ^ x83 ;
  assign n15282 = n15280 & ~n15281 ;
  assign n15283 = n15282 ^ x83 ;
  assign n15287 = n15286 ^ n15283 ;
  assign n15288 = n15286 ^ x84 ;
  assign n15289 = n15287 & ~n15288 ;
  assign n15290 = n15289 ^ x84 ;
  assign n15294 = n15293 ^ n15290 ;
  assign n15295 = n15293 ^ x85 ;
  assign n15296 = n15294 & ~n15295 ;
  assign n15297 = n15296 ^ x85 ;
  assign n15342 = n15341 ^ n15297 ;
  assign n15343 = n15341 ^ x86 ;
  assign n15344 = n15342 & ~n15343 ;
  assign n15345 = n15344 ^ x86 ;
  assign n15349 = n15348 ^ n15345 ;
  assign n15350 = n15348 ^ x87 ;
  assign n15351 = n15349 & ~n15350 ;
  assign n15352 = n15351 ^ x87 ;
  assign n15356 = n15355 ^ n15352 ;
  assign n15357 = n15355 ^ x88 ;
  assign n15358 = n15356 & ~n15357 ;
  assign n15359 = n15358 ^ x88 ;
  assign n15363 = n15362 ^ n15359 ;
  assign n15364 = n15362 ^ x89 ;
  assign n15365 = n15363 & ~n15364 ;
  assign n15366 = n15365 ^ x89 ;
  assign n15370 = n15369 ^ n15366 ;
  assign n15371 = n15369 ^ x90 ;
  assign n15372 = n15370 & ~n15371 ;
  assign n15373 = n15372 ^ x90 ;
  assign n15377 = n15376 ^ n15373 ;
  assign n15378 = n15376 ^ x91 ;
  assign n15379 = n15377 & ~n15378 ;
  assign n15380 = n15379 ^ x91 ;
  assign n15384 = n15383 ^ n15380 ;
  assign n15385 = n15383 ^ x92 ;
  assign n15386 = n15384 & ~n15385 ;
  assign n15387 = n15386 ^ x92 ;
  assign n15391 = n15390 ^ n15387 ;
  assign n15392 = n15390 ^ x93 ;
  assign n15393 = n15391 & ~n15392 ;
  assign n15394 = n15393 ^ x93 ;
  assign n15398 = n15397 ^ n15394 ;
  assign n15399 = n15397 ^ x94 ;
  assign n15400 = n15398 & ~n15399 ;
  assign n15401 = n15400 ^ x94 ;
  assign n15404 = n15403 ^ n15401 ;
  assign n15405 = n15403 ^ x95 ;
  assign n15406 = n15404 & ~n15405 ;
  assign n15407 = n15406 ^ x95 ;
  assign n15411 = n15410 ^ n15407 ;
  assign n15412 = n15410 ^ x96 ;
  assign n15413 = n15411 & ~n15412 ;
  assign n15414 = n15413 ^ x96 ;
  assign n15418 = n15417 ^ n15414 ;
  assign n15419 = n15417 ^ x97 ;
  assign n15420 = n15418 & ~n15419 ;
  assign n15421 = n15420 ^ x97 ;
  assign n15425 = n15424 ^ n15421 ;
  assign n15426 = n15424 ^ x98 ;
  assign n15427 = n15425 & ~n15426 ;
  assign n15428 = n15427 ^ x98 ;
  assign n15432 = n15431 ^ n15428 ;
  assign n15433 = n15431 ^ x99 ;
  assign n15434 = n15432 & ~n15433 ;
  assign n15435 = n15434 ^ x99 ;
  assign n15439 = n15438 ^ n15435 ;
  assign n15440 = n15438 ^ x100 ;
  assign n15441 = n15439 & ~n15440 ;
  assign n15442 = n15441 ^ x100 ;
  assign n15454 = n15453 ^ n15442 ;
  assign n15455 = n15453 ^ x101 ;
  assign n15456 = n15454 & ~n15455 ;
  assign n15457 = n15456 ^ x101 ;
  assign n15461 = n15460 ^ n15457 ;
  assign n15462 = n15460 ^ x102 ;
  assign n15463 = n15461 & ~n15462 ;
  assign n15464 = n15463 ^ x102 ;
  assign n15465 = n15464 ^ n15337 ;
  assign n15466 = ~n15338 & n15465 ;
  assign n15467 = n15466 ^ x103 ;
  assign n15468 = n15467 ^ n15333 ;
  assign n15469 = ~n15334 & n15468 ;
  assign n15470 = n15469 ^ x104 ;
  assign n15474 = n15473 ^ n15470 ;
  assign n15475 = n15473 ^ x105 ;
  assign n15476 = n15474 & ~n15475 ;
  assign n15477 = n15476 ^ x105 ;
  assign n15481 = n15480 ^ n15477 ;
  assign n15482 = n15480 ^ x106 ;
  assign n15483 = n15481 & ~n15482 ;
  assign n15484 = n15483 ^ x106 ;
  assign n15488 = n15487 ^ n15484 ;
  assign n15489 = n15487 ^ x107 ;
  assign n15490 = n15488 & ~n15489 ;
  assign n15491 = n15490 ^ x107 ;
  assign n15495 = n15494 ^ n15491 ;
  assign n15496 = n15494 ^ x108 ;
  assign n15497 = n15495 & ~n15496 ;
  assign n15498 = n15497 ^ x108 ;
  assign n15502 = n15501 ^ n15498 ;
  assign n15503 = n15501 ^ x109 ;
  assign n15504 = n15502 & ~n15503 ;
  assign n15505 = n15504 ^ x109 ;
  assign n15509 = n15508 ^ n15505 ;
  assign n15510 = n15508 ^ x110 ;
  assign n15511 = n15509 & ~n15510 ;
  assign n15512 = n15511 ^ x110 ;
  assign n15516 = n15515 ^ n15512 ;
  assign n15517 = n15515 ^ x111 ;
  assign n15518 = n15516 & ~n15517 ;
  assign n15519 = n15518 ^ x111 ;
  assign n15523 = n15522 ^ n15519 ;
  assign n15524 = n15522 ^ x112 ;
  assign n15525 = n15523 & ~n15524 ;
  assign n15526 = n15525 ^ x112 ;
  assign n15527 = n15526 ^ n15315 ;
  assign n15528 = n15527 ^ n15321 ;
  assign n15529 = ~n15322 & n15528 ;
  assign n15530 = n15529 ^ n15321 ;
  assign n15531 = ~n15316 & n15530 ;
  assign n15532 = n15531 ^ x114 ;
  assign n15536 = n15535 ^ n15532 ;
  assign n15537 = n15535 ^ x115 ;
  assign n15538 = n15536 & ~n15537 ;
  assign n15539 = n15538 ^ x115 ;
  assign n15543 = n15542 ^ n15539 ;
  assign n15544 = n15542 ^ x116 ;
  assign n15545 = n15543 & ~n15544 ;
  assign n15546 = n15545 ^ x116 ;
  assign n15558 = n15557 ^ n15546 ;
  assign n15559 = n15557 ^ x117 ;
  assign n15560 = n15558 & ~n15559 ;
  assign n15561 = n15560 ^ x117 ;
  assign n15562 = n15561 ^ n15305 ;
  assign n15563 = n15562 ^ n15311 ;
  assign n15564 = ~n15312 & n15563 ;
  assign n15565 = n15564 ^ n15311 ;
  assign n15566 = ~n15306 & n15565 ;
  assign n15567 = n15566 ^ x119 ;
  assign n15571 = n15570 ^ n15567 ;
  assign n15572 = n15570 ^ x120 ;
  assign n15573 = n15571 & ~n15572 ;
  assign n15574 = n15573 ^ x120 ;
  assign n15578 = n15577 ^ n15574 ;
  assign n15579 = n15577 ^ x121 ;
  assign n15580 = n15578 & ~n15579 ;
  assign n15581 = n15580 ^ x121 ;
  assign n15585 = n15584 ^ n15581 ;
  assign n15586 = n15584 ^ x122 ;
  assign n15587 = n15585 & ~n15586 ;
  assign n15588 = n15587 ^ x122 ;
  assign n15592 = n15591 ^ n15588 ;
  assign n15593 = n15591 ^ x123 ;
  assign n15594 = n15592 & ~n15593 ;
  assign n15595 = n15594 ^ x123 ;
  assign n15599 = n15598 ^ n15595 ;
  assign n15600 = n15598 ^ x124 ;
  assign n15601 = n15599 & ~n15600 ;
  assign n15602 = n15601 ^ x124 ;
  assign n15606 = n15605 ^ n15602 ;
  assign n16080 = n15602 ^ x125 ;
  assign n15610 = n15606 & n16080 ;
  assign n15607 = x126 ^ x125 ;
  assign n15611 = n15610 ^ n15607 ;
  assign n15614 = ~n15302 & n15611 ;
  assign n15615 = n15614 ^ x126 ;
  assign n15616 = ~x127 & ~n15615 ;
  assign n16081 = n15616 & n16080 ;
  assign n16082 = n16081 ^ n15605 ;
  assign n16073 = n15595 ^ x124 ;
  assign n16074 = n15616 & n16073 ;
  assign n16075 = n16074 ^ n15598 ;
  assign n16066 = n15588 ^ x123 ;
  assign n16067 = n15616 & n16066 ;
  assign n16068 = n16067 ^ n15591 ;
  assign n16059 = n15581 ^ x122 ;
  assign n16060 = n15616 & n16059 ;
  assign n16061 = n16060 ^ n15584 ;
  assign n16052 = n15574 ^ x121 ;
  assign n16053 = n15616 & n16052 ;
  assign n16054 = n16053 ^ n15577 ;
  assign n16045 = n15567 ^ x120 ;
  assign n16046 = n15616 & n16045 ;
  assign n16047 = n16046 ^ n15570 ;
  assign n16030 = n15309 ^ x119 ;
  assign n16031 = n16030 ^ n15561 ;
  assign n16032 = n16031 ^ x118 ;
  assign n16033 = n16032 ^ n16030 ;
  assign n16035 = n15561 ^ x119 ;
  assign n16036 = n16035 ^ n16030 ;
  assign n16037 = ~n16033 & ~n16036 ;
  assign n16038 = n16037 ^ n16030 ;
  assign n16039 = n15616 & ~n16038 ;
  assign n16040 = n16039 ^ n15305 ;
  assign n16023 = n15561 ^ x118 ;
  assign n16024 = n15616 & n16023 ;
  assign n16025 = n16024 ^ n15309 ;
  assign n16016 = n15546 ^ x117 ;
  assign n16017 = n15616 & n16016 ;
  assign n16018 = n16017 ^ n15557 ;
  assign n16009 = n15539 ^ x116 ;
  assign n16010 = n15616 & n16009 ;
  assign n16011 = n16010 ^ n15542 ;
  assign n16002 = n15532 ^ x115 ;
  assign n16003 = n15616 & n16002 ;
  assign n16004 = n16003 ^ n15535 ;
  assign n15987 = n15319 ^ x114 ;
  assign n15988 = n15987 ^ n15526 ;
  assign n15989 = n15988 ^ x113 ;
  assign n15990 = n15989 ^ n15987 ;
  assign n15992 = n15526 ^ x114 ;
  assign n15993 = n15992 ^ n15987 ;
  assign n15994 = ~n15990 & ~n15993 ;
  assign n15995 = n15994 ^ n15987 ;
  assign n15996 = n15616 & ~n15995 ;
  assign n15997 = n15996 ^ n15315 ;
  assign n15980 = n15526 ^ x113 ;
  assign n15981 = n15616 & n15980 ;
  assign n15982 = n15981 ^ n15319 ;
  assign n15973 = n15519 ^ x112 ;
  assign n15974 = n15616 & n15973 ;
  assign n15975 = n15974 ^ n15522 ;
  assign n15966 = n15512 ^ x111 ;
  assign n15967 = n15616 & n15966 ;
  assign n15968 = n15967 ^ n15515 ;
  assign n15959 = n15505 ^ x110 ;
  assign n15960 = n15616 & n15959 ;
  assign n15961 = n15960 ^ n15508 ;
  assign n15952 = n15498 ^ x109 ;
  assign n15953 = n15616 & n15952 ;
  assign n15954 = n15953 ^ n15501 ;
  assign n15945 = n15491 ^ x108 ;
  assign n15946 = n15616 & n15945 ;
  assign n15947 = n15946 ^ n15494 ;
  assign n15938 = n15484 ^ x107 ;
  assign n15939 = n15616 & n15938 ;
  assign n15940 = n15939 ^ n15487 ;
  assign n15931 = n15477 ^ x106 ;
  assign n15932 = n15616 & n15931 ;
  assign n15933 = n15932 ^ n15480 ;
  assign n15924 = n15470 ^ x105 ;
  assign n15925 = n15616 & n15924 ;
  assign n15926 = n15925 ^ n15473 ;
  assign n15917 = n15467 ^ x104 ;
  assign n15918 = n15616 & n15917 ;
  assign n15919 = n15918 ^ n15333 ;
  assign n15910 = n15464 ^ x103 ;
  assign n15911 = n15616 & n15910 ;
  assign n15912 = n15911 ^ n15337 ;
  assign n15903 = n15457 ^ x102 ;
  assign n15904 = n15616 & n15903 ;
  assign n15905 = n15904 ^ n15460 ;
  assign n15896 = n15442 ^ x101 ;
  assign n15897 = n15616 & n15896 ;
  assign n15898 = n15897 ^ n15453 ;
  assign n15889 = n15435 ^ x100 ;
  assign n15890 = n15616 & n15889 ;
  assign n15891 = n15890 ^ n15438 ;
  assign n15882 = n15428 ^ x99 ;
  assign n15883 = n15616 & n15882 ;
  assign n15884 = n15883 ^ n15431 ;
  assign n15875 = n15421 ^ x98 ;
  assign n15876 = n15616 & n15875 ;
  assign n15877 = n15876 ^ n15424 ;
  assign n15868 = n15414 ^ x97 ;
  assign n15869 = n15616 & n15868 ;
  assign n15870 = n15869 ^ n15417 ;
  assign n15861 = n15407 ^ x96 ;
  assign n15862 = n15616 & n15861 ;
  assign n15863 = n15862 ^ n15410 ;
  assign n15854 = n15401 ^ x95 ;
  assign n15855 = n15616 & n15854 ;
  assign n15856 = n15855 ^ n15403 ;
  assign n15847 = n15394 ^ x94 ;
  assign n15848 = n15616 & n15847 ;
  assign n15849 = n15848 ^ n15397 ;
  assign n15840 = n15387 ^ x93 ;
  assign n15841 = n15616 & n15840 ;
  assign n15842 = n15841 ^ n15390 ;
  assign n15833 = n15380 ^ x92 ;
  assign n15834 = n15616 & n15833 ;
  assign n15835 = n15834 ^ n15383 ;
  assign n15826 = n15373 ^ x91 ;
  assign n15827 = n15616 & n15826 ;
  assign n15828 = n15827 ^ n15376 ;
  assign n15819 = n15366 ^ x90 ;
  assign n15820 = n15616 & n15819 ;
  assign n15821 = n15820 ^ n15369 ;
  assign n15812 = n15359 ^ x89 ;
  assign n15813 = n15616 & n15812 ;
  assign n15814 = n15813 ^ n15362 ;
  assign n15805 = n15352 ^ x88 ;
  assign n15806 = n15616 & n15805 ;
  assign n15807 = n15806 ^ n15355 ;
  assign n15798 = n15345 ^ x87 ;
  assign n15799 = n15616 & n15798 ;
  assign n15800 = n15799 ^ n15348 ;
  assign n15298 = n15297 ^ x86 ;
  assign n15617 = n15298 & n15616 ;
  assign n15618 = n15617 ^ n15341 ;
  assign n15619 = n15618 ^ x87 ;
  assign n15624 = n15618 ^ x86 ;
  assign n15620 = n15290 ^ x85 ;
  assign n15621 = n15616 & n15620 ;
  assign n15622 = n15621 ^ n15293 ;
  assign n15623 = n15622 ^ n15618 ;
  assign n15625 = n15624 ^ n15623 ;
  assign n15785 = n15283 ^ x84 ;
  assign n15786 = n15616 & n15785 ;
  assign n15787 = n15786 ^ n15286 ;
  assign n15778 = n15276 ^ x83 ;
  assign n15779 = n15616 & n15778 ;
  assign n15780 = n15779 ^ n15279 ;
  assign n15771 = n15269 ^ x82 ;
  assign n15772 = n15616 & n15771 ;
  assign n15773 = n15772 ^ n15272 ;
  assign n15764 = n15262 ^ x81 ;
  assign n15765 = n15616 & n15764 ;
  assign n15766 = n15765 ^ n15265 ;
  assign n15757 = n15255 ^ x80 ;
  assign n15758 = n15616 & n15757 ;
  assign n15759 = n15758 ^ n15258 ;
  assign n15750 = n15248 ^ x79 ;
  assign n15751 = n15616 & n15750 ;
  assign n15752 = n15751 ^ n15251 ;
  assign n15743 = n15241 ^ x78 ;
  assign n15744 = n15616 & n15743 ;
  assign n15745 = n15744 ^ n15244 ;
  assign n15736 = n15234 ^ x77 ;
  assign n15737 = n15616 & n15736 ;
  assign n15738 = n15737 ^ n15237 ;
  assign n15626 = n15227 ^ x76 ;
  assign n15627 = n15616 & n15626 ;
  assign n15628 = n15627 ^ n15230 ;
  assign n15629 = n15628 ^ x77 ;
  assign n15634 = n15628 ^ x76 ;
  assign n15630 = n15220 ^ x75 ;
  assign n15631 = n15616 & n15630 ;
  assign n15632 = n15631 ^ n15223 ;
  assign n15633 = n15632 ^ n15628 ;
  assign n15635 = n15634 ^ n15633 ;
  assign n15723 = n15214 ^ x74 ;
  assign n15724 = n15616 & n15723 ;
  assign n15725 = n15724 ^ n15216 ;
  assign n15716 = n15207 ^ x73 ;
  assign n15717 = n15616 & n15716 ;
  assign n15718 = n15717 ^ n15210 ;
  assign n15709 = n15192 ^ x72 ;
  assign n15710 = n15616 & n15709 ;
  assign n15711 = n15710 ^ n15203 ;
  assign n15636 = n15185 ^ x71 ;
  assign n15637 = n15616 & n15636 ;
  assign n15638 = n15637 ^ n15188 ;
  assign n15639 = n15638 ^ x72 ;
  assign n15640 = n15178 ^ x70 ;
  assign n15641 = n15616 & n15640 ;
  assign n15642 = n15641 ^ n15181 ;
  assign n15643 = n15642 ^ x71 ;
  assign n15688 = n15128 ^ x69 ;
  assign n15689 = n15688 ^ n15172 ;
  assign n15690 = n15689 ^ x68 ;
  assign n15691 = n15690 ^ n15688 ;
  assign n15693 = n15172 ^ x69 ;
  assign n15694 = n15693 ^ n15688 ;
  assign n15695 = ~n15691 & ~n15694 ;
  assign n15696 = n15695 ^ n15688 ;
  assign n15697 = n15616 & ~n15696 ;
  assign n15698 = n15697 ^ n15125 ;
  assign n15681 = n15172 ^ x68 ;
  assign n15682 = n15616 & n15681 ;
  assign n15683 = n15682 ^ n15128 ;
  assign n15674 = n15151 ^ x67 ;
  assign n15675 = n15616 & n15674 ;
  assign n15676 = n15675 ^ n15168 ;
  assign n15661 = x1 & x65 ;
  assign n15658 = x65 ^ x0 ;
  assign n15654 = x64 ^ x1 ;
  assign n15655 = n15654 ^ x65 ;
  assign n15659 = n15655 ^ n15616 ;
  assign n15660 = ~n15658 & n15659 ;
  assign n15662 = n15661 ^ n15660 ;
  assign n15663 = x64 & n15662 ;
  assign n15664 = n15663 ^ n15661 ;
  assign n15665 = n15664 ^ x65 ;
  assign n15652 = x64 & n15123 ;
  assign n15648 = ~x1 & x64 ;
  assign n15649 = n15648 ^ x65 ;
  assign n15650 = n15616 & n15649 ;
  assign n15651 = n15650 ^ x2 ;
  assign n15653 = n15652 ^ n15651 ;
  assign n15666 = n15665 ^ n15653 ;
  assign n15667 = n15665 ^ x66 ;
  assign n15668 = n15666 & n15667 ;
  assign n15669 = n15668 ^ x66 ;
  assign n15644 = n15143 ^ x66 ;
  assign n15645 = n15616 & n15644 ;
  assign n15646 = n15645 ^ n15147 ;
  assign n15670 = n15669 ^ n15646 ;
  assign n15671 = n15669 ^ x67 ;
  assign n15672 = n15670 & n15671 ;
  assign n15673 = n15672 ^ x67 ;
  assign n15677 = n15676 ^ n15673 ;
  assign n15678 = n15676 ^ x68 ;
  assign n15679 = n15677 & ~n15678 ;
  assign n15680 = n15679 ^ x68 ;
  assign n15684 = n15683 ^ n15680 ;
  assign n15685 = n15683 ^ x69 ;
  assign n15686 = n15684 & ~n15685 ;
  assign n15687 = n15686 ^ x69 ;
  assign n15699 = n15698 ^ n15687 ;
  assign n15700 = n15698 ^ x70 ;
  assign n15701 = n15699 & ~n15700 ;
  assign n15702 = n15701 ^ x70 ;
  assign n15703 = n15702 ^ n15642 ;
  assign n15704 = ~n15643 & n15703 ;
  assign n15705 = n15704 ^ x71 ;
  assign n15706 = n15705 ^ n15638 ;
  assign n15707 = ~n15639 & n15706 ;
  assign n15708 = n15707 ^ x72 ;
  assign n15712 = n15711 ^ n15708 ;
  assign n15713 = n15711 ^ x73 ;
  assign n15714 = n15712 & ~n15713 ;
  assign n15715 = n15714 ^ x73 ;
  assign n15719 = n15718 ^ n15715 ;
  assign n15720 = n15718 ^ x74 ;
  assign n15721 = n15719 & ~n15720 ;
  assign n15722 = n15721 ^ x74 ;
  assign n15726 = n15725 ^ n15722 ;
  assign n15727 = n15725 ^ x75 ;
  assign n15728 = n15726 & ~n15727 ;
  assign n15729 = n15728 ^ x75 ;
  assign n15730 = n15729 ^ n15628 ;
  assign n15731 = n15730 ^ n15634 ;
  assign n15732 = ~n15635 & n15731 ;
  assign n15733 = n15732 ^ n15634 ;
  assign n15734 = ~n15629 & n15733 ;
  assign n15735 = n15734 ^ x77 ;
  assign n15739 = n15738 ^ n15735 ;
  assign n15740 = n15738 ^ x78 ;
  assign n15741 = n15739 & ~n15740 ;
  assign n15742 = n15741 ^ x78 ;
  assign n15746 = n15745 ^ n15742 ;
  assign n15747 = n15745 ^ x79 ;
  assign n15748 = n15746 & ~n15747 ;
  assign n15749 = n15748 ^ x79 ;
  assign n15753 = n15752 ^ n15749 ;
  assign n15754 = n15752 ^ x80 ;
  assign n15755 = n15753 & ~n15754 ;
  assign n15756 = n15755 ^ x80 ;
  assign n15760 = n15759 ^ n15756 ;
  assign n15761 = n15759 ^ x81 ;
  assign n15762 = n15760 & ~n15761 ;
  assign n15763 = n15762 ^ x81 ;
  assign n15767 = n15766 ^ n15763 ;
  assign n15768 = n15766 ^ x82 ;
  assign n15769 = n15767 & ~n15768 ;
  assign n15770 = n15769 ^ x82 ;
  assign n15774 = n15773 ^ n15770 ;
  assign n15775 = n15773 ^ x83 ;
  assign n15776 = n15774 & ~n15775 ;
  assign n15777 = n15776 ^ x83 ;
  assign n15781 = n15780 ^ n15777 ;
  assign n15782 = n15780 ^ x84 ;
  assign n15783 = n15781 & ~n15782 ;
  assign n15784 = n15783 ^ x84 ;
  assign n15788 = n15787 ^ n15784 ;
  assign n15789 = n15787 ^ x85 ;
  assign n15790 = n15788 & ~n15789 ;
  assign n15791 = n15790 ^ x85 ;
  assign n15792 = n15791 ^ n15618 ;
  assign n15793 = n15792 ^ n15624 ;
  assign n15794 = ~n15625 & n15793 ;
  assign n15795 = n15794 ^ n15624 ;
  assign n15796 = ~n15619 & n15795 ;
  assign n15797 = n15796 ^ x87 ;
  assign n15801 = n15800 ^ n15797 ;
  assign n15802 = n15800 ^ x88 ;
  assign n15803 = n15801 & ~n15802 ;
  assign n15804 = n15803 ^ x88 ;
  assign n15808 = n15807 ^ n15804 ;
  assign n15809 = n15807 ^ x89 ;
  assign n15810 = n15808 & ~n15809 ;
  assign n15811 = n15810 ^ x89 ;
  assign n15815 = n15814 ^ n15811 ;
  assign n15816 = n15814 ^ x90 ;
  assign n15817 = n15815 & ~n15816 ;
  assign n15818 = n15817 ^ x90 ;
  assign n15822 = n15821 ^ n15818 ;
  assign n15823 = n15821 ^ x91 ;
  assign n15824 = n15822 & ~n15823 ;
  assign n15825 = n15824 ^ x91 ;
  assign n15829 = n15828 ^ n15825 ;
  assign n15830 = n15828 ^ x92 ;
  assign n15831 = n15829 & ~n15830 ;
  assign n15832 = n15831 ^ x92 ;
  assign n15836 = n15835 ^ n15832 ;
  assign n15837 = n15835 ^ x93 ;
  assign n15838 = n15836 & ~n15837 ;
  assign n15839 = n15838 ^ x93 ;
  assign n15843 = n15842 ^ n15839 ;
  assign n15844 = n15842 ^ x94 ;
  assign n15845 = n15843 & ~n15844 ;
  assign n15846 = n15845 ^ x94 ;
  assign n15850 = n15849 ^ n15846 ;
  assign n15851 = n15849 ^ x95 ;
  assign n15852 = n15850 & ~n15851 ;
  assign n15853 = n15852 ^ x95 ;
  assign n15857 = n15856 ^ n15853 ;
  assign n15858 = n15856 ^ x96 ;
  assign n15859 = n15857 & ~n15858 ;
  assign n15860 = n15859 ^ x96 ;
  assign n15864 = n15863 ^ n15860 ;
  assign n15865 = n15863 ^ x97 ;
  assign n15866 = n15864 & ~n15865 ;
  assign n15867 = n15866 ^ x97 ;
  assign n15871 = n15870 ^ n15867 ;
  assign n15872 = n15870 ^ x98 ;
  assign n15873 = n15871 & ~n15872 ;
  assign n15874 = n15873 ^ x98 ;
  assign n15878 = n15877 ^ n15874 ;
  assign n15879 = n15877 ^ x99 ;
  assign n15880 = n15878 & ~n15879 ;
  assign n15881 = n15880 ^ x99 ;
  assign n15885 = n15884 ^ n15881 ;
  assign n15886 = n15884 ^ x100 ;
  assign n15887 = n15885 & ~n15886 ;
  assign n15888 = n15887 ^ x100 ;
  assign n15892 = n15891 ^ n15888 ;
  assign n15893 = n15891 ^ x101 ;
  assign n15894 = n15892 & ~n15893 ;
  assign n15895 = n15894 ^ x101 ;
  assign n15899 = n15898 ^ n15895 ;
  assign n15900 = n15898 ^ x102 ;
  assign n15901 = n15899 & ~n15900 ;
  assign n15902 = n15901 ^ x102 ;
  assign n15906 = n15905 ^ n15902 ;
  assign n15907 = n15905 ^ x103 ;
  assign n15908 = n15906 & ~n15907 ;
  assign n15909 = n15908 ^ x103 ;
  assign n15913 = n15912 ^ n15909 ;
  assign n15914 = n15912 ^ x104 ;
  assign n15915 = n15913 & ~n15914 ;
  assign n15916 = n15915 ^ x104 ;
  assign n15920 = n15919 ^ n15916 ;
  assign n15921 = n15919 ^ x105 ;
  assign n15922 = n15920 & ~n15921 ;
  assign n15923 = n15922 ^ x105 ;
  assign n15927 = n15926 ^ n15923 ;
  assign n15928 = n15926 ^ x106 ;
  assign n15929 = n15927 & ~n15928 ;
  assign n15930 = n15929 ^ x106 ;
  assign n15934 = n15933 ^ n15930 ;
  assign n15935 = n15933 ^ x107 ;
  assign n15936 = n15934 & ~n15935 ;
  assign n15937 = n15936 ^ x107 ;
  assign n15941 = n15940 ^ n15937 ;
  assign n15942 = n15940 ^ x108 ;
  assign n15943 = n15941 & ~n15942 ;
  assign n15944 = n15943 ^ x108 ;
  assign n15948 = n15947 ^ n15944 ;
  assign n15949 = n15947 ^ x109 ;
  assign n15950 = n15948 & ~n15949 ;
  assign n15951 = n15950 ^ x109 ;
  assign n15955 = n15954 ^ n15951 ;
  assign n15956 = n15954 ^ x110 ;
  assign n15957 = n15955 & ~n15956 ;
  assign n15958 = n15957 ^ x110 ;
  assign n15962 = n15961 ^ n15958 ;
  assign n15963 = n15961 ^ x111 ;
  assign n15964 = n15962 & ~n15963 ;
  assign n15965 = n15964 ^ x111 ;
  assign n15969 = n15968 ^ n15965 ;
  assign n15970 = n15968 ^ x112 ;
  assign n15971 = n15969 & ~n15970 ;
  assign n15972 = n15971 ^ x112 ;
  assign n15976 = n15975 ^ n15972 ;
  assign n15977 = n15975 ^ x113 ;
  assign n15978 = n15976 & ~n15977 ;
  assign n15979 = n15978 ^ x113 ;
  assign n15983 = n15982 ^ n15979 ;
  assign n15984 = n15982 ^ x114 ;
  assign n15985 = n15983 & ~n15984 ;
  assign n15986 = n15985 ^ x114 ;
  assign n15998 = n15997 ^ n15986 ;
  assign n15999 = n15997 ^ x115 ;
  assign n16000 = n15998 & ~n15999 ;
  assign n16001 = n16000 ^ x115 ;
  assign n16005 = n16004 ^ n16001 ;
  assign n16006 = n16004 ^ x116 ;
  assign n16007 = n16005 & ~n16006 ;
  assign n16008 = n16007 ^ x116 ;
  assign n16012 = n16011 ^ n16008 ;
  assign n16013 = n16011 ^ x117 ;
  assign n16014 = n16012 & ~n16013 ;
  assign n16015 = n16014 ^ x117 ;
  assign n16019 = n16018 ^ n16015 ;
  assign n16020 = n16018 ^ x118 ;
  assign n16021 = n16019 & ~n16020 ;
  assign n16022 = n16021 ^ x118 ;
  assign n16026 = n16025 ^ n16022 ;
  assign n16027 = n16025 ^ x119 ;
  assign n16028 = n16026 & ~n16027 ;
  assign n16029 = n16028 ^ x119 ;
  assign n16041 = n16040 ^ n16029 ;
  assign n16042 = n16040 ^ x120 ;
  assign n16043 = n16041 & ~n16042 ;
  assign n16044 = n16043 ^ x120 ;
  assign n16048 = n16047 ^ n16044 ;
  assign n16049 = n16047 ^ x121 ;
  assign n16050 = n16048 & ~n16049 ;
  assign n16051 = n16050 ^ x121 ;
  assign n16055 = n16054 ^ n16051 ;
  assign n16056 = n16054 ^ x122 ;
  assign n16057 = n16055 & ~n16056 ;
  assign n16058 = n16057 ^ x122 ;
  assign n16062 = n16061 ^ n16058 ;
  assign n16063 = n16061 ^ x123 ;
  assign n16064 = n16062 & ~n16063 ;
  assign n16065 = n16064 ^ x123 ;
  assign n16069 = n16068 ^ n16065 ;
  assign n16070 = n16068 ^ x124 ;
  assign n16071 = n16069 & ~n16070 ;
  assign n16072 = n16071 ^ x124 ;
  assign n16076 = n16075 ^ n16072 ;
  assign n16077 = n16075 ^ x125 ;
  assign n16078 = n16076 & ~n16077 ;
  assign n16079 = n16078 ^ x125 ;
  assign n16083 = n16082 ^ n16079 ;
  assign n16084 = n16082 ^ x126 ;
  assign n16085 = n16083 & ~n16084 ;
  assign n16086 = n16085 ^ x126 ;
  assign n16087 = n16086 ^ x127 ;
  assign n16090 = n15301 & ~n15611 ;
  assign n16091 = n16090 ^ n14080 ;
  assign n16092 = n16086 & ~n16091 ;
  assign n16093 = n16092 ^ n14080 ;
  assign n16094 = n16087 & ~n16093 ;
  assign n16095 = n16094 ^ n16086 ;
  assign n16096 = n267 ^ n220 ;
  assign n16097 = ~x63 & x64 ;
  assign n16098 = ~x65 & ~x66 ;
  assign n16099 = ~n16097 & n16098 ;
  assign n16100 = n194 & n16099 ;
  assign n16101 = x64 & ~n16095 ;
  assign n16102 = n16101 ^ x0 ;
  assign n16108 = x64 & n15616 ;
  assign n16104 = ~x0 & x64 ;
  assign n16105 = n16104 ^ x65 ;
  assign n16106 = ~n16095 & n16105 ;
  assign n16107 = n16106 ^ x1 ;
  assign n16109 = n16108 ^ n16107 ;
  assign n16110 = n15667 & ~n16095 ;
  assign n16111 = n16110 ^ n15653 ;
  assign n16112 = n15671 & ~n16095 ;
  assign n16113 = n16112 ^ n15646 ;
  assign n16114 = n15673 ^ x68 ;
  assign n16115 = ~n16095 & n16114 ;
  assign n16116 = n16115 ^ n15676 ;
  assign n16117 = n15680 ^ x69 ;
  assign n16118 = ~n16095 & n16117 ;
  assign n16119 = n16118 ^ n15683 ;
  assign n16120 = n15687 ^ x70 ;
  assign n16121 = ~n16095 & n16120 ;
  assign n16122 = n16121 ^ n15698 ;
  assign n16123 = n15702 ^ x71 ;
  assign n16124 = ~n16095 & n16123 ;
  assign n16125 = n16124 ^ n15642 ;
  assign n16126 = n15705 ^ x72 ;
  assign n16127 = ~n16095 & n16126 ;
  assign n16128 = n16127 ^ n15638 ;
  assign n16129 = n15708 ^ x73 ;
  assign n16130 = ~n16095 & n16129 ;
  assign n16131 = n16130 ^ n15711 ;
  assign n16132 = n15715 ^ x74 ;
  assign n16133 = ~n16095 & n16132 ;
  assign n16134 = n16133 ^ n15718 ;
  assign n16135 = n15722 ^ x75 ;
  assign n16136 = ~n16095 & n16135 ;
  assign n16137 = n16136 ^ n15725 ;
  assign n16138 = n15729 ^ x76 ;
  assign n16139 = ~n16095 & n16138 ;
  assign n16140 = n16139 ^ n15632 ;
  assign n16141 = n15632 ^ x77 ;
  assign n16142 = n16141 ^ x76 ;
  assign n16143 = n16142 ^ n15729 ;
  assign n16144 = n16143 ^ n16141 ;
  assign n16146 = x77 ^ x76 ;
  assign n16147 = n16146 ^ n16141 ;
  assign n16148 = ~n16144 & ~n16147 ;
  assign n16149 = n16148 ^ n16141 ;
  assign n16150 = ~n16095 & ~n16149 ;
  assign n16151 = n16150 ^ n15628 ;
  assign n16152 = n15735 ^ x78 ;
  assign n16153 = ~n16095 & n16152 ;
  assign n16154 = n16153 ^ n15738 ;
  assign n16155 = n15742 ^ x79 ;
  assign n16156 = ~n16095 & n16155 ;
  assign n16157 = n16156 ^ n15745 ;
  assign n16158 = n15749 ^ x80 ;
  assign n16159 = ~n16095 & n16158 ;
  assign n16160 = n16159 ^ n15752 ;
  assign n16161 = n15756 ^ x81 ;
  assign n16162 = ~n16095 & n16161 ;
  assign n16163 = n16162 ^ n15759 ;
  assign n16164 = n15763 ^ x82 ;
  assign n16165 = ~n16095 & n16164 ;
  assign n16166 = n16165 ^ n15766 ;
  assign n16167 = n15770 ^ x83 ;
  assign n16168 = ~n16095 & n16167 ;
  assign n16169 = n16168 ^ n15773 ;
  assign n16170 = n15777 ^ x84 ;
  assign n16171 = ~n16095 & n16170 ;
  assign n16172 = n16171 ^ n15780 ;
  assign n16173 = n15784 ^ x85 ;
  assign n16174 = ~n16095 & n16173 ;
  assign n16175 = n16174 ^ n15787 ;
  assign n16176 = n15791 ^ x86 ;
  assign n16177 = ~n16095 & n16176 ;
  assign n16178 = n16177 ^ n15622 ;
  assign n16179 = n15622 ^ x87 ;
  assign n16180 = n16179 ^ x86 ;
  assign n16181 = n16180 ^ n15791 ;
  assign n16182 = n16181 ^ n16179 ;
  assign n16185 = n16179 ^ n2532 ;
  assign n16186 = ~n16182 & ~n16185 ;
  assign n16187 = n16186 ^ n16179 ;
  assign n16188 = ~n16095 & ~n16187 ;
  assign n16189 = n16188 ^ n15618 ;
  assign n16190 = n15797 ^ x88 ;
  assign n16191 = ~n16095 & n16190 ;
  assign n16192 = n16191 ^ n15800 ;
  assign n16193 = n15804 ^ x89 ;
  assign n16194 = ~n16095 & n16193 ;
  assign n16195 = n16194 ^ n15807 ;
  assign n16196 = n15811 ^ x90 ;
  assign n16197 = ~n16095 & n16196 ;
  assign n16198 = n16197 ^ n15814 ;
  assign n16199 = n15818 ^ x91 ;
  assign n16200 = ~n16095 & n16199 ;
  assign n16201 = n16200 ^ n15821 ;
  assign n16202 = n15825 ^ x92 ;
  assign n16203 = ~n16095 & n16202 ;
  assign n16204 = n16203 ^ n15828 ;
  assign n16205 = n15832 ^ x93 ;
  assign n16206 = ~n16095 & n16205 ;
  assign n16207 = n16206 ^ n15835 ;
  assign n16208 = n15839 ^ x94 ;
  assign n16209 = ~n16095 & n16208 ;
  assign n16210 = n16209 ^ n15842 ;
  assign n16211 = n15846 ^ x95 ;
  assign n16212 = ~n16095 & n16211 ;
  assign n16213 = n16212 ^ n15849 ;
  assign n16214 = n15853 ^ x96 ;
  assign n16215 = ~n16095 & n16214 ;
  assign n16216 = n16215 ^ n15856 ;
  assign n16217 = n15860 ^ x97 ;
  assign n16218 = ~n16095 & n16217 ;
  assign n16219 = n16218 ^ n15863 ;
  assign n16220 = n15867 ^ x98 ;
  assign n16221 = ~n16095 & n16220 ;
  assign n16222 = n16221 ^ n15870 ;
  assign n16223 = n15874 ^ x99 ;
  assign n16224 = ~n16095 & n16223 ;
  assign n16225 = n16224 ^ n15877 ;
  assign n16226 = n15881 ^ x100 ;
  assign n16227 = ~n16095 & n16226 ;
  assign n16228 = n16227 ^ n15884 ;
  assign n16229 = n15888 ^ x101 ;
  assign n16230 = ~n16095 & n16229 ;
  assign n16231 = n16230 ^ n15891 ;
  assign n16232 = n15895 ^ x102 ;
  assign n16233 = ~n16095 & n16232 ;
  assign n16234 = n16233 ^ n15898 ;
  assign n16235 = n15902 ^ x103 ;
  assign n16236 = ~n16095 & n16235 ;
  assign n16237 = n16236 ^ n15905 ;
  assign n16238 = n15909 ^ x104 ;
  assign n16239 = ~n16095 & n16238 ;
  assign n16240 = n16239 ^ n15912 ;
  assign n16241 = n15916 ^ x105 ;
  assign n16242 = ~n16095 & n16241 ;
  assign n16243 = n16242 ^ n15919 ;
  assign n16244 = n15923 ^ x106 ;
  assign n16245 = ~n16095 & n16244 ;
  assign n16246 = n16245 ^ n15926 ;
  assign n16247 = n15930 ^ x107 ;
  assign n16248 = ~n16095 & n16247 ;
  assign n16249 = n16248 ^ n15933 ;
  assign n16250 = n15937 ^ x108 ;
  assign n16251 = ~n16095 & n16250 ;
  assign n16252 = n16251 ^ n15940 ;
  assign n16253 = n15944 ^ x109 ;
  assign n16254 = ~n16095 & n16253 ;
  assign n16255 = n16254 ^ n15947 ;
  assign n16256 = n15951 ^ x110 ;
  assign n16257 = ~n16095 & n16256 ;
  assign n16258 = n16257 ^ n15954 ;
  assign n16259 = n15958 ^ x111 ;
  assign n16260 = ~n16095 & n16259 ;
  assign n16261 = n16260 ^ n15961 ;
  assign n16262 = n15965 ^ x112 ;
  assign n16263 = ~n16095 & n16262 ;
  assign n16264 = n16263 ^ n15968 ;
  assign n16265 = n15972 ^ x113 ;
  assign n16266 = ~n16095 & n16265 ;
  assign n16267 = n16266 ^ n15975 ;
  assign n16268 = n15979 ^ x114 ;
  assign n16269 = ~n16095 & n16268 ;
  assign n16270 = n16269 ^ n15982 ;
  assign n16271 = n15986 ^ x115 ;
  assign n16272 = ~n16095 & n16271 ;
  assign n16273 = n16272 ^ n15997 ;
  assign n16274 = n16001 ^ x116 ;
  assign n16275 = ~n16095 & n16274 ;
  assign n16276 = n16275 ^ n16004 ;
  assign n16277 = n16008 ^ x117 ;
  assign n16278 = ~n16095 & n16277 ;
  assign n16279 = n16278 ^ n16011 ;
  assign n16280 = n16015 ^ x118 ;
  assign n16281 = ~n16095 & n16280 ;
  assign n16282 = n16281 ^ n16018 ;
  assign n16283 = n16022 ^ x119 ;
  assign n16284 = ~n16095 & n16283 ;
  assign n16285 = n16284 ^ n16025 ;
  assign n16286 = n16029 ^ x120 ;
  assign n16287 = ~n16095 & n16286 ;
  assign n16288 = n16287 ^ n16040 ;
  assign n16289 = n16044 ^ x121 ;
  assign n16290 = ~n16095 & n16289 ;
  assign n16291 = n16290 ^ n16047 ;
  assign n16292 = n16051 ^ x122 ;
  assign n16293 = ~n16095 & n16292 ;
  assign n16294 = n16293 ^ n16054 ;
  assign n16295 = n16058 ^ x123 ;
  assign n16296 = ~n16095 & n16295 ;
  assign n16297 = n16296 ^ n16061 ;
  assign n16298 = n16065 ^ x124 ;
  assign n16299 = ~n16095 & n16298 ;
  assign n16300 = n16299 ^ n16068 ;
  assign n16301 = n16072 ^ x125 ;
  assign n16302 = ~n16095 & n16301 ;
  assign n16303 = n16302 ^ n16075 ;
  assign n16304 = n16079 ^ x126 ;
  assign n16305 = ~n16095 & n16304 ;
  assign n16306 = n16305 ^ n16082 ;
  assign n16307 = n15301 & ~n16087 ;
  assign n16308 = n15611 & n16307 ;
  assign n16309 = ~n16086 & n16308 ;
  assign n16310 = n16309 ^ n16307 ;
  assign y0 = ~n16095 ;
  assign y1 = n15616 ;
  assign y2 = n15123 ;
  assign y3 = n14632 ;
  assign y4 = n14165 ;
  assign y5 = n13710 ;
  assign y6 = n13277 ;
  assign y7 = n12847 ;
  assign y8 = n12413 ;
  assign y9 = n11973 ;
  assign y10 = n11508 ;
  assign y11 = n11106 ;
  assign y12 = n10662 ;
  assign y13 = n10273 ;
  assign y14 = n9852 ;
  assign y15 = n9479 ;
  assign y16 = n9100 ;
  assign y17 = n8723 ;
  assign y18 = n8360 ;
  assign y19 = ~n8010 ;
  assign y20 = n7650 ;
  assign y21 = n7295 ;
  assign y22 = n6935 ;
  assign y23 = n6618 ;
  assign y24 = n6316 ;
  assign y25 = n6015 ;
  assign y26 = n5697 ;
  assign y27 = n5377 ;
  assign y28 = n5079 ;
  assign y29 = n4818 ;
  assign y30 = n4569 ;
  assign y31 = n4324 ;
  assign y32 = n4069 ;
  assign y33 = n3834 ;
  assign y34 = n3583 ;
  assign y35 = n3350 ;
  assign y36 = n3145 ;
  assign y37 = n2941 ;
  assign y38 = n2735 ;
  assign y39 = n2548 ;
  assign y40 = n2372 ;
  assign y41 = n2194 ;
  assign y42 = n2032 ;
  assign y43 = n1882 ;
  assign y44 = n1726 ;
  assign y45 = n1581 ;
  assign y46 = n1456 ;
  assign y47 = n1327 ;
  assign y48 = n1212 ;
  assign y49 = n1111 ;
  assign y50 = n1004 ;
  assign y51 = n908 ;
  assign y52 = n816 ;
  assign y53 = n727 ;
  assign y54 = n639 ;
  assign y55 = n555 ;
  assign y56 = n486 ;
  assign y57 = n431 ;
  assign y58 = n372 ;
  assign y59 = n330 ;
  assign y60 = n284 ;
  assign y61 = n254 ;
  assign y62 = n16096 ;
  assign y63 = n16100 ;
  assign y64 = n16102 ;
  assign y65 = n16109 ;
  assign y66 = n16111 ;
  assign y67 = n16113 ;
  assign y68 = n16116 ;
  assign y69 = n16119 ;
  assign y70 = n16122 ;
  assign y71 = n16125 ;
  assign y72 = n16128 ;
  assign y73 = n16131 ;
  assign y74 = n16134 ;
  assign y75 = n16137 ;
  assign y76 = n16140 ;
  assign y77 = n16151 ;
  assign y78 = n16154 ;
  assign y79 = n16157 ;
  assign y80 = n16160 ;
  assign y81 = n16163 ;
  assign y82 = n16166 ;
  assign y83 = n16169 ;
  assign y84 = n16172 ;
  assign y85 = n16175 ;
  assign y86 = n16178 ;
  assign y87 = n16189 ;
  assign y88 = n16192 ;
  assign y89 = n16195 ;
  assign y90 = n16198 ;
  assign y91 = n16201 ;
  assign y92 = n16204 ;
  assign y93 = n16207 ;
  assign y94 = n16210 ;
  assign y95 = n16213 ;
  assign y96 = n16216 ;
  assign y97 = n16219 ;
  assign y98 = n16222 ;
  assign y99 = n16225 ;
  assign y100 = n16228 ;
  assign y101 = n16231 ;
  assign y102 = n16234 ;
  assign y103 = n16237 ;
  assign y104 = n16240 ;
  assign y105 = n16243 ;
  assign y106 = n16246 ;
  assign y107 = n16249 ;
  assign y108 = n16252 ;
  assign y109 = n16255 ;
  assign y110 = n16258 ;
  assign y111 = n16261 ;
  assign y112 = n16264 ;
  assign y113 = n16267 ;
  assign y114 = n16270 ;
  assign y115 = n16273 ;
  assign y116 = n16276 ;
  assign y117 = n16279 ;
  assign y118 = n16282 ;
  assign y119 = n16285 ;
  assign y120 = n16288 ;
  assign y121 = n16291 ;
  assign y122 = n16294 ;
  assign y123 = n16297 ;
  assign y124 = n16300 ;
  assign y125 = n16303 ;
  assign y126 = n16306 ;
  assign y127 = n16310 ;
endmodule
