module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n168 , n169 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3518 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3980 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4401 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4433 , n4434 , n4435 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4655 , n4656 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4882 , n4883 , n4884 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4992 , n4993 , n4994 , n4995 , n4996 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5220 , n5221 , n5224 , n5225 , n5226 , n5232 , n5233 , n5234 , n5235 , n5239 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5888 , n5889 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6015 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6145 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6736 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6846 , n6847 , n6848 , n6849 , n6850 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6870 , n6871 , n6872 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7157 , n7158 , n7159 , n7160 , n7161 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7310 , n7311 , n7312 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7433 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7688 , n7691 , n7692 , n7693 , n7694 , n7695 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7824 , n7825 , n7826 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8484 , n8485 , n8486 , n8487 , n8489 , n8490 , n8491 , n8492 , n8493 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8583 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8835 , n8836 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8860 , n8861 , n8862 , n8863 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8976 , n8977 , n8978 , n8979 , n8980 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9067 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9400 , n9401 , n9402 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9611 , n9612 , n9613 , n9615 , n9616 , n9617 , n9619 , n9620 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9645 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9811 , n9812 , n9813 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9896 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10407 , n10408 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10662 , n10672 , n10674 , n10677 , n10678 , n10679 , n10680 , n10682 , n10684 , n10688 , n10698 , n10699 , n10700 , n10701 , n10703 , n10706 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10742 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11029 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11152 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11235 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11310 , n11311 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11330 , n11331 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11349 , n11350 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11667 , n11671 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11709 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12020 , n12021 , n12022 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12192 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12413 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12434 , n12435 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12805 , n12806 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12939 , n12940 , n12941 , n12942 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13084 , n13085 , n13086 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13119 , n13120 , n13121 , n13125 , n13126 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13197 , n13201 , n13202 , n13203 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13214 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14095 , n14096 , n14097 , n14098 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14435 , n14436 , n14437 , n14438 , n14439 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14554 , n14555 , n14556 , n14557 , n14558 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15798 , n15799 , n15800 , n15801 , n15802 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17125 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17178 , n17179 , n17180 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17260 , n17261 , n17262 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17328 , n17329 , n17330 , n17334 , n17335 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17353 , n17359 , n17360 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17604 , n17609 , n17610 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19042 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19289 , n19290 , n19291 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19342 , n19343 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19399 , n19400 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19472 , n19473 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19490 , n19491 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19506 , n19507 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19546 , n19547 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19587 , n19588 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19621 , n19622 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19726 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19882 , n19883 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20432 , n20433 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20649 , n20650 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20662 , n20663 , n20664 , n20665 , n20667 , n20668 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20788 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20922 , n20924 , n20925 , n20926 , n20927 , n20929 , n20930 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20943 , n20944 , n20946 , n20947 , n20948 , n20949 , n20951 , n20952 , n20953 , n20955 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20984 , n20985 , n20986 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21044 , n21045 , n21046 , n21049 , n21050 , n21051 , n21052 , n21053 , n21055 , n21058 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21257 , n21258 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21751 , n21752 , n21753 , n21754 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24104 , n24105 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24158 , n24159 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24268 , n24269 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24367 , n24368 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24447 , n24448 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25780 , n25781 , n25782 , n25783 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26780 , n26781 , n26782 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27741 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27890 , n27891 , n27892 , n27893 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28489 , n28490 , n28491 , n28492 , n28493 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29178 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29434 , n29435 , n29436 , n29437 , n29438 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 ;
  assign n52 = ~x29 & ~x30 ;
  assign n53 = x27 & x28 ;
  assign n54 = n53 ^ x27 ;
  assign n55 = n52 & n54 ;
  assign n72 = ~x23 & ~x24 ;
  assign n86 = ~x25 & n72 ;
  assign n75 = x25 ^ x24 ;
  assign n74 = x24 & x25 ;
  assign n76 = n75 ^ n74 ;
  assign n87 = n86 ^ n76 ;
  assign n154 = n87 ^ x24 ;
  assign n155 = n154 ^ n72 ;
  assign n203 = n155 ^ n74 ;
  assign n365 = ~x26 & ~n203 ;
  assign n366 = n55 & n365 ;
  assign n56 = ~x28 & n52 ;
  assign n57 = n56 ^ n55 ;
  assign n367 = n366 ^ n57 ;
  assign n48 = x25 & ~x26 ;
  assign n110 = x23 & n48 ;
  assign n102 = ~x24 & ~x26 ;
  assign n103 = n102 ^ x26 ;
  assign n79 = n76 ^ x26 ;
  assign n80 = n79 ^ n48 ;
  assign n77 = x26 & n76 ;
  assign n78 = n77 ^ x26 ;
  assign n81 = n80 ^ n78 ;
  assign n104 = n103 ^ n81 ;
  assign n96 = x24 ^ x23 ;
  assign n97 = x26 & ~n96 ;
  assign n98 = n97 ^ x26 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n99 ^ x26 ;
  assign n95 = ~x26 & n72 ;
  assign n101 = n100 ^ n95 ;
  assign n105 = n104 ^ n101 ;
  assign n88 = ~x23 & ~x25 ;
  assign n89 = n88 ^ n87 ;
  assign n49 = n48 ^ x25 ;
  assign n50 = n49 ^ x26 ;
  assign n83 = n72 ^ x24 ;
  assign n84 = n83 ^ x23 ;
  assign n85 = n50 & n84 ;
  assign n90 = n89 ^ n85 ;
  assign n51 = n50 ^ x25 ;
  assign n91 = n90 ^ n51 ;
  assign n106 = n105 ^ n91 ;
  assign n107 = n106 ^ n104 ;
  assign n111 = n110 ^ n107 ;
  assign n156 = n155 ^ n111 ;
  assign n299 = n52 & n53 ;
  assign n362 = ~n156 & n299 ;
  assign n146 = n74 ^ x26 ;
  assign n147 = n146 ^ n104 ;
  assign n132 = n89 ^ x25 ;
  assign n133 = n132 ^ n84 ;
  assign n134 = n133 ^ x26 ;
  assign n135 = n134 ^ n107 ;
  assign n148 = n147 ^ n135 ;
  assign n347 = n55 & ~n148 ;
  assign n20601 = n135 ^ n86 ;
  assign n20600 = ~n86 & ~n135 ;
  assign n20602 = n20601 ^ n20600 ;
  assign n212 = ~n20602 ^ n78 ;
  assign n346 = n212 & n299 ;
  assign n348 = n347 ^ n346 ;
  assign n332 = n299 ^ n52 ;
  assign n333 = n332 ^ n56 ;
  assign n344 = ~n101 & n333 ;
  assign n190 = n77 ^ n49 ;
  assign n343 = n190 & n333 ;
  assign n345 = n344 ^ n343 ;
  assign n349 = n348 ^ n345 ;
  assign n139 = n95 ^ n72 ;
  assign n141 = ~n20602 ^ n139 ;
  assign n340 = n55 & n141 ;
  assign n152 = n85 ^ n50 ;
  assign n339 = n55 & n152 ;
  assign n341 = n340 ^ n339 ;
  assign n335 = ~n111 & n333 ;
  assign n115 = n102 ^ n95 ;
  assign n334 = n115 & n333 ;
  assign n336 = n335 ^ n334 ;
  assign n116 = n115 ^ n111 ;
  assign n331 = ~n116 & n299 ;
  assign n337 = n336 ^ n331 ;
  assign n191 = n190 ^ n152 ;
  assign n306 = n191 ^ n139 ;
  assign n305 = n132 ^ n48 ;
  assign n307 = n306 ^ n305 ;
  assign n308 = n299 & n307 ;
  assign n338 = n337 ^ n308 ;
  assign n342 = n341 ^ n338 ;
  assign n350 = n349 ^ n342 ;
  assign n354 = n55 & ~n156 ;
  assign n353 = ~n148 & n333 ;
  assign n355 = n354 ^ n353 ;
  assign n351 = ~x23 & ~n51 ;
  assign n352 = n299 & n351 ;
  assign n356 = n355 ^ n352 ;
  assign n136 = n135 ^ x26 ;
  assign n357 = n55 & n136 ;
  assign n358 = n357 ^ n345 ;
  assign n359 = n358 ^ n333 ;
  assign n360 = ~n356 & ~n359 ;
  assign n361 = ~n350 & n360 ;
  assign n363 = n362 ^ n361 ;
  assign n328 = n104 ^ n85 ;
  assign n329 = n55 & ~n328 ;
  assign n327 = n55 & ~n111 ;
  assign n330 = n329 ^ n327 ;
  assign n364 = n363 ^ n330 ;
  assign n368 = n367 ^ n364 ;
  assign n112 = n104 ^ n48 ;
  assign n113 = n112 ^ n111 ;
  assign n60 = n52 ^ x29 ;
  assign n131 = n53 & ~n60 ;
  assign n199 = n113 & n131 ;
  assign n197 = ~n111 & n131 ;
  assign n195 = n78 & n131 ;
  assign n182 = n106 & n131 ;
  assign n196 = n195 ^ n182 ;
  assign n198 = n197 ^ n196 ;
  assign n200 = n199 ^ n198 ;
  assign n192 = n131 & n191 ;
  assign n189 = n91 & n131 ;
  assign n193 = n192 ^ n189 ;
  assign n73 = n72 ^ x23 ;
  assign n82 = n81 ^ n73 ;
  assign n92 = n91 ^ n82 ;
  assign n93 = n92 ^ n73 ;
  assign n188 = n93 & n131 ;
  assign n194 = n193 ^ n188 ;
  assign n201 = n200 ^ n194 ;
  assign n59 = n53 ^ x28 ;
  assign n176 = n59 & ~n60 ;
  assign n174 = n54 & ~n60 ;
  assign n175 = n90 & n174 ;
  assign n177 = n176 ^ n175 ;
  assign n184 = n93 & n176 ;
  assign n181 = ~n104 & n131 ;
  assign n183 = n182 ^ n181 ;
  assign n185 = n184 ^ n183 ;
  assign n179 = n91 & n176 ;
  assign n178 = n93 & n174 ;
  assign n180 = n179 ^ n178 ;
  assign n186 = n185 ^ n180 ;
  assign n187 = ~n177 & ~n186 ;
  assign n202 = n201 ^ n187 ;
  assign n123 = n113 ^ n95 ;
  assign n215 = n123 & n131 ;
  assign n214 = ~n116 & n174 ;
  assign n216 = n215 ^ n214 ;
  assign n213 = n176 & n212 ;
  assign n217 = n216 ^ n213 ;
  assign n211 = n113 & n176 ;
  assign n218 = n217 ^ n211 ;
  assign n209 = ~n116 & n131 ;
  assign n204 = n102 ^ x24 ;
  assign n205 = ~n20602 ^ n204 ;
  assign n206 = n205 ^ x26 ;
  assign n207 = ~n203 & n206 ;
  assign n208 = n176 & ~n207 ;
  assign n210 = n209 ^ n208 ;
  assign n219 = n218 ^ n210 ;
  assign n220 = n202 & ~n219 ;
  assign n231 = n57 & n110 ;
  assign n1239 = x24 & n231 ;
  assign n61 = n60 ^ x30 ;
  assign n66 = n53 & ~n61 ;
  assign n171 = n66 & n106 ;
  assign n172 = n1239 ^ n171 ;
  assign n162 = x26 & ~n88 ;
  assign n165 = n66 & n92 ;
  assign n168 = n162 & n165 ;
  assign n67 = n66 ^ n61 ;
  assign n63 = ~x27 & ~n61 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = ~n49 & ~n68 ;
  assign n163 = n69 ^ n68 ;
  assign n62 = n59 & ~n61 ;
  assign n127 = n68 ^ n62 ;
  assign n128 = n49 & ~n127 ;
  assign n164 = n163 ^ n128 ;
  assign n166 = n165 ^ n164 ;
  assign n169 = n168 ^ n166 ;
  assign n173 = n172 ^ n169 ;
  assign n221 = n220 ^ n173 ;
  assign n157 = n131 & ~n156 ;
  assign n153 = n131 & n152 ;
  assign n158 = n157 ^ n153 ;
  assign n149 = n131 & ~n148 ;
  assign n64 = n63 ^ n62 ;
  assign n145 = n64 & n113 ;
  assign n150 = n149 ^ n145 ;
  assign n142 = n131 & n141 ;
  assign n138 = n64 & ~n111 ;
  assign n143 = n142 ^ n138 ;
  assign n137 = n131 & n136 ;
  assign n144 = n143 ^ n137 ;
  assign n151 = n150 ^ n144 ;
  assign n159 = n158 ^ n151 ;
  assign n129 = n128 ^ n62 ;
  assign n125 = n64 & n106 ;
  assign n124 = n64 & n123 ;
  assign n126 = n125 ^ n124 ;
  assign n130 = n129 ^ n126 ;
  assign n160 = n159 ^ n130 ;
  assign n118 = n64 & n91 ;
  assign n117 = n64 & ~n116 ;
  assign n119 = n118 ^ n117 ;
  assign n114 = n57 & n113 ;
  assign n120 = n119 ^ n114 ;
  assign n108 = n64 & ~n107 ;
  assign n94 = n64 & n93 ;
  assign n109 = n108 ^ n94 ;
  assign n121 = n120 ^ n109 ;
  assign n65 = x26 & n64 ;
  assign n70 = n69 ^ n65 ;
  assign n58 = ~n51 & n57 ;
  assign n71 = n70 ^ n58 ;
  assign n122 = n121 ^ n71 ;
  assign n161 = n160 ^ n122 ;
  assign n222 = n221 ^ n161 ;
  assign n1689 = x25 & n344 ;
  assign n403 = n354 ^ n341 ;
  assign n300 = x26 & n299 ;
  assign n301 = n74 & n300 ;
  assign n223 = n61 ^ x29 ;
  assign n227 = n59 ^ x27 ;
  assign n298 = ~n223 & ~n227 ;
  assign n302 = n301 ^ n298 ;
  assign n260 = n54 & ~n223 ;
  assign n380 = n91 & n260 ;
  assign n267 = n81 & n260 ;
  assign n390 = n380 ^ n267 ;
  assign n389 = n113 & n260 ;
  assign n391 = n390 ^ n389 ;
  assign n387 = n347 ^ n336 ;
  assign n385 = n123 & n333 ;
  assign n386 = n385 ^ n357 ;
  assign n388 = n387 ^ n386 ;
  assign n392 = n391 ^ n388 ;
  assign n382 = ~n148 & n298 ;
  assign n296 = n123 & n260 ;
  assign n383 = n382 ^ n296 ;
  assign n378 = ~n116 & n260 ;
  assign n377 = n93 & n333 ;
  assign n379 = n378 ^ n377 ;
  assign n381 = n380 ^ n379 ;
  assign n384 = n383 ^ n381 ;
  assign n393 = n392 ^ n384 ;
  assign n394 = ~n302 & ~n393 ;
  assign n399 = n113 & n333 ;
  assign n398 = n106 & n333 ;
  assign n400 = n399 ^ n398 ;
  assign n395 = n191 & n298 ;
  assign n396 = n395 ^ n335 ;
  assign n369 = n91 & n333 ;
  assign n397 = n396 ^ n369 ;
  assign n401 = n400 ^ n397 ;
  assign n402 = n394 & ~n401 ;
  assign n404 = n403 ^ n402 ;
  assign n405 = n404 ^ n329 ;
  assign n252 = n62 & ~n148 ;
  assign n251 = n62 & n141 ;
  assign n253 = n252 ^ n251 ;
  assign n232 = n1239 ^ n231 ;
  assign n373 = n253 ^ n232 ;
  assign n270 = n110 & n260 ;
  assign n374 = n373 ^ n270 ;
  assign n234 = n57 & n106 ;
  assign n375 = n374 ^ n234 ;
  assign n371 = n147 ^ n106 ;
  assign n372 = n260 & ~n371 ;
  assign n376 = n375 ^ n372 ;
  assign n406 = n405 ^ n376 ;
  assign n407 = n1689 ^ n406 ;
  assign n408 = ~n222 & n407 ;
  assign n446 = ~n148 & n260 ;
  assign n447 = n446 ^ n403 ;
  assign n264 = n59 & ~n223 ;
  assign n444 = ~n116 & n264 ;
  assign n445 = n444 ^ n189 ;
  assign n448 = n447 ^ n445 ;
  assign n322 = n57 & n123 ;
  assign n224 = n53 & ~n223 ;
  assign n320 = n93 & n224 ;
  assign n318 = ~n116 & n224 ;
  assign n317 = n91 & n224 ;
  assign n319 = n318 ^ n317 ;
  assign n321 = n320 ^ n319 ;
  assign n323 = n322 ^ n321 ;
  assign n449 = n448 ^ n323 ;
  assign n440 = n123 & n264 ;
  assign n256 = n57 & ~n20602 ;
  assign n441 = n440 ^ n256 ;
  assign n409 = n136 & n299 ;
  assign n437 = n409 ^ n301 ;
  assign n436 = ~n116 & n298 ;
  assign n438 = n437 ^ n436 ;
  assign n434 = n136 & n260 ;
  assign n435 = n434 ^ n199 ;
  assign n439 = n438 ^ n435 ;
  assign n442 = n441 ^ n439 ;
  assign n430 = n57 & ~n116 ;
  assign n429 = n57 & ~n148 ;
  assign n431 = n430 ^ n429 ;
  assign n432 = n431 ^ n177 ;
  assign n265 = n93 & n264 ;
  assign n427 = n265 ^ n183 ;
  assign n426 = n214 ^ n178 ;
  assign n428 = n427 ^ n426 ;
  assign n433 = n432 ^ n428 ;
  assign n443 = n442 ^ n433 ;
  assign n450 = n449 ^ n443 ;
  assign n422 = n57 & n190 ;
  assign n419 = n136 & n264 ;
  assign n275 = n113 & n224 ;
  assign n273 = n95 & n224 ;
  assign n274 = n273 ^ n224 ;
  assign n276 = n275 ^ n274 ;
  assign n277 = n276 ^ n224 ;
  assign n420 = n419 ^ n277 ;
  assign n243 = n57 & n212 ;
  assign n421 = n420 ^ n243 ;
  assign n423 = n422 ^ n421 ;
  assign n416 = n113 & n298 ;
  assign n415 = n95 & n298 ;
  assign n417 = n416 ^ n415 ;
  assign n413 = n56 & n141 ;
  assign n414 = n413 ^ n340 ;
  assign n418 = n417 ^ n414 ;
  assign n424 = n423 ^ n418 ;
  assign n411 = n57 & ~n156 ;
  assign n410 = n409 ^ n198 ;
  assign n412 = n411 ^ n410 ;
  assign n425 = n424 ^ n412 ;
  assign n451 = n450 ^ n425 ;
  assign n533 = n123 & n299 ;
  assign n484 = n264 & ~n20602 ;
  assign n534 = n533 ^ n484 ;
  assign n248 = n66 & ~n148 ;
  assign n535 = n534 ^ n248 ;
  assign n519 = n152 & n264 ;
  assign n536 = n535 ^ n519 ;
  assign n530 = n416 ^ n188 ;
  assign n279 = x23 & n264 ;
  assign n527 = ~n104 & n279 ;
  assign n526 = n152 & n298 ;
  assign n528 = n527 ^ n526 ;
  assign n529 = n528 ^ n215 ;
  assign n531 = n530 ^ n529 ;
  assign n523 = n55 & n106 ;
  assign n522 = ~n156 & n264 ;
  assign n524 = n523 ^ n522 ;
  assign n518 = n132 & n264 ;
  assign n520 = n519 ^ n518 ;
  assign n517 = n106 & n264 ;
  assign n521 = n520 ^ n517 ;
  assign n525 = n524 ^ n521 ;
  assign n532 = n531 ^ n525 ;
  assign n537 = n536 ^ n532 ;
  assign n513 = n141 & n298 ;
  assign n514 = n513 ^ n395 ;
  assign n511 = n212 & n298 ;
  assign n510 = n353 ^ n184 ;
  assign n512 = n511 ^ n510 ;
  assign n515 = n514 ^ n512 ;
  assign n1209 = x23 & n343 ;
  assign n507 = n1209 ^ n343 ;
  assign n506 = n136 & n333 ;
  assign n508 = n507 ^ n506 ;
  assign n504 = n55 & ~n20602 ;
  assign n505 = n504 ^ n211 ;
  assign n509 = n508 ^ n505 ;
  assign n516 = n515 ^ n509 ;
  assign n538 = n537 ^ n516 ;
  assign n269 = n139 & n264 ;
  assign n485 = n484 ^ n269 ;
  assign n480 = n55 & n212 ;
  assign n478 = n212 & n333 ;
  assign n247 = n66 & n212 ;
  assign n479 = n478 ^ n247 ;
  assign n481 = n480 ^ n479 ;
  assign n483 = n1209 ^ n481 ;
  assign n486 = n485 ^ n483 ;
  assign n476 = n91 & n298 ;
  assign n240 = n66 & n136 ;
  assign n239 = n66 & n152 ;
  assign n241 = n240 ^ n239 ;
  assign n237 = n66 & n191 ;
  assign n236 = n66 & n141 ;
  assign n238 = n237 ^ n236 ;
  assign n242 = n241 ^ n238 ;
  assign n477 = n476 ^ n242 ;
  assign n487 = n486 ^ n477 ;
  assign n471 = ~n148 & n264 ;
  assign n470 = n113 & n264 ;
  assign n472 = n471 ^ n470 ;
  assign n468 = n191 & n264 ;
  assign n469 = n468 ^ n213 ;
  assign n473 = n472 ^ n469 ;
  assign n465 = ~n111 & n264 ;
  assign n464 = n212 & n264 ;
  assign n466 = n465 ^ n464 ;
  assign n462 = n93 & n298 ;
  assign n250 = n66 & ~n156 ;
  assign n463 = n462 ^ n250 ;
  assign n467 = n466 ^ n463 ;
  assign n474 = n473 ^ n467 ;
  assign n459 = ~n107 & n176 ;
  assign n457 = n86 & n333 ;
  assign n458 = n457 ^ n385 ;
  assign n460 = n459 ^ n458 ;
  assign n455 = n55 & ~n107 ;
  assign n453 = n298 & ~n20602 ;
  assign n452 = n141 & n333 ;
  assign n454 = n453 ^ n452 ;
  assign n456 = n455 ^ n454 ;
  assign n461 = n460 ^ n456 ;
  assign n475 = n474 ^ n461 ;
  assign n488 = n487 ^ n475 ;
  assign n501 = n141 & n176 ;
  assign n498 = ~n156 & n333 ;
  assign n495 = ~n111 & n298 ;
  assign n493 = n106 & n298 ;
  assign n494 = n493 ^ n331 ;
  assign n496 = n495 ^ n494 ;
  assign n490 = n55 & n191 ;
  assign n489 = ~n107 & n298 ;
  assign n491 = n490 ^ n489 ;
  assign n492 = n491 ^ n179 ;
  assign n497 = n496 ^ n492 ;
  assign n499 = n498 ^ n497 ;
  assign n500 = n499 ^ n210 ;
  assign n502 = n501 ^ n500 ;
  assign n503 = ~n488 & ~n502 ;
  assign n539 = n538 ^ n503 ;
  assign n540 = ~n451 & n539 ;
  assign n577 = n55 & ~n116 ;
  assign n575 = n57 & n136 ;
  assign n576 = n575 ^ n114 ;
  assign n578 = n577 ^ n576 ;
  assign n579 = n578 ^ n192 ;
  assign n580 = n579 ^ n426 ;
  assign n571 = ~n133 & n298 ;
  assign n572 = n571 ^ n489 ;
  assign n570 = ~n68 & n113 ;
  assign n573 = n572 ^ n570 ;
  assign n567 = n93 & n299 ;
  assign n566 = ~n107 & n299 ;
  assign n568 = n567 ^ n566 ;
  assign n569 = n568 ^ n527 ;
  assign n574 = n573 ^ n569 ;
  assign n581 = n580 ^ n574 ;
  assign n563 = ~n156 & n298 ;
  assign n562 = n55 & n123 ;
  assign n564 = n563 ^ n562 ;
  assign n558 = n57 & ~n77 ;
  assign n559 = n558 ^ n58 ;
  assign n312 = n57 & n79 ;
  assign n560 = n559 ^ n312 ;
  assign n556 = n91 & n299 ;
  assign n555 = n113 & n299 ;
  assign n557 = n556 ^ n555 ;
  assign n561 = n560 ^ n557 ;
  assign n565 = n564 ^ n561 ;
  assign n582 = n581 ^ n565 ;
  assign n550 = ~n111 & n299 ;
  assign n551 = n550 ^ n465 ;
  assign n547 = n106 & n299 ;
  assign n546 = ~n68 & n91 ;
  assign n548 = n547 ^ n546 ;
  assign n549 = n548 ^ n484 ;
  assign n552 = n551 ^ n549 ;
  assign n228 = ~n60 & ~n227 ;
  assign n542 = ~n111 & n228 ;
  assign n541 = n115 & n228 ;
  assign n543 = n542 ^ n541 ;
  assign n544 = n543 ^ n470 ;
  assign n545 = n544 ^ n521 ;
  assign n553 = n552 ^ n545 ;
  assign n554 = n553 ^ n393 ;
  assign n583 = n582 ^ n554 ;
  assign n690 = n110 & n224 ;
  assign n691 = n690 ^ n481 ;
  assign n688 = n110 & n174 ;
  assign n225 = x26 & n224 ;
  assign n915 = ~n87 & n225 ;
  assign n687 = n915 ^ n446 ;
  assign n689 = n688 ^ n687 ;
  assign n692 = n691 ^ n689 ;
  assign n684 = n174 & n212 ;
  assign n682 = n64 & ~n148 ;
  assign n680 = ~n68 & n123 ;
  assign n681 = n680 ^ n125 ;
  assign n683 = n682 ^ n681 ;
  assign n685 = n684 ^ n683 ;
  assign n693 = n692 ^ n685 ;
  assign n677 = n64 & ~n20602 ;
  assign n678 = n677 ^ n438 ;
  assign n675 = n132 & n225 ;
  assign n676 = n675 ^ n343 ;
  assign n679 = n678 ^ n676 ;
  assign n694 = n693 ^ n679 ;
  assign n670 = n256 ^ n124 ;
  assign n671 = n670 ^ n137 ;
  assign n672 = n671 ^ n434 ;
  assign n667 = n64 & ~n133 ;
  assign n668 = n667 ^ n108 ;
  assign n664 = n123 & n228 ;
  assign n663 = n123 & n176 ;
  assign n665 = n664 ^ n663 ;
  assign n666 = n665 ^ n142 ;
  assign n669 = n668 ^ n666 ;
  assign n673 = n672 ^ n669 ;
  assign n659 = n64 & n191 ;
  assign n660 = n659 ^ n243 ;
  assign n657 = n113 & n174 ;
  assign n658 = n657 ^ n250 ;
  assign n661 = n660 ^ n658 ;
  assign n655 = ~n156 & n174 ;
  assign n653 = n91 & n174 ;
  assign n654 = n653 ^ n149 ;
  assign n656 = n655 ^ n654 ;
  assign n662 = n661 ^ n656 ;
  assign n674 = n673 ^ n662 ;
  assign n695 = n694 ^ n674 ;
  assign n649 = n191 & n224 ;
  assign n647 = n504 ^ n145 ;
  assign n645 = n64 & n152 ;
  assign n646 = n645 ^ n240 ;
  assign n648 = n647 ^ n646 ;
  assign n650 = n649 ^ n648 ;
  assign n641 = n174 & n191 ;
  assign n640 = n136 & n224 ;
  assign n642 = n641 ^ n640 ;
  assign n643 = n642 ^ n476 ;
  assign n644 = n643 ^ n109 ;
  assign n651 = n650 ^ n644 ;
  assign n637 = n141 & n174 ;
  assign n636 = n239 ^ n184 ;
  assign n638 = n637 ^ n636 ;
  assign n634 = ~n156 & n224 ;
  assign n635 = n634 ^ n455 ;
  assign n639 = n638 ^ n635 ;
  assign n652 = n651 ^ n639 ;
  assign n696 = n695 ^ n652 ;
  assign n628 = ~n68 & ~n116 ;
  assign n1179 = n64 & n212 ;
  assign n627 = n1179 ^ n157 ;
  assign n629 = n628 ^ n627 ;
  assign n622 = n174 & ~n20602 ;
  assign n623 = n622 ^ n409 ;
  assign n624 = n623 ^ n523 ;
  assign n630 = n629 ^ n624 ;
  assign n975 = x23 & n422 ;
  assign n618 = n975 ^ n422 ;
  assign n619 = n618 ^ n462 ;
  assign n620 = n619 ^ n444 ;
  assign n621 = n620 ^ n238 ;
  assign n631 = n630 ^ n621 ;
  assign n615 = n106 & n224 ;
  assign n610 = n64 & n141 ;
  assign n609 = n106 & n174 ;
  assign n611 = n610 ^ n609 ;
  assign n612 = n611 ^ n248 ;
  assign n613 = n612 ^ n440 ;
  assign n614 = n613 ^ n265 ;
  assign n616 = n615 ^ n614 ;
  assign n632 = n631 ^ n616 ;
  assign n603 = n141 & n224 ;
  assign n602 = ~n148 & n224 ;
  assign n604 = n603 ^ n602 ;
  assign n600 = ~n68 & n93 ;
  assign n598 = n152 & n174 ;
  assign n226 = ~n86 & n225 ;
  assign n596 = n226 ^ n225 ;
  assign n597 = n596 ^ n275 ;
  assign n599 = n598 ^ n597 ;
  assign n601 = n600 ^ n599 ;
  assign n605 = n604 ^ n601 ;
  assign n594 = n138 ^ n118 ;
  assign n595 = n594 ^ n458 ;
  assign n606 = n605 ^ n595 ;
  assign n592 = n64 & ~n156 ;
  assign n589 = ~n148 & n174 ;
  assign n590 = n589 ^ n153 ;
  assign n591 = n590 ^ n117 ;
  assign n593 = n592 ^ n591 ;
  assign n607 = n606 ^ n593 ;
  assign n585 = n136 & n174 ;
  assign n584 = ~n116 & n176 ;
  assign n586 = n585 ^ n584 ;
  assign n587 = n586 ^ n452 ;
  assign n588 = n587 ^ n415 ;
  assign n608 = n607 ^ n588 ;
  assign n633 = n632 ^ n608 ;
  assign n697 = n696 ^ n633 ;
  assign n698 = ~n583 & ~n697 ;
  assign n755 = n414 ^ n339 ;
  assign n753 = n55 & n91 ;
  assign n754 = n753 ^ n192 ;
  assign n756 = n755 ^ n754 ;
  assign n750 = n62 & n93 ;
  assign n751 = n750 ^ n399 ;
  assign n752 = n751 ^ n241 ;
  assign n757 = n756 ^ n752 ;
  assign n747 = n493 ^ n250 ;
  assign n746 = n485 ^ n265 ;
  assign n748 = n747 ^ n746 ;
  assign n743 = n62 & n91 ;
  assign n744 = n743 ^ n490 ;
  assign n741 = n62 & n123 ;
  assign n742 = n741 ^ n434 ;
  assign n745 = n744 ^ n742 ;
  assign n749 = n748 ^ n745 ;
  assign n758 = n757 ^ n749 ;
  assign n737 = n55 & n93 ;
  assign n738 = n737 ^ n687 ;
  assign n735 = n58 & ~n73 ;
  assign n734 = n426 ^ n248 ;
  assign n736 = n735 ^ n734 ;
  assign n739 = n738 ^ n736 ;
  assign n730 = n191 & n299 ;
  assign n731 = n730 ^ n383 ;
  assign n732 = n731 ^ n440 ;
  assign n733 = n975 ^ n732 ;
  assign n740 = n739 ^ n733 ;
  assign n759 = n758 ^ n740 ;
  assign n725 = n57 & n91 ;
  assign n722 = n299 & ~n20602 ;
  assign n721 = n62 & n113 ;
  assign n723 = n722 ^ n721 ;
  assign n724 = n723 ^ n179 ;
  assign n726 = n725 ^ n724 ;
  assign n719 = n62 & ~n116 ;
  assign n716 = ~n111 & n176 ;
  assign n717 = n716 ^ n444 ;
  assign n718 = n717 ^ n211 ;
  assign n720 = n719 ^ n718 ;
  assign n727 = n726 ^ n720 ;
  assign n714 = n468 ^ n236 ;
  assign n712 = n353 ^ n243 ;
  assign n707 = ~n68 & ~n84 ;
  assign n709 = n707 ^ n546 ;
  assign n285 = x26 ^ x25 ;
  assign n708 = n285 & n707 ;
  assign n710 = n709 ^ n708 ;
  assign n706 = n62 & ~n111 ;
  assign n711 = n710 ^ n706 ;
  assign n713 = n712 ^ n711 ;
  assign n715 = n714 ^ n713 ;
  assign n728 = n727 ^ n715 ;
  assign n703 = n522 ^ n498 ;
  assign n701 = n571 ^ n519 ;
  assign n702 = n701 ^ n346 ;
  assign n704 = n703 ^ n702 ;
  assign n699 = n495 ^ n369 ;
  assign n700 = n699 ^ n649 ;
  assign n705 = n704 ^ n700 ;
  assign n729 = n728 ^ n705 ;
  assign n760 = n759 ^ n729 ;
  assign n847 = ~n68 & n106 ;
  assign n848 = n847 ^ n213 ;
  assign n791 = ~n107 & n224 ;
  assign n849 = n848 ^ n791 ;
  assign n845 = n91 & n228 ;
  assign n846 = n845 ^ n94 ;
  assign n850 = n849 ^ n846 ;
  assign n842 = n48 & n707 ;
  assign n843 = n842 ^ n542 ;
  assign n844 = n843 ^ n322 ;
  assign n851 = n850 ^ n844 ;
  assign n838 = ~n68 & ~n156 ;
  assign n839 = n838 ^ n458 ;
  assign n840 = n839 ^ n409 ;
  assign n836 = n176 & ~n20602 ;
  assign n837 = n836 ^ n158 ;
  assign n841 = n840 ^ n837 ;
  assign n852 = n851 ^ n841 ;
  assign n831 = n176 & n191 ;
  assign n832 = n831 ^ n464 ;
  assign n830 = n453 ^ n275 ;
  assign n833 = n832 ^ n830 ;
  assign n272 = n212 & n260 ;
  assign n829 = n272 ^ n118 ;
  assign n834 = n833 ^ n829 ;
  assign n825 = n113 & n228 ;
  assign n826 = n825 ^ n455 ;
  assign n827 = n826 ^ n622 ;
  assign n828 = n827 ^ n564 ;
  assign n835 = n834 ^ n828 ;
  assign n853 = n852 ^ n835 ;
  assign n820 = ~n68 & ~n148 ;
  assign n821 = n820 ^ n684 ;
  assign n822 = n821 ^ n256 ;
  assign n818 = n106 & n176 ;
  assign n819 = n818 ^ n556 ;
  assign n823 = n822 ^ n819 ;
  assign n815 = n106 & n260 ;
  assign n816 = n815 ^ n347 ;
  assign n813 = ~n68 & n152 ;
  assign n814 = n813 ^ n615 ;
  assign n817 = n816 ^ n814 ;
  assign n824 = n823 ^ n817 ;
  assign n854 = n853 ^ n824 ;
  assign n805 = ~n68 & n141 ;
  assign n806 = n805 ^ n501 ;
  assign n807 = n806 ^ n232 ;
  assign n808 = n807 ^ n575 ;
  assign n803 = n260 & ~n20602 ;
  assign n769 = ~n104 & n174 ;
  assign n770 = n769 ^ n609 ;
  assign n801 = n770 ^ n688 ;
  assign n800 = ~n156 & n176 ;
  assign n802 = n801 ^ n800 ;
  assign n804 = n803 ^ n802 ;
  assign n809 = n808 ^ n804 ;
  assign n798 = n234 ^ n117 ;
  assign n799 = n798 ^ n609 ;
  assign n810 = n809 ^ n799 ;
  assign n794 = n653 ^ n459 ;
  assign n795 = n794 ^ n479 ;
  assign n991 = ~x24 & n690 ;
  assign n793 = n991 ^ n417 ;
  assign n796 = n795 ^ n793 ;
  assign n788 = ~n68 & n212 ;
  assign n789 = n788 ^ n438 ;
  assign n784 = ~n68 & ~n111 ;
  assign n785 = n784 ^ n237 ;
  assign n786 = n785 ^ n270 ;
  assign n787 = n786 ^ n386 ;
  assign n790 = n789 ^ n787 ;
  assign n797 = n796 ^ n790 ;
  assign n811 = n810 ^ n797 ;
  assign n778 = n228 & ~n20602 ;
  assign n779 = n778 ^ n596 ;
  assign n776 = ~n68 & n191 ;
  assign n777 = n776 ^ n124 ;
  assign n780 = n779 ^ n777 ;
  assign n773 = ~n68 & ~n20602 ;
  assign n772 = n106 & n228 ;
  assign n774 = n773 ^ n772 ;
  assign n771 = n770 ^ n555 ;
  assign n775 = n774 ^ n771 ;
  assign n781 = n780 ^ n775 ;
  assign n782 = n781 ^ n151 ;
  assign n766 = n152 & n176 ;
  assign n764 = ~n107 & n228 ;
  assign n765 = n764 ^ n657 ;
  assign n767 = n766 ^ n765 ;
  assign n761 = n93 & n228 ;
  assign n762 = n761 ^ n567 ;
  assign n763 = n762 ^ n523 ;
  assign n768 = n767 ^ n763 ;
  assign n783 = n782 ^ n768 ;
  assign n812 = n811 ^ n783 ;
  assign n855 = n854 ^ n812 ;
  assign n856 = ~n760 & ~n855 ;
  assign n1040 = n610 ^ n153 ;
  assign n1041 = n1040 ^ n567 ;
  assign n1038 = n677 ^ n335 ;
  assign n1036 = n152 & n260 ;
  assign n1037 = n1036 ^ n815 ;
  assign n1039 = n1038 ^ n1037 ;
  assign n1042 = n1041 ^ n1039 ;
  assign n1034 = n659 ^ n637 ;
  assign n1032 = n975 ^ n178 ;
  assign n1033 = n1032 ^ n395 ;
  assign n1035 = n1034 ^ n1033 ;
  assign n1043 = n1042 ^ n1035 ;
  assign n956 = n62 & n152 ;
  assign n1028 = n956 ^ n722 ;
  assign n1027 = n550 ^ n237 ;
  assign n1029 = n1028 ^ n1027 ;
  assign n1026 = n825 ^ n813 ;
  assign n1030 = n1029 ^ n1026 ;
  assign n1024 = n603 ^ n188 ;
  assign n1020 = n55 & n113 ;
  assign n1021 = n1020 ^ n575 ;
  assign n1022 = n1021 ^ n179 ;
  assign n1023 = n1022 ^ n655 ;
  assign n1025 = n1024 ^ n1023 ;
  assign n1031 = n1030 ^ n1025 ;
  assign n1044 = n1043 ^ n1031 ;
  assign n1015 = n437 ^ n125 ;
  assign n1016 = n1015 ^ n340 ;
  assign n1014 = n62 & ~n156 ;
  assign n1017 = n1016 ^ n1014 ;
  assign n1011 = n465 ^ n214 ;
  assign n1012 = n1011 ^ n598 ;
  assign n1013 = n1012 ^ n533 ;
  assign n1018 = n1017 ^ n1013 ;
  assign n1008 = n141 & n299 ;
  assign n1009 = n1008 ^ n149 ;
  assign n1010 = n1009 ^ n508 ;
  assign n1019 = n1018 ^ n1010 ;
  assign n1045 = n1044 ^ n1019 ;
  assign n1001 = n791 ^ n471 ;
  assign n1000 = n520 ^ n275 ;
  assign n1002 = n1001 ^ n1000 ;
  assign n999 = n191 & n260 ;
  assign n1003 = n1002 ^ n999 ;
  assign n998 = n470 ^ n193 ;
  assign n1004 = n1003 ^ n998 ;
  assign n995 = n419 ^ n378 ;
  assign n996 = n995 ^ n387 ;
  assign n994 = n615 ^ n446 ;
  assign n997 = n996 ^ n994 ;
  assign n1005 = n1004 ^ n997 ;
  assign n254 = n253 ^ n250 ;
  assign n249 = n248 ^ n247 ;
  assign n255 = n254 ^ n249 ;
  assign n257 = n256 ^ n255 ;
  assign n1006 = n1005 ^ n257 ;
  assign n992 = n498 ^ n232 ;
  assign n993 = n992 ^ n991 ;
  assign n1007 = n1006 ^ n993 ;
  assign n1046 = n1045 ^ n1007 ;
  assign n1111 = n845 ^ n788 ;
  assign n908 = ~n148 & n176 ;
  assign n1110 = n908 ^ n493 ;
  assign n1112 = n1111 ^ n1110 ;
  assign n1108 = n440 ^ n277 ;
  assign n1106 = n62 & n191 ;
  assign n1107 = n1106 ^ n618 ;
  assign n1109 = n1108 ^ n1107 ;
  assign n1113 = n1112 ^ n1109 ;
  assign n1103 = n589 ^ n142 ;
  assign n903 = n152 & n228 ;
  assign n1104 = n1103 ^ n903 ;
  assign n1105 = n1104 ^ n346 ;
  assign n1114 = n1113 ^ n1105 ;
  assign n1099 = n836 ^ n794 ;
  assign n1100 = n1099 ^ n737 ;
  assign n943 = n62 & ~n107 ;
  assign n944 = n943 ^ n240 ;
  assign n1098 = n944 ^ n490 ;
  assign n1101 = n1100 ^ n1098 ;
  assign n1095 = n476 ^ n215 ;
  assign n1096 = n1095 ^ n511 ;
  assign n1092 = n634 ^ n409 ;
  assign n1093 = n1092 ^ n209 ;
  assign n1094 = n1093 ^ n495 ;
  assign n1097 = n1096 ^ n1094 ;
  assign n1102 = n1101 ^ n1097 ;
  assign n1115 = n1114 ^ n1102 ;
  assign n876 = n212 & n228 ;
  assign n1087 = n876 ^ n641 ;
  assign n1088 = n1087 ^ n773 ;
  assign n867 = ~n107 & n260 ;
  assign n900 = n867 ^ n270 ;
  assign n1089 = n1088 ^ n900 ;
  assign n1086 = n657 ^ n382 ;
  assign n1090 = n1089 ^ n1086 ;
  assign n1084 = n62 & n212 ;
  assign n1085 = n1084 ^ n556 ;
  assign n1091 = n1090 ^ n1085 ;
  assign n1116 = n1115 ^ n1091 ;
  assign n1078 = n805 ^ n776 ;
  assign n1077 = n136 & n176 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1080 = n1079 ^ n645 ;
  assign n1076 = n842 ^ n675 ;
  assign n1081 = n1080 ^ n1076 ;
  assign n1075 = n818 ^ n236 ;
  assign n1082 = n1081 ^ n1075 ;
  assign n873 = n152 & n299 ;
  assign n1073 = n873 ^ n390 ;
  assign n1074 = n1179 ^ n1073 ;
  assign n1083 = n1082 ^ n1074 ;
  assign n1117 = n1116 ^ n1083 ;
  assign n1066 = n62 & ~n20602 ;
  assign n1067 = n1066 ^ n592 ;
  assign n1068 = n1067 ^ n505 ;
  assign n1064 = n191 & n228 ;
  assign n1065 = n1064 ^ n468 ;
  assign n1069 = n1068 ^ n1065 ;
  assign n1062 = n523 ^ n137 ;
  assign n1060 = n735 ^ n369 ;
  assign n1061 = n1060 ^ n847 ;
  assign n1063 = n1062 ^ n1061 ;
  assign n1070 = n1069 ^ n1063 ;
  assign n1058 = n464 ^ n458 ;
  assign n1056 = n761 ^ n411 ;
  assign n1057 = n1056 ^ n462 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1071 = n1070 ^ n1059 ;
  assign n1052 = n141 & n228 ;
  assign n950 = n62 & n106 ;
  assign n1050 = n950 ^ n563 ;
  assign n1051 = n1050 ^ n239 ;
  assign n1053 = n1052 ^ n1051 ;
  assign n1048 = n784 ^ n519 ;
  assign n1049 = n1048 ^ n434 ;
  assign n1054 = n1053 ^ n1049 ;
  assign n926 = n157 ^ n108 ;
  assign n1047 = n926 ^ n716 ;
  assign n1055 = n1054 ^ n1047 ;
  assign n1072 = n1071 ^ n1055 ;
  assign n1118 = n1117 ^ n1072 ;
  assign n1119 = ~n1046 & ~n1118 ;
  assign n918 = ~n156 & n228 ;
  assign n919 = n918 ^ n213 ;
  assign n920 = n919 ^ n764 ;
  assign n917 = n645 ^ n600 ;
  assign n921 = n920 ^ n917 ;
  assign n262 = n141 & n260 ;
  assign n916 = n915 ^ n262 ;
  assign n922 = n921 ^ n916 ;
  assign n910 = n66 & n123 ;
  assign n911 = n910 ^ n437 ;
  assign n909 = n908 ^ n847 ;
  assign n912 = n911 ^ n909 ;
  assign n905 = n136 & n228 ;
  assign n906 = n905 ^ n409 ;
  assign n904 = n903 ^ n183 ;
  assign n907 = n906 ^ n904 ;
  assign n913 = n912 ^ n907 ;
  assign n898 = n520 ^ n468 ;
  assign n899 = n898 ^ n682 ;
  assign n901 = n900 ^ n899 ;
  assign n895 = n66 & ~n111 ;
  assign n896 = n895 ^ n577 ;
  assign n897 = n896 ^ n493 ;
  assign n902 = n901 ^ n897 ;
  assign n914 = n913 ^ n902 ;
  assign n923 = n922 ^ n914 ;
  assign n890 = n354 ^ n243 ;
  assign n891 = n890 ^ n517 ;
  assign n888 = n743 ^ n211 ;
  assign n889 = n888 ^ n192 ;
  assign n892 = n891 ^ n889 ;
  assign n886 = n753 ^ n506 ;
  assign n887 = n886 ^ n318 ;
  assign n893 = n892 ^ n887 ;
  assign n884 = n776 ^ n585 ;
  assign n883 = n761 ^ n489 ;
  assign n885 = n884 ^ n883 ;
  assign n894 = n893 ^ n885 ;
  assign n924 = n923 ^ n894 ;
  assign n877 = n876 ^ n584 ;
  assign n875 = n566 ^ n331 ;
  assign n878 = n877 ^ n875 ;
  assign n874 = n873 ^ n801 ;
  assign n879 = n878 ^ n874 ;
  assign n871 = n179 ^ n171 ;
  assign n872 = n871 ^ n251 ;
  assign n880 = n879 ^ n872 ;
  assign n868 = n1239 ^ n867 ;
  assign n869 = n868 ^ n737 ;
  assign n866 = n659 ^ n369 ;
  assign n870 = n869 ^ n866 ;
  assign n881 = n880 ^ n870 ;
  assign n861 = n66 & ~n116 ;
  assign n862 = n861 ^ n527 ;
  assign n863 = n862 ^ n818 ;
  assign n864 = n863 ^ n398 ;
  assign n858 = n730 ^ n239 ;
  assign n857 = n845 ^ n380 ;
  assign n859 = n858 ^ n857 ;
  assign n860 = n859 ^ n416 ;
  assign n865 = n864 ^ n860 ;
  assign n882 = n881 ^ n865 ;
  assign n925 = n924 ^ n882 ;
  assign n982 = n664 ^ n501 ;
  assign n983 = n982 ^ n478 ;
  assign n981 = n622 ^ n145 ;
  assign n984 = n983 ^ n981 ;
  assign n980 = n641 ^ n273 ;
  assign n985 = n984 ^ n980 ;
  assign n977 = n317 ^ n237 ;
  assign n978 = n977 ^ n703 ;
  assign n974 = ~n84 & ~n164 ;
  assign n976 = n975 ^ n974 ;
  assign n979 = n978 ^ n976 ;
  assign n986 = n985 ^ n979 ;
  assign n969 = n66 & n113 ;
  assign n970 = n969 ^ n788 ;
  assign n968 = n322 ^ n214 ;
  assign n971 = n970 ^ n968 ;
  assign n965 = n430 ^ n265 ;
  assign n966 = n965 ^ n444 ;
  assign n967 = n966 ^ n357 ;
  assign n972 = n971 ^ n967 ;
  assign n963 = n615 ^ n453 ;
  assign n962 = n1209 ^ n628 ;
  assign n964 = n963 ^ n962 ;
  assign n973 = n972 ^ n964 ;
  assign n987 = n986 ^ n973 ;
  assign n958 = n209 ^ n126 ;
  assign n957 = n956 ^ n820 ;
  assign n959 = n958 ^ n957 ;
  assign n955 = n547 ^ n182 ;
  assign n960 = n959 ^ n955 ;
  assign n951 = n950 ^ n118 ;
  assign n952 = n951 ^ n347 ;
  assign n953 = n952 ^ n390 ;
  assign n948 = n429 ^ n114 ;
  assign n949 = n948 ^ n495 ;
  assign n954 = n953 ^ n949 ;
  assign n961 = n960 ^ n954 ;
  assign n988 = n987 ^ n961 ;
  assign n941 = n838 ^ n247 ;
  assign n942 = n941 ^ n604 ;
  assign n945 = n944 ^ n942 ;
  assign n938 = n815 ^ n471 ;
  assign n937 = n784 ^ n653 ;
  assign n939 = n938 ^ n937 ;
  assign n935 = n750 ^ n199 ;
  assign n934 = n766 ^ n377 ;
  assign n936 = n935 ^ n934 ;
  assign n940 = n939 ^ n936 ;
  assign n946 = n945 ^ n940 ;
  assign n261 = ~n156 & n260 ;
  assign n930 = n637 ^ n261 ;
  assign n931 = n930 ^ n389 ;
  assign n928 = n675 ^ n555 ;
  assign n929 = n928 ^ n542 ;
  assign n932 = n931 ^ n929 ;
  assign n927 = n926 ^ n446 ;
  assign n933 = n932 ^ n927 ;
  assign n947 = n946 ^ n933 ;
  assign n989 = n988 ^ n947 ;
  assign n990 = ~n925 & ~n989 ;
  assign n1120 = n1119 ^ n990 ;
  assign n1189 = n66 & n91 ;
  assign n1190 = n1189 ^ n142 ;
  assign n1188 = n908 ^ n125 ;
  assign n1191 = n1190 ^ n1188 ;
  assign n1187 = n974 ^ n178 ;
  assign n1192 = n1191 ^ n1187 ;
  assign n1184 = n737 ^ n462 ;
  assign n1185 = n1184 ^ n347 ;
  assign n1183 = n675 ^ n197 ;
  assign n1186 = n1185 ^ n1183 ;
  assign n1193 = n1192 ^ n1186 ;
  assign n1180 = n1179 ^ n517 ;
  assign n1176 = n1077 ^ n94 ;
  assign n1177 = n1176 ^ n470 ;
  assign n1178 = n1177 ^ n716 ;
  assign n1181 = n1180 ^ n1178 ;
  assign n1175 = n975 ^ n873 ;
  assign n1182 = n1181 ^ n1175 ;
  assign n1194 = n1193 ^ n1182 ;
  assign n1170 = n663 ^ n434 ;
  assign n1171 = n1170 ^ n327 ;
  assign n1172 = n1171 ^ n991 ;
  assign n1173 = n1172 ^ n354 ;
  assign n1167 = n598 ^ n411 ;
  assign n1168 = n1167 ^ n419 ;
  assign n1169 = n1168 ^ n1106 ;
  assign n1174 = n1173 ^ n1169 ;
  assign n1195 = n1194 ^ n1174 ;
  assign n1162 = n437 ^ n341 ;
  assign n1163 = n1162 ^ n236 ;
  assign n1160 = n66 & n93 ;
  assign n1161 = n1160 ^ n262 ;
  assign n1164 = n1163 ^ n1161 ;
  assign n1158 = n682 ^ n153 ;
  assign n1159 = n1158 ^ n1066 ;
  assign n1165 = n1164 ^ n1159 ;
  assign n1156 = n1084 ^ n761 ;
  assign n1155 = n357 ^ n114 ;
  assign n1157 = n1156 ^ n1155 ;
  assign n1166 = n1165 ^ n1157 ;
  assign n1196 = n1195 ^ n1166 ;
  assign n1148 = n950 ^ n722 ;
  assign n1149 = n1148 ^ n464 ;
  assign n1150 = n1149 ^ n774 ;
  assign n1146 = n446 ^ n124 ;
  assign n1147 = n1146 ^ n602 ;
  assign n1151 = n1150 ^ n1147 ;
  assign n1143 = n577 ^ n550 ;
  assign n1142 = n250 ^ n179 ;
  assign n1144 = n1143 ^ n1142 ;
  assign n1140 = n668 ^ n526 ;
  assign n1139 = n380 ^ n239 ;
  assign n1141 = n1140 ^ n1139 ;
  assign n1145 = n1144 ^ n1141 ;
  assign n1152 = n1151 ^ n1145 ;
  assign n1136 = n504 ^ n417 ;
  assign n1135 = n803 ^ n444 ;
  assign n1137 = n1136 ^ n1135 ;
  assign n1133 = n609 ^ n256 ;
  assign n1134 = n1133 ^ n563 ;
  assign n1138 = n1137 ^ n1134 ;
  assign n1153 = n1152 ^ n1138 ;
  assign n1129 = n910 ^ n455 ;
  assign n1130 = n1129 ^ n471 ;
  assign n1127 = n770 ^ n567 ;
  assign n1128 = n1127 ^ n490 ;
  assign n1131 = n1130 ^ n1128 ;
  assign n1124 = n918 ^ n640 ;
  assign n1125 = n1124 ^ n1020 ;
  assign n1122 = n847 ^ n820 ;
  assign n1121 = n430 ^ n192 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1126 = n1125 ^ n1123 ;
  assign n1132 = n1131 ^ n1126 ;
  assign n1154 = n1153 ^ n1132 ;
  assign n1197 = n1196 ^ n1154 ;
  assign n1240 = n1239 ^ n213 ;
  assign n1241 = n1240 ^ n485 ;
  assign n1242 = n1241 ^ n867 ;
  assign n1236 = ~n148 & n228 ;
  assign n1237 = n1236 ^ n108 ;
  assign n1238 = n1237 ^ n735 ;
  assign n1243 = n1242 ^ n1238 ;
  assign n1233 = n831 ^ n320 ;
  assign n1234 = n1233 ^ n843 ;
  assign n1235 = n1234 ^ n1038 ;
  assign n1244 = n1243 ^ n1235 ;
  assign n1229 = n876 ^ n199 ;
  assign n1230 = n1229 ^ n1064 ;
  assign n1228 = n801 ^ n680 ;
  assign n1231 = n1230 ^ n1228 ;
  assign n1226 = n571 ^ n248 ;
  assign n1225 = n999 ^ n785 ;
  assign n1227 = n1226 ^ n1225 ;
  assign n1232 = n1231 ^ n1227 ;
  assign n1245 = n1244 ^ n1232 ;
  assign n1221 = n941 ^ n362 ;
  assign n1220 = n400 ^ n117 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1216 = n378 ^ n353 ;
  assign n1217 = n1216 ^ n511 ;
  assign n1218 = n1217 ^ n547 ;
  assign n1214 = n900 ^ n520 ;
  assign n1215 = n1214 ^ n585 ;
  assign n1219 = n1218 ^ n1215 ;
  assign n1223 = n1222 ^ n1219 ;
  assign n1210 = n1209 ^ n943 ;
  assign n1211 = n1210 ^ n523 ;
  assign n1212 = n1211 ^ n741 ;
  assign n1213 = n1212 ^ n887 ;
  assign n1224 = n1223 ^ n1213 ;
  assign n1246 = n1245 ^ n1224 ;
  assign n1204 = n719 ^ n480 ;
  assign n1205 = n1204 ^ n232 ;
  assign n1206 = n1205 ^ n414 ;
  assign n1201 = n710 ^ n641 ;
  assign n1202 = n1201 ^ n507 ;
  assign n1203 = n1202 ^ n861 ;
  assign n1207 = n1206 ^ n1203 ;
  assign n1198 = n495 ^ n211 ;
  assign n1199 = n1198 ^ n216 ;
  assign n1200 = n1199 ^ n597 ;
  assign n1208 = n1207 ^ n1200 ;
  assign n1247 = n1246 ^ n1208 ;
  assign n1248 = ~n1197 & ~n1247 ;
  assign n1249 = n1248 ^ n990 ;
  assign n1250 = ~n1120 & n1249 ;
  assign n1251 = n1045 ^ n794 ;
  assign n1291 = n974 ^ n464 ;
  assign n1292 = n1291 ^ n446 ;
  assign n1293 = n1292 ^ n240 ;
  assign n1289 = n778 ^ n275 ;
  assign n230 = n123 & n174 ;
  assign n1288 = n230 ^ n197 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1294 = n1293 ^ n1290 ;
  assign n1285 = n416 ^ n357 ;
  assign n1284 = n721 ^ n520 ;
  assign n1286 = n1285 ^ n1284 ;
  assign n1283 = n950 ^ n801 ;
  assign n1287 = n1286 ^ n1283 ;
  assign n1295 = n1294 ^ n1287 ;
  assign n1276 = n66 & ~n104 ;
  assign n1277 = n1276 ^ n171 ;
  assign n1278 = n1277 ^ n725 ;
  assign n1279 = n1278 ^ n495 ;
  assign n1280 = n1279 ^ n546 ;
  assign n1281 = n1280 ^ n969 ;
  assign n1274 = n868 ^ n471 ;
  assign n1273 = n563 ^ n138 ;
  assign n1275 = n1274 ^ n1273 ;
  assign n1282 = n1281 ^ n1275 ;
  assign n1296 = n1295 ^ n1282 ;
  assign n1268 = n526 ^ n513 ;
  assign n1269 = n1268 ^ n124 ;
  assign n1265 = n845 ^ n766 ;
  assign n1266 = n1265 ^ n184 ;
  assign n1263 = ~n51 & n333 ;
  assign n1264 = x23 & n1263 ;
  assign n1267 = n1266 ^ n1264 ;
  assign n1270 = n1269 ^ n1267 ;
  assign n1260 = n991 ^ n382 ;
  assign n1261 = n1260 ^ n839 ;
  assign n1258 = n1077 ^ n322 ;
  assign n1257 = n910 ^ n596 ;
  assign n1259 = n1258 ^ n1257 ;
  assign n1262 = n1261 ^ n1259 ;
  assign n1271 = n1270 ^ n1262 ;
  assign n1254 = n511 ^ n247 ;
  assign n1255 = n1254 ^ n772 ;
  assign n1252 = n1052 ^ n876 ;
  assign n1253 = n1252 ^ n750 ;
  assign n1256 = n1255 ^ n1253 ;
  assign n1272 = n1271 ^ n1256 ;
  assign n1297 = n1296 ^ n1272 ;
  assign n1337 = n1075 ^ n331 ;
  assign n1338 = n1337 ^ n905 ;
  assign n1335 = n1209 ^ n118 ;
  assign n1336 = n1335 ^ n440 ;
  assign n1339 = n1338 ^ n1336 ;
  assign n1332 = n788 ^ n584 ;
  assign n1333 = n1332 ^ n896 ;
  assign n1330 = n478 ^ n378 ;
  assign n1329 = n628 ^ n572 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1334 = n1333 ^ n1331 ;
  assign n1340 = n1339 ^ n1334 ;
  assign n1327 = n765 ^ n527 ;
  assign n1328 = n1327 ^ n843 ;
  assign n1341 = n1340 ^ n1328 ;
  assign n1324 = n915 ^ n485 ;
  assign n1323 = n798 ^ n327 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1321 = n1064 ^ n430 ;
  assign n1322 = n1321 ^ n417 ;
  assign n1326 = n1325 ^ n1322 ;
  assign n1342 = n1341 ^ n1326 ;
  assign n1317 = n755 ^ n668 ;
  assign n1314 = n730 ^ n682 ;
  assign n1315 = n1314 ^ n182 ;
  assign n1316 = n1315 ^ n602 ;
  assign n1318 = n1317 ^ n1316 ;
  assign n1312 = n903 ^ n634 ;
  assign n1313 = n1312 ^ n1066 ;
  assign n1319 = n1318 ^ n1313 ;
  assign n1307 = n131 & ~n20602 ;
  assign n1308 = n1307 ^ n1160 ;
  assign n1306 = n436 ^ n261 ;
  assign n1309 = n1308 ^ n1306 ;
  assign n1304 = n710 ^ n318 ;
  assign n1303 = n918 ^ n609 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1310 = n1309 ^ n1305 ;
  assign n1300 = n784 ^ n296 ;
  assign n1299 = n999 ^ n908 ;
  assign n1301 = n1300 ^ n1299 ;
  assign n1298 = n1236 ^ n547 ;
  assign n1302 = n1301 ^ n1298 ;
  assign n1311 = n1310 ^ n1302 ;
  assign n1320 = n1319 ^ n1311 ;
  assign n1343 = n1342 ^ n1320 ;
  assign n1344 = ~n1297 & ~n1343 ;
  assign n1345 = ~n1251 & n1344 ;
  assign n1694 = n1133 ^ n1085 ;
  assign n1693 = n1142 ^ n188 ;
  assign n1695 = n1694 ^ n1693 ;
  assign n1690 = n1689 ^ n498 ;
  assign n1691 = n1690 ^ n1058 ;
  assign n1687 = n778 ^ n157 ;
  assign n1688 = n1687 ^ n723 ;
  assign n1692 = n1691 ^ n1688 ;
  assign n1696 = n1695 ^ n1692 ;
  assign n1683 = n550 ^ n125 ;
  assign n1684 = n1683 ^ n262 ;
  assign n1685 = n1684 ^ n645 ;
  assign n1680 = n1160 ^ n766 ;
  assign n1681 = n1680 ^ n563 ;
  assign n1682 = n1681 ^ n452 ;
  assign n1686 = n1685 ^ n1682 ;
  assign n1697 = n1696 ^ n1686 ;
  assign n1676 = n1187 ^ n604 ;
  assign n1674 = n1307 ^ n357 ;
  assign n1675 = n1674 ^ n1277 ;
  assign n1677 = n1676 ^ n1675 ;
  assign n1673 = n1037 ^ n240 ;
  assign n1678 = n1677 ^ n1673 ;
  assign n1679 = n1678 ^ n1223 ;
  assign n1698 = n1697 ^ n1679 ;
  assign n1743 = n522 ^ n346 ;
  assign n1744 = n1743 ^ n197 ;
  assign n1745 = n1744 ^ n618 ;
  assign n314 = n57 & ~n87 ;
  assign n1742 = n737 ^ n314 ;
  assign n1746 = n1745 ^ n1742 ;
  assign n1653 = n513 ^ n184 ;
  assign n1740 = n1653 ^ n108 ;
  assign n1741 = n1740 ^ n507 ;
  assign n1747 = n1746 ^ n1741 ;
  assign n1735 = n706 ^ n380 ;
  assign n1736 = n1735 ^ n831 ;
  assign n1737 = n1736 ^ n628 ;
  assign n1738 = n1737 ^ n429 ;
  assign n1733 = n641 ^ n317 ;
  assign n1734 = n1733 ^ n772 ;
  assign n1739 = n1738 ^ n1734 ;
  assign n1748 = n1747 ^ n1739 ;
  assign n1729 = n764 ^ n137 ;
  assign n1728 = n491 ^ n265 ;
  assign n1730 = n1729 ^ n1728 ;
  assign n1726 = n820 ^ n600 ;
  assign n1727 = n1726 ^ n567 ;
  assign n1731 = n1730 ^ n1727 ;
  assign n1376 = n417 ^ n320 ;
  assign n1725 = n1376 ^ n640 ;
  assign n1732 = n1731 ^ n1725 ;
  assign n1749 = n1748 ^ n1732 ;
  assign n1719 = n637 ^ n434 ;
  assign n1720 = n1719 ^ n468 ;
  assign n1718 = n845 ^ n825 ;
  assign n1721 = n1720 ^ n1718 ;
  assign n1716 = n710 ^ n437 ;
  assign n1717 = n1716 ^ n382 ;
  assign n1722 = n1721 ^ n1717 ;
  assign n1723 = n1722 ^ n801 ;
  assign n1711 = n543 ^ n251 ;
  assign n1710 = n523 ^ n239 ;
  assign n1712 = n1711 ^ n1710 ;
  assign n1709 = n214 ^ n213 ;
  assign n1713 = n1712 ^ n1709 ;
  assign n1499 = n1014 ^ n419 ;
  assign n1708 = n1499 ^ n928 ;
  assign n1714 = n1713 ^ n1708 ;
  assign n1704 = n969 ^ n153 ;
  assign n1705 = n1704 ^ n981 ;
  assign n1702 = n680 ^ n209 ;
  assign n1703 = n1702 ^ n668 ;
  assign n1706 = n1705 ^ n1703 ;
  assign n1699 = n455 ^ n182 ;
  assign n1700 = n1699 ^ n741 ;
  assign n1701 = n1700 ^ n659 ;
  assign n1707 = n1706 ^ n1701 ;
  assign n1715 = n1714 ^ n1707 ;
  assign n1724 = n1723 ^ n1715 ;
  assign n1750 = n1749 ^ n1724 ;
  assign n1751 = ~n1698 & ~n1750 ;
  assign n1793 = n908 ^ n378 ;
  assign n1794 = n1793 ^ n613 ;
  assign n1790 = n750 ^ n677 ;
  assign n1791 = n1790 ^ n564 ;
  assign n1362 = n813 ^ n618 ;
  assign n1792 = n1791 ^ n1362 ;
  assign n1795 = n1794 ^ n1792 ;
  assign n1786 = n818 ^ n805 ;
  assign n1787 = n1786 ^ n585 ;
  assign n1785 = n861 ^ n197 ;
  assign n1788 = n1787 ^ n1785 ;
  assign n1783 = n791 ^ n416 ;
  assign n1784 = n1783 ^ n550 ;
  assign n1789 = n1788 ^ n1784 ;
  assign n1796 = n1795 ^ n1789 ;
  assign n1778 = n680 ^ n485 ;
  assign n1779 = n1778 ^ n1298 ;
  assign n1776 = n764 ^ n434 ;
  assign n1377 = n603 ^ n470 ;
  assign n1777 = n1776 ^ n1377 ;
  assign n1780 = n1779 ^ n1777 ;
  assign n1774 = n876 ^ n395 ;
  assign n1772 = n763 ^ n211 ;
  assign n1773 = n1772 ^ n1277 ;
  assign n1775 = n1774 ^ n1773 ;
  assign n1781 = n1780 ^ n1775 ;
  assign n1770 = n1313 ^ n948 ;
  assign n1768 = n517 ^ n385 ;
  assign n1769 = n1768 ^ n975 ;
  assign n1771 = n1770 ^ n1769 ;
  assign n1782 = n1781 ^ n1771 ;
  assign n1797 = n1796 ^ n1782 ;
  assign n1762 = n436 ^ n125 ;
  assign n1763 = n1762 ^ n675 ;
  assign n1764 = n1763 ^ n722 ;
  assign n1760 = n1189 ^ n230 ;
  assign n1761 = n1760 ^ n743 ;
  assign n1765 = n1764 ^ n1761 ;
  assign n1757 = n533 ^ n179 ;
  assign n1756 = n820 ^ n655 ;
  assign n1758 = n1757 ^ n1756 ;
  assign n1754 = n1014 ^ n918 ;
  assign n1755 = n1754 ^ n344 ;
  assign n1759 = n1758 ^ n1755 ;
  assign n1766 = n1765 ^ n1759 ;
  assign n1752 = n801 ^ n182 ;
  assign n1753 = n1752 ^ n277 ;
  assign n1767 = n1766 ^ n1753 ;
  assign n1798 = n1797 ^ n1767 ;
  assign n1811 = n493 ^ n480 ;
  assign n1812 = n1811 ^ n171 ;
  assign n1813 = n1812 ^ n741 ;
  assign n1814 = n1813 ^ n453 ;
  assign n1810 = n1184 ^ n831 ;
  assign n1815 = n1814 ^ n1810 ;
  assign n1389 = n560 ^ n256 ;
  assign n1808 = n1389 ^ n592 ;
  assign n1807 = n1052 ^ n251 ;
  assign n1809 = n1808 ^ n1807 ;
  assign n1816 = n1815 ^ n1809 ;
  assign n1817 = n1816 ^ n651 ;
  assign n1404 = n943 ^ n596 ;
  assign n1803 = n1404 ^ n353 ;
  assign n1804 = n1803 ^ n1268 ;
  assign n1661 = n663 ^ n213 ;
  assign n1662 = n1661 ^ n772 ;
  assign n1660 = n668 ^ n215 ;
  assign n1663 = n1662 ^ n1660 ;
  assign n1805 = n1804 ^ n1663 ;
  assign n1498 = n382 ^ n327 ;
  assign n1800 = n1674 ^ n1498 ;
  assign n1422 = n974 ^ n209 ;
  assign n1799 = n1422 ^ n994 ;
  assign n1801 = n1800 ^ n1799 ;
  assign n1590 = n1265 ^ n546 ;
  assign n1591 = n1590 ^ n754 ;
  assign n1802 = n1801 ^ n1591 ;
  assign n1806 = n1805 ^ n1802 ;
  assign n1818 = n1817 ^ n1806 ;
  assign n1819 = ~n1798 & ~n1818 ;
  assign n1820 = n1751 & n1819 ;
  assign n1378 = n1377 ^ n1376 ;
  assign n1374 = n1066 ^ n566 ;
  assign n1375 = n1374 ^ n270 ;
  assign n1379 = n1378 ^ n1375 ;
  assign n1372 = n1123 ^ n275 ;
  assign n1371 = n609 ^ n498 ;
  assign n1373 = n1372 ^ n1371 ;
  assign n1380 = n1379 ^ n1373 ;
  assign n1367 = n542 ^ n296 ;
  assign n1368 = n1367 ^ n272 ;
  assign n1369 = n1368 ^ n628 ;
  assign n1366 = n948 ^ n577 ;
  assign n1370 = n1369 ^ n1366 ;
  assign n1381 = n1380 ^ n1370 ;
  assign n1363 = n1362 ^ n1176 ;
  assign n1364 = n1363 ^ n1047 ;
  assign n1360 = n66 & ~n20602 ;
  assign n1361 = n1360 ^ n396 ;
  assign n1365 = n1364 ^ n1361 ;
  assign n1382 = n1381 ^ n1365 ;
  assign n1354 = n562 ^ n471 ;
  assign n1355 = n1354 ^ n831 ;
  assign n1356 = n1355 ^ n480 ;
  assign n1353 = n657 ^ n555 ;
  assign n1357 = n1356 ^ n1353 ;
  assign n1350 = n546 ^ n179 ;
  assign n1351 = n1350 ^ n641 ;
  assign n1352 = n1351 ^ n1180 ;
  assign n1358 = n1357 ^ n1352 ;
  assign n1347 = n615 ^ n490 ;
  assign n1348 = n1347 ^ n567 ;
  assign n1346 = n1036 ^ n649 ;
  assign n1349 = n1348 ^ n1346 ;
  assign n1359 = n1358 ^ n1349 ;
  assign n1383 = n1382 ^ n1359 ;
  assign n1441 = n575 ^ n236 ;
  assign n1442 = n1441 ^ n741 ;
  assign n1443 = n1442 ^ n527 ;
  assign n1440 = n825 ^ n452 ;
  assign n1444 = n1443 ^ n1440 ;
  assign n1437 = n640 ^ n318 ;
  assign n1438 = n1437 ^ n784 ;
  assign n1439 = n1438 ^ n547 ;
  assign n1445 = n1444 ^ n1439 ;
  assign n1434 = n747 ^ n712 ;
  assign n1432 = n1020 ^ n484 ;
  assign n1433 = n1432 ^ n665 ;
  assign n1435 = n1434 ^ n1433 ;
  assign n1436 = n1435 ^ n1185 ;
  assign n1446 = n1445 ^ n1436 ;
  assign n1428 = n460 ^ n117 ;
  assign n1427 = n1189 ^ n681 ;
  assign n1429 = n1428 ^ n1427 ;
  assign n1424 = n773 ^ n416 ;
  assign n1425 = n1424 ^ n573 ;
  assign n1426 = n1425 ^ n802 ;
  assign n1430 = n1429 ^ n1426 ;
  assign n1423 = n1422 ^ n776 ;
  assign n1431 = n1430 ^ n1423 ;
  assign n1447 = n1446 ^ n1431 ;
  assign n1418 = n504 ^ n252 ;
  assign n1419 = n1418 ^ n523 ;
  assign n1417 = n842 ^ n182 ;
  assign n1420 = n1419 ^ n1417 ;
  assign n1414 = n634 ^ n398 ;
  assign n1415 = n1414 ^ n340 ;
  assign n1416 = n1415 ^ n655 ;
  assign n1421 = n1420 ^ n1416 ;
  assign n1448 = n1447 ^ n1421 ;
  assign n1408 = n684 ^ n414 ;
  assign n1407 = n511 ^ n455 ;
  assign n1409 = n1408 ^ n1407 ;
  assign n1405 = n389 ^ n234 ;
  assign n1406 = n1405 ^ n1404 ;
  assign n1410 = n1409 ^ n1406 ;
  assign n1401 = n845 ^ n199 ;
  assign n1402 = n1401 ^ n446 ;
  assign n1400 = n898 ^ n677 ;
  assign n1403 = n1402 ^ n1400 ;
  assign n1411 = n1410 ^ n1403 ;
  assign n1397 = n479 ^ n331 ;
  assign n1398 = n1397 ^ n466 ;
  assign n1395 = n1084 ^ n805 ;
  assign n1396 = n1395 ^ n427 ;
  assign n1399 = n1398 ^ n1396 ;
  assign n1412 = n1411 ^ n1399 ;
  assign n1390 = n1389 ^ n1140 ;
  assign n1391 = n1390 ^ n419 ;
  assign n1392 = n1391 ^ n409 ;
  assign n1388 = n838 ^ n600 ;
  assign n1393 = n1392 ^ n1388 ;
  assign n1386 = n970 ^ n654 ;
  assign n1384 = n710 ^ n378 ;
  assign n1385 = n1384 ^ n951 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1394 = n1393 ^ n1387 ;
  assign n1413 = n1412 ^ n1394 ;
  assign n1449 = n1448 ^ n1413 ;
  assign n1450 = ~n1383 & ~n1449 ;
  assign n1472 = n213 ^ n171 ;
  assign n1471 = n556 ^ n398 ;
  assign n1473 = n1472 ^ n1471 ;
  assign n1469 = n659 ^ n211 ;
  assign n1470 = n1469 ^ n1015 ;
  assign n1474 = n1473 ^ n1470 ;
  assign n1467 = n1299 ^ n1176 ;
  assign n1465 = n772 ^ n543 ;
  assign n1466 = n1465 ^ n1329 ;
  assign n1468 = n1467 ^ n1466 ;
  assign n1475 = n1474 ^ n1468 ;
  assign n1461 = n1300 ^ n241 ;
  assign n1462 = n1461 ^ n566 ;
  assign n1459 = n1689 ^ n517 ;
  assign n1460 = n1459 ^ n513 ;
  assign n1463 = n1462 ^ n1460 ;
  assign n1464 = n1463 ^ n1402 ;
  assign n1476 = n1475 ^ n1464 ;
  assign n1456 = n956 ^ n479 ;
  assign n1454 = n867 ^ n354 ;
  assign n1455 = n1454 ^ n1020 ;
  assign n1457 = n1456 ^ n1455 ;
  assign n1451 = n577 ^ n138 ;
  assign n1452 = n1451 ^ n721 ;
  assign n1453 = n1452 ^ n533 ;
  assign n1458 = n1457 ^ n1453 ;
  assign n1477 = n1476 ^ n1458 ;
  assign n1533 = n1066 ^ n250 ;
  assign n1534 = n1533 ^ n318 ;
  assign n1532 = n1236 ^ n188 ;
  assign n1535 = n1534 ^ n1532 ;
  assign n1536 = n1535 ^ n184 ;
  assign n1531 = n1306 ^ n1128 ;
  assign n1537 = n1536 ^ n1531 ;
  assign n1528 = n1179 ^ n189 ;
  assign n1526 = n680 ^ n522 ;
  assign n1525 = ~n96 & n1263 ;
  assign n1527 = n1526 ^ n1525 ;
  assign n1529 = n1528 ^ n1527 ;
  assign n1523 = n484 ^ n434 ;
  assign n1522 = n831 ^ n444 ;
  assign n1524 = n1523 ^ n1522 ;
  assign n1530 = n1529 ^ n1524 ;
  assign n1538 = n1537 ^ n1530 ;
  assign n1518 = n637 ^ n570 ;
  assign n1519 = n1518 ^ n422 ;
  assign n1517 = n1209 ^ n153 ;
  assign n1520 = n1519 ^ n1517 ;
  assign n1514 = n1360 ^ n776 ;
  assign n1515 = n1514 ^ n238 ;
  assign n1512 = n955 ^ n641 ;
  assign n1513 = n1512 ^ n458 ;
  assign n1516 = n1515 ^ n1513 ;
  assign n1521 = n1520 ^ n1516 ;
  assign n1539 = n1538 ^ n1521 ;
  assign n1506 = n649 ^ n452 ;
  assign n1507 = n1506 ^ n480 ;
  assign n1508 = n1507 ^ n335 ;
  assign n1503 = n943 ^ n585 ;
  assign n1504 = n1503 ^ n506 ;
  assign n1505 = n1504 ^ n767 ;
  assign n1509 = n1508 ^ n1505 ;
  assign n1500 = n1499 ^ n1498 ;
  assign n1501 = n1500 ^ n341 ;
  assign n1495 = n664 ^ n440 ;
  assign n1496 = n1495 ^ n216 ;
  assign n1494 = n1184 ^ n825 ;
  assign n1497 = n1496 ^ n1494 ;
  assign n1502 = n1501 ^ n1497 ;
  assign n1510 = n1509 ^ n1502 ;
  assign n1489 = n584 ^ n453 ;
  assign n1490 = n1489 ^ n1008 ;
  assign n1491 = n1490 ^ n805 ;
  assign n1486 = n493 ^ n117 ;
  assign n1487 = n1486 ^ n411 ;
  assign n1485 = n597 ^ n389 ;
  assign n1488 = n1487 ^ n1485 ;
  assign n1492 = n1491 ^ n1488 ;
  assign n1481 = n750 ^ n232 ;
  assign n1482 = n1481 ^ n592 ;
  assign n1483 = n1482 ^ n969 ;
  assign n1478 = n730 ^ n609 ;
  assign n1479 = n1478 ^ n459 ;
  assign n1480 = n1479 ^ n800 ;
  assign n1484 = n1483 ^ n1480 ;
  assign n1493 = n1492 ^ n1484 ;
  assign n1511 = n1510 ^ n1493 ;
  assign n1540 = n1539 ^ n1511 ;
  assign n1541 = ~n1477 & ~n1540 ;
  assign n1549 = n570 ^ n511 ;
  assign n1550 = n1549 ^ n842 ;
  assign n1551 = n1550 ^ n417 ;
  assign n1547 = n831 ^ n275 ;
  assign n1548 = n1547 ^ n1360 ;
  assign n1552 = n1551 ^ n1548 ;
  assign n1544 = n730 ^ n188 ;
  assign n1545 = n1544 ^ n249 ;
  assign n1542 = n905 ^ n230 ;
  assign n1543 = n1542 ^ n1258 ;
  assign n1546 = n1545 ^ n1543 ;
  assign n1553 = n1552 ^ n1546 ;
  assign n1593 = n238 ^ n211 ;
  assign n1594 = n1593 ^ n262 ;
  assign n1592 = n1239 ^ n480 ;
  assign n1595 = n1594 ^ n1592 ;
  assign n1596 = n1595 ^ n1591 ;
  assign n1588 = n1021 ^ n999 ;
  assign n1587 = n440 ^ n250 ;
  assign n1589 = n1588 ^ n1587 ;
  assign n1597 = n1596 ^ n1589 ;
  assign n1581 = n741 ^ n722 ;
  assign n1582 = n1581 ^ n649 ;
  assign n1583 = n1582 ^ n153 ;
  assign n1580 = n1300 ^ n142 ;
  assign n1584 = n1583 ^ n1580 ;
  assign n1577 = n861 ^ n438 ;
  assign n1578 = n1577 ^ n956 ;
  assign n1576 = n1008 ^ n347 ;
  assign n1579 = n1578 ^ n1576 ;
  assign n1585 = n1584 ^ n1579 ;
  assign n1572 = n788 ^ n114 ;
  assign n1571 = n452 ^ n265 ;
  assign n1573 = n1572 ^ n1571 ;
  assign n1569 = n495 ^ n256 ;
  assign n1568 = n395 ^ n182 ;
  assign n1570 = n1569 ^ n1568 ;
  assign n1574 = n1573 ^ n1570 ;
  assign n1565 = n542 ^ n533 ;
  assign n1566 = n1565 ^ n472 ;
  assign n1564 = n991 ^ n711 ;
  assign n1567 = n1566 ^ n1564 ;
  assign n1575 = n1574 ^ n1567 ;
  assign n1586 = n1585 ^ n1575 ;
  assign n1598 = n1597 ^ n1586 ;
  assign n1558 = n716 ^ n610 ;
  assign n1559 = n1558 ^ n446 ;
  assign n1560 = n1559 ^ n813 ;
  assign n1556 = n847 ^ n677 ;
  assign n1557 = n1556 ^ n876 ;
  assign n1561 = n1560 ^ n1557 ;
  assign n1554 = n1277 ^ n577 ;
  assign n1555 = n1554 ^ n712 ;
  assign n1562 = n1561 ^ n1555 ;
  assign n1563 = n1562 ^ n873 ;
  assign n1599 = n1598 ^ n1563 ;
  assign n278 = n277 ^ n272 ;
  assign n1664 = n1663 ^ n278 ;
  assign n1658 = n803 ^ n239 ;
  assign n1659 = n1658 ^ n1486 ;
  assign n1665 = n1664 ^ n1659 ;
  assign n1654 = n1653 ^ n655 ;
  assign n1655 = n1654 ^ n761 ;
  assign n1656 = n1655 ^ n504 ;
  assign n1650 = n1273 ^ n498 ;
  assign n1651 = n1650 ^ n603 ;
  assign n1652 = n1651 ^ n1032 ;
  assign n1657 = n1656 ^ n1652 ;
  assign n1666 = n1665 ^ n1657 ;
  assign n1646 = n465 ^ n414 ;
  assign n1645 = n1499 ^ n382 ;
  assign n1647 = n1646 ^ n1645 ;
  assign n1643 = n900 ^ n137 ;
  assign n1644 = n1643 ^ n527 ;
  assign n1648 = n1647 ^ n1644 ;
  assign n1641 = n1167 ^ n1078 ;
  assign n1639 = n773 ^ n125 ;
  assign n1638 = n398 ^ n320 ;
  assign n1640 = n1639 ^ n1638 ;
  assign n1642 = n1641 ^ n1640 ;
  assign n1649 = n1648 ^ n1642 ;
  assign n1667 = n1666 ^ n1649 ;
  assign n1631 = n1066 ^ n199 ;
  assign n1632 = n1631 ^ n183 ;
  assign n1630 = n684 ^ n240 ;
  assign n1633 = n1632 ^ n1630 ;
  assign n1628 = n609 ^ n566 ;
  assign n1629 = n1628 ^ n770 ;
  assign n1634 = n1633 ^ n1629 ;
  assign n1625 = n171 ^ n124 ;
  assign n1626 = n1625 ^ n269 ;
  assign n1624 = n339 ^ n157 ;
  assign n1627 = n1626 ^ n1624 ;
  assign n1635 = n1634 ^ n1627 ;
  assign n1620 = n915 ^ n468 ;
  assign n1619 = n657 ^ n409 ;
  assign n1621 = n1620 ^ n1619 ;
  assign n1616 = n618 ^ n327 ;
  assign n1617 = n1616 ^ n523 ;
  assign n1618 = n1617 ^ n458 ;
  assign n1622 = n1621 ^ n1618 ;
  assign n1614 = n1084 ^ n252 ;
  assign n1615 = n1614 ^ n664 ;
  assign n1623 = n1622 ^ n1615 ;
  assign n1636 = n1635 ^ n1623 ;
  assign n1609 = n1064 ^ n637 ;
  assign n1610 = n1609 ^ n1160 ;
  assign n1607 = n867 ^ n522 ;
  assign n1608 = n1607 ^ n149 ;
  assign n1611 = n1610 ^ n1608 ;
  assign n1603 = n659 ^ n94 ;
  assign n1604 = n1603 ^ n640 ;
  assign n1605 = n1604 ^ n547 ;
  assign n1602 = n744 ^ n543 ;
  assign n1606 = n1605 ^ n1602 ;
  assign n1612 = n1611 ^ n1606 ;
  assign n1600 = n622 ^ n489 ;
  assign n1601 = n1600 ^ n434 ;
  assign n1613 = n1612 ^ n1601 ;
  assign n1637 = n1636 ^ n1613 ;
  assign n1668 = n1667 ^ n1637 ;
  assign n1669 = ~n1599 & ~n1668 ;
  assign n1670 = ~n1553 & n1669 ;
  assign n1671 = n1541 & n1670 ;
  assign n1672 = n1450 & n1671 ;
  assign n1821 = n1820 ^ n1672 ;
  assign n1928 = n1811 ^ n873 ;
  assign n1929 = n1928 ^ n1239 ;
  assign n1925 = n575 ^ n498 ;
  assign n1926 = n1925 ^ n905 ;
  assign n1927 = n1926 ^ n572 ;
  assign n1930 = n1929 ^ n1927 ;
  assign n1923 = n848 ^ n252 ;
  assign n1883 = n564 ^ n444 ;
  assign n1924 = n1923 ^ n1883 ;
  assign n1931 = n1930 ^ n1924 ;
  assign n1919 = n1209 ^ n464 ;
  assign n1920 = n1919 ^ n567 ;
  assign n1917 = n682 ^ n339 ;
  assign n1915 = n1036 ^ n753 ;
  assign n1916 = n1915 ^ n570 ;
  assign n1918 = n1917 ^ n1916 ;
  assign n1921 = n1920 ^ n1918 ;
  assign n1912 = n336 ^ n317 ;
  assign n1913 = n1912 ^ n1544 ;
  assign n1914 = n1913 ^ n1465 ;
  assign n1922 = n1921 ^ n1914 ;
  assign n1932 = n1931 ^ n1922 ;
  assign n1908 = n1179 ^ n277 ;
  assign n1906 = n589 ^ n566 ;
  assign n1907 = n1906 ^ n399 ;
  assign n1909 = n1908 ^ n1907 ;
  assign n1903 = n526 ^ n192 ;
  assign n1904 = n1903 ^ n216 ;
  assign n1905 = n1904 ^ n1190 ;
  assign n1910 = n1909 ^ n1905 ;
  assign n1900 = n1106 ^ n800 ;
  assign n1901 = n1900 ^ n803 ;
  assign n1898 = n390 ^ n265 ;
  assign n1899 = n1898 ^ n766 ;
  assign n1902 = n1901 ^ n1899 ;
  assign n1911 = n1910 ^ n1902 ;
  assign n1933 = n1932 ^ n1911 ;
  assign n1849 = n484 ^ n145 ;
  assign n1850 = n1849 ^ n118 ;
  assign n1851 = n1850 ^ n546 ;
  assign n1848 = n771 ^ n506 ;
  assign n1852 = n1851 ^ n1848 ;
  assign n1845 = n716 ^ n615 ;
  assign n1846 = n1845 ^ n1653 ;
  assign n1844 = n519 ^ n453 ;
  assign n1847 = n1846 ^ n1844 ;
  assign n1853 = n1852 ^ n1847 ;
  assign n1840 = n346 ^ n117 ;
  assign n1839 = n641 ^ n452 ;
  assign n1841 = n1840 ^ n1839 ;
  assign n1837 = n628 ^ n550 ;
  assign n1838 = n1837 ^ n687 ;
  assign n1842 = n1841 ^ n1838 ;
  assign n1834 = n489 ^ n124 ;
  assign n1833 = n584 ^ n250 ;
  assign n1835 = n1834 ^ n1833 ;
  assign n1831 = n943 ^ n178 ;
  assign n1832 = n1831 ^ n664 ;
  assign n1836 = n1835 ^ n1832 ;
  assign n1843 = n1842 ^ n1836 ;
  assign n1854 = n1853 ^ n1843 ;
  assign n1855 = n1854 ^ n1771 ;
  assign n1934 = n1933 ^ n1855 ;
  assign n1968 = n764 ^ n230 ;
  assign n1962 = n1008 ^ n999 ;
  assign n1963 = n1962 ^ n622 ;
  assign n1960 = n501 ^ n261 ;
  assign n1961 = n1960 ^ n533 ;
  assign n1964 = n1963 ^ n1961 ;
  assign n1957 = n818 ^ n610 ;
  assign n1958 = n1957 ^ n659 ;
  assign n1956 = n838 ^ n199 ;
  assign n1959 = n1958 ^ n1956 ;
  assign n1965 = n1964 ^ n1959 ;
  assign n1953 = n1360 ^ n125 ;
  assign n1954 = n1953 ^ n1689 ;
  assign n1952 = n1002 ^ n417 ;
  assign n1955 = n1954 ^ n1952 ;
  assign n1966 = n1965 ^ n1955 ;
  assign n1948 = n735 ^ n272 ;
  assign n1947 = n1616 ^ n655 ;
  assign n1949 = n1948 ^ n1947 ;
  assign n1945 = n340 ^ n189 ;
  assign n1944 = n1702 ^ n108 ;
  assign n1946 = n1945 ^ n1944 ;
  assign n1950 = n1949 ^ n1946 ;
  assign n1940 = n1184 ^ n719 ;
  assign n1941 = n1940 ^ n653 ;
  assign n1939 = n867 ^ n331 ;
  assign n1942 = n1941 ^ n1939 ;
  assign n1937 = n1405 ^ n1303 ;
  assign n1938 = n1937 ^ n396 ;
  assign n1943 = n1942 ^ n1938 ;
  assign n1951 = n1950 ^ n1943 ;
  assign n1967 = n1966 ^ n1951 ;
  assign n1969 = n1968 ^ n1967 ;
  assign n1936 = n788 ^ n314 ;
  assign n1970 = n1969 ^ n1936 ;
  assign n1935 = n640 ^ n440 ;
  assign n1971 = n1970 ^ n1935 ;
  assign n1972 = ~n1934 & ~n1971 ;
  assign n1827 = n956 ^ n340 ;
  assign n1828 = n1827 ^ n485 ;
  assign n1825 = n618 ^ n183 ;
  assign n1826 = n1825 ^ n478 ;
  assign n1829 = n1828 ^ n1826 ;
  assign n1823 = n706 ^ n602 ;
  assign n1822 = n867 ^ n857 ;
  assign n1824 = n1823 ^ n1822 ;
  assign n1830 = n1829 ^ n1824 ;
  assign n1856 = n1855 ^ n1830 ;
  assign n1889 = n459 ^ n399 ;
  assign n1890 = n1889 ^ n441 ;
  assign n1887 = n818 ^ n592 ;
  assign n1885 = ~x23 & n49 ;
  assign n1886 = n228 & n1885 ;
  assign n1888 = n1887 ^ n1886 ;
  assign n1891 = n1890 ^ n1888 ;
  assign n1892 = n1891 ^ n1595 ;
  assign n1884 = n1883 ^ n737 ;
  assign n1893 = n1892 ^ n1884 ;
  assign n1879 = n1179 ^ n108 ;
  assign n1880 = n1879 ^ n1757 ;
  assign n1878 = n1299 ^ n779 ;
  assign n1881 = n1880 ^ n1878 ;
  assign n1876 = n766 ^ n437 ;
  assign n1875 = n567 ^ n317 ;
  assign n1877 = n1876 ^ n1875 ;
  assign n1882 = n1881 ^ n1877 ;
  assign n1894 = n1893 ^ n1882 ;
  assign n1895 = n1894 ^ n1553 ;
  assign n1869 = n1704 ^ n1689 ;
  assign n1870 = n1869 ^ n680 ;
  assign n1868 = n609 ^ n357 ;
  assign n1871 = n1870 ^ n1868 ;
  assign n1866 = n1554 ^ n816 ;
  assign n1864 = n436 ^ n362 ;
  assign n1865 = n1864 ^ n826 ;
  assign n1867 = n1866 ^ n1865 ;
  assign n1872 = n1871 ^ n1867 ;
  assign n1861 = n1783 ^ n520 ;
  assign n1862 = n1861 ^ n1160 ;
  assign n1858 = n600 ^ n377 ;
  assign n1859 = n1858 ^ n354 ;
  assign n1857 = n974 ^ n462 ;
  assign n1860 = n1859 ^ n1857 ;
  assign n1863 = n1862 ^ n1860 ;
  assign n1873 = n1872 ^ n1863 ;
  assign n1874 = n1873 ^ n1649 ;
  assign n1896 = n1895 ^ n1874 ;
  assign n1897 = ~n1856 & ~n1896 ;
  assign n1973 = n1972 ^ n1897 ;
  assign n1974 = n1897 ^ n1541 ;
  assign n2043 = n788 ^ n94 ;
  assign n2042 = n1277 ^ n637 ;
  assign n2044 = n2043 ^ n2042 ;
  assign n2045 = n2044 ^ n570 ;
  assign n2046 = n2045 ^ n527 ;
  assign n2040 = n604 ^ n555 ;
  assign n2041 = n2040 ^ n504 ;
  assign n2047 = n2046 ^ n2041 ;
  assign n2035 = n1052 ^ n138 ;
  assign n2036 = n2035 ^ n1350 ;
  assign n2033 = n770 ^ n663 ;
  assign n2032 = n1014 ^ n618 ;
  assign n2034 = n2033 ^ n2032 ;
  assign n2037 = n2036 ^ n2034 ;
  assign n2038 = n2037 ^ n1627 ;
  assign n2028 = n564 ^ n230 ;
  assign n2029 = n2028 ^ n498 ;
  assign n2030 = n2029 ^ n680 ;
  assign n2025 = n1236 ^ n800 ;
  assign n2026 = n2025 ^ n389 ;
  assign n2024 = n867 ^ n145 ;
  assign n2027 = n2026 ^ n2024 ;
  assign n2031 = n2030 ^ n2027 ;
  assign n2039 = n2038 ^ n2031 ;
  assign n2048 = n2047 ^ n2039 ;
  assign n2021 = n1254 ^ n820 ;
  assign n2019 = n239 ^ n199 ;
  assign n2018 = n596 ^ n517 ;
  assign n2020 = n2019 ^ n2018 ;
  assign n2022 = n2021 ^ n2020 ;
  assign n2015 = n513 ^ n458 ;
  assign n2014 = n706 ^ n575 ;
  assign n2016 = n2015 ^ n2014 ;
  assign n2012 = n675 ^ n256 ;
  assign n2010 = n1209 ^ n188 ;
  assign n2011 = n2010 ^ n362 ;
  assign n2013 = n2012 ^ n2011 ;
  assign n2017 = n2016 ^ n2013 ;
  assign n2023 = n2022 ^ n2017 ;
  assign n2049 = n2048 ^ n2023 ;
  assign n2004 = n1581 ^ n764 ;
  assign n2005 = n2004 ^ n117 ;
  assign n2002 = n1095 ^ n682 ;
  assign n2003 = n2002 ^ n585 ;
  assign n2006 = n2005 ^ n2003 ;
  assign n2000 = n1469 ^ n937 ;
  assign n1998 = n999 ^ n801 ;
  assign n1997 = n815 ^ n465 ;
  assign n1999 = n1998 ^ n1997 ;
  assign n2001 = n2000 ^ n1999 ;
  assign n2007 = n2006 ^ n2001 ;
  assign n1994 = n900 ^ n380 ;
  assign n1995 = n1994 ^ n335 ;
  assign n1992 = n737 ^ n183 ;
  assign n1993 = n1992 ^ n615 ;
  assign n1996 = n1995 ^ n1993 ;
  assign n2008 = n2007 ^ n1996 ;
  assign n1987 = n773 ^ n272 ;
  assign n1988 = n1987 ^ n197 ;
  assign n1985 = n813 ^ n452 ;
  assign n1986 = n1985 ^ n873 ;
  assign n1989 = n1988 ^ n1986 ;
  assign n1983 = n1837 ^ n275 ;
  assign n1981 = n721 ^ n523 ;
  assign n1982 = n1981 ^ n440 ;
  assign n1984 = n1983 ^ n1982 ;
  assign n1990 = n1989 ^ n1984 ;
  assign n1978 = n1155 ^ n915 ;
  assign n1979 = n1978 ^ n836 ;
  assign n1975 = n842 ^ n556 ;
  assign n1976 = n1975 ^ n251 ;
  assign n1977 = n1976 ^ n1189 ;
  assign n1980 = n1979 ^ n1977 ;
  assign n1991 = n1990 ^ n1980 ;
  assign n2009 = n2008 ^ n1991 ;
  assign n2050 = n2049 ^ n2009 ;
  assign n2088 = n848 ^ n462 ;
  assign n2089 = n2088 ^ n655 ;
  assign n2086 = n1084 ^ n592 ;
  assign n2087 = n2086 ^ n385 ;
  assign n2090 = n2089 ^ n2087 ;
  assign n2084 = n1313 ^ n895 ;
  assign n2082 = n1307 ^ n195 ;
  assign n2083 = n2082 ^ n778 ;
  assign n2085 = n2084 ^ n2083 ;
  assign n2091 = n2090 ^ n2085 ;
  assign n2079 = n1075 ^ n346 ;
  assign n2078 = n1020 ^ n436 ;
  assign n2080 = n2079 ^ n2078 ;
  assign n2076 = n1906 ^ n1321 ;
  assign n2077 = n2076 ^ n1233 ;
  assign n2081 = n2080 ^ n2077 ;
  assign n2092 = n2091 ^ n2081 ;
  assign n2072 = n716 ^ n331 ;
  assign n2073 = n2072 ^ n641 ;
  assign n2070 = n898 ^ n209 ;
  assign n2068 = n1106 ^ n750 ;
  assign n2069 = n2068 ^ n153 ;
  assign n2071 = n2070 ^ n2069 ;
  assign n2074 = n2073 ^ n2071 ;
  assign n2065 = n955 ^ n354 ;
  assign n2066 = n2065 ^ n507 ;
  assign n2064 = n735 ^ n382 ;
  assign n2067 = n2066 ^ n2064 ;
  assign n2075 = n2074 ^ n2067 ;
  assign n2093 = n2092 ^ n2075 ;
  assign n2059 = n1124 ^ n243 ;
  assign n2060 = n2059 ^ n265 ;
  assign n2058 = n471 ^ n409 ;
  assign n2061 = n2060 ^ n2058 ;
  assign n2057 = n1601 ^ n395 ;
  assign n2062 = n2061 ^ n2057 ;
  assign n2054 = n725 ^ n277 ;
  assign n2053 = n327 ^ n252 ;
  assign n2055 = n2054 ^ n2053 ;
  assign n2051 = n533 ^ n318 ;
  assign n2052 = n2051 ^ n231 ;
  assign n2056 = n2055 ^ n2052 ;
  assign n2063 = n2062 ^ n2056 ;
  assign n2094 = n2093 ^ n2063 ;
  assign n2095 = ~n2050 & ~n2094 ;
  assign n2127 = n637 ^ n269 ;
  assign n2125 = n1160 ^ n189 ;
  assign n2126 = n2125 ^ n1189 ;
  assign n2128 = n2127 ^ n2126 ;
  assign n2129 = n2128 ^ n1813 ;
  assign n2120 = n215 ^ n94 ;
  assign n2121 = n2120 ^ n495 ;
  assign n2122 = n2121 ^ n108 ;
  assign n2117 = n719 ^ n275 ;
  assign n2118 = n2117 ^ n622 ;
  assign n2119 = n2118 ^ n585 ;
  assign n2123 = n2122 ^ n2119 ;
  assign n2115 = n2025 ^ n1565 ;
  assign n2114 = n1837 ^ n400 ;
  assign n2116 = n2115 ^ n2114 ;
  assign n2124 = n2123 ^ n2116 ;
  assign n2130 = n2129 ^ n2124 ;
  assign n2110 = n1576 ^ n600 ;
  assign n2111 = n2110 ^ n634 ;
  assign n2107 = n584 ^ n262 ;
  assign n2108 = n2107 ^ n252 ;
  assign n2105 = n649 ^ n277 ;
  assign n2106 = n2105 ^ n340 ;
  assign n2109 = n2108 ^ n2106 ;
  assign n2112 = n2111 ^ n2109 ;
  assign n2102 = n1953 ^ n969 ;
  assign n2103 = n2102 ^ n556 ;
  assign n2100 = n478 ^ n251 ;
  assign n2101 = n2100 ^ n436 ;
  assign n2104 = n2103 ^ n2101 ;
  assign n2113 = n2112 ^ n2104 ;
  assign n2131 = n2130 ^ n2113 ;
  assign n2132 = n2131 ^ n948 ;
  assign n2192 = n660 ^ n248 ;
  assign n2193 = n2192 ^ n663 ;
  assign n2190 = n1233 ^ n465 ;
  assign n2191 = n2190 ^ n825 ;
  assign n2194 = n2193 ^ n2191 ;
  assign n2187 = n362 ^ n296 ;
  assign n2188 = n2187 ^ n911 ;
  assign n2185 = n570 ^ n336 ;
  assign n2186 = n2185 ^ n2019 ;
  assign n2189 = n2188 ^ n2186 ;
  assign n2195 = n2194 ^ n2189 ;
  assign n2183 = n382 ^ n346 ;
  assign n2182 = n546 ^ n504 ;
  assign n2184 = n2183 ^ n2182 ;
  assign n2196 = n2195 ^ n2184 ;
  assign n2176 = n803 ^ n339 ;
  assign n2177 = n2176 ^ n943 ;
  assign n2178 = n2177 ^ n459 ;
  assign n2175 = n592 ^ n343 ;
  assign n2179 = n2178 ^ n2175 ;
  assign n2173 = n1441 ^ n378 ;
  assign n2172 = n1790 ^ n788 ;
  assign n2174 = n2173 ^ n2172 ;
  assign n2180 = n2179 ^ n2174 ;
  assign n2168 = n722 ^ n142 ;
  assign n2169 = n2168 ^ n417 ;
  assign n2166 = n250 ^ n231 ;
  assign n2167 = n2166 ^ n522 ;
  assign n2170 = n2169 ^ n2167 ;
  assign n2163 = n838 ^ n240 ;
  assign n2162 = n861 ^ n675 ;
  assign n2164 = n2163 ^ n2162 ;
  assign n2161 = n1643 ^ n905 ;
  assign n2165 = n2164 ^ n2161 ;
  assign n2171 = n2170 ^ n2165 ;
  assign n2181 = n2180 ^ n2171 ;
  assign n2197 = n2196 ^ n2181 ;
  assign n2155 = n1052 ^ n327 ;
  assign n2156 = n2155 ^ n1307 ;
  assign n2153 = n778 ^ n470 ;
  assign n2154 = n2153 ^ n1689 ;
  assign n2157 = n2156 ^ n2154 ;
  assign n2150 = n836 ^ n389 ;
  assign n2151 = n2150 ^ n1273 ;
  assign n2152 = n2151 ^ n857 ;
  assign n2158 = n2157 ^ n2152 ;
  assign n2145 = n322 ^ n197 ;
  assign n2144 = n770 ^ n411 ;
  assign n2146 = n2145 ^ n2144 ;
  assign n2147 = n2146 ^ n903 ;
  assign n2143 = n458 ^ n192 ;
  assign n2148 = n2147 ^ n2143 ;
  assign n2139 = n434 ^ n118 ;
  assign n2140 = n2139 ^ n265 ;
  assign n2141 = n2140 ^ n386 ;
  assign n2137 = n776 ^ n589 ;
  assign n2138 = n2137 ^ n668 ;
  assign n2142 = n2141 ^ n2138 ;
  assign n2149 = n2148 ^ n2142 ;
  assign n2159 = n2158 ^ n2149 ;
  assign n2134 = n957 ^ n543 ;
  assign n2135 = n2134 ^ n1654 ;
  assign n2133 = n1844 ^ n815 ;
  assign n2136 = n2135 ^ n2133 ;
  assign n2160 = n2159 ^ n2136 ;
  assign n2198 = n2197 ^ n2160 ;
  assign n2199 = ~n2132 & ~n2198 ;
  assign n2251 = n610 ^ n462 ;
  assign n2250 = n1360 ^ n1277 ;
  assign n2252 = n2251 ^ n2250 ;
  assign n2248 = n2051 ^ n585 ;
  assign n2249 = n2248 ^ n743 ;
  assign n2253 = n2252 ^ n2249 ;
  assign n2246 = n317 ^ n142 ;
  assign n2247 = n2246 ^ n505 ;
  assign n2254 = n2253 ^ n2247 ;
  assign n2243 = n805 ^ n480 ;
  assign n2242 = n950 ^ n915 ;
  assign n2244 = n2243 ^ n2242 ;
  assign n2241 = n1189 ^ n380 ;
  assign n2245 = n2244 ^ n2241 ;
  assign n2255 = n2254 ^ n2245 ;
  assign n2236 = n452 ^ n336 ;
  assign n2237 = n2236 ^ n1064 ;
  assign n2238 = n2237 ^ n1306 ;
  assign n2233 = n861 ^ n395 ;
  assign n2234 = n2233 ^ n444 ;
  assign n2235 = n2234 ^ n900 ;
  assign n2239 = n2238 ^ n2235 ;
  assign n2240 = n2239 ^ n2157 ;
  assign n2256 = n2255 ^ n2240 ;
  assign n2230 = n1528 ^ n526 ;
  assign n2229 = n592 ^ n485 ;
  assign n2231 = n2230 ^ n2229 ;
  assign n2227 = n507 ^ n357 ;
  assign n2226 = n838 ^ n335 ;
  assign n2228 = n2227 ^ n2226 ;
  assign n2232 = n2231 ^ n2228 ;
  assign n2257 = n2256 ^ n2232 ;
  assign n2220 = n774 ^ n240 ;
  assign n2221 = n2220 ^ n320 ;
  assign n2219 = n2107 ^ n721 ;
  assign n2222 = n2221 ^ n2219 ;
  assign n2215 = n1845 ^ n419 ;
  assign n2216 = n2215 ^ n753 ;
  assign n2217 = n2216 ^ n478 ;
  assign n2214 = n1354 ^ n455 ;
  assign n2218 = n2217 ^ n2214 ;
  assign n2223 = n2222 ^ n2218 ;
  assign n2224 = n2223 ^ n2023 ;
  assign n2210 = n1898 ^ n604 ;
  assign n2209 = n1935 ^ n1095 ;
  assign n2211 = n2210 ^ n2209 ;
  assign n2205 = n659 ^ n234 ;
  assign n2206 = n2205 ^ n571 ;
  assign n2207 = n2206 ^ n1556 ;
  assign n2204 = n999 ^ n668 ;
  assign n2208 = n2207 ^ n2204 ;
  assign n2212 = n2211 ^ n2208 ;
  assign n2201 = n813 ^ n340 ;
  assign n2202 = n2201 ^ n399 ;
  assign n2200 = n493 ^ n252 ;
  assign n2203 = n2202 ^ n2200 ;
  assign n2213 = n2212 ^ n2203 ;
  assign n2225 = n2224 ^ n2213 ;
  assign n2258 = n2257 ^ n2225 ;
  assign n2283 = n1479 ^ n466 ;
  assign n2281 = n896 ^ n184 ;
  assign n2282 = n2281 ^ n1060 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2285 = n2284 ^ n1723 ;
  assign n2277 = n663 ^ n331 ;
  assign n2278 = n2277 ^ n114 ;
  assign n2279 = n2278 ^ n1037 ;
  assign n2276 = n1327 ^ n354 ;
  assign n2280 = n2279 ^ n2276 ;
  assign n2286 = n2285 ^ n2280 ;
  assign n2271 = n903 ^ n836 ;
  assign n2272 = n2271 ^ n2105 ;
  assign n2270 = n378 ^ n118 ;
  assign n2273 = n2272 ^ n2270 ;
  assign n2267 = n1077 ^ n867 ;
  assign n2268 = n2267 ^ n555 ;
  assign n2265 = n1683 ^ n171 ;
  assign n2266 = n2265 ^ n761 ;
  assign n2269 = n2268 ^ n2266 ;
  assign n2274 = n2273 ^ n2269 ;
  assign n2261 = n831 ^ n430 ;
  assign n2262 = n2261 ^ n737 ;
  assign n2263 = n2262 ^ n389 ;
  assign n2259 = n417 ^ n192 ;
  assign n2260 = n2259 ^ n974 ;
  assign n2264 = n2263 ^ n2260 ;
  assign n2275 = n2274 ^ n2264 ;
  assign n2287 = n2286 ^ n2275 ;
  assign n2288 = ~n2258 & ~n2287 ;
  assign n2325 = n1254 ^ n417 ;
  assign n2323 = n1188 ^ n240 ;
  assign n2324 = n2323 ^ n737 ;
  assign n2326 = n2325 ^ n2324 ;
  assign n2320 = n577 ^ n178 ;
  assign n2321 = n2320 ^ n1362 ;
  assign n2319 = n1160 ^ n248 ;
  assign n2322 = n2321 ^ n2319 ;
  assign n2327 = n2326 ^ n2322 ;
  assign n2316 = n390 ^ n357 ;
  assign n2315 = n2068 ^ n1065 ;
  assign n2317 = n2316 ^ n2315 ;
  assign n2318 = n2317 ^ n2059 ;
  assign n2328 = n2327 ^ n2318 ;
  assign n2310 = n1277 ^ n836 ;
  assign n2311 = n2310 ^ n251 ;
  assign n2312 = n2311 ^ n436 ;
  assign n2309 = n905 ^ n555 ;
  assign n2313 = n2312 ^ n2309 ;
  assign n2306 = n1209 ^ n803 ;
  assign n2305 = n831 ^ n721 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2303 = n507 ^ n230 ;
  assign n2304 = n2303 ^ n668 ;
  assign n2308 = n2307 ^ n2304 ;
  assign n2314 = n2313 ^ n2308 ;
  assign n2329 = n2328 ^ n2314 ;
  assign n2297 = n609 ^ n556 ;
  assign n2298 = n2297 ^ n2107 ;
  assign n2295 = n1036 ^ n895 ;
  assign n2296 = n2295 ^ n1273 ;
  assign n2299 = n2298 ^ n2296 ;
  assign n2294 = n1582 ^ n319 ;
  assign n2300 = n2299 ^ n2294 ;
  assign n2291 = n1139 ^ n331 ;
  assign n2292 = n2291 ^ n1040 ;
  assign n2289 = n1175 ^ n214 ;
  assign n2290 = n2289 ^ n623 ;
  assign n2293 = n2292 ^ n2290 ;
  assign n2301 = n2300 ^ n2293 ;
  assign n2302 = n2301 ^ n1575 ;
  assign n2330 = n2329 ^ n2302 ;
  assign n2363 = n1052 ^ n465 ;
  assign n2364 = n2363 ^ n818 ;
  assign n2365 = n2364 ^ n910 ;
  assign n2362 = n703 ^ n527 ;
  assign n2366 = n2365 ^ n2362 ;
  assign n2359 = n1360 ^ n493 ;
  assign n2358 = n459 ^ n362 ;
  assign n2360 = n2359 ^ n2358 ;
  assign n2356 = n820 ^ n725 ;
  assign n2357 = n2356 ^ n1170 ;
  assign n2361 = n2360 ^ n2357 ;
  assign n2367 = n2366 ^ n2361 ;
  assign n2352 = n680 ^ n657 ;
  assign n2353 = n2352 ^ n339 ;
  assign n2354 = n2353 ^ n969 ;
  assign n2349 = n399 ^ n189 ;
  assign n2350 = n2349 ^ n504 ;
  assign n2348 = n1329 ^ n188 ;
  assign n2351 = n2350 ^ n2348 ;
  assign n2355 = n2354 ^ n2351 ;
  assign n2368 = n2367 ^ n2355 ;
  assign n2344 = n429 ^ n278 ;
  assign n2345 = n2344 ^ n1313 ;
  assign n2343 = n826 ^ n762 ;
  assign n2346 = n2345 ^ n2343 ;
  assign n2341 = n382 ^ n213 ;
  assign n2340 = n2270 ^ n377 ;
  assign n2342 = n2341 ^ n2340 ;
  assign n2347 = n2346 ^ n2342 ;
  assign n2369 = n2368 ^ n2347 ;
  assign n2337 = n1289 ^ n354 ;
  assign n2336 = n543 ^ n320 ;
  assign n2338 = n2337 ^ n2336 ;
  assign n2334 = n2082 ^ n562 ;
  assign n2331 = n523 ^ n444 ;
  assign n2332 = n2331 ^ n145 ;
  assign n2333 = n2332 ^ n974 ;
  assign n2335 = n2334 ^ n2333 ;
  assign n2339 = n2338 ^ n2335 ;
  assign n2370 = n2369 ^ n2339 ;
  assign n2371 = ~n2330 & ~n2370 ;
  assign n2415 = n876 ^ n458 ;
  assign n2416 = n2415 ^ n265 ;
  assign n2417 = n2416 ^ n2082 ;
  assign n2414 = n636 ^ n429 ;
  assign n2418 = n2417 ^ n2414 ;
  assign n2413 = n1209 ^ n815 ;
  assign n2419 = n2418 ^ n2413 ;
  assign n2410 = n2040 ^ n903 ;
  assign n2409 = n845 ^ n716 ;
  assign n2411 = n2410 ^ n2409 ;
  assign n2408 = n680 ^ n347 ;
  assign n2412 = n2411 ^ n2408 ;
  assign n2420 = n2419 ^ n2412 ;
  assign n2403 = n722 ^ n437 ;
  assign n2404 = n2403 ^ n1549 ;
  assign n2405 = n2404 ^ n2297 ;
  assign n2401 = n906 ^ n779 ;
  assign n2400 = n1783 ^ n1236 ;
  assign n2402 = n2401 ^ n2400 ;
  assign n2406 = n2405 ^ n2402 ;
  assign n2397 = n2246 ^ n567 ;
  assign n2398 = n2397 ^ n411 ;
  assign n2396 = n1066 ^ n522 ;
  assign n2399 = n2398 ^ n2396 ;
  assign n2407 = n2406 ^ n2399 ;
  assign n2421 = n2420 ^ n2407 ;
  assign n2391 = n2177 ^ n197 ;
  assign n2390 = n1762 ^ n641 ;
  assign n2392 = n2391 ^ n2390 ;
  assign n2388 = n243 ^ n188 ;
  assign n2389 = n2388 ^ n214 ;
  assign n2393 = n2392 ^ n2389 ;
  assign n2384 = n1106 ^ n1014 ;
  assign n2385 = n2384 ^ n1300 ;
  assign n2383 = n547 ^ n145 ;
  assign n2386 = n2385 ^ n2383 ;
  assign n2387 = n2386 ^ n497 ;
  assign n2394 = n2393 ^ n2387 ;
  assign n2379 = n788 ^ n453 ;
  assign n2378 = n1160 ^ n838 ;
  assign n2380 = n2379 ^ n2378 ;
  assign n2376 = n563 ^ n252 ;
  assign n2377 = n2376 ^ n658 ;
  assign n2381 = n2380 ^ n2377 ;
  assign n2373 = n772 ^ n506 ;
  assign n2374 = n2373 ^ n501 ;
  assign n2372 = n800 ^ n320 ;
  assign n2375 = n2374 ^ n2372 ;
  assign n2382 = n2381 ^ n2375 ;
  assign n2395 = n2394 ^ n2382 ;
  assign n2422 = n2421 ^ n2395 ;
  assign n2457 = n336 ^ n318 ;
  assign n2458 = n2457 ^ n470 ;
  assign n2459 = n2458 ^ n895 ;
  assign n2460 = n2459 ^ n991 ;
  assign n2461 = n2460 ^ n725 ;
  assign n2454 = n766 ^ n117 ;
  assign n2455 = n2454 ^ n610 ;
  assign n2453 = n710 ^ n248 ;
  assign n2456 = n2455 ^ n2453 ;
  assign n2462 = n2461 ^ n2456 ;
  assign n2449 = n1189 ^ n149 ;
  assign n2450 = n2449 ^ n362 ;
  assign n2448 = n655 ^ n353 ;
  assign n2451 = n2450 ^ n2448 ;
  assign n2445 = n649 ^ n183 ;
  assign n2446 = n2445 ^ n1000 ;
  assign n2444 = n598 ^ n322 ;
  assign n2447 = n2446 ^ n2444 ;
  assign n2452 = n2451 ^ n2447 ;
  assign n2463 = n2462 ^ n2452 ;
  assign n2464 = n2463 ^ n1083 ;
  assign n2439 = n1660 ^ n615 ;
  assign n2440 = n2439 ^ n459 ;
  assign n2438 = n663 ^ n480 ;
  assign n2441 = n2440 ^ n2438 ;
  assign n2437 = n753 ^ n382 ;
  assign n2442 = n2441 ^ n2437 ;
  assign n2434 = n1768 ^ n1414 ;
  assign n2432 = n910 ^ n192 ;
  assign n2433 = n2432 ^ n1689 ;
  assign n2435 = n2434 ^ n2433 ;
  assign n2436 = n2435 ^ n2263 ;
  assign n2443 = n2442 ^ n2436 ;
  assign n2465 = n2464 ^ n2443 ;
  assign n2428 = n542 ^ n414 ;
  assign n2426 = n585 ^ n237 ;
  assign n2427 = n2426 ^ n659 ;
  assign n2429 = n2428 ^ n2427 ;
  assign n2425 = n566 ^ n256 ;
  assign n2430 = n2429 ^ n2425 ;
  assign n2423 = n1925 ^ n1026 ;
  assign n2424 = n2423 ^ n2233 ;
  assign n2431 = n2430 ^ n2424 ;
  assign n2466 = n2465 ^ n2431 ;
  assign n2467 = ~n2422 & ~n2466 ;
  assign n2493 = n637 ^ n232 ;
  assign n2494 = n2493 ^ n399 ;
  assign n2495 = n2494 ^ n800 ;
  assign n2491 = n670 ^ n108 ;
  assign n2492 = n2491 ^ n876 ;
  assign n2496 = n2495 ^ n2492 ;
  assign n2486 = n842 ^ n471 ;
  assign n2487 = n2486 ^ n275 ;
  assign n2488 = n2487 ^ n1106 ;
  assign n2484 = n719 ^ n462 ;
  assign n2485 = n2484 ^ n784 ;
  assign n2489 = n2488 ^ n2485 ;
  assign n2481 = n566 ^ n248 ;
  assign n2482 = n2481 ^ n1142 ;
  assign n2479 = n455 ^ n389 ;
  assign n2480 = n2479 ^ n2457 ;
  assign n2483 = n2482 ^ n2480 ;
  assign n2490 = n2489 ^ n2483 ;
  assign n2497 = n2496 ^ n2490 ;
  assign n2475 = n1687 ^ n514 ;
  assign n2476 = n2475 ^ n427 ;
  assign n2473 = n884 ^ n252 ;
  assign n2474 = n2473 ^ n339 ;
  assign n2477 = n2476 ^ n2474 ;
  assign n2470 = n741 ^ n215 ;
  assign n2469 = n1175 ^ n770 ;
  assign n2471 = n2470 ^ n2469 ;
  assign n2468 = n1092 ^ n815 ;
  assign n2472 = n2471 ^ n2468 ;
  assign n2478 = n2477 ^ n2472 ;
  assign n2498 = n2497 ^ n2478 ;
  assign n2499 = n2498 ^ n1710 ;
  assign n2543 = n655 ^ n262 ;
  assign n2544 = n2543 ^ n1066 ;
  assign n2545 = n2544 ^ n357 ;
  assign n2546 = n2545 ^ n556 ;
  assign n2542 = n943 ^ n847 ;
  assign n2547 = n2546 ^ n2542 ;
  assign n2548 = n2547 ^ n591 ;
  assign n2540 = n1811 ^ n142 ;
  assign n2539 = n1858 ^ n506 ;
  assign n2541 = n2540 ^ n2539 ;
  assign n2549 = n2548 ^ n2541 ;
  assign n2532 = n895 ^ n825 ;
  assign n2533 = n2532 ^ n470 ;
  assign n2534 = n2533 ^ n1307 ;
  assign n2531 = n765 ^ n436 ;
  assign n2535 = n2534 ^ n2531 ;
  assign n2529 = n1495 ^ n571 ;
  assign n2528 = n1542 ^ n546 ;
  assign n2530 = n2529 ^ n2528 ;
  assign n2536 = n2535 ^ n2530 ;
  assign n2525 = n791 ^ n622 ;
  assign n2526 = n2525 ^ n716 ;
  assign n2523 = n956 ^ n417 ;
  assign n2524 = n2523 ^ n788 ;
  assign n2527 = n2526 ^ n2524 ;
  assign n2537 = n2536 ^ n2527 ;
  assign n2519 = n317 ^ n171 ;
  assign n2520 = n2519 ^ n1422 ;
  assign n2521 = n2520 ^ n899 ;
  assign n2522 = n2521 ^ n954 ;
  assign n2538 = n2537 ^ n2522 ;
  assign n2550 = n2549 ^ n2538 ;
  assign n2514 = n1395 ^ n668 ;
  assign n2513 = n991 ^ n750 ;
  assign n2515 = n2514 ^ n2513 ;
  assign n2510 = n603 ^ n476 ;
  assign n2509 = n766 ^ n94 ;
  assign n2511 = n2510 ^ n2509 ;
  assign n2507 = n562 ^ n251 ;
  assign n2506 = n861 ^ n801 ;
  assign n2508 = n2507 ^ n2506 ;
  assign n2512 = n2511 ^ n2508 ;
  assign n2516 = n2515 ^ n2512 ;
  assign n2503 = n968 ^ n838 ;
  assign n2504 = n2503 ^ n1397 ;
  assign n2500 = n398 ^ n340 ;
  assign n2501 = n2500 ^ n327 ;
  assign n2502 = n2501 ^ n1021 ;
  assign n2505 = n2504 ^ n2502 ;
  assign n2517 = n2516 ^ n2505 ;
  assign n2518 = n2517 ^ n1530 ;
  assign n2551 = n2550 ^ n2518 ;
  assign n2552 = ~n2499 & ~n2551 ;
  assign n2553 = n2009 ^ n1539 ;
  assign n2582 = n905 ^ n414 ;
  assign n2581 = n743 ^ n592 ;
  assign n2583 = n2582 ^ n2581 ;
  assign n2584 = n2583 ^ n430 ;
  assign n2580 = n526 ^ n248 ;
  assign n2585 = n2584 ^ n2580 ;
  assign n2576 = n1008 ^ n429 ;
  assign n2577 = n2576 ^ n1239 ;
  assign n2575 = n719 ^ n209 ;
  assign n2578 = n2577 ^ n2575 ;
  assign n2573 = n2072 ^ n542 ;
  assign n2574 = n2573 ^ n803 ;
  assign n2579 = n2578 ^ n2574 ;
  assign n2586 = n2585 ^ n2579 ;
  assign n2569 = n677 ^ n645 ;
  assign n2567 = n766 ^ n234 ;
  assign n2568 = n2567 ^ n2295 ;
  assign n2570 = n2569 ^ n2568 ;
  assign n2566 = n657 ^ n137 ;
  assign n2571 = n2570 ^ n2566 ;
  assign n2572 = n2571 ^ n1863 ;
  assign n2587 = n2586 ^ n2572 ;
  assign n2562 = n991 ^ n684 ;
  assign n2561 = n610 ^ n464 ;
  assign n2563 = n2562 ^ n2561 ;
  assign n2558 = n1188 ^ n108 ;
  assign n2559 = n2558 ^ n589 ;
  assign n2557 = n903 ^ n725 ;
  assign n2560 = n2559 ^ n2557 ;
  assign n2564 = n2563 ^ n2560 ;
  assign n2554 = n572 ^ n262 ;
  assign n2555 = n2554 ^ n1709 ;
  assign n2556 = n2555 ^ n2233 ;
  assign n2565 = n2564 ^ n2556 ;
  assign n2588 = n2587 ^ n2565 ;
  assign n2589 = ~n2553 & ~n2588 ;
  assign n2622 = n684 ^ n239 ;
  assign n2623 = n2622 ^ n546 ;
  assign n2624 = n2623 ^ n563 ;
  assign n2621 = n710 ^ n213 ;
  assign n2625 = n2624 ^ n2621 ;
  assign n2619 = n420 ^ n272 ;
  assign n2620 = n2619 ^ n716 ;
  assign n2626 = n2625 ^ n2620 ;
  assign n2616 = n1189 ^ n511 ;
  assign n2617 = n2616 ^ n1879 ;
  assign n2618 = n2617 ^ n1811 ;
  assign n2627 = n2626 ^ n2618 ;
  assign n2611 = n1960 ^ n440 ;
  assign n2610 = n743 ^ n336 ;
  assign n2612 = n2611 ^ n2610 ;
  assign n2608 = n778 ^ n236 ;
  assign n2607 = n761 ^ n753 ;
  assign n2609 = n2608 ^ n2607 ;
  assign n2613 = n2612 ^ n2609 ;
  assign n2604 = n1236 ^ n1176 ;
  assign n2603 = n1785 ^ n398 ;
  assign n2605 = n2604 ^ n2603 ;
  assign n2600 = n682 ^ n572 ;
  assign n2601 = n2600 ^ n429 ;
  assign n2599 = n915 ^ n741 ;
  assign n2602 = n2601 ^ n2599 ;
  assign n2606 = n2605 ^ n2602 ;
  assign n2614 = n2613 ^ n2606 ;
  assign n2596 = n495 ^ n479 ;
  assign n2593 = n600 ^ n124 ;
  assign n2594 = n2593 ^ n1360 ;
  assign n2595 = n2594 ^ n380 ;
  assign n2597 = n2596 ^ n2595 ;
  assign n2591 = n2315 ^ n1171 ;
  assign n2590 = n2479 ^ n1353 ;
  assign n2592 = n2591 ^ n2590 ;
  assign n2598 = n2597 ^ n2592 ;
  assign n2615 = n2614 ^ n2598 ;
  assign n2628 = n2627 ^ n2615 ;
  assign n2648 = n1512 ^ n322 ;
  assign n2649 = n2648 ^ n820 ;
  assign n2650 = n2649 ^ n527 ;
  assign n2651 = n2650 ^ n1209 ;
  assign n2646 = n2259 ^ n416 ;
  assign n2647 = n2646 ^ n1084 ;
  assign n2652 = n2651 ^ n2647 ;
  assign n2644 = n1793 ^ n622 ;
  assign n2645 = n2644 ^ n2219 ;
  assign n2653 = n2652 ^ n2645 ;
  assign n2639 = n730 ^ n377 ;
  assign n2640 = n2639 ^ n596 ;
  assign n2641 = n2640 ^ n1506 ;
  assign n2638 = n1459 ^ n602 ;
  assign n2642 = n2641 ^ n2638 ;
  assign n2634 = n1887 ^ n1277 ;
  assign n2635 = n2634 ^ n369 ;
  assign n2636 = n2635 ^ n411 ;
  assign n2631 = n444 ^ n138 ;
  assign n2632 = n2631 ^ n390 ;
  assign n2630 = n560 ^ n117 ;
  assign n2633 = n2632 ^ n2630 ;
  assign n2637 = n2636 ^ n2633 ;
  assign n2643 = n2642 ^ n2637 ;
  assign n2654 = n2653 ^ n2643 ;
  assign n2629 = n1105 ^ n430 ;
  assign n2655 = n2654 ^ n2629 ;
  assign n2656 = n2655 ^ n1045 ;
  assign n2657 = ~n2628 & ~n2656 ;
  assign n2658 = n2347 ^ n900 ;
  assign n2659 = n2658 ^ n2301 ;
  assign n2705 = n1898 ^ n1879 ;
  assign n2704 = n1790 ^ n1229 ;
  assign n2706 = n2705 ^ n2704 ;
  assign n2701 = n1008 ^ n189 ;
  assign n2702 = n2701 ^ n520 ;
  assign n2700 = n730 ^ n114 ;
  assign n2703 = n2702 ^ n2700 ;
  assign n2707 = n2706 ^ n2703 ;
  assign n2697 = n1465 ^ n322 ;
  assign n2698 = n2697 ^ n1283 ;
  assign n2699 = n2698 ^ n1063 ;
  assign n2708 = n2707 ^ n2699 ;
  assign n2693 = n1084 ^ n663 ;
  assign n2694 = n2693 ^ n2486 ;
  assign n2691 = n555 ^ n438 ;
  assign n2692 = n2691 ^ n956 ;
  assign n2695 = n2694 ^ n2692 ;
  assign n2689 = n1064 ^ n640 ;
  assign n2690 = n2689 ^ n969 ;
  assign n2696 = n2695 ^ n2690 ;
  assign n2709 = n2708 ^ n2696 ;
  assign n2684 = n1441 ^ n791 ;
  assign n2685 = n2684 ^ n395 ;
  assign n2682 = n1900 ^ n572 ;
  assign n2683 = n2682 ^ n493 ;
  assign n2686 = n2685 ^ n2683 ;
  assign n2679 = n485 ^ n327 ;
  assign n2678 = n589 ^ n519 ;
  assign n2680 = n2679 ^ n2678 ;
  assign n2677 = n1689 ^ n598 ;
  assign n2681 = n2680 ^ n2677 ;
  assign n2687 = n2686 ^ n2681 ;
  assign n2676 = n1408 ^ n551 ;
  assign n2688 = n2687 ^ n2676 ;
  assign n2710 = n2709 ^ n2688 ;
  assign n2670 = n788 ^ n600 ;
  assign n2671 = n2670 ^ n653 ;
  assign n2672 = n2671 ^ n1020 ;
  assign n2673 = n2672 ^ n2451 ;
  assign n2667 = n2432 ^ n930 ;
  assign n2668 = n2667 ^ n2507 ;
  assign n2665 = n2267 ^ n1095 ;
  assign n2664 = n1198 ^ n619 ;
  assign n2666 = n2665 ^ n2664 ;
  assign n2669 = n2668 ^ n2666 ;
  assign n2674 = n2673 ^ n2669 ;
  assign n2661 = n2427 ^ n498 ;
  assign n2662 = n2661 ^ n602 ;
  assign n2660 = n886 ^ n517 ;
  assign n2663 = n2662 ^ n2660 ;
  assign n2675 = n2674 ^ n2663 ;
  assign n2711 = n2710 ^ n2675 ;
  assign n2712 = ~n2659 & ~n2711 ;
  assign n2742 = n2082 ^ n770 ;
  assign n2741 = n836 ^ n138 ;
  assign n2743 = n2742 ^ n2741 ;
  assign n2744 = n2743 ^ n2585 ;
  assign n2737 = n1844 ^ n501 ;
  assign n2738 = n2737 ^ n417 ;
  assign n2736 = n975 ^ n247 ;
  assign n2739 = n2738 ^ n2736 ;
  assign n2735 = n389 ^ n150 ;
  assign n2740 = n2739 ^ n2735 ;
  assign n2745 = n2744 ^ n2740 ;
  assign n2732 = n1179 ^ n179 ;
  assign n2733 = n2732 ^ n1284 ;
  assign n2734 = n2733 ^ n1996 ;
  assign n2746 = n2745 ^ n2734 ;
  assign n2727 = n1156 ^ n847 ;
  assign n2728 = n2727 ^ n547 ;
  assign n2724 = n951 ^ n355 ;
  assign n2725 = n2724 ^ n523 ;
  assign n2726 = n2725 ^ n1252 ;
  assign n2729 = n2728 ^ n2726 ;
  assign n2720 = n419 ^ n239 ;
  assign n2721 = n2720 ^ n2432 ;
  assign n2719 = n2072 ^ n1362 ;
  assign n2722 = n2721 ^ n2719 ;
  assign n2723 = n2722 ^ n1589 ;
  assign n2730 = n2729 ^ n2723 ;
  assign n2715 = n687 ^ n238 ;
  assign n2716 = n2715 ^ n1544 ;
  assign n2717 = n2716 ^ n1730 ;
  assign n2713 = n2568 ^ n1014 ;
  assign n2714 = n2713 ^ n1040 ;
  assign n2718 = n2717 ^ n2714 ;
  assign n2731 = n2730 ^ n2718 ;
  assign n2747 = n2746 ^ n2731 ;
  assign n2748 = ~n2132 & ~n2747 ;
  assign n2755 = n1052 ^ n546 ;
  assign n2756 = n2755 ^ n813 ;
  assign n2754 = n645 ^ n275 ;
  assign n2757 = n2756 ^ n2754 ;
  assign n2752 = n791 ^ n770 ;
  assign n2753 = n2752 ^ n414 ;
  assign n2758 = n2757 ^ n2753 ;
  assign n2749 = n1239 ^ n668 ;
  assign n2750 = n2749 ^ n1210 ;
  assign n2751 = n2750 ^ n1143 ;
  assign n2759 = n2758 ^ n2751 ;
  assign n2760 = n2759 ^ n1946 ;
  assign n2784 = n628 ^ n243 ;
  assign n2783 = n750 ^ n622 ;
  assign n2785 = n2784 ^ n2783 ;
  assign n2781 = n589 ^ n236 ;
  assign n2780 = n716 ^ n506 ;
  assign n2782 = n2781 ^ n2780 ;
  assign n2786 = n2785 ^ n2782 ;
  assign n2787 = n2786 ^ n1618 ;
  assign n2778 = n957 ^ n838 ;
  assign n2779 = n2778 ^ n872 ;
  assign n2788 = n2787 ^ n2779 ;
  assign n2773 = n655 ^ n94 ;
  assign n2774 = n2773 ^ n142 ;
  assign n2775 = n2774 ^ n1264 ;
  assign n2771 = n2634 ^ n452 ;
  assign n2770 = n909 ^ n114 ;
  assign n2772 = n2771 ^ n2770 ;
  assign n2776 = n2775 ^ n2772 ;
  assign n2766 = n455 ^ n157 ;
  assign n2767 = n2766 ^ n773 ;
  assign n2765 = n766 ^ n761 ;
  assign n2768 = n2767 ^ n2765 ;
  assign n2762 = n794 ^ n347 ;
  assign n2763 = n2762 ^ n1236 ;
  assign n2761 = n707 ^ n557 ;
  assign n2764 = n2763 ^ n2761 ;
  assign n2769 = n2768 ^ n2764 ;
  assign n2777 = n2776 ^ n2769 ;
  assign n2789 = n2788 ^ n2777 ;
  assign n2790 = ~n2760 & ~n2789 ;
  assign n2832 = n543 ^ n247 ;
  assign n2830 = n888 ^ n296 ;
  assign n2831 = n2830 ^ n301 ;
  assign n2833 = n2832 ^ n2831 ;
  assign n2828 = n504 ^ n362 ;
  assign n2829 = n2828 ^ n1077 ;
  assign n2834 = n2833 ^ n2829 ;
  assign n2835 = n2834 ^ n2067 ;
  assign n2824 = n1709 ^ n682 ;
  assign n2825 = n2824 ^ n805 ;
  assign n2823 = n2481 ^ n649 ;
  assign n2826 = n2825 ^ n2823 ;
  assign n2821 = n1718 ^ n1229 ;
  assign n2819 = n918 ^ n395 ;
  assign n291 = n110 ^ n86 ;
  assign n292 = n291 ^ n104 ;
  assign n283 = x26 ^ x24 ;
  assign n293 = n292 ^ n283 ;
  assign n294 = n260 & n293 ;
  assign n284 = n283 ^ n97 ;
  assign n286 = n285 ^ x23 ;
  assign n287 = n286 ^ n97 ;
  assign n288 = n284 & ~n287 ;
  assign n289 = n288 ^ n97 ;
  assign n290 = n264 & ~n289 ;
  assign n295 = n294 ^ n290 ;
  assign n2818 = n991 ^ n295 ;
  assign n2820 = n2819 ^ n2818 ;
  assign n2822 = n2821 ^ n2820 ;
  assign n2827 = n2826 ^ n2822 ;
  assign n2836 = n2835 ^ n2827 ;
  assign n2811 = n584 ^ n533 ;
  assign n2812 = n2811 ^ n335 ;
  assign n2813 = n2812 ^ n905 ;
  assign n2810 = n594 ^ n188 ;
  assign n2814 = n2813 ^ n2810 ;
  assign n2807 = n1106 ^ n567 ;
  assign n2808 = n2807 ^ n124 ;
  assign n2809 = n2808 ^ n501 ;
  assign n2815 = n2814 ^ n2809 ;
  assign n2805 = n2277 ^ n150 ;
  assign n2806 = n2805 ^ n884 ;
  assign n2816 = n2815 ^ n2806 ;
  assign n2801 = n764 ^ n677 ;
  assign n2802 = n2801 ^ n1160 ;
  assign n2803 = n2802 ^ n642 ;
  assign n2798 = n753 ^ n741 ;
  assign n2797 = n873 ^ n232 ;
  assign n2799 = n2798 ^ n2797 ;
  assign n2796 = n1020 ^ n664 ;
  assign n2800 = n2799 ^ n2796 ;
  assign n2804 = n2803 ^ n2800 ;
  assign n2817 = n2816 ^ n2804 ;
  assign n2837 = n2836 ^ n2817 ;
  assign n2792 = n306 ^ x23 ;
  assign n2793 = n2792 ^ n86 ;
  assign n2791 = n147 ^ n78 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2795 = n298 & ~n2794 ;
  assign n2838 = n2837 ^ n2795 ;
  assign n2839 = n2790 & ~n2838 ;
  assign n2872 = n2801 ^ n411 ;
  assign n2873 = n2872 ^ n975 ;
  assign n2870 = n910 ^ n791 ;
  assign n2871 = n2870 ^ n398 ;
  assign n2874 = n2873 ^ n2871 ;
  assign n2868 = n511 ^ n183 ;
  assign n2869 = n2868 ^ n714 ;
  assign n2875 = n2874 ^ n2869 ;
  assign n2865 = n1236 ^ n861 ;
  assign n2866 = n2865 ^ n1857 ;
  assign n2867 = n2866 ^ n2028 ;
  assign n2876 = n2875 ^ n2867 ;
  assign n2862 = n1646 ^ n441 ;
  assign n2859 = n476 ^ n192 ;
  assign n2860 = n2859 ^ n788 ;
  assign n2857 = n530 ^ n124 ;
  assign n2858 = n2857 ^ n478 ;
  assign n2861 = n2860 ^ n2858 ;
  assign n2863 = n2862 ^ n2861 ;
  assign n2855 = n2457 ^ n2058 ;
  assign n2854 = n634 ^ n335 ;
  assign n2856 = n2855 ^ n2854 ;
  assign n2864 = n2863 ^ n2856 ;
  assign n2877 = n2876 ^ n2864 ;
  assign n2849 = n1014 ^ n348 ;
  assign n2850 = n2849 ^ n490 ;
  assign n2851 = n2850 ^ n1314 ;
  assign n2847 = n589 ^ n377 ;
  assign n2848 = n2847 ^ n836 ;
  assign n2852 = n2851 ^ n2848 ;
  assign n2843 = n2082 ^ n1689 ;
  assign n2844 = n2843 ^ n470 ;
  assign n2845 = n2844 ^ n555 ;
  assign n2840 = n838 ^ n645 ;
  assign n2841 = n2840 ^ n453 ;
  assign n2842 = n2841 ^ n992 ;
  assign n2846 = n2845 ^ n2842 ;
  assign n2853 = n2852 ^ n2846 ;
  assign n2878 = n2877 ^ n2853 ;
  assign n2928 = n1180 ^ n818 ;
  assign n2929 = n2928 ^ n603 ;
  assign n2926 = n721 ^ n247 ;
  assign n2927 = n2926 ^ n380 ;
  assign n2930 = n2929 ^ n2927 ;
  assign n2924 = n969 ^ n182 ;
  assign n2925 = n2924 ^ n642 ;
  assign n2931 = n2930 ^ n2925 ;
  assign n2919 = n340 ^ n261 ;
  assign n2920 = n2919 ^ n357 ;
  assign n2921 = n2920 ^ n157 ;
  assign n2917 = n362 ^ n137 ;
  assign n2918 = n2917 ^ n275 ;
  assign n2922 = n2921 ^ n2918 ;
  assign n2916 = n1811 ^ n519 ;
  assign n2923 = n2922 ^ n2916 ;
  assign n2932 = n2931 ^ n2923 ;
  assign n2912 = n437 ^ n118 ;
  assign n2910 = n2784 ^ n1360 ;
  assign n2909 = n1052 ^ n214 ;
  assign n2911 = n2910 ^ n2909 ;
  assign n2913 = n2912 ^ n2911 ;
  assign n2907 = ~x29 & n113 ;
  assign n2908 = n54 & n2907 ;
  assign n2914 = n2913 ^ n2908 ;
  assign n2905 = n772 ^ n610 ;
  assign n2906 = n2905 ^ n1299 ;
  assign n2915 = n2914 ^ n2906 ;
  assign n2933 = n2932 ^ n2915 ;
  assign n2898 = n903 ^ n464 ;
  assign n2899 = n2898 ^ n211 ;
  assign n2900 = n2899 ^ n895 ;
  assign n2897 = n1307 ^ n149 ;
  assign n2901 = n2900 ^ n2897 ;
  assign n2894 = n991 ^ n663 ;
  assign n2895 = n2894 ^ n524 ;
  assign n2896 = n2895 ^ n1517 ;
  assign n2902 = n2901 ^ n2896 ;
  assign n2891 = n1084 ^ n884 ;
  assign n2892 = n2891 ^ n2216 ;
  assign n2889 = n1027 ^ n543 ;
  assign n2890 = n2889 ^ n1226 ;
  assign n2893 = n2892 ^ n2890 ;
  assign n2903 = n2902 ^ n2893 ;
  assign n2884 = n847 ^ n215 ;
  assign n2885 = n2884 ^ n2127 ;
  assign n2886 = n2885 ^ n708 ;
  assign n2883 = n1832 ^ n390 ;
  assign n2887 = n2886 ^ n2883 ;
  assign n2881 = n1160 ^ n399 ;
  assign n2879 = n735 ^ n548 ;
  assign n2880 = n2879 ^ n900 ;
  assign n2882 = n2881 ^ n2880 ;
  assign n2888 = n2887 ^ n2882 ;
  assign n2904 = n2903 ^ n2888 ;
  assign n2934 = n2933 ^ n2904 ;
  assign n2935 = ~n2878 & ~n2934 ;
  assign n2975 = n419 ^ n317 ;
  assign n2976 = n2975 ^ n919 ;
  assign n2973 = n867 ^ n773 ;
  assign n2972 = n430 ^ n395 ;
  assign n2974 = n2973 ^ n2972 ;
  assign n2977 = n2976 ^ n2974 ;
  assign n2971 = n992 ^ n842 ;
  assign n2978 = n2977 ^ n2971 ;
  assign n2969 = n1052 ^ n252 ;
  assign n2970 = n2969 ^ n1591 ;
  assign n2979 = n2978 ^ n2970 ;
  assign n2965 = n788 ^ n272 ;
  assign n2966 = n2965 ^ n566 ;
  assign n2964 = n1037 ^ n353 ;
  assign n2967 = n2966 ^ n2964 ;
  assign n2962 = n1471 ^ n261 ;
  assign n2963 = n2962 ^ n1021 ;
  assign n2968 = n2967 ^ n2963 ;
  assign n2980 = n2979 ^ n2968 ;
  assign n2956 = n677 ^ n417 ;
  assign n2957 = n2956 ^ n322 ;
  assign n2955 = n858 ^ n171 ;
  assign n2958 = n2957 ^ n2955 ;
  assign n2953 = n1992 ^ n1689 ;
  assign n2954 = n2953 ^ n722 ;
  assign n2959 = n2958 ^ n2954 ;
  assign n2951 = n1040 ^ n725 ;
  assign n2949 = n975 ^ n563 ;
  assign n2950 = n2949 ^ n1832 ;
  assign n2952 = n2951 ^ n2950 ;
  assign n2960 = n2959 ^ n2952 ;
  assign n2946 = n900 ^ n262 ;
  assign n2944 = n2847 ^ n145 ;
  assign n2945 = n2944 ^ n550 ;
  assign n2947 = n2946 ^ n2945 ;
  assign n2940 = n719 ^ n182 ;
  assign n2941 = n2940 ^ n908 ;
  assign n2938 = n667 ^ n320 ;
  assign n2939 = n2938 ^ n1064 ;
  assign n2942 = n2941 ^ n2939 ;
  assign n2936 = n2072 ^ n710 ;
  assign n2937 = n2936 ^ n1525 ;
  assign n2943 = n2942 ^ n2937 ;
  assign n2948 = n2947 ^ n2943 ;
  assign n2961 = n2960 ^ n2948 ;
  assign n2981 = n2980 ^ n2961 ;
  assign n3013 = n2082 ^ n506 ;
  assign n3014 = n3013 ^ n347 ;
  assign n3015 = n3014 ^ n411 ;
  assign n3012 = n2600 ^ n784 ;
  assign n3016 = n3015 ^ n3012 ;
  assign n3010 = n2773 ^ n746 ;
  assign n3008 = n490 ^ n340 ;
  assign n3009 = n3008 ^ n438 ;
  assign n3011 = n3010 ^ n3009 ;
  assign n3017 = n3016 ^ n3011 ;
  assign n3005 = n1312 ^ n761 ;
  assign n3006 = n3005 ^ n765 ;
  assign n3007 = n3006 ^ n630 ;
  assign n3018 = n3017 ^ n3007 ;
  assign n3019 = n3018 ^ n1295 ;
  assign n3001 = n645 ^ n522 ;
  assign n3002 = n3001 ^ n847 ;
  assign n2998 = n547 ^ n380 ;
  assign n2999 = n2998 ^ n237 ;
  assign n3000 = n2999 ^ n465 ;
  assign n3003 = n3002 ^ n3000 ;
  assign n3004 = n3003 ^ n562 ;
  assign n3020 = n3019 ^ n3004 ;
  assign n2993 = n501 ^ n354 ;
  assign n2994 = n2993 ^ n1277 ;
  assign n2995 = n2994 ^ n463 ;
  assign n2990 = n1077 ^ n124 ;
  assign n2991 = n2990 ^ n1260 ;
  assign n2988 = n1236 ^ n389 ;
  assign n2989 = n2988 ^ n1889 ;
  assign n2992 = n2991 ^ n2989 ;
  assign n2996 = n2995 ^ n2992 ;
  assign n2984 = n1323 ^ n277 ;
  assign n2985 = n2984 ^ n743 ;
  assign n2983 = n1084 ^ n444 ;
  assign n2986 = n2985 ^ n2983 ;
  assign n2982 = n1811 ^ n1711 ;
  assign n2987 = n2986 ^ n2982 ;
  assign n2997 = n2996 ^ n2987 ;
  assign n3021 = n3020 ^ n2997 ;
  assign n3022 = ~n2981 & ~n3021 ;
  assign n3048 = n1040 ^ n385 ;
  assign n3049 = n3048 ^ n895 ;
  assign n3050 = n3049 ^ n1699 ;
  assign n3046 = n2100 ^ n918 ;
  assign n3047 = n3046 ^ n355 ;
  assign n3051 = n3050 ^ n3047 ;
  assign n3044 = n2854 ^ n471 ;
  assign n3043 = n645 ^ n209 ;
  assign n3045 = n3044 ^ n3043 ;
  assign n3052 = n3051 ^ n3045 ;
  assign n3038 = n800 ^ n142 ;
  assign n3039 = n3038 ^ n2150 ;
  assign n3036 = n950 ^ n682 ;
  assign n3037 = n3036 ^ n2778 ;
  assign n3040 = n3039 ^ n3037 ;
  assign n3033 = n1459 ^ n145 ;
  assign n3034 = n3033 ^ n2576 ;
  assign n3031 = n675 ^ n462 ;
  assign n3032 = n3031 ^ n2798 ;
  assign n3035 = n3034 ^ n3032 ;
  assign n3041 = n3040 ^ n3035 ;
  assign n3027 = n1718 ^ n232 ;
  assign n3028 = n3027 ^ n296 ;
  assign n3026 = n699 ^ n261 ;
  assign n3029 = n3028 ^ n3026 ;
  assign n3024 = n910 ^ n710 ;
  assign n3023 = n1209 ^ n974 ;
  assign n3025 = n3024 ^ n3023 ;
  assign n3030 = n3029 ^ n3025 ;
  assign n3042 = n3041 ^ n3030 ;
  assign n3053 = n3052 ^ n3042 ;
  assign n3054 = n3053 ^ n1637 ;
  assign n3055 = ~n1895 & ~n3054 ;
  assign n3072 = n2146 ^ n453 ;
  assign n3071 = n805 ^ n495 ;
  assign n3073 = n3072 ^ n3071 ;
  assign n3069 = n435 ^ n377 ;
  assign n3067 = n772 ^ n719 ;
  assign n3068 = n3067 ^ n543 ;
  assign n3070 = n3069 ^ n3068 ;
  assign n3074 = n3073 ^ n3070 ;
  assign n3075 = n3074 ^ n2914 ;
  assign n3063 = n779 ^ n534 ;
  assign n3061 = n895 ^ n602 ;
  assign n3062 = n3061 ^ n654 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3060 = n773 ^ n391 ;
  assign n3065 = n3064 ^ n3060 ;
  assign n3058 = n1268 ^ n399 ;
  assign n3057 = n1917 ^ n1209 ;
  assign n3059 = n3058 ^ n3057 ;
  assign n3066 = n3065 ^ n3059 ;
  assign n3076 = n3075 ^ n3066 ;
  assign n3056 = n2543 ^ n1879 ;
  assign n3077 = n3076 ^ n3056 ;
  assign n3118 = n2344 ^ n1900 ;
  assign n3117 = n637 ^ n317 ;
  assign n3119 = n3118 ^ n3117 ;
  assign n3115 = n3008 ^ n1768 ;
  assign n3116 = n3115 ^ n2383 ;
  assign n3120 = n3119 ^ n3116 ;
  assign n3111 = n1036 ^ n125 ;
  assign n3112 = n3111 ^ n261 ;
  assign n3113 = n3112 ^ n512 ;
  assign n3110 = n2690 ^ n1225 ;
  assign n3114 = n3113 ^ n3110 ;
  assign n3121 = n3120 ^ n3114 ;
  assign n3122 = n3121 ^ n2171 ;
  assign n3105 = n1778 ^ n452 ;
  assign n3104 = n2741 ^ n555 ;
  assign n3106 = n3105 ^ n3104 ;
  assign n3102 = n476 ^ n248 ;
  assign n3101 = n1014 ^ n252 ;
  assign n3103 = n3102 ^ n3101 ;
  assign n3107 = n3106 ^ n3103 ;
  assign n3099 = n3013 ^ n915 ;
  assign n3097 = n791 ^ n362 ;
  assign n3098 = n3097 ^ n189 ;
  assign n3100 = n3099 ^ n3098 ;
  assign n3108 = n3107 ^ n3100 ;
  assign n3090 = n95 ^ n91 ;
  assign n3091 = n3090 ^ n78 ;
  assign n3092 = n62 & n3091 ;
  assign n3093 = n3092 ^ n710 ;
  assign n3094 = n3093 ^ n2899 ;
  assign n3085 = n618 ^ n419 ;
  assign n3086 = n3085 ^ n239 ;
  assign n3087 = n3086 ^ n382 ;
  assign n3084 = n816 ^ n318 ;
  assign n3088 = n3087 ^ n3084 ;
  assign n3083 = n1883 ^ n1832 ;
  assign n3089 = n3088 ^ n3083 ;
  assign n3095 = n3094 ^ n3089 ;
  assign n3081 = n3046 ^ n2770 ;
  assign n3079 = n876 ^ n440 ;
  assign n3078 = n730 ^ n409 ;
  assign n3080 = n3079 ^ n3078 ;
  assign n3082 = n3081 ^ n3080 ;
  assign n3096 = n3095 ^ n3082 ;
  assign n3109 = n3108 ^ n3096 ;
  assign n3123 = n3122 ^ n3109 ;
  assign n3124 = ~n3077 & ~n3123 ;
  assign n3153 = n346 ^ n138 ;
  assign n3154 = n3153 ^ n419 ;
  assign n3151 = n434 ^ n149 ;
  assign n3150 = n690 ^ n598 ;
  assign n3152 = n3151 ^ n3150 ;
  assign n3155 = n3154 ^ n3152 ;
  assign n3148 = n935 ^ n820 ;
  assign n3149 = n3148 ^ n2507 ;
  assign n3156 = n3155 ^ n3149 ;
  assign n3157 = n3156 ^ n1080 ;
  assign n4722 = n975 ^ n622 ;
  assign n3144 = n4722 ^ n1660 ;
  assign n3145 = n3144 ^ n518 ;
  assign n3140 = n498 ^ n209 ;
  assign n3141 = n3140 ^ n737 ;
  assign n3142 = n3141 ^ n1014 ;
  assign n3146 = n3145 ^ n3142 ;
  assign n3138 = n2363 ^ n555 ;
  assign n3135 = n735 ^ n409 ;
  assign n3136 = n3135 ^ n550 ;
  assign n3137 = n3136 ^ n801 ;
  assign n3139 = n3138 ^ n3137 ;
  assign n3147 = n3146 ^ n3139 ;
  assign n3158 = n3157 ^ n3147 ;
  assign n3131 = n2641 ^ n414 ;
  assign n625 = n63 & n212 ;
  assign n3130 = n857 ^ n625 ;
  assign n3132 = n3131 ^ n3130 ;
  assign n3129 = n762 ^ n495 ;
  assign n3133 = n3132 ^ n3129 ;
  assign n3126 = n2843 ^ n468 ;
  assign n3127 = n3126 ^ n653 ;
  assign n3125 = n670 ^ n296 ;
  assign n3128 = n3127 ^ n3125 ;
  assign n3134 = n3133 ^ n3128 ;
  assign n3159 = n3158 ^ n3134 ;
  assign n3188 = n663 ^ n247 ;
  assign n3189 = n3188 ^ n462 ;
  assign n3190 = n3189 ^ n230 ;
  assign n3185 = n873 ^ n803 ;
  assign n3186 = n3185 ^ n182 ;
  assign n3187 = n3186 ^ n179 ;
  assign n3191 = n3190 ^ n3187 ;
  assign n3182 = n1307 ^ n369 ;
  assign n3183 = n3182 ^ n458 ;
  assign n3181 = n1277 ^ n684 ;
  assign n3184 = n3183 ^ n3181 ;
  assign n3192 = n3191 ^ n3184 ;
  assign n3178 = n867 ^ n213 ;
  assign n3177 = n2261 ^ n575 ;
  assign n3179 = n3178 ^ n3177 ;
  assign n3175 = n1160 ^ n493 ;
  assign n3176 = n3175 ^ n769 ;
  assign n3180 = n3179 ^ n3176 ;
  assign n3193 = n3192 ^ n3180 ;
  assign n3170 = n2993 ^ n183 ;
  assign n3171 = n3170 ^ n534 ;
  assign n3169 = n1414 ^ n603 ;
  assign n3172 = n3171 ^ n3169 ;
  assign n3166 = n453 ^ n416 ;
  assign n3167 = n3166 ^ n438 ;
  assign n3165 = n1465 ^ n396 ;
  assign n3168 = n3167 ^ n3165 ;
  assign n3173 = n3172 ^ n3168 ;
  assign n3162 = n1327 ^ n1130 ;
  assign n3163 = n3162 ^ n585 ;
  assign n3160 = n716 ^ n157 ;
  assign n3161 = n3160 ^ n600 ;
  assign n3164 = n3163 ^ n3161 ;
  assign n3174 = n3173 ^ n3164 ;
  assign n3194 = n3193 ^ n3174 ;
  assign n3195 = n3194 ^ n3122 ;
  assign n3196 = ~n3159 & ~n3195 ;
  assign n3197 = ~n3124 & ~n3196 ;
  assign n3198 = n3055 & ~n3197 ;
  assign n3199 = ~n3022 & ~n3198 ;
  assign n3226 = n1239 ^ n272 ;
  assign n3227 = n3226 ^ n400 ;
  assign n3228 = n3227 ^ n964 ;
  assign n3224 = n1423 ^ n820 ;
  assign n3223 = n1066 ^ n380 ;
  assign n3225 = n3224 ^ n3223 ;
  assign n3229 = n3228 ^ n3225 ;
  assign n3221 = n2243 ^ n883 ;
  assign n3219 = n446 ^ n434 ;
  assign n3220 = n3219 ^ n896 ;
  assign n3222 = n3221 ^ n3220 ;
  assign n3230 = n3229 ^ n3222 ;
  assign n3213 = n825 ^ n188 ;
  assign n3214 = n3213 ^ n275 ;
  assign n3212 = n903 ^ n250 ;
  assign n3215 = n3214 ^ n3212 ;
  assign n3209 = n743 ^ n706 ;
  assign n3210 = n3209 ^ n567 ;
  assign n3207 = n234 ^ n179 ;
  assign n3208 = n3207 ^ n675 ;
  assign n3211 = n3210 ^ n3208 ;
  assign n3216 = n3215 ^ n3211 ;
  assign n3206 = n56 & ~n20602 ;
  assign n3217 = n3216 ^ n3206 ;
  assign n3202 = n803 ^ n411 ;
  assign n3203 = n3202 ^ n818 ;
  assign n3200 = n468 ^ n314 ;
  assign n3201 = n3200 ^ n318 ;
  assign n3204 = n3203 ^ n3201 ;
  assign n3205 = n3204 ^ n334 ;
  assign n3218 = n3217 ^ n3205 ;
  assign n3231 = n3230 ^ n3218 ;
  assign n3232 = n3231 ^ n2961 ;
  assign n3243 = n842 ^ n536 ;
  assign n3244 = n3243 ^ n735 ;
  assign n3245 = n3244 ^ n1256 ;
  assign n3239 = n214 ^ n143 ;
  assign n3240 = n3239 ^ n378 ;
  assign n3237 = n557 ^ n94 ;
  assign n3238 = n3237 ^ n684 ;
  assign n3241 = n3240 ^ n3238 ;
  assign n3234 = n815 ^ n184 ;
  assign n3235 = n3234 ^ n2576 ;
  assign n3236 = n3235 ^ n2153 ;
  assign n3242 = n3241 ^ n3236 ;
  assign n3246 = n3245 ^ n3242 ;
  assign n3233 = n2675 ^ n649 ;
  assign n3247 = n3246 ^ n3233 ;
  assign n3248 = ~n3232 & ~n3247 ;
  assign n3249 = ~n3199 & n3248 ;
  assign n3250 = ~n2935 & ~n3249 ;
  assign n3251 = n2839 & ~n3250 ;
  assign n3252 = ~n2748 & ~n3251 ;
  assign n3282 = n1528 ^ n520 ;
  assign n3283 = n3282 ^ n1252 ;
  assign n3284 = n3283 ^ n1377 ;
  assign n3279 = n610 ^ n178 ;
  assign n3280 = n3279 ^ n317 ;
  assign n3277 = n1273 ^ n240 ;
  assign n3278 = n3277 ^ n369 ;
  assign n3281 = n3280 ^ n3278 ;
  assign n3285 = n3284 ^ n3281 ;
  assign n3273 = n3219 ^ n243 ;
  assign n3274 = n3273 ^ n800 ;
  assign n3272 = n600 ^ n414 ;
  assign n3275 = n3274 ^ n3272 ;
  assign n3276 = n3275 ^ n2080 ;
  assign n3286 = n3285 ^ n3276 ;
  assign n3270 = n805 ^ n183 ;
  assign n3271 = n3270 ^ n2356 ;
  assign n3287 = n3286 ^ n3271 ;
  assign n3265 = n1397 ^ n362 ;
  assign n3266 = n3265 ^ n771 ;
  assign n3263 = n1603 ^ n150 ;
  assign n3262 = n1027 ^ n108 ;
  assign n3264 = n3263 ^ n3262 ;
  assign n3267 = n3266 ^ n3264 ;
  assign n3268 = n3267 ^ n3217 ;
  assign n3257 = n2058 ^ n542 ;
  assign n3255 = n2068 ^ n918 ;
  assign n3256 = n3255 ^ n493 ;
  assign n3258 = n3257 ^ n3256 ;
  assign n3259 = n3258 ^ n664 ;
  assign n3260 = n3259 ^ n710 ;
  assign n3253 = n1753 ^ n591 ;
  assign n3254 = n3253 ^ n3060 ;
  assign n3261 = n3260 ^ n3254 ;
  assign n3269 = n3268 ^ n3261 ;
  assign n3288 = n3287 ^ n3269 ;
  assign n3317 = n956 ^ n895 ;
  assign n3318 = n3317 ^ n2576 ;
  assign n3315 = n813 ^ n784 ;
  assign n3316 = n3315 ^ n199 ;
  assign n3319 = n3318 ^ n3316 ;
  assign n3314 = n1156 ^ n886 ;
  assign n3320 = n3319 ^ n3314 ;
  assign n3313 = n2737 ^ n2307 ;
  assign n3321 = n3320 ^ n3313 ;
  assign n3310 = n2840 ^ n1526 ;
  assign n3311 = n3310 ^ n2102 ;
  assign n3307 = n1307 ^ n653 ;
  assign n3306 = n585 ^ n339 ;
  assign n3308 = n3307 ^ n3306 ;
  assign n3304 = n641 ^ n137 ;
  assign n3303 = n950 ^ n507 ;
  assign n3305 = n3304 ^ n3303 ;
  assign n3309 = n3308 ^ n3305 ;
  assign n3312 = n3311 ^ n3309 ;
  assign n3322 = n3321 ^ n3312 ;
  assign n3297 = n637 ^ n322 ;
  assign n3296 = n1845 ^ n1077 ;
  assign n3298 = n3297 ^ n3296 ;
  assign n3295 = n592 ^ n419 ;
  assign n3299 = n3298 ^ n3295 ;
  assign n3292 = n2749 ^ n778 ;
  assign n3293 = n3292 ^ n340 ;
  assign n3290 = n943 ^ n353 ;
  assign n3291 = n3290 ^ n437 ;
  assign n3294 = n3293 ^ n3291 ;
  assign n3300 = n3299 ^ n3294 ;
  assign n3289 = n4722 ^ n2894 ;
  assign n3301 = n3300 ^ n3289 ;
  assign n3302 = n3301 ^ n2484 ;
  assign n3323 = n3322 ^ n3302 ;
  assign n3324 = ~n3288 & ~n3323 ;
  assign n3325 = ~n3252 & n3324 ;
  assign n3326 = ~n2712 & ~n3325 ;
  assign n3327 = n2657 & ~n3326 ;
  assign n3328 = ~n2589 & ~n3327 ;
  assign n3329 = n2552 & ~n3328 ;
  assign n3330 = ~n2467 & ~n3329 ;
  assign n3331 = n2371 & ~n3330 ;
  assign n3332 = ~n2288 & ~n3331 ;
  assign n3333 = n2199 & ~n3332 ;
  assign n3334 = ~n2095 & ~n3333 ;
  assign n3335 = n3334 ^ n1897 ;
  assign n2096 = n2095 ^ n1897 ;
  assign n3336 = n3335 ^ n2096 ;
  assign n3337 = ~n1972 & ~n3336 ;
  assign n3338 = n3337 ^ n2096 ;
  assign n3339 = ~n1974 & ~n3338 ;
  assign n3340 = n3339 ^ n1541 ;
  assign n3371 = n2500 ^ n2054 ;
  assign n3370 = n243 ^ n117 ;
  assign n3372 = n3371 ^ n3370 ;
  assign n3366 = n609 ^ n230 ;
  assign n3367 = n3366 ^ n195 ;
  assign n3368 = n3367 ^ n737 ;
  assign n3365 = n1404 ^ n480 ;
  assign n3369 = n3368 ^ n3365 ;
  assign n3373 = n3372 ^ n3369 ;
  assign n3362 = n213 ^ n138 ;
  assign n3363 = n3362 ^ n773 ;
  assign n3364 = n3363 ^ n1440 ;
  assign n3374 = n3373 ^ n3364 ;
  assign n3358 = n1129 ^ n427 ;
  assign n3359 = n3358 ^ n645 ;
  assign n3357 = n2998 ^ n517 ;
  assign n3360 = n3359 ^ n3357 ;
  assign n3355 = n1702 ^ n389 ;
  assign n3356 = n3355 ^ n3203 ;
  assign n3361 = n3360 ^ n3356 ;
  assign n3375 = n3374 ^ n3361 ;
  assign n3351 = n1630 ^ n562 ;
  assign n3352 = n3351 ^ n845 ;
  assign n3349 = n861 ^ n261 ;
  assign n3350 = n3349 ^ n668 ;
  assign n3353 = n3352 ^ n3350 ;
  assign n3346 = n1844 ^ n950 ;
  assign n3345 = n3209 ^ n876 ;
  assign n3347 = n3346 ^ n3345 ;
  assign n3344 = n791 ^ n426 ;
  assign n3348 = n3347 ^ n3344 ;
  assign n3354 = n3353 ^ n3348 ;
  assign n3376 = n3375 ^ n3354 ;
  assign n3421 = n2107 ^ n369 ;
  assign n3422 = n3421 ^ n199 ;
  assign n3423 = n3422 ^ n501 ;
  assign n3420 = n677 ^ n526 ;
  assign n3424 = n3423 ^ n3420 ;
  assign n3418 = n2363 ^ n1653 ;
  assign n3417 = n2975 ^ n1517 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n3425 = n3424 ^ n3419 ;
  assign n3414 = n2425 ^ n1064 ;
  assign n3415 = n3414 ^ n1644 ;
  assign n3413 = n1285 ^ n476 ;
  assign n3416 = n3415 ^ n3413 ;
  assign n3426 = n3425 ^ n3416 ;
  assign n3409 = n898 ^ n742 ;
  assign n3407 = n1106 ^ n179 ;
  assign n3408 = n3407 ^ n926 ;
  assign n3410 = n3409 ^ n3408 ;
  assign n3405 = n437 ^ n337 ;
  assign n3404 = n379 ^ n150 ;
  assign n3406 = n3405 ^ n3404 ;
  assign n3411 = n3410 ^ n3406 ;
  assign n3402 = n3315 ^ n2828 ;
  assign n3401 = n572 ^ n322 ;
  assign n3403 = n3402 ^ n3401 ;
  assign n3412 = n3411 ^ n3403 ;
  assign n3427 = n3426 ^ n3412 ;
  assign n3395 = n788 ^ n211 ;
  assign n3396 = n3395 ^ n471 ;
  assign n3393 = n570 ^ n189 ;
  assign n3392 = n522 ^ n171 ;
  assign n3394 = n3393 ^ n3392 ;
  assign n3397 = n3396 ^ n3394 ;
  assign n3389 = n642 ^ n484 ;
  assign n3390 = n3389 ^ n722 ;
  assign n3387 = n489 ^ n347 ;
  assign n3386 = n546 ^ n495 ;
  assign n3388 = n3387 ^ n3386 ;
  assign n3391 = n3390 ^ n3388 ;
  assign n3398 = n3397 ^ n3391 ;
  assign n3383 = n2359 ^ n928 ;
  assign n3384 = n3383 ^ n414 ;
  assign n3382 = n2924 ^ n873 ;
  assign n3385 = n3384 ^ n3382 ;
  assign n3399 = n3398 ^ n3385 ;
  assign n3380 = n2964 ^ n1456 ;
  assign n3378 = n2781 ^ n2025 ;
  assign n3377 = n1176 ^ n523 ;
  assign n3379 = n3378 ^ n3377 ;
  assign n3381 = n3380 ^ n3379 ;
  assign n3400 = n3399 ^ n3381 ;
  assign n3428 = n3427 ^ n3400 ;
  assign n3429 = ~n3376 & ~n3428 ;
  assign n3430 = n3124 & n3429 ;
  assign n3431 = n3430 ^ n3429 ;
  assign n3432 = n3431 ^ n3124 ;
  assign n3433 = n3196 & n3432 ;
  assign n3434 = ~n3055 & ~n3433 ;
  assign n3435 = n3022 & ~n3434 ;
  assign n3436 = ~n3249 & ~n3435 ;
  assign n3437 = n3436 ^ n3248 ;
  assign n3438 = n2935 & n3437 ;
  assign n3439 = n3438 ^ n3249 ;
  assign n3440 = ~n2839 & ~n3439 ;
  assign n3343 = n3251 ^ n3250 ;
  assign n3441 = n3440 ^ n3343 ;
  assign n3442 = n2748 & n3441 ;
  assign n3443 = ~n3324 & ~n3442 ;
  assign n3444 = n2712 & ~n3443 ;
  assign n3445 = ~n2657 & ~n3444 ;
  assign n3446 = n2589 & ~n3445 ;
  assign n3447 = ~n2552 & ~n3446 ;
  assign n3448 = n2467 & ~n3447 ;
  assign n3449 = ~n2371 & ~n3448 ;
  assign n3450 = n2288 & ~n3449 ;
  assign n3451 = ~n2199 & ~n3450 ;
  assign n3456 = ~n1897 & n3451 ;
  assign n3457 = ~n3340 & n3456 ;
  assign n3458 = n3457 ^ n3340 ;
  assign n3459 = n3458 ^ n1541 ;
  assign n3460 = n1973 & n3459 ;
  assign n3461 = n3460 ^ n1972 ;
  assign n3462 = n1821 & n3461 ;
  assign n3463 = n1751 ^ n1670 ;
  assign n3464 = n1670 ^ n1450 ;
  assign n3465 = n1819 ^ n1670 ;
  assign n3466 = ~n3464 & n3465 ;
  assign n3474 = ~n1541 & n3466 ;
  assign n3475 = n1751 & n3474 ;
  assign n3476 = n3475 ^ n1751 ;
  assign n3467 = n3466 ^ n3464 ;
  assign n3468 = n3467 ^ n1751 ;
  assign n3477 = n3476 ^ n3468 ;
  assign n3478 = n3463 & n3477 ;
  assign n3479 = n3478 ^ n1670 ;
  assign n3480 = ~n3462 & ~n3479 ;
  assign n3483 = n3480 ^ n1450 ;
  assign n3481 = ~n1450 & n3480 ;
  assign n3484 = n3483 ^ n3481 ;
  assign n3485 = ~n1345 & ~n3484 ;
  assign n3482 = n1345 & ~n3481 ;
  assign n3486 = n3485 ^ n3482 ;
  assign n3487 = n3485 ^ n1248 ;
  assign n3488 = n3487 ^ n3485 ;
  assign n3489 = n3486 & n3488 ;
  assign n3490 = n3489 ^ n3485 ;
  assign n3491 = n1250 & ~n3490 ;
  assign n3492 = n3491 ^ n1248 ;
  assign n3493 = n3492 ^ n1119 ;
  assign n3494 = n1119 ^ n856 ;
  assign n3495 = ~n3493 & n3494 ;
  assign n3496 = n856 & ~n3495 ;
  assign n3497 = n3496 ^ n3495 ;
  assign n3498 = n698 & n3497 ;
  assign n3499 = ~n540 & ~n3498 ;
  assign n3500 = n408 & ~n3499 ;
  assign n3502 = n276 ^ n228 ;
  assign n280 = n279 ^ n278 ;
  assign n271 = n270 ^ n269 ;
  assign n281 = n280 ^ n271 ;
  assign n263 = n262 ^ n261 ;
  assign n266 = n265 ^ n263 ;
  assign n268 = n267 ^ n266 ;
  assign n282 = n281 ^ n268 ;
  assign n297 = n296 ^ n295 ;
  assign n303 = n302 ^ n297 ;
  assign n304 = ~n282 & ~n303 ;
  assign n3503 = n3502 ^ n304 ;
  assign n3504 = n3503 ^ n327 ;
  assign n3501 = n367 ^ n230 ;
  assign n3505 = n3504 ^ n3501 ;
  assign n3506 = ~n698 & ~n3496 ;
  assign n3507 = n540 & ~n3506 ;
  assign n3508 = ~n408 & ~n3507 ;
  assign n3509 = n3505 & ~n3508 ;
  assign n3510 = ~n3500 & ~n3509 ;
  assign n3511 = n3510 ^ n3509 ;
  assign n3512 = n3511 ^ n3505 ;
  assign n3513 = n3512 ^ n3509 ;
  assign n3514 = n368 & n3513 ;
  assign n3515 = n3514 ^ n3509 ;
  assign n6141 = x15 ^ x14 ;
  assign n23445 = x16 & n6141 ;
  assign n16849 = x17 & n6141 ;
  assign n6147 = n16849 ^ n6141 ;
  assign n6148 = n23445 ^ n6147 ;
  assign n6163 = n6148 ^ n6141 ;
  assign n6386 = n3515 & n6163 ;
  assign n3930 = n3495 ^ n698 ;
  assign n5212 = ~x17 & x18 ;
  assign n5214 = n5212 ^ x17 ;
  assign n5213 = n5212 ^ x18 ;
  assign n5215 = n5214 ^ n5213 ;
  assign n27193 = x20 & n5215 ;
  assign n5216 = x19 & n5215 ;
  assign n5217 = n5216 ^ n5215 ;
  assign n5220 = n27193 ^ n5217 ;
  assign n5221 = n5220 ^ n5215 ;
  assign n5980 = ~n3930 & n5221 ;
  assign n5978 = ~n698 & n5220 ;
  assign n5425 = n5216 ^ x19 ;
  assign n5426 = n5425 ^ n5213 ;
  assign n5975 = ~n856 & n5426 ;
  assign n13431 = n5216 ^ n5214 ;
  assign n5224 = x20 ^ x19 ;
  assign n5218 = x20 & ~n5215 ;
  assign n5225 = n5218 ^ n5214 ;
  assign n5226 = ~n5224 & n5225 ;
  assign n13432 = n13431 ^ n5226 ;
  assign n13433 = n13432 ^ x20 ;
  assign n5974 = ~n1119 & n13433 ;
  assign n5976 = n5975 ^ n5974 ;
  assign n5977 = n5976 ^ x20 ;
  assign n5979 = n5978 ^ n5977 ;
  assign n5981 = n5980 ^ n5979 ;
  assign n4025 = n598 ^ n480 ;
  assign n4235 = n4025 ^ n470 ;
  assign n5564 = n4235 ^ n1307 ;
  assign n5563 = n1975 ^ n634 ;
  assign n5565 = n5564 ^ n5563 ;
  assign n5560 = n1276 ^ n265 ;
  assign n5561 = n5560 ^ n999 ;
  assign n5562 = n5561 ^ n1095 ;
  assign n5566 = n5565 ^ n5562 ;
  assign n3565 = n1064 ^ n546 ;
  assign n5557 = n3565 ^ n1518 ;
  assign n3767 = n845 ^ n507 ;
  assign n5556 = n3767 ^ n590 ;
  assign n5558 = n5557 ^ n5556 ;
  assign n5554 = n2425 ^ n618 ;
  assign n5551 = n416 ^ n395 ;
  assign n5552 = n5551 ^ n369 ;
  assign n5553 = n5552 ^ n2990 ;
  assign n5555 = n5554 ^ n5553 ;
  assign n5559 = n5558 ^ n5555 ;
  assign n5567 = n5566 ^ n5559 ;
  assign n5499 = n2379 ^ n236 ;
  assign n5500 = n5499 ^ n382 ;
  assign n5496 = n719 ^ n452 ;
  assign n5497 = n5496 ^ n730 ;
  assign n5498 = n5497 ^ n335 ;
  assign n5501 = n5500 ^ n5498 ;
  assign n5494 = n836 ^ n528 ;
  assign n5495 = n5494 ^ n346 ;
  assign n5502 = n5501 ^ n5495 ;
  assign n5492 = n2025 ^ n926 ;
  assign n5491 = n1699 ^ n1690 ;
  assign n5493 = n5492 ^ n5491 ;
  assign n5503 = n5502 ^ n5493 ;
  assign n5568 = n5567 ^ n5503 ;
  assign n4763 = n684 ^ n230 ;
  assign n4764 = n4763 ^ n150 ;
  assign n4761 = n641 ^ n331 ;
  assign n4762 = n4761 ^ n1735 ;
  assign n4765 = n4764 ^ n4762 ;
  assign n4766 = n4765 ^ n3031 ;
  assign n5549 = n4766 ^ n2355 ;
  assign n5545 = n3226 ^ n1465 ;
  assign n5543 = n721 ^ n430 ;
  assign n3571 = n773 ^ n490 ;
  assign n5544 = n5543 ^ n3571 ;
  assign n5546 = n5545 ^ n5544 ;
  assign n5542 = n1935 ^ n209 ;
  assign n5547 = n5546 ^ n5542 ;
  assign n5539 = n436 ^ n142 ;
  assign n5540 = n5539 ^ n1603 ;
  assign n5537 = n1106 ^ n1036 ;
  assign n5538 = n5537 ^ n806 ;
  assign n5541 = n5540 ^ n5538 ;
  assign n5548 = n5547 ^ n5541 ;
  assign n5550 = n5549 ^ n5548 ;
  assign n5569 = n5568 ^ n5550 ;
  assign n5570 = ~n924 & ~n5569 ;
  assign n5487 = n2105 ^ n1000 ;
  assign n3573 = n680 ^ n377 ;
  assign n5486 = n3573 ^ n385 ;
  assign n5488 = n5487 ^ n5486 ;
  assign n5485 = n1176 ^ n794 ;
  assign n5489 = n5488 ^ n5485 ;
  assign n5483 = n943 ^ n399 ;
  assign n3560 = n398 ^ n234 ;
  assign n3559 = n369 ^ n171 ;
  assign n3561 = n3560 ^ n3559 ;
  assign n3562 = n3561 ^ n3001 ;
  assign n5484 = n5483 ^ n3562 ;
  assign n5490 = n5489 ^ n5484 ;
  assign n5504 = n5503 ^ n5490 ;
  assign n4058 = n1609 ^ n555 ;
  assign n5506 = n4058 ^ n2724 ;
  assign n4908 = n1898 ^ n577 ;
  assign n5505 = n4908 ^ n2161 ;
  assign n5507 = n5506 ^ n5505 ;
  assign n4193 = n2082 ^ n468 ;
  assign n4192 = n1187 ^ n511 ;
  assign n4194 = n4193 ^ n4192 ;
  assign n233 = n232 ^ n230 ;
  assign n4190 = n842 ^ n233 ;
  assign n4191 = n4190 ^ n845 ;
  assign n4195 = n4194 ^ n4191 ;
  assign n3740 = n956 ^ n411 ;
  assign n4188 = n3740 ^ n975 ;
  assign n4189 = n4188 ^ n1556 ;
  assign n4196 = n4195 ^ n4189 ;
  assign n5508 = n5507 ^ n4196 ;
  assign n4100 = n1157 ^ n1011 ;
  assign n4098 = n784 ^ n533 ;
  assign n4099 = n4098 ^ n3370 ;
  assign n4101 = n4100 ^ n4099 ;
  assign n4095 = n941 ^ n903 ;
  assign n4096 = n4095 ^ n1279 ;
  assign n4093 = n2162 ^ n209 ;
  assign n4094 = n4093 ^ n825 ;
  assign n4097 = n4096 ^ n4094 ;
  assign n4102 = n4101 ^ n4097 ;
  assign n5509 = n5508 ^ n4102 ;
  assign n5527 = n684 ^ n211 ;
  assign n5526 = n640 ^ n430 ;
  assign n5528 = n5527 ^ n5526 ;
  assign n5529 = n5528 ^ n409 ;
  assign n5525 = n1514 ^ n188 ;
  assign n5530 = n5529 ^ n5525 ;
  assign n5524 = n2982 ^ n1727 ;
  assign n5531 = n5530 ^ n5524 ;
  assign n5532 = n5531 ^ n1739 ;
  assign n5520 = n1252 ^ n1020 ;
  assign n3753 = n1495 ^ n570 ;
  assign n5521 = n5520 ^ n3753 ;
  assign n5517 = n778 ^ n657 ;
  assign n5518 = n5517 ^ n458 ;
  assign n5515 = n2457 ^ n395 ;
  assign n5514 = n436 ^ n215 ;
  assign n5516 = n5515 ^ n5514 ;
  assign n5519 = n5518 ^ n5516 ;
  assign n5522 = n5521 ^ n5519 ;
  assign n5511 = n2432 ^ n213 ;
  assign n5512 = n5511 ^ n688 ;
  assign n3604 = n753 ^ n296 ;
  assign n5510 = n3604 ^ n149 ;
  assign n5513 = n5512 ^ n5510 ;
  assign n5523 = n5522 ^ n5513 ;
  assign n5533 = n5532 ^ n5523 ;
  assign n5534 = ~n5509 & ~n5533 ;
  assign n5535 = ~n5504 & n5534 ;
  assign n5771 = n5570 ^ n5535 ;
  assign n5772 = n5570 ^ x11 ;
  assign n5773 = ~n5771 & n5772 ;
  assign n5774 = n5773 ^ x11 ;
  assign n5762 = ~n61 & ~n2199 ;
  assign n3518 = x30 ^ x29 ;
  assign n5381 = ~n2095 & n3518 ;
  assign n5763 = n5762 ^ n5381 ;
  assign n5468 = ~n61 & ~n2288 ;
  assign n5764 = n5763 ^ n5468 ;
  assign n5386 = n52 & ~n2199 ;
  assign n5765 = n5764 ^ n5386 ;
  assign n5759 = n3451 ^ n3333 ;
  assign n5760 = n5759 ^ n2095 ;
  assign n5761 = n3518 & n5760 ;
  assign n5766 = n5765 ^ n5761 ;
  assign n5767 = x31 & n5766 ;
  assign n5768 = n5767 ^ n5763 ;
  assign n5794 = n5774 ^ n5768 ;
  assign n4716 = n485 ^ n234 ;
  assign n4717 = n4716 ^ n240 ;
  assign n4718 = n4717 ^ n2569 ;
  assign n4113 = n480 ^ n251 ;
  assign n4714 = n4113 ^ n845 ;
  assign n4519 = n411 ^ n153 ;
  assign n4713 = n4519 ^ n124 ;
  assign n4715 = n4714 ^ n4713 ;
  assign n4719 = n4718 ^ n4715 ;
  assign n4710 = n773 ^ n248 ;
  assign n4711 = n4710 ^ n431 ;
  assign n4712 = n4711 ^ n2363 ;
  assign n4720 = n4719 ^ n4712 ;
  assign n4742 = n905 ^ n390 ;
  assign n4743 = n4742 ^ n970 ;
  assign n4744 = n4743 ^ n3061 ;
  assign n4740 = n1489 ^ n108 ;
  assign n4738 = n776 ^ n507 ;
  assign n4739 = n4738 ^ n555 ;
  assign n4741 = n4740 ^ n4739 ;
  assign n4745 = n4744 ^ n4741 ;
  assign n4735 = n1518 ^ n142 ;
  assign n4736 = n4735 ^ n1304 ;
  assign n4734 = n1347 ^ n610 ;
  assign n4737 = n4736 ^ n4734 ;
  assign n4746 = n4745 ^ n4737 ;
  assign n4731 = n938 ^ n742 ;
  assign n4730 = n2025 ^ n1525 ;
  assign n4732 = n4731 ^ n4730 ;
  assign n4728 = n653 ^ n117 ;
  assign n4727 = n1544 ^ n813 ;
  assign n4729 = n4728 ^ n4727 ;
  assign n4733 = n4732 ^ n4729 ;
  assign n4747 = n4746 ^ n4733 ;
  assign n4723 = n4722 ^ n320 ;
  assign n4724 = n4723 ^ n993 ;
  assign n4721 = n1506 ^ n495 ;
  assign n4725 = n4724 ^ n4721 ;
  assign n4726 = n4725 ^ n3006 ;
  assign n4748 = n4747 ^ n4726 ;
  assign n4782 = n659 ^ n484 ;
  assign n4783 = n4782 ^ n3013 ;
  assign n3742 = n908 ^ n791 ;
  assign n4781 = n3742 ^ n1209 ;
  assign n4784 = n4783 ^ n4781 ;
  assign n4087 = n1307 ^ n341 ;
  assign n4785 = n4784 ^ n4087 ;
  assign n4778 = n900 ^ n197 ;
  assign n4777 = n1239 ^ n335 ;
  assign n4779 = n4778 ^ n4777 ;
  assign n3563 = n3112 ^ n184 ;
  assign n4780 = n4779 ^ n3563 ;
  assign n4786 = n4785 ^ n4780 ;
  assign n4773 = n663 ^ n511 ;
  assign n3713 = n600 ^ n519 ;
  assign n4771 = n3713 ^ n409 ;
  assign n4772 = n4771 ^ n237 ;
  assign n4774 = n4773 ^ n4772 ;
  assign n4769 = n721 ^ n446 ;
  assign n4770 = n4769 ^ n1277 ;
  assign n4775 = n4774 ^ n4770 ;
  assign n4776 = n4775 ^ n1138 ;
  assign n4787 = n4786 ^ n4776 ;
  assign n4758 = n779 ^ n520 ;
  assign n4759 = n4758 ^ n1645 ;
  assign n4760 = n4759 ^ n862 ;
  assign n4767 = n4766 ^ n4760 ;
  assign n4754 = n1085 ^ n594 ;
  assign n4755 = n4754 ^ n524 ;
  assign n4752 = n603 ^ n426 ;
  assign n4753 = n4752 ^ n348 ;
  assign n4756 = n4755 ^ n4753 ;
  assign n4749 = n493 ^ n199 ;
  assign n4750 = n4749 ^ n1020 ;
  assign n4751 = n4750 ^ n1533 ;
  assign n4757 = n4756 ^ n4751 ;
  assign n4768 = n4767 ^ n4757 ;
  assign n4788 = n4787 ^ n4768 ;
  assign n4789 = ~n4748 & ~n4788 ;
  assign n4790 = ~n4720 & n4789 ;
  assign n5795 = n5794 ^ n4790 ;
  assign n3833 = x27 ^ x26 ;
  assign n3834 = ~x28 & n3833 ;
  assign n3829 = x26 & x27 ;
  assign n3832 = n3829 ^ x28 ;
  assign n3835 = n3834 ^ n3832 ;
  assign n3836 = x29 & n3835 ;
  assign n3830 = x28 & n3829 ;
  assign n3831 = n3830 ^ x29 ;
  assign n3837 = n3836 ^ n3831 ;
  assign n5757 = ~n1897 & n3837 ;
  assign n3985 = n3835 ^ n3833 ;
  assign n5755 = ~n1972 & n3985 ;
  assign n4883 = n2095 & ~n3451 ;
  assign n4884 = n4883 ^ n3334 ;
  assign n4887 = n3334 ^ n1972 ;
  assign n4888 = n4887 ^ n3334 ;
  assign n4889 = n4884 & n4888 ;
  assign n4890 = n4889 ^ n3334 ;
  assign n4891 = n1973 & ~n4890 ;
  assign n5065 = x29 ^ x28 ;
  assign n5751 = n4891 & n5065 ;
  assign n5752 = n5751 ^ n1541 ;
  assign n5753 = n3833 & ~n5752 ;
  assign n5754 = n5753 ^ x29 ;
  assign n5756 = n5755 ^ n5754 ;
  assign n5758 = n5757 ^ n5756 ;
  assign n5536 = n5535 ^ x11 ;
  assign n5571 = n5570 ^ n5536 ;
  assign n5479 = n3450 ^ n3332 ;
  assign n5480 = n5479 ^ n2199 ;
  assign n3801 = n61 ^ x31 ;
  assign n3802 = ~n3518 & n3801 ;
  assign n22543 = x31 & n3802 ;
  assign n3799 = ~x31 & n52 ;
  assign n3800 = n3799 ^ x31 ;
  assign n5280 = n3800 ^ n52 ;
  assign n22005 = n22543 ^ n5280 ;
  assign n5481 = n5480 & n22005 ;
  assign n5474 = ~n2199 & n3518 ;
  assign n5467 = ~n61 & ~n2371 ;
  assign n5469 = n5468 ^ n5467 ;
  assign n5475 = n5474 ^ n5469 ;
  assign n5476 = ~x31 & n5475 ;
  assign n5477 = n5476 ^ n5467 ;
  assign n5465 = n5280 ^ x31 ;
  assign n5466 = ~n2288 & n5465 ;
  assign n5478 = n5477 ^ n5466 ;
  assign n5482 = n5481 ^ n5478 ;
  assign n5572 = n5571 ^ n5482 ;
  assign n5593 = n3117 ^ n562 ;
  assign n5592 = n547 ^ n211 ;
  assign n5594 = n5593 ^ n5592 ;
  assign n5590 = n1014 ^ n322 ;
  assign n5591 = n5590 ^ n908 ;
  assign n5595 = n5594 ^ n5591 ;
  assign n4034 = n1307 ^ n114 ;
  assign n4035 = n4034 ^ n320 ;
  assign n5596 = n5595 ^ n4035 ;
  assign n5587 = n2201 ^ n462 ;
  assign n5586 = n544 ^ n434 ;
  assign n5588 = n5587 ^ n5586 ;
  assign n5589 = n5588 ^ n2883 ;
  assign n5597 = n5596 ^ n5589 ;
  assign n5581 = n346 ^ n232 ;
  assign n5582 = n5581 ^ n506 ;
  assign n5583 = n5582 ^ n2766 ;
  assign n4930 = n476 ^ n240 ;
  assign n5579 = n4930 ^ n867 ;
  assign n5580 = n5579 ^ n751 ;
  assign n5584 = n5583 ^ n5580 ;
  assign n5576 = n1161 ^ n459 ;
  assign n5573 = n847 ^ n533 ;
  assign n5574 = n5573 ^ n431 ;
  assign n5575 = n5574 ^ n846 ;
  assign n5577 = n5576 ^ n5575 ;
  assign n5578 = n5577 ^ n1535 ;
  assign n5585 = n5584 ^ n5578 ;
  assign n5598 = n5597 ^ n5585 ;
  assign n5629 = n4763 ^ n1384 ;
  assign n4012 = n741 ^ n247 ;
  assign n5628 = n4012 ^ n2828 ;
  assign n5630 = n5629 ^ n5628 ;
  assign n4181 = n831 ^ n446 ;
  assign n5626 = n4181 ^ n4025 ;
  assign n5625 = n2532 ^ n1653 ;
  assign n5627 = n5626 ^ n5625 ;
  assign n5631 = n5630 ^ n5627 ;
  assign n4159 = n2082 ^ n640 ;
  assign n4836 = n4159 ^ n820 ;
  assign n3555 = n1260 ^ n615 ;
  assign n3556 = n3555 ^ n542 ;
  assign n4835 = n3556 ^ n398 ;
  assign n4837 = n4836 ^ n4835 ;
  assign n5632 = n5631 ^ n4837 ;
  assign n5621 = n1252 ^ n354 ;
  assign n5622 = n5621 ^ n784 ;
  assign n5619 = n485 ^ n239 ;
  assign n5620 = n5619 ^ n773 ;
  assign n5623 = n5622 ^ n5620 ;
  assign n5624 = n5623 ^ n2133 ;
  assign n5633 = n5632 ^ n5624 ;
  assign n5615 = n2819 ^ n806 ;
  assign n4535 = n600 ^ n117 ;
  assign n5613 = n4535 ^ n903 ;
  assign n5614 = n5613 ^ n3067 ;
  assign n5616 = n5615 ^ n5614 ;
  assign n3533 = n440 ^ n243 ;
  assign n3534 = n3533 ^ n2018 ;
  assign n3532 = n1405 ^ n1135 ;
  assign n3535 = n3534 ^ n3532 ;
  assign n3529 = n343 ^ n197 ;
  assign n3530 = n3529 ^ n468 ;
  assign n3528 = n369 ^ n331 ;
  assign n3531 = n3530 ^ n3528 ;
  assign n3536 = n3535 ^ n3531 ;
  assign n5617 = n5616 ^ n3536 ;
  assign n3890 = n649 ^ n570 ;
  assign n5609 = n3890 ^ n723 ;
  assign n5608 = n5537 ^ n2352 ;
  assign n5610 = n5609 ^ n5608 ;
  assign n5605 = n928 ^ n153 ;
  assign n5606 = n5605 ^ n585 ;
  assign n5603 = n883 ^ n215 ;
  assign n5604 = n5603 ^ n275 ;
  assign n5607 = n5606 ^ n5604 ;
  assign n5611 = n5610 ^ n5607 ;
  assign n5314 = n577 ^ n149 ;
  assign n5600 = n5314 ^ n193 ;
  assign n5599 = n2949 ^ n974 ;
  assign n5601 = n5600 ^ n5599 ;
  assign n5602 = n5601 ^ n2527 ;
  assign n5612 = n5611 ^ n5602 ;
  assign n5618 = n5617 ^ n5612 ;
  assign n5634 = n5633 ^ n5618 ;
  assign n5635 = ~n5598 & ~n5634 ;
  assign n5636 = n5635 ^ x8 ;
  assign n5657 = n755 ^ n179 ;
  assign n5656 = n1125 ^ n327 ;
  assign n5658 = n5657 ^ n5656 ;
  assign n4503 = n1389 ^ n489 ;
  assign n4504 = n4503 ^ n1886 ;
  assign n5659 = n5658 ^ n4504 ;
  assign n4814 = n446 ^ n137 ;
  assign n5652 = n4814 ^ n803 ;
  assign n5653 = n5652 ^ n484 ;
  assign n4942 = n1689 ^ n905 ;
  assign n5651 = n4942 ^ n511 ;
  assign n5654 = n5653 ^ n5651 ;
  assign n5655 = n5654 ^ n2069 ;
  assign n5660 = n5659 ^ n5655 ;
  assign n5647 = n1936 ^ n840 ;
  assign n5648 = n5647 ^ n2349 ;
  assign n3626 = n895 ^ n250 ;
  assign n5644 = n3626 ^ n184 ;
  assign n5645 = n5644 ^ n527 ;
  assign n5643 = n1906 ^ n157 ;
  assign n5646 = n5645 ^ n5643 ;
  assign n5649 = n5648 ^ n5646 ;
  assign n5639 = n3890 ^ n379 ;
  assign n5640 = n5639 ^ n874 ;
  assign n5638 = n495 ^ n172 ;
  assign n5641 = n5640 ^ n5638 ;
  assign n5637 = n1187 ^ n663 ;
  assign n5642 = n5641 ^ n5637 ;
  assign n5650 = n5649 ^ n5642 ;
  assign n5661 = n5660 ^ n5650 ;
  assign n4547 = n1581 ^ n634 ;
  assign n4548 = n4547 ^ n272 ;
  assign n4549 = n4548 ^ n505 ;
  assign n4546 = n1129 ^ n602 ;
  assign n4550 = n4549 ^ n4546 ;
  assign n3762 = n493 ^ n429 ;
  assign n4543 = n3762 ^ n1362 ;
  assign n4541 = n1189 ^ n550 ;
  assign n4542 = n4541 ^ n2205 ;
  assign n4544 = n4543 ^ n4542 ;
  assign n4545 = n4544 ^ n1804 ;
  assign n4551 = n4550 ^ n4545 ;
  assign n4537 = n2242 ^ n664 ;
  assign n4538 = n4537 ^ n2720 ;
  assign n4536 = n4535 ^ n2742 ;
  assign n4539 = n4538 ^ n4536 ;
  assign n4532 = n1577 ^ n389 ;
  assign n4533 = n4532 ^ n657 ;
  assign n4530 = n975 ^ n232 ;
  assign n4531 = n4530 ^ n385 ;
  assign n4534 = n4533 ^ n4531 ;
  assign n4540 = n4539 ^ n4534 ;
  assign n4552 = n4551 ^ n4540 ;
  assign n5662 = n5661 ^ n4552 ;
  assign n5684 = n2243 ^ n762 ;
  assign n5685 = n5684 ^ n836 ;
  assign n5682 = n2303 ^ n1161 ;
  assign n5683 = n5682 ^ n1953 ;
  assign n5686 = n5685 ^ n5683 ;
  assign n5687 = n5686 ^ n616 ;
  assign n5679 = n1037 ^ n296 ;
  assign n3663 = n478 ^ n348 ;
  assign n5680 = n5679 ^ n3663 ;
  assign n5678 = n1844 ^ n335 ;
  assign n5681 = n5680 ^ n5678 ;
  assign n5688 = n5687 ^ n5681 ;
  assign n4816 = n876 ^ n825 ;
  assign n5674 = n4816 ^ n390 ;
  assign n5675 = n5674 ^ n578 ;
  assign n5671 = n1077 ^ n653 ;
  assign n5672 = n5671 ^ n886 ;
  assign n5669 = n592 ^ n320 ;
  assign n5670 = n5669 ^ n667 ;
  assign n5673 = n5672 ^ n5670 ;
  assign n5676 = n5675 ^ n5673 ;
  assign n5665 = n928 ^ n603 ;
  assign n3655 = n318 ^ n118 ;
  assign n5663 = n3655 ^ n730 ;
  assign n5664 = n5663 ^ n564 ;
  assign n5666 = n5665 ^ n5664 ;
  assign n5667 = n5666 ^ n1064 ;
  assign n5668 = n5667 ^ n1711 ;
  assign n5677 = n5676 ^ n5668 ;
  assign n5689 = n5688 ^ n5677 ;
  assign n5690 = ~n5662 & ~n5689 ;
  assign n5691 = n5690 ^ n5635 ;
  assign n5692 = n5636 & ~n5691 ;
  assign n5693 = n5692 ^ x8 ;
  assign n5694 = n5693 ^ n5570 ;
  assign n5707 = ~n61 & ~n2467 ;
  assign n5708 = n5707 ^ n2371 ;
  assign n5695 = n3448 ^ n3330 ;
  assign n5696 = n5695 ^ n2371 ;
  assign n5698 = n5696 ^ n2467 ;
  assign n5697 = n5696 ^ n2552 ;
  assign n5699 = n5698 ^ n5697 ;
  assign n5702 = x30 & n5699 ;
  assign n5703 = n5702 ^ n5698 ;
  assign n5704 = ~n3518 & ~n5703 ;
  assign n5705 = n5704 ^ n5696 ;
  assign n5706 = n5705 ^ n5467 ;
  assign n5709 = n5708 ^ n5706 ;
  assign n5710 = n5709 ^ n5705 ;
  assign n5713 = ~n52 & ~n5710 ;
  assign n5714 = n5713 ^ n5705 ;
  assign n5715 = ~x31 & n5714 ;
  assign n5716 = n5715 ^ n5705 ;
  assign n5717 = n5716 ^ n5693 ;
  assign n5718 = ~n5694 & n5717 ;
  assign n5734 = n1879 ^ n653 ;
  assign n5732 = n838 ^ n484 ;
  assign n5733 = n5732 ^ n550 ;
  assign n5735 = n5734 ^ n5733 ;
  assign n5730 = n416 ^ n346 ;
  assign n5731 = n5730 ^ n1960 ;
  assign n5736 = n5735 ^ n5731 ;
  assign n5727 = n3008 ^ n1076 ;
  assign n5726 = n2988 ^ n1095 ;
  assign n5728 = n5727 ^ n5726 ;
  assign n5724 = n2205 ^ n615 ;
  assign n5725 = n5724 ^ n915 ;
  assign n5729 = n5728 ^ n5725 ;
  assign n5737 = n5736 ^ n5729 ;
  assign n5722 = n1084 ^ n871 ;
  assign n5721 = n2677 ^ n1060 ;
  assign n5723 = n5722 ^ n5721 ;
  assign n5738 = n5737 ^ n5723 ;
  assign n4106 = n2373 ^ n462 ;
  assign n4105 = n547 ^ n336 ;
  assign n4107 = n4106 ^ n4105 ;
  assign n4103 = n1014 ^ n664 ;
  assign n4104 = n4103 ^ n1037 ;
  assign n4108 = n4107 ^ n4104 ;
  assign n5739 = n5738 ^ n4108 ;
  assign n5740 = ~n1599 & ~n5739 ;
  assign n5741 = ~n2370 & n5740 ;
  assign n5742 = n5741 ^ n5570 ;
  assign n5743 = n5718 & ~n5742 ;
  assign n5719 = n5570 ^ n5482 ;
  assign n5744 = n5743 ^ n5719 ;
  assign n5745 = ~n5572 & ~n5744 ;
  assign n5746 = n5745 ^ n5571 ;
  assign n5781 = n5758 ^ n5746 ;
  assign n5796 = n5795 ^ n5781 ;
  assign n35 = x21 ^ x20 ;
  assign n38 = x22 & n35 ;
  assign n39 = n38 ^ x22 ;
  assign n33 = ~x20 & ~x21 ;
  assign n37 = n35 ^ n33 ;
  assign n40 = n39 ^ n37 ;
  assign n34 = ~x22 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n34 ^ x23 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n42 & n44 ;
  assign n4651 = n45 ^ n34 ;
  assign n5445 = ~n1345 & n4651 ;
  assign n5444 = ~n40 & ~n990 ;
  assign n5446 = n5445 ^ n5444 ;
  assign n4332 = n990 & ~n3485 ;
  assign n4331 = ~n990 & ~n3482 ;
  assign n4333 = n4332 ^ n4331 ;
  assign n5437 = n1248 ^ x23 ;
  assign n5438 = n5437 ^ x22 ;
  assign n5439 = n5438 ^ n1248 ;
  assign n5440 = ~n4333 & n5439 ;
  assign n5441 = n5440 ^ n1248 ;
  assign n5442 = n35 & ~n5441 ;
  assign n5443 = n5442 ^ x23 ;
  assign n5447 = n5446 ^ n5443 ;
  assign n5843 = n5796 ^ n5447 ;
  assign n4433 = n97 ^ n88 ;
  assign n4434 = n4433 ^ n79 ;
  assign n4435 = n4434 ^ n96 ;
  assign n4488 = n3461 ^ n1541 ;
  assign n4485 = n1541 & n3461 ;
  assign n4489 = n4488 ^ n4485 ;
  assign n4490 = n1819 & n4489 ;
  assign n4491 = ~n1670 & ~n4490 ;
  assign n4486 = ~n1819 & ~n4485 ;
  assign n4487 = n1670 & ~n4486 ;
  assign n4492 = n4491 ^ n4487 ;
  assign n4690 = n4492 ^ n1751 ;
  assign n5792 = ~n4435 & n4690 ;
  assign n4600 = n203 ^ n89 ;
  assign n5790 = ~n1670 & n4600 ;
  assign n20603 = n20602 ^ n107 ;
  assign n5787 = ~n1819 & n20603 ;
  assign n5786 = ~n1751 & ~n4434 ;
  assign n5788 = n5787 ^ n5786 ;
  assign n5789 = n5788 ^ x26 ;
  assign n5791 = n5790 ^ n5789 ;
  assign n5793 = n5792 ^ n5791 ;
  assign n5797 = n5796 ^ n5793 ;
  assign n5809 = ~n2095 & n3837 ;
  assign n5807 = ~n1897 & n3985 ;
  assign n5285 = ~n1897 & n4884 ;
  assign n5286 = n5285 ^ n3334 ;
  assign n5803 = n5065 & n5286 ;
  assign n5804 = n5803 ^ n1972 ;
  assign n5805 = n3833 & ~n5804 ;
  assign n5806 = n5805 ^ x29 ;
  assign n5808 = n5807 ^ n5806 ;
  assign n5810 = n5809 ^ n5808 ;
  assign n5840 = n5810 ^ n5796 ;
  assign n5798 = n5744 ^ n5571 ;
  assign n5811 = n5810 ^ n5798 ;
  assign n3805 = n22543 ^ n61 ;
  assign n3806 = n3805 ^ x31 ;
  assign n3807 = n3806 ^ n3799 ;
  assign n5814 = n3449 ^ n3331 ;
  assign n5815 = n5814 ^ n2371 ;
  assign n5818 = n3807 & n5815 ;
  assign n5816 = n5815 ^ n2288 ;
  assign n5817 = n3518 & ~n5816 ;
  assign n5819 = n5818 ^ n5817 ;
  assign n5820 = n5819 ^ n2371 ;
  assign n5813 = n3801 & ~n5708 ;
  assign n5821 = n5820 ^ n5813 ;
  assign n5812 = n5741 ^ n5718 ;
  assign n5822 = n5821 ^ n5812 ;
  assign n5833 = ~n2095 & n3985 ;
  assign n5831 = n5821 ^ x29 ;
  assign n5828 = ~n4884 & n5065 ;
  assign n5829 = n5828 ^ n1897 ;
  assign n5830 = n3833 & ~n5829 ;
  assign n5832 = n5831 ^ n5830 ;
  assign n5834 = n5833 ^ n5832 ;
  assign n5823 = ~n2199 & n3837 ;
  assign n5835 = n5834 ^ n5823 ;
  assign n5836 = n5822 & ~n5835 ;
  assign n5837 = n5836 ^ n5821 ;
  assign n5838 = n5837 ^ n5810 ;
  assign n5839 = ~n5811 & ~n5838 ;
  assign n5841 = n5840 ^ n5839 ;
  assign n5842 = n5797 & n5841 ;
  assign n5844 = n5843 ^ n5842 ;
  assign n5769 = n5768 ^ n5758 ;
  assign n5782 = ~n5769 & n5781 ;
  assign n5770 = n5769 ^ n5746 ;
  assign n5775 = n5774 ^ n5770 ;
  assign n5385 = x31 & n3451 ;
  assign n5387 = n5386 ^ n5381 ;
  assign n5388 = n5385 & ~n5387 ;
  assign n5382 = x31 & ~n3333 ;
  assign n5383 = n5381 & n5382 ;
  assign n5375 = ~n3333 & n3450 ;
  assign n5376 = ~n61 & n5375 ;
  assign n5377 = n5376 ^ n61 ;
  assign n5367 = n2095 ^ x31 ;
  assign n5378 = n5377 ^ n5367 ;
  assign n5379 = n3801 & ~n5378 ;
  assign n5297 = n1600 ^ n153 ;
  assign n5296 = n600 ^ n188 ;
  assign n5298 = n5297 ^ n5296 ;
  assign n5294 = n452 ^ n213 ;
  assign n5295 = n5294 ^ n230 ;
  assign n5299 = n5298 ^ n5295 ;
  assign n5300 = n5299 ^ n2629 ;
  assign n3887 = n1136 ^ n547 ;
  assign n5337 = n3887 ^ n137 ;
  assign n5338 = n5337 ^ n2965 ;
  assign n5336 = n1175 ^ n592 ;
  assign n5339 = n5338 ^ n5336 ;
  assign n5333 = n2068 ^ n910 ;
  assign n5334 = n5333 ^ n1363 ;
  assign n5335 = n5334 ^ n1569 ;
  assign n5340 = n5339 ^ n5335 ;
  assign n5327 = n735 ^ n437 ;
  assign n5328 = n5327 ^ n522 ;
  assign n5326 = n815 ^ n663 ;
  assign n5329 = n5328 ^ n5326 ;
  assign n5330 = n5329 ^ n2125 ;
  assign n5325 = n3140 ^ n1754 ;
  assign n5331 = n5330 ^ n5325 ;
  assign n5322 = n1185 ^ n353 ;
  assign n5323 = n5322 ^ n382 ;
  assign n5321 = n842 ^ n339 ;
  assign n5324 = n5323 ^ n5321 ;
  assign n5332 = n5331 ^ n5324 ;
  assign n5341 = n5340 ^ n5332 ;
  assign n5316 = n826 ^ n714 ;
  assign n4857 = n1189 ^ n645 ;
  assign n5315 = n5314 ^ n4857 ;
  assign n5317 = n5316 ^ n5315 ;
  assign n5318 = n5317 ^ n1270 ;
  assign n5312 = n464 ^ n320 ;
  assign n5311 = n957 ^ n357 ;
  assign n5313 = n5312 ^ n5311 ;
  assign n5319 = n5318 ^ n5313 ;
  assign n5307 = n4098 ^ n261 ;
  assign n5308 = n5307 ^ n2481 ;
  assign n5306 = n1793 ^ n1689 ;
  assign n5309 = n5308 ^ n5306 ;
  assign n5302 = n741 ^ n476 ;
  assign n5303 = n5302 ^ n335 ;
  assign n5304 = n5303 ^ n484 ;
  assign n5301 = n597 ^ n435 ;
  assign n5305 = n5304 ^ n5301 ;
  assign n5310 = n5309 ^ n5305 ;
  assign n5320 = n5319 ^ n5310 ;
  assign n5342 = n5341 ^ n5320 ;
  assign n3685 = n801 ^ n546 ;
  assign n5354 = n3685 ^ n2493 ;
  assign n5355 = n5354 ^ n411 ;
  assign n5353 = n716 ^ n664 ;
  assign n5356 = n5355 ^ n5353 ;
  assign n5351 = n1768 ^ n550 ;
  assign n4173 = n1354 ^ n1284 ;
  assign n5352 = n5351 ^ n4173 ;
  assign n5357 = n5356 ^ n5352 ;
  assign n3880 = n1066 ^ n501 ;
  assign n3881 = n3880 ^ n465 ;
  assign n3882 = n3881 ^ n655 ;
  assign n3877 = n458 ^ n440 ;
  assign n3878 = n3877 ^ n684 ;
  assign n3876 = n2741 ^ n800 ;
  assign n3879 = n3878 ^ n3876 ;
  assign n3883 = n3882 ^ n3879 ;
  assign n5358 = n5357 ^ n3883 ;
  assign n5347 = n872 ^ n575 ;
  assign n5348 = n5347 ^ n586 ;
  assign n5349 = n5348 ^ n3655 ;
  assign n5343 = n861 ^ n557 ;
  assign n5344 = n5343 ^ n1360 ;
  assign n3645 = n969 ^ n572 ;
  assign n5345 = n5344 ^ n3645 ;
  assign n5346 = n5345 ^ n2679 ;
  assign n5350 = n5349 ^ n5346 ;
  assign n5359 = n5358 ^ n5350 ;
  assign n5360 = n5359 ^ n999 ;
  assign n5361 = ~n5342 & ~n5360 ;
  assign n5362 = ~n5300 & n5361 ;
  assign n5366 = n5362 ^ n52 ;
  assign n5368 = n5367 ^ n5366 ;
  assign n5380 = n5379 ^ n5368 ;
  assign n5384 = n5383 ^ n5380 ;
  assign n5389 = n5388 ^ n5384 ;
  assign n5365 = n1897 & n3518 ;
  assign n5390 = n5389 ^ n5365 ;
  assign n5776 = n5390 ^ n4790 ;
  assign n5777 = n5776 ^ n5390 ;
  assign n5778 = n5777 ^ n5774 ;
  assign n5779 = n5775 & n5778 ;
  assign n5780 = n5779 ^ n5776 ;
  assign n5783 = n5782 ^ n5780 ;
  assign n5463 = ~n1972 & n3837 ;
  assign n5460 = ~n1541 & n3985 ;
  assign n3976 = n3834 ^ n3833 ;
  assign n3977 = n3976 ^ x29 ;
  assign n3982 = n5065 ^ n3977 ;
  assign n3978 = x29 & ~n3833 ;
  assign n28382 = x29 & ~n3978 ;
  assign n3980 = n28382 ^ x28 ;
  assign n3983 = n3982 ^ n3980 ;
  assign n5154 = n4488 ^ n1819 ;
  assign n5458 = n3983 & ~n5154 ;
  assign n4493 = n1751 & n4492 ;
  assign n4494 = n4493 ^ n4487 ;
  assign n4495 = n4494 ^ n1450 ;
  assign n5455 = ~n4435 & ~n4495 ;
  assign n5453 = ~n1670 & n20603 ;
  assign n5450 = ~n1450 & ~n4434 ;
  assign n5449 = ~n1751 & n4600 ;
  assign n5451 = n5450 ^ n5449 ;
  assign n5452 = n5451 ^ x26 ;
  assign n5454 = n5453 ^ n5452 ;
  assign n5456 = n5455 ^ n5454 ;
  assign n5457 = n5456 ^ x29 ;
  assign n5459 = n5458 ^ n5457 ;
  assign n5461 = n5460 ^ n5459 ;
  assign n4368 = n28382 ^ n3833 ;
  assign n4369 = n4368 ^ n3976 ;
  assign n5448 = ~n1819 & n4369 ;
  assign n5462 = n5461 ^ n5448 ;
  assign n5464 = n5463 ^ n5462 ;
  assign n5784 = n5783 ^ n5464 ;
  assign n5973 = n5844 ^ n5784 ;
  assign n5982 = n5981 ^ n5973 ;
  assign n5992 = n5841 ^ n5793 ;
  assign n4307 = n3486 ^ n990 ;
  assign n13743 = x23 & ~n35 ;
  assign n13744 = n13743 ^ x23 ;
  assign n13745 = n13744 ^ n35 ;
  assign n4655 = n13745 ^ n38 ;
  assign n4656 = n4655 ^ n35 ;
  assign n5987 = n4307 & n4656 ;
  assign n5986 = ~n1450 & n4651 ;
  assign n5988 = n5987 ^ n5986 ;
  assign n5989 = n5988 ^ x23 ;
  assign n5984 = ~n40 & ~n1345 ;
  assign n5983 = ~n990 & n4655 ;
  assign n5985 = n5984 ^ n5983 ;
  assign n5990 = n5989 ^ n5985 ;
  assign n5993 = n5992 ^ n5990 ;
  assign n4985 = n4490 ^ n4486 ;
  assign n4986 = n4985 ^ n1670 ;
  assign n6120 = ~n4435 & n4986 ;
  assign n6118 = ~n1670 & ~n4434 ;
  assign n6115 = ~n1819 & n4600 ;
  assign n6114 = ~n1541 & n20603 ;
  assign n6116 = n6115 ^ n6114 ;
  assign n6117 = n6116 ^ x26 ;
  assign n6119 = n6118 ^ n6117 ;
  assign n6121 = n6120 ^ n6119 ;
  assign n6002 = n5835 ^ n5812 ;
  assign n6000 = ~n4435 & ~n5154 ;
  assign n5998 = ~n1972 & n20603 ;
  assign n5995 = ~n1819 & ~n4434 ;
  assign n5994 = ~n1541 & n4600 ;
  assign n5996 = n5995 ^ n5994 ;
  assign n5997 = n5996 ^ x26 ;
  assign n5999 = n5998 ^ n5997 ;
  assign n6001 = n6000 ^ n5999 ;
  assign n6003 = n6002 ^ n6001 ;
  assign n6022 = n5690 ^ n5636 ;
  assign n6015 = x31 ^ x30 ;
  assign n6018 = ~n2552 & n6015 ;
  assign n6007 = n3447 ^ n3329 ;
  assign n6008 = n6007 ^ n2467 ;
  assign n6009 = n6008 & n22005 ;
  assign n6006 = ~n2589 & n22543 ;
  assign n6010 = n6009 ^ n6006 ;
  assign n6005 = ~x31 & ~n2467 ;
  assign n6011 = n6010 ^ n6005 ;
  assign n6012 = n6011 ^ n6010 ;
  assign n6019 = n6018 ^ n6012 ;
  assign n6020 = ~n3518 & n6019 ;
  assign n6021 = n6020 ^ n6011 ;
  assign n6023 = n6022 ^ n6021 ;
  assign n4018 = n680 ^ n459 ;
  assign n4267 = n4018 ^ n1324 ;
  assign n3867 = n1209 ^ n296 ;
  assign n4266 = n3867 ^ n1021 ;
  assign n4268 = n4267 ^ n4266 ;
  assign n4263 = n1998 ^ n506 ;
  assign n4264 = n4263 ^ n956 ;
  assign n4262 = n1401 ^ n725 ;
  assign n4265 = n4264 ^ n4262 ;
  assign n4269 = n4268 ^ n4265 ;
  assign n4270 = n4269 ^ n2280 ;
  assign n4259 = n2891 ^ n976 ;
  assign n4257 = n1239 ^ n911 ;
  assign n4256 = n1404 ^ n189 ;
  assign n4258 = n4257 ^ n4256 ;
  assign n4260 = n4259 ^ n4258 ;
  assign n4254 = n1581 ^ n197 ;
  assign n4252 = n825 ^ n584 ;
  assign n4253 = n4252 ^ n2058 ;
  assign n4255 = n4254 ^ n4253 ;
  assign n4261 = n4260 ^ n4255 ;
  assign n4271 = n4270 ^ n4261 ;
  assign n6045 = n2303 ^ n2153 ;
  assign n6046 = n6045 ^ n1089 ;
  assign n4242 = n770 ^ n416 ;
  assign n6041 = n4242 ^ n317 ;
  assign n6042 = n6041 ^ n1008 ;
  assign n6043 = n6042 ^ n398 ;
  assign n6040 = n735 ^ n377 ;
  assign n6044 = n6043 ^ n6040 ;
  assign n6047 = n6046 ^ n6044 ;
  assign n6037 = n5669 ^ n717 ;
  assign n6038 = n6037 ^ n1506 ;
  assign n6035 = n2053 ^ n898 ;
  assign n6036 = n6035 ^ n1142 ;
  assign n6039 = n6038 ^ n6036 ;
  assign n6048 = n6047 ^ n6039 ;
  assign n6049 = n6048 ^ n1613 ;
  assign n6031 = n5671 ^ n1221 ;
  assign n4197 = n895 ^ n125 ;
  assign n6030 = n4197 ^ n1565 ;
  assign n6032 = n6031 ^ n6030 ;
  assign n6027 = n1052 ^ n510 ;
  assign n6028 = n6027 ^ n431 ;
  assign n6025 = n1185 ^ n380 ;
  assign n6026 = n6025 ^ n969 ;
  assign n6029 = n6028 ^ n6026 ;
  assign n6033 = n6032 ^ n6029 ;
  assign n6024 = n5666 ^ n5616 ;
  assign n6034 = n6033 ^ n6024 ;
  assign n6050 = n6049 ^ n6034 ;
  assign n6051 = ~n4271 & ~n6050 ;
  assign n6052 = n6051 ^ n5635 ;
  assign n6053 = x5 ^ x2 ;
  assign n4807 = n1786 ^ n149 ;
  assign n4808 = n4807 ^ n677 ;
  assign n4805 = n2236 ^ n1689 ;
  assign n4806 = n4805 ^ n1020 ;
  assign n4809 = n4808 ^ n4806 ;
  assign n3647 = n905 ^ n527 ;
  assign n4803 = n3647 ^ n530 ;
  assign n4804 = n4803 ^ n3645 ;
  assign n4810 = n4809 ^ n4804 ;
  assign n4811 = n4810 ^ n3282 ;
  assign n4798 = n1355 ^ n1036 ;
  assign n4799 = n4798 ^ n453 ;
  assign n4796 = n2277 ^ n813 ;
  assign n4795 = n327 ^ n318 ;
  assign n4797 = n4796 ^ n4795 ;
  assign n4800 = n4799 ^ n4797 ;
  assign n4793 = n1136 ^ n1085 ;
  assign n4792 = n1454 ^ n158 ;
  assign n4794 = n4793 ^ n4792 ;
  assign n4801 = n4800 ^ n4794 ;
  assign n4802 = n4801 ^ n728 ;
  assign n4812 = n4811 ^ n4802 ;
  assign n6066 = n1675 ^ n434 ;
  assign n6065 = n596 ^ n339 ;
  assign n6067 = n6066 ^ n6065 ;
  assign n6062 = n602 ^ n458 ;
  assign n3870 = n847 ^ n634 ;
  assign n6063 = n6062 ^ n3870 ;
  assign n3909 = n320 ^ n197 ;
  assign n6061 = n3909 ^ n216 ;
  assign n6064 = n6063 ^ n6061 ;
  assign n6068 = n6067 ^ n6064 ;
  assign n6060 = n3358 ^ n932 ;
  assign n6069 = n6068 ^ n6060 ;
  assign n6056 = n2561 ^ n489 ;
  assign n6057 = n6056 ^ n3135 ;
  assign n6055 = n1143 ^ n743 ;
  assign n6058 = n6057 ^ n6055 ;
  assign n6059 = n6058 ^ n908 ;
  assign n6070 = n6069 ^ n6059 ;
  assign n6054 = n986 ^ n761 ;
  assign n6071 = n6070 ^ n6054 ;
  assign n3722 = n1240 ^ n124 ;
  assign n3723 = n3722 ^ n825 ;
  assign n3719 = n655 ^ n567 ;
  assign n3720 = n3719 ^ n543 ;
  assign n3721 = n3720 ^ n2025 ;
  assign n3724 = n3723 ^ n3721 ;
  assign n3716 = n398 ^ n178 ;
  assign n3717 = n3716 ^ n1300 ;
  assign n3714 = n3713 ^ n495 ;
  assign n3715 = n3714 ^ n1503 ;
  assign n3718 = n3717 ^ n3715 ;
  assign n3725 = n3724 ^ n3718 ;
  assign n3711 = n2562 ^ n385 ;
  assign n3710 = n1680 ^ n829 ;
  assign n3712 = n3711 ^ n3710 ;
  assign n3726 = n3725 ^ n3712 ;
  assign n3705 = n1077 ^ n526 ;
  assign n3706 = n3705 ^ n490 ;
  assign n3707 = n3706 ^ n382 ;
  assign n3704 = n3317 ^ n592 ;
  assign n3708 = n3707 ^ n3704 ;
  assign n3701 = n598 ^ n232 ;
  assign n3702 = n3701 ^ n1568 ;
  assign n3703 = n3702 ^ n1968 ;
  assign n3709 = n3708 ^ n3703 ;
  assign n3727 = n3726 ^ n3709 ;
  assign n6072 = n6071 ^ n3727 ;
  assign n6073 = ~n4812 & ~n6072 ;
  assign n6074 = n6073 ^ x5 ;
  assign n6075 = n6053 & ~n6074 ;
  assign n6076 = n6075 ^ x2 ;
  assign n6077 = n6076 ^ n5635 ;
  assign n6089 = ~n2712 & n22543 ;
  assign n3849 = n3805 ^ n52 ;
  assign n3850 = n3849 ^ n3799 ;
  assign n6088 = ~n2657 & ~n3850 ;
  assign n6090 = n6089 ^ n6088 ;
  assign n6078 = n3445 ^ n3327 ;
  assign n6085 = x31 & ~n6078 ;
  assign n6086 = n6085 ^ n2589 ;
  assign n6087 = n3518 & ~n6086 ;
  assign n6091 = n6090 ^ n6087 ;
  assign n6092 = n6091 ^ n6076 ;
  assign n6093 = ~n6077 & n6092 ;
  assign n6094 = ~n6052 & n6093 ;
  assign n6095 = n6094 ^ n5635 ;
  assign n6096 = n6095 ^ n6021 ;
  assign n6097 = ~n6023 & n6096 ;
  assign n6098 = n6097 ^ n6021 ;
  assign n6110 = n6098 ^ n6002 ;
  assign n6004 = n5716 ^ n5694 ;
  assign n6099 = n6098 ^ n6004 ;
  assign n6103 = ~n2095 & n4369 ;
  assign n6102 = ~n2288 & n3837 ;
  assign n6104 = n6103 ^ n6102 ;
  assign n6105 = n6104 ^ x29 ;
  assign n6101 = n3983 & n5760 ;
  assign n6106 = n6105 ^ n6101 ;
  assign n6100 = ~n2199 & n3985 ;
  assign n6107 = n6106 ^ n6100 ;
  assign n6108 = n6107 ^ n6098 ;
  assign n6109 = ~n6099 & n6108 ;
  assign n6111 = n6110 ^ n6109 ;
  assign n6112 = n6003 & n6111 ;
  assign n6113 = n6112 ^ n6002 ;
  assign n6122 = n6121 ^ n6113 ;
  assign n6123 = n5837 ^ n5811 ;
  assign n6124 = n6123 ^ n6121 ;
  assign n6125 = n6122 & n6124 ;
  assign n6126 = n6125 ^ n6121 ;
  assign n6127 = n6126 ^ n5990 ;
  assign n6128 = n5993 & n6127 ;
  assign n5991 = n5990 ^ n5981 ;
  assign n6129 = n6128 ^ n5991 ;
  assign n6130 = ~n5982 & n6129 ;
  assign n6131 = n6130 ^ n5981 ;
  assign n6132 = n6131 ^ x20 ;
  assign n5972 = ~n856 & n13433 ;
  assign n6133 = n6132 ^ n5972 ;
  assign n5971 = ~n540 & n5220 ;
  assign n6134 = n6133 ^ n5971 ;
  assign n5970 = ~n698 & n5426 ;
  assign n6135 = n6134 ^ n5970 ;
  assign n3955 = n3506 ^ n3498 ;
  assign n3968 = n3955 ^ n540 ;
  assign n5969 = n3968 & n5221 ;
  assign n6136 = n6135 ^ n5969 ;
  assign n4475 = n3483 ^ n1345 ;
  assign n5927 = ~n4435 & n4475 ;
  assign n5924 = ~n1345 & ~n4434 ;
  assign n5922 = ~n1450 & n4600 ;
  assign n5876 = ~n4790 & n5768 ;
  assign n5877 = ~n5746 & n5758 ;
  assign n5878 = ~n5774 & n5877 ;
  assign n5879 = n5876 & n5878 ;
  assign n5880 = n5879 ^ n4790 ;
  assign n5881 = n5774 ^ n5769 ;
  assign n5882 = ~n5770 & ~n5881 ;
  assign n5883 = n5882 ^ n5769 ;
  assign n5884 = ~n5880 & ~n5883 ;
  assign n5885 = n5884 ^ n5880 ;
  assign n5888 = n5885 ^ n5758 ;
  assign n5889 = n5888 ^ n5885 ;
  assign n5892 = n5884 & n5889 ;
  assign n5893 = n5768 & n5892 ;
  assign n5894 = n5893 ^ n5768 ;
  assign n5886 = n5885 ^ n5768 ;
  assign n5895 = n5894 ^ n5886 ;
  assign n5896 = n5390 & ~n5895 ;
  assign n5897 = n5896 ^ n5880 ;
  assign n5898 = n4790 & n5390 ;
  assign n5899 = n5898 ^ n5758 ;
  assign n5900 = n5899 ^ n5898 ;
  assign n5901 = n5898 ^ n5768 ;
  assign n5902 = n5901 ^ n5898 ;
  assign n5903 = ~n5900 & ~n5902 ;
  assign n5904 = n5903 ^ n5898 ;
  assign n5912 = n5902 ^ n5900 ;
  assign n5913 = n5912 ^ n5898 ;
  assign n5906 = n5898 ^ n5774 ;
  assign n5905 = n5898 ^ n5746 ;
  assign n5907 = n5906 ^ n5905 ;
  assign n5908 = n5905 ^ n5899 ;
  assign n5909 = n5908 ^ n5901 ;
  assign n5910 = n5909 ^ n5898 ;
  assign n5911 = ~n5907 & n5910 ;
  assign n5914 = n5913 ^ n5911 ;
  assign n5915 = n5904 & n5914 ;
  assign n5916 = n5915 ^ n5898 ;
  assign n5919 = n5897 & ~n5916 ;
  assign n5874 = ~n1541 & n3837 ;
  assign n5872 = ~n1819 & n3985 ;
  assign n5867 = n5362 ^ n4790 ;
  assign n5868 = ~n5390 & ~n5867 ;
  assign n4846 = n795 ^ n659 ;
  assign n4845 = n802 ^ n506 ;
  assign n4847 = n4846 ^ n4845 ;
  assign n4843 = n1549 ^ n377 ;
  assign n4844 = n4843 ^ n2035 ;
  assign n4848 = n4847 ^ n4844 ;
  assign n4840 = n1576 ^ n1321 ;
  assign n4838 = n730 ^ n493 ;
  assign n4839 = n4838 ^ n3085 ;
  assign n4841 = n4840 ^ n4839 ;
  assign n4295 = n1472 ^ n908 ;
  assign n4842 = n4841 ^ n4295 ;
  assign n4849 = n4848 ^ n4842 ;
  assign n4850 = n4849 ^ n4837 ;
  assign n4831 = n2920 ^ n682 ;
  assign n4154 = n956 ^ n322 ;
  assign n4830 = n4154 ^ n918 ;
  assign n4832 = n4831 ^ n4830 ;
  assign n4833 = n4832 ^ n1835 ;
  assign n4827 = n743 ^ n346 ;
  assign n4828 = n4827 ^ n1495 ;
  assign n4829 = n4828 ^ n2271 ;
  assign n4834 = n4833 ^ n4829 ;
  assign n4851 = n4850 ^ n4834 ;
  assign n4822 = n1408 ^ n145 ;
  assign n4823 = n4822 ^ n362 ;
  assign n4820 = n2840 ^ n269 ;
  assign n4821 = n4820 ^ n465 ;
  assign n4824 = n4823 ^ n4821 ;
  assign n4817 = n4816 ^ n1095 ;
  assign n4815 = n4814 ^ n241 ;
  assign n4818 = n4817 ^ n4815 ;
  assign n4819 = n4818 ^ n1676 ;
  assign n4825 = n4824 ^ n4819 ;
  assign n4813 = n4534 ^ n2882 ;
  assign n4826 = n4825 ^ n4813 ;
  assign n4852 = n4851 ^ n4826 ;
  assign n4853 = ~n4812 & ~n4852 ;
  assign n5292 = n4853 ^ x14 ;
  assign n4878 = x31 & ~n1897 ;
  assign n5281 = ~n4878 & ~n5280 ;
  assign n5279 = n2095 & n22543 ;
  assign n5282 = n5281 ^ n5279 ;
  assign n5287 = n5286 ^ n1972 ;
  assign n5288 = n3518 & n5287 ;
  assign n5289 = ~n5282 & n5288 ;
  assign n5276 = ~n61 & n1973 ;
  assign n5277 = n5276 ^ n1972 ;
  assign n5278 = ~n3800 & ~n5277 ;
  assign n5283 = n5282 ^ n5278 ;
  assign n5290 = n5289 ^ n5283 ;
  assign n5866 = n5292 ^ n5290 ;
  assign n5869 = n5868 ^ n5866 ;
  assign n5870 = n5869 ^ x29 ;
  assign n5863 = ~n4985 & n5065 ;
  assign n5864 = n5863 ^ n1670 ;
  assign n5865 = n3833 & ~n5864 ;
  assign n5871 = n5870 ^ n5865 ;
  assign n5873 = n5872 ^ n5871 ;
  assign n5875 = n5874 ^ n5873 ;
  assign n5920 = n5919 ^ n5875 ;
  assign n5921 = n5920 ^ x26 ;
  assign n5923 = n5922 ^ n5921 ;
  assign n5925 = n5924 ^ n5923 ;
  assign n5859 = ~n1751 & n20603 ;
  assign n5926 = n5925 ^ n5859 ;
  assign n5928 = n5927 ^ n5926 ;
  assign n5856 = n5783 ^ n5456 ;
  assign n5857 = ~n5464 & ~n5856 ;
  assign n5858 = n5857 ^ n5783 ;
  assign n5929 = n5928 ^ n5858 ;
  assign n5854 = ~n990 & n4651 ;
  assign n5852 = ~n1119 & n4655 ;
  assign n5850 = ~n40 & ~n1248 ;
  assign n4334 = n1248 & n4333 ;
  assign n4335 = n4334 ^ n4332 ;
  assign n4336 = n4335 ^ n1119 ;
  assign n5848 = ~n4336 & n4656 ;
  assign n5785 = n5784 ^ n5447 ;
  assign n5845 = ~n5785 & ~n5844 ;
  assign n5846 = n5845 ^ n5784 ;
  assign n5847 = n5846 ^ x23 ;
  assign n5849 = n5848 ^ n5847 ;
  assign n5851 = n5850 ^ n5849 ;
  assign n5853 = n5852 ^ n5851 ;
  assign n5855 = n5854 ^ n5853 ;
  assign n5968 = n5929 ^ n5855 ;
  assign n6380 = n6131 ^ n5968 ;
  assign n6381 = ~n6136 & n6380 ;
  assign n6382 = n6381 ^ n5968 ;
  assign n6383 = n6382 ^ x17 ;
  assign n6142 = x16 ^ x15 ;
  assign n6143 = ~n6141 & n6142 ;
  assign n6379 = ~n368 & n6143 ;
  assign n6384 = n6383 ^ n6379 ;
  assign n6154 = n6143 ^ n6141 ;
  assign n6139 = x14 & x15 ;
  assign n6153 = x16 & n6139 ;
  assign n20432 = n6153 ^ x17 ;
  assign n6155 = n6154 ^ n6153 ;
  assign n20433 = n20432 ^ n6155 ;
  assign n20436 = ~n6154 & n20433 ;
  assign n20437 = n20436 ^ n6153 ;
  assign n6378 = ~n3505 & n20437 ;
  assign n6385 = n6384 ^ n6378 ;
  assign n6387 = n6386 ^ n6385 ;
  assign n5961 = n5920 ^ n5858 ;
  assign n5962 = n5928 & ~n5961 ;
  assign n5963 = n5962 ^ n5920 ;
  assign n5959 = ~n856 & n4655 ;
  assign n5956 = ~n40 & ~n1119 ;
  assign n4359 = n3493 ^ n856 ;
  assign n5954 = ~n4359 & n4656 ;
  assign n5950 = n4307 & ~n4435 ;
  assign n5947 = ~n990 & ~n4434 ;
  assign n5945 = ~n1345 & n4600 ;
  assign n5405 = ~n1819 & n3837 ;
  assign n5403 = ~n1751 & n4369 ;
  assign n5400 = n3983 & n4690 ;
  assign n5399 = ~n1670 & n3985 ;
  assign n5401 = n5400 ^ n5399 ;
  assign n5402 = n5401 ^ x29 ;
  assign n5404 = n5403 ^ n5402 ;
  assign n5406 = n5405 ^ n5404 ;
  assign n5291 = n5290 ^ n4790 ;
  assign n5293 = n5292 ^ n5291 ;
  assign n5363 = n5362 ^ n5290 ;
  assign n5364 = n5363 ^ n5292 ;
  assign n5393 = n5364 & ~n5390 ;
  assign n5394 = n5393 ^ n5292 ;
  assign n5395 = n5293 & n5394 ;
  assign n5396 = n5395 ^ n5290 ;
  assign n3747 = n3275 ^ n2886 ;
  assign n3746 = n1498 ^ n803 ;
  assign n3748 = n3747 ^ n3746 ;
  assign n3743 = n3742 ^ n1614 ;
  assign n3741 = n3740 ^ n3571 ;
  assign n3744 = n3743 ^ n3741 ;
  assign n3735 = n655 ^ n137 ;
  assign n3736 = n3735 ^ n468 ;
  assign n3737 = n3736 ^ n766 ;
  assign n3738 = n3737 ^ n1422 ;
  assign n3734 = n2678 ^ n1300 ;
  assign n3739 = n3738 ^ n3734 ;
  assign n3745 = n3744 ^ n3739 ;
  assign n3749 = n3748 ^ n3745 ;
  assign n3750 = n3749 ^ n2816 ;
  assign n4905 = n3750 ^ n873 ;
  assign n4934 = n4503 ^ n2930 ;
  assign n4931 = n4930 ^ n1108 ;
  assign n4932 = n4931 ^ n2616 ;
  assign n4929 = n3112 ^ n377 ;
  assign n4933 = n4932 ^ n4929 ;
  assign n4935 = n4934 ^ n4933 ;
  assign n4925 = n3013 ^ n1405 ;
  assign n4923 = n2378 ^ n831 ;
  assign n4924 = n4923 ^ n820 ;
  assign n4926 = n4925 ^ n4924 ;
  assign n4922 = n2519 ^ n347 ;
  assign n4927 = n4926 ^ n4922 ;
  assign n4928 = n4927 ^ n3059 ;
  assign n4936 = n4935 ^ n4928 ;
  assign n4917 = n1040 ^ n636 ;
  assign n4916 = n868 ^ n830 ;
  assign n4918 = n4917 ^ n4916 ;
  assign n4919 = n4918 ^ n2703 ;
  assign n4912 = n653 ^ n562 ;
  assign n4913 = n4912 ^ n480 ;
  assign n4911 = n504 ^ n478 ;
  assign n4914 = n4913 ^ n4911 ;
  assign n4909 = n4908 ^ n734 ;
  assign n4906 = n772 ^ n556 ;
  assign n4907 = n4906 ^ n1066 ;
  assign n4910 = n4909 ^ n4907 ;
  assign n4915 = n4914 ^ n4910 ;
  assign n4920 = n4919 ^ n4915 ;
  assign n4921 = n4920 ^ n4726 ;
  assign n4937 = n4936 ^ n4921 ;
  assign n4938 = ~n4905 & ~n4937 ;
  assign n4791 = n4790 ^ x14 ;
  assign n4854 = n4853 ^ n4790 ;
  assign n4855 = n4791 & ~n4854 ;
  assign n4856 = n4855 ^ x14 ;
  assign n4939 = n4938 ^ n4856 ;
  assign n4899 = x31 & ~n1972 ;
  assign n4892 = n4891 ^ n1541 ;
  assign n4893 = x31 & ~n4892 ;
  assign n4882 = ~n1541 & ~n22005 ;
  assign n4894 = n4893 ^ n4882 ;
  assign n4900 = n4899 ^ n4894 ;
  assign n4901 = ~n3518 & n4900 ;
  assign n4902 = n4901 ^ n4894 ;
  assign n4879 = n4878 ^ n1972 ;
  assign n4880 = ~n61 & ~n4879 ;
  assign n4903 = n4902 ^ n4880 ;
  assign n5271 = n4939 ^ n4903 ;
  assign n5397 = n5396 ^ n5271 ;
  assign n5943 = n5406 ^ n5397 ;
  assign n5944 = n5943 ^ x26 ;
  assign n5946 = n5945 ^ n5944 ;
  assign n5948 = n5947 ^ n5946 ;
  assign n5942 = ~n1450 & n20603 ;
  assign n5949 = n5948 ^ n5942 ;
  assign n5951 = n5950 ^ n5949 ;
  assign n5939 = n5919 ^ n5869 ;
  assign n5940 = ~n5875 & n5939 ;
  assign n5941 = n5940 ^ n5919 ;
  assign n5952 = n5951 ^ n5941 ;
  assign n5953 = n5952 ^ x23 ;
  assign n5955 = n5954 ^ n5953 ;
  assign n5957 = n5956 ^ n5955 ;
  assign n5938 = ~n1248 & n4651 ;
  assign n5958 = n5957 ^ n5938 ;
  assign n5960 = n5959 ^ n5958 ;
  assign n5964 = n5963 ^ n5960 ;
  assign n5930 = n5929 ^ n5846 ;
  assign n5931 = n5855 & n5930 ;
  assign n5932 = n5931 ^ n5929 ;
  assign n5933 = n5932 ^ x20 ;
  assign n5436 = ~n408 & n5220 ;
  assign n5934 = n5933 ^ n5436 ;
  assign n5435 = ~n540 & n5426 ;
  assign n5935 = n5934 ^ n5435 ;
  assign n5434 = ~n698 & n13433 ;
  assign n5936 = n5935 ^ n5434 ;
  assign n3811 = n3507 ^ n3499 ;
  assign n3812 = n3811 ^ n408 ;
  assign n5433 = n3812 & n5221 ;
  assign n5937 = n5936 ^ n5433 ;
  assign n6377 = n5964 ^ n5937 ;
  assign n6388 = n6387 ^ n6377 ;
  assign n6137 = n6136 ^ n5968 ;
  assign n3839 = n3508 ^ n3500 ;
  assign n3840 = n3839 ^ n3505 ;
  assign n6164 = n3840 & n6163 ;
  assign n6161 = ~n540 & n20437 ;
  assign n6150 = ~n408 & n6143 ;
  assign n6149 = ~n3505 & n6148 ;
  assign n6151 = n6150 ^ n6149 ;
  assign n6152 = n6151 ^ x17 ;
  assign n6162 = n6161 ^ n6152 ;
  assign n6165 = n6164 ^ n6162 ;
  assign n6138 = n6129 ^ n5973 ;
  assign n6166 = n6165 ^ n6138 ;
  assign n6174 = ~n4359 & n5221 ;
  assign n6172 = ~n1248 & n13433 ;
  assign n6169 = ~n856 & n5220 ;
  assign n6168 = ~n1119 & n5426 ;
  assign n6170 = n6169 ^ n6168 ;
  assign n6171 = n6170 ^ x20 ;
  assign n6173 = n6172 ^ n6171 ;
  assign n6175 = n6174 ^ n6173 ;
  assign n6167 = n6126 ^ n5993 ;
  assign n6176 = n6175 ^ n6167 ;
  assign n6356 = n6124 ^ n6113 ;
  assign n6368 = n6356 ^ n6175 ;
  assign n6185 = n6111 ^ n6001 ;
  assign n6181 = ~n4495 & n4656 ;
  assign n6180 = ~n1670 & n4651 ;
  assign n6182 = n6181 ^ n6180 ;
  assign n6183 = n6182 ^ x23 ;
  assign n6178 = ~n1450 & n4655 ;
  assign n6177 = ~n40 & ~n1751 ;
  assign n6179 = n6178 ^ n6177 ;
  assign n6184 = n6183 ^ n6179 ;
  assign n6186 = n6185 ^ n6184 ;
  assign n6194 = ~n4435 & ~n4892 ;
  assign n6192 = ~n1541 & ~n4434 ;
  assign n6189 = ~n1897 & n20603 ;
  assign n6188 = ~n1972 & n4600 ;
  assign n6190 = n6189 ^ n6188 ;
  assign n6191 = n6190 ^ x26 ;
  assign n6193 = n6192 ^ n6191 ;
  assign n6195 = n6194 ^ n6193 ;
  assign n6187 = n6107 ^ n6099 ;
  assign n6196 = n6195 ^ n6187 ;
  assign n6201 = ~n2199 & n4369 ;
  assign n6200 = ~n2371 & n3837 ;
  assign n6202 = n6201 ^ n6200 ;
  assign n6203 = n6202 ^ x29 ;
  assign n6199 = n3983 & n5480 ;
  assign n6204 = n6203 ^ n6199 ;
  assign n6198 = ~n2288 & n3985 ;
  assign n6205 = n6204 ^ n6198 ;
  assign n6197 = n6095 ^ n6023 ;
  assign n6206 = n6205 ^ n6197 ;
  assign n6216 = n6093 ^ n6051 ;
  assign n6211 = n3446 ^ n3328 ;
  assign n6212 = n6211 ^ n2552 ;
  assign n6213 = n6212 & n22005 ;
  assign n6210 = ~n2657 & n22543 ;
  assign n6214 = n6213 ^ n6210 ;
  assign n6208 = ~n2552 & n3807 ;
  assign n6207 = ~n2589 & ~n3850 ;
  assign n6209 = n6208 ^ n6207 ;
  assign n6215 = n6214 ^ n6209 ;
  assign n6217 = n6216 ^ n6215 ;
  assign n6226 = n6091 ^ n6077 ;
  assign n6343 = n6226 ^ n6215 ;
  assign n6221 = ~n2552 & n3837 ;
  assign n6220 = ~n2371 & n4369 ;
  assign n6222 = n6221 ^ n6220 ;
  assign n6223 = n6222 ^ x29 ;
  assign n6219 = n3983 & n5696 ;
  assign n6224 = n6223 ^ n6219 ;
  assign n6218 = ~n2467 & n3985 ;
  assign n6225 = n6224 ^ n6218 ;
  assign n6227 = n6226 ^ n6225 ;
  assign n6243 = n6073 ^ n6053 ;
  assign n6239 = ~n3324 & n22543 ;
  assign n6238 = ~n2712 & ~n3850 ;
  assign n6240 = n6239 ^ n6238 ;
  assign n6228 = n3444 ^ n3326 ;
  assign n6235 = x31 & ~n6228 ;
  assign n6236 = n6235 ^ n2657 ;
  assign n6237 = n3518 & ~n6236 ;
  assign n6241 = n6240 ^ n6237 ;
  assign n6244 = n6243 ^ n6241 ;
  assign n6283 = n604 ^ n470 ;
  assign n6284 = n6283 ^ n501 ;
  assign n6281 = n556 ^ n237 ;
  assign n6282 = n6281 ^ n873 ;
  assign n6285 = n6284 ^ n6282 ;
  assign n6278 = n5732 ^ n493 ;
  assign n6279 = n6278 ^ n387 ;
  assign n6277 = n2561 ^ n637 ;
  assign n6280 = n6279 ^ n6277 ;
  assign n6286 = n6285 ^ n6280 ;
  assign n3686 = n3685 ^ n1036 ;
  assign n6275 = n3686 ^ n3413 ;
  assign n3646 = n3645 ^ n1889 ;
  assign n6276 = n6275 ^ n3646 ;
  assign n6287 = n6286 ^ n6276 ;
  assign n3615 = n2319 ^ n145 ;
  assign n3616 = n3615 ^ n788 ;
  assign n3613 = n682 ^ n188 ;
  assign n3614 = n3613 ^ n444 ;
  assign n3617 = n3616 ^ n3614 ;
  assign n3618 = n3617 ^ n3421 ;
  assign n6288 = n6287 ^ n3618 ;
  assign n6289 = n6288 ^ n3354 ;
  assign n6270 = n1191 ^ n784 ;
  assign n6271 = n6270 ^ n829 ;
  assign n6269 = n1324 ^ n1128 ;
  assign n6272 = n6271 ^ n6269 ;
  assign n6267 = n2639 ^ n1236 ;
  assign n6268 = n6267 ^ n948 ;
  assign n6273 = n6272 ^ n6268 ;
  assign n6264 = n5724 ^ n3068 ;
  assign n6265 = n6264 ^ n2428 ;
  assign n6266 = n6265 ^ n5601 ;
  assign n6274 = n6273 ^ n6266 ;
  assign n6290 = n6289 ^ n6274 ;
  assign n6291 = ~n2094 & ~n6290 ;
  assign n6256 = n1581 ^ n948 ;
  assign n6257 = n6256 ^ n339 ;
  assign n6255 = n476 ^ n262 ;
  assign n6258 = n6257 ^ n6255 ;
  assign n3548 = n659 ^ n504 ;
  assign n6253 = n3740 ^ n3548 ;
  assign n6252 = n1362 ^ n1037 ;
  assign n6254 = n6253 ^ n6252 ;
  assign n6259 = n6258 ^ n6254 ;
  assign n3695 = n1360 ^ n1204 ;
  assign n3696 = n3695 ^ n1020 ;
  assign n3693 = n1374 ^ n157 ;
  assign n3694 = n3693 ^ n547 ;
  assign n3697 = n3696 ^ n3694 ;
  assign n3690 = n873 ^ n94 ;
  assign n3691 = n3690 ^ n2408 ;
  assign n3692 = n3691 ^ n2331 ;
  assign n3698 = n3697 ^ n3692 ;
  assign n6260 = n6259 ^ n3698 ;
  assign n6248 = n5669 ^ n400 ;
  assign n6249 = n6248 ^ n2150 ;
  assign n6250 = n6249 ^ n4737 ;
  assign n6245 = n4098 ^ n1709 ;
  assign n4182 = n556 ^ n188 ;
  assign n6246 = n6245 ^ n4182 ;
  assign n6247 = n6246 ^ n892 ;
  assign n6251 = n6250 ^ n6247 ;
  assign n6261 = n6260 ^ n6251 ;
  assign n6262 = n6261 ^ n1342 ;
  assign n6263 = ~n3159 & ~n6262 ;
  assign n6292 = n6291 ^ n6263 ;
  assign n6293 = n6291 ^ x2 ;
  assign n6301 = n3441 ^ n3251 ;
  assign n6302 = n6301 ^ n2748 ;
  assign n6303 = ~n6302 & n22005 ;
  assign n6300 = ~n2839 & n5465 ;
  assign n6304 = n6303 ^ n6300 ;
  assign n6305 = n6304 ^ n2935 ;
  assign n6297 = ~n61 & ~n2839 ;
  assign n6298 = n6297 ^ n2748 ;
  assign n6299 = ~n3800 & ~n6298 ;
  assign n6306 = n6305 ^ n6299 ;
  assign n6294 = ~n61 & ~n2748 ;
  assign n6295 = n6294 ^ n2935 ;
  assign n6296 = ~n6295 & ~n22543 ;
  assign n6307 = n6306 ^ n6296 ;
  assign n6308 = n6307 ^ n6291 ;
  assign n6309 = ~n6293 & ~n6308 ;
  assign n6310 = ~n6292 & n6309 ;
  assign n6311 = n2961 ^ n1007 ;
  assign n6328 = n1440 ^ n188 ;
  assign n6329 = n6328 ^ n751 ;
  assign n6330 = n6329 ^ n541 ;
  assign n6325 = n596 ^ n265 ;
  assign n6326 = n6325 ^ n1095 ;
  assign n6327 = n6326 ^ n2506 ;
  assign n6331 = n6330 ^ n6327 ;
  assign n6332 = n6331 ^ n1949 ;
  assign n6321 = n1324 ^ n682 ;
  assign n3756 = n566 ^ n495 ;
  assign n3757 = n3756 ^ n1014 ;
  assign n6320 = n3757 ^ n489 ;
  assign n6322 = n6321 ^ n6320 ;
  assign n6319 = n1183 ^ n1073 ;
  assign n6323 = n6322 ^ n6319 ;
  assign n6316 = n1709 ^ n548 ;
  assign n6317 = n6316 ^ n5528 ;
  assign n6314 = n1066 ^ n526 ;
  assign n6312 = n1128 ^ n261 ;
  assign n6313 = n6312 ^ n598 ;
  assign n6315 = n6314 ^ n6313 ;
  assign n6318 = n6317 ^ n6315 ;
  assign n6324 = n6323 ^ n6318 ;
  assign n6333 = n6332 ^ n6324 ;
  assign n6334 = n6333 ^ n3322 ;
  assign n6335 = ~n6311 & ~n6334 ;
  assign n6336 = n6335 ^ n6263 ;
  assign n6337 = n6310 & ~n6336 ;
  assign n6338 = n6337 ^ x2 ;
  assign n6339 = n6338 ^ n6241 ;
  assign n6340 = ~n6244 & n6339 ;
  assign n6242 = n6241 ^ n6225 ;
  assign n6341 = n6340 ^ n6242 ;
  assign n6342 = ~n6227 & ~n6341 ;
  assign n6344 = n6343 ^ n6342 ;
  assign n6345 = ~n6217 & n6344 ;
  assign n6346 = n6345 ^ n6216 ;
  assign n6347 = n6346 ^ n6205 ;
  assign n6348 = ~n6206 & ~n6347 ;
  assign n6349 = n6348 ^ n6205 ;
  assign n6350 = n6349 ^ n6195 ;
  assign n6351 = ~n6196 & n6350 ;
  assign n6352 = n6351 ^ n6195 ;
  assign n6353 = n6352 ^ n6184 ;
  assign n6354 = n6186 & n6353 ;
  assign n6355 = n6354 ^ n6184 ;
  assign n6357 = n6356 ^ n6355 ;
  assign n6365 = ~n1751 & n4651 ;
  assign n6361 = n6356 ^ x23 ;
  assign n6360 = n4475 & n4656 ;
  assign n6362 = n6361 ^ n6360 ;
  assign n6359 = ~n40 & ~n1450 ;
  assign n6363 = n6362 ^ n6359 ;
  assign n6358 = ~n1345 & n4655 ;
  assign n6364 = n6363 ^ n6358 ;
  assign n6366 = n6365 ^ n6364 ;
  assign n6367 = n6357 & n6366 ;
  assign n6369 = n6368 ^ n6367 ;
  assign n6370 = n6176 & n6369 ;
  assign n6371 = n6370 ^ n6175 ;
  assign n6372 = n6371 ^ n6165 ;
  assign n6373 = ~n6166 & n6372 ;
  assign n6374 = n6373 ^ n6165 ;
  assign n6375 = n6374 ^ n6137 ;
  assign n6376 = ~n6137 & ~n6375 ;
  assign n6389 = n6388 ^ n6376 ;
  assign n6410 = n6371 ^ n6166 ;
  assign n6391 = x12 ^ x11 ;
  assign n6390 = ~x11 & ~x12 ;
  assign n6392 = n6391 ^ n6390 ;
  assign n6397 = ~x13 & ~n368 ;
  assign n6398 = n6397 ^ x14 ;
  assign n6399 = ~n3509 & ~n6398 ;
  assign n6400 = n6399 ^ x14 ;
  assign n6401 = n6392 & ~n6400 ;
  assign n6402 = n6390 ^ x14 ;
  assign n6403 = n6390 ^ x13 ;
  assign n6404 = ~n6402 & n6403 ;
  assign n6407 = ~n368 & n6404 ;
  assign n6408 = n6407 ^ x14 ;
  assign n6409 = ~n6401 & n6408 ;
  assign n6411 = n6410 ^ n6409 ;
  assign n6491 = ~n698 & n20437 ;
  assign n6490 = ~n540 & n6143 ;
  assign n6492 = n6491 ^ n6490 ;
  assign n6145 = x17 & ~n6141 ;
  assign n6493 = n6492 ^ n6145 ;
  assign n6496 = n408 ^ x16 ;
  assign n6494 = n6147 ^ x16 ;
  assign n6495 = n3811 & ~n6494 ;
  assign n6497 = n6496 ^ n6495 ;
  assign n6498 = n6497 ^ n6492 ;
  assign n6499 = n6498 ^ x17 ;
  assign n6502 = ~n6147 & ~n6496 ;
  assign n6503 = n6502 ^ n408 ;
  assign n6504 = ~n3811 & n6503 ;
  assign n6505 = n6504 ^ n408 ;
  assign n6506 = ~n6499 & n6505 ;
  assign n6507 = n6506 ^ n6497 ;
  assign n6508 = ~n6493 & n6507 ;
  assign n6420 = ~n4336 & n5221 ;
  assign n6417 = ~n1119 & n5220 ;
  assign n6415 = ~n1248 & n5426 ;
  assign n6413 = n6366 ^ n6355 ;
  assign n6414 = n6413 ^ x20 ;
  assign n6416 = n6415 ^ n6414 ;
  assign n6418 = n6417 ^ n6416 ;
  assign n6412 = ~n990 & n13433 ;
  assign n6419 = n6418 ^ n6412 ;
  assign n6421 = n6420 ^ n6419 ;
  assign n4580 = n4333 ^ n1248 ;
  assign n6429 = n4580 & n5221 ;
  assign n6427 = ~n990 & n5426 ;
  assign n6424 = ~n1345 & n13433 ;
  assign n6423 = ~n1248 & n5220 ;
  assign n6425 = n6424 ^ n6423 ;
  assign n6426 = n6425 ^ x20 ;
  assign n6428 = n6427 ^ n6426 ;
  assign n6430 = n6429 ^ n6428 ;
  assign n6422 = n6352 ^ n6186 ;
  assign n6431 = n6430 ^ n6422 ;
  assign n6442 = ~n40 & ~n1670 ;
  assign n6441 = ~n1819 & n4651 ;
  assign n6443 = n6442 ^ n6441 ;
  assign n6434 = n1751 ^ x23 ;
  assign n6435 = n6434 ^ x22 ;
  assign n6436 = n6435 ^ n1751 ;
  assign n6437 = ~n4492 & n6436 ;
  assign n6438 = n6437 ^ n1751 ;
  assign n6439 = n35 & ~n6438 ;
  assign n6440 = n6439 ^ x23 ;
  assign n6444 = n6443 ^ n6440 ;
  assign n6483 = n6444 ^ n6422 ;
  assign n6432 = n6349 ^ n6196 ;
  assign n6445 = n6444 ^ n6432 ;
  assign n5824 = n4884 ^ n1897 ;
  assign n6463 = ~n4435 & n5824 ;
  assign n6461 = ~n1897 & ~n4434 ;
  assign n6458 = ~n2095 & n4600 ;
  assign n6457 = ~n2199 & n20603 ;
  assign n6459 = n6458 ^ n6457 ;
  assign n6460 = n6459 ^ x26 ;
  assign n6462 = n6461 ^ n6460 ;
  assign n6464 = n6463 ^ n6462 ;
  assign n6452 = ~n2467 & n3837 ;
  assign n6451 = ~n2288 & n4369 ;
  assign n6453 = n6452 ^ n6451 ;
  assign n6454 = n6453 ^ x29 ;
  assign n6449 = n5814 ^ n2288 ;
  assign n6450 = n3983 & n6449 ;
  assign n6455 = n6454 ^ n6450 ;
  assign n6448 = ~n2371 & n3985 ;
  assign n6456 = n6455 ^ n6448 ;
  assign n6465 = n6464 ^ n6456 ;
  assign n6466 = n6344 ^ n6216 ;
  assign n6467 = n6466 ^ n6456 ;
  assign n6468 = n6465 & ~n6467 ;
  assign n6469 = n6468 ^ n6464 ;
  assign n6446 = n6346 ^ n6206 ;
  assign n6470 = n6469 ^ n6446 ;
  assign n6478 = ~n4435 & ~n5287 ;
  assign n6474 = n6446 ^ x26 ;
  assign n6473 = ~n1897 & n4600 ;
  assign n6475 = n6474 ^ n6473 ;
  assign n6472 = ~n1972 & ~n4434 ;
  assign n6476 = n6475 ^ n6472 ;
  assign n6471 = ~n2095 & n20603 ;
  assign n6477 = n6476 ^ n6471 ;
  assign n6479 = n6478 ^ n6477 ;
  assign n6480 = n6470 & n6479 ;
  assign n6447 = n6446 ^ n6444 ;
  assign n6481 = n6480 ^ n6447 ;
  assign n6482 = ~n6445 & n6481 ;
  assign n6484 = n6483 ^ n6482 ;
  assign n6485 = n6431 & ~n6484 ;
  assign n6486 = n6485 ^ n6430 ;
  assign n6487 = n6486 ^ n6413 ;
  assign n6488 = n6421 & n6487 ;
  assign n6489 = n6488 ^ n6413 ;
  assign n6509 = n6508 ^ n6489 ;
  assign n6510 = n6369 ^ n6167 ;
  assign n6511 = n6510 ^ n6508 ;
  assign n6512 = ~n6509 & ~n6511 ;
  assign n6513 = n6512 ^ n6508 ;
  assign n6514 = n6513 ^ n6410 ;
  assign n6515 = ~n6411 & n6514 ;
  assign n6516 = n6515 ^ n6410 ;
  assign n6524 = ~n3513 & n6148 ;
  assign n6520 = n6516 ^ x17 ;
  assign n6519 = ~n408 & n20437 ;
  assign n6521 = n6520 ^ n6519 ;
  assign n6518 = ~n3505 & n6143 ;
  assign n6522 = n6521 ^ n6518 ;
  assign n4398 = n3513 ^ n368 ;
  assign n6517 = n4398 & n6141 ;
  assign n6523 = n6522 ^ n6517 ;
  assign n6525 = n6524 ^ n6523 ;
  assign n6526 = ~n6516 & n6525 ;
  assign n7022 = n6513 ^ n6411 ;
  assign n6531 = n6392 ^ x13 ;
  assign n6528 = ~x13 & n6391 ;
  assign n6532 = n6531 ^ n6528 ;
  assign n20347 = n6532 ^ x14 ;
  assign n6534 = x13 & ~n6392 ;
  assign n6535 = n6534 ^ n6532 ;
  assign n6537 = x14 & n6391 ;
  assign n6536 = n6391 ^ x14 ;
  assign n6538 = n6537 ^ n6536 ;
  assign n6541 = ~x12 & ~x13 ;
  assign n6540 = x13 ^ x12 ;
  assign n6542 = n6541 ^ n6540 ;
  assign n6543 = ~n6538 & n6542 ;
  assign n6544 = n6543 ^ n6534 ;
  assign n6539 = n6538 ^ x14 ;
  assign n6545 = n6544 ^ n6539 ;
  assign n6546 = ~n6535 & n6545 ;
  assign n6547 = n20347 ^ n6546 ;
  assign n6548 = ~n3505 & ~n6547 ;
  assign n6529 = n6528 ^ n6403 ;
  assign n6530 = ~n368 & ~n6529 ;
  assign n6549 = n6548 ^ n6530 ;
  assign n6550 = n6549 ^ x14 ;
  assign n6551 = n6550 ^ x13 ;
  assign n6552 = n3515 & n6391 ;
  assign n6553 = n6551 & n6552 ;
  assign n6554 = n6553 ^ n6550 ;
  assign n6527 = n6511 ^ n6489 ;
  assign n6555 = n6554 ^ n6527 ;
  assign n6564 = n3968 & n6163 ;
  assign n6559 = n6486 ^ n6421 ;
  assign n6560 = n6559 ^ x17 ;
  assign n6558 = ~n856 & n20437 ;
  assign n6561 = n6560 ^ n6558 ;
  assign n6557 = ~n540 & n6148 ;
  assign n6562 = n6561 ^ n6557 ;
  assign n6556 = ~n698 & n6143 ;
  assign n6563 = n6562 ^ n6556 ;
  assign n6565 = n6564 ^ n6563 ;
  assign n6576 = ~n3930 & n6163 ;
  assign n6573 = ~n1119 & n20437 ;
  assign n6571 = ~n698 & n6148 ;
  assign n6569 = n6484 ^ n6430 ;
  assign n6570 = n6569 ^ x17 ;
  assign n6572 = n6571 ^ n6570 ;
  assign n6574 = n6573 ^ n6572 ;
  assign n6568 = ~n856 & n6143 ;
  assign n6575 = n6574 ^ n6568 ;
  assign n6577 = n6576 ^ n6575 ;
  assign n6586 = n4307 & n5221 ;
  assign n6583 = ~n990 & n5220 ;
  assign n6581 = ~n1345 & n5426 ;
  assign n6579 = n6481 ^ n6432 ;
  assign n6580 = n6579 ^ x20 ;
  assign n6582 = n6581 ^ n6580 ;
  assign n6584 = n6583 ^ n6582 ;
  assign n6578 = ~n1450 & n13433 ;
  assign n6585 = n6584 ^ n6578 ;
  assign n6587 = n6586 ^ n6585 ;
  assign n6597 = ~n40 & ~n1541 ;
  assign n6594 = ~n1972 & n4651 ;
  assign n6592 = n4656 & ~n5154 ;
  assign n6590 = n6467 ^ n6464 ;
  assign n6591 = n6590 ^ x23 ;
  assign n6593 = n6592 ^ n6591 ;
  assign n6595 = n6594 ^ n6593 ;
  assign n6589 = ~n1819 & n4655 ;
  assign n6596 = n6595 ^ n6589 ;
  assign n6598 = n6597 ^ n6596 ;
  assign n6610 = n6341 ^ n6226 ;
  assign n6606 = ~n2199 & n4600 ;
  assign n6605 = ~n2288 & n20603 ;
  assign n6607 = n6606 ^ n6605 ;
  assign n6608 = n6607 ^ x26 ;
  assign n6602 = n285 & ~n5759 ;
  assign n6603 = n6602 ^ n2095 ;
  assign n6604 = n96 & ~n6603 ;
  assign n6609 = n6608 ^ n6604 ;
  assign n6611 = n6610 ^ n6609 ;
  assign n6616 = ~n2467 & n4369 ;
  assign n6615 = ~n2589 & n3837 ;
  assign n6617 = n6616 ^ n6615 ;
  assign n6618 = n6617 ^ x29 ;
  assign n6614 = n3983 & n6008 ;
  assign n6619 = n6618 ^ n6614 ;
  assign n6613 = ~n2552 & n3985 ;
  assign n6620 = n6619 ^ n6613 ;
  assign n6612 = n6338 ^ n6244 ;
  assign n6621 = n6620 ^ n6612 ;
  assign n6627 = n6307 ^ n6263 ;
  assign n6628 = n6309 & ~n6627 ;
  assign n6629 = n6628 ^ n6335 ;
  assign n6630 = n6629 ^ n6294 ;
  assign n6631 = n6630 ^ n6629 ;
  assign n6632 = n6631 ^ n3324 ;
  assign n6633 = n6632 ^ n6631 ;
  assign n6634 = n6631 ^ n3806 ;
  assign n6635 = n6634 ^ n6631 ;
  assign n6636 = ~n6633 & ~n6635 ;
  assign n6637 = n6636 ^ n6631 ;
  assign n6638 = ~n3849 & n6637 ;
  assign n6639 = n6638 ^ n6630 ;
  assign n6622 = n3443 ^ n3325 ;
  assign n6625 = n3807 & ~n6622 ;
  assign n6623 = n6622 ^ n2712 ;
  assign n6624 = n3518 & n6623 ;
  assign n6626 = n6625 ^ n6624 ;
  assign n6640 = n6639 ^ n6626 ;
  assign n6643 = n3442 ^ n3252 ;
  assign n6644 = n6643 ^ n2748 ;
  assign n6647 = n3807 & n6644 ;
  assign n6645 = n6644 ^ n3324 ;
  assign n6646 = n3518 & ~n6645 ;
  assign n6648 = n6647 ^ n6646 ;
  assign n6649 = n6648 ^ n2748 ;
  assign n6642 = n3801 & ~n6298 ;
  assign n6650 = n6649 ^ n6642 ;
  assign n6641 = n6309 ^ n6263 ;
  assign n6651 = n6650 ^ n6641 ;
  assign n6661 = n6307 ^ n6293 ;
  assign n6655 = ~n3324 & n3837 ;
  assign n6654 = ~n2657 & n4369 ;
  assign n6656 = n6655 ^ n6654 ;
  assign n6657 = n6656 ^ x29 ;
  assign n6229 = n6228 ^ n2657 ;
  assign n6653 = n3983 & n6229 ;
  assign n6658 = n6657 ^ n6653 ;
  assign n6652 = ~n2712 & n3985 ;
  assign n6659 = n6658 ^ n6652 ;
  assign n6662 = n6661 ^ n6659 ;
  assign n6700 = ~n3248 & n22543 ;
  assign n6699 = ~n2935 & ~n3850 ;
  assign n6701 = n6700 ^ n6699 ;
  assign n6697 = n3439 & n3807 ;
  assign n6695 = n3439 ^ n2839 ;
  assign n6696 = n3518 & ~n6695 ;
  assign n6698 = n6697 ^ n6696 ;
  assign n6702 = n6701 ^ n6698 ;
  assign n6672 = n1919 ^ n517 ;
  assign n6673 = n6672 ^ n1554 ;
  assign n6671 = n2567 ^ n1360 ;
  assign n6674 = n6673 ^ n6671 ;
  assign n6668 = n335 ^ n185 ;
  assign n6669 = n6668 ^ n915 ;
  assign n3621 = n1189 ^ n778 ;
  assign n3622 = n3621 ^ n721 ;
  assign n6670 = n6669 ^ n3622 ;
  assign n6675 = n6674 ^ n6670 ;
  assign n6666 = n977 ^ n761 ;
  assign n6667 = n6666 ^ n2384 ;
  assign n6676 = n6675 ^ n6667 ;
  assign n6663 = n2425 ^ n710 ;
  assign n6664 = n6663 ^ n3706 ;
  assign n6665 = n6664 ^ n6256 ;
  assign n6677 = n6676 ^ n6665 ;
  assign n6678 = n6677 ^ n4811 ;
  assign n6687 = n1099 ^ n592 ;
  assign n6688 = n6687 ^ n609 ;
  assign n6686 = n820 ^ n504 ;
  assign n6689 = n6688 ^ n6686 ;
  assign n6684 = n1661 ^ n126 ;
  assign n6682 = n725 ^ n409 ;
  assign n6683 = n6682 ^ n1837 ;
  assign n6685 = n6684 ^ n6683 ;
  assign n6690 = n6689 ^ n6685 ;
  assign n6679 = n4827 ^ n2144 ;
  assign n6680 = n6679 ^ n1793 ;
  assign n6681 = n6680 ^ n4741 ;
  assign n6691 = n6690 ^ n6681 ;
  assign n6692 = n6691 ^ n2549 ;
  assign n6693 = n6692 ^ n4826 ;
  assign n6694 = ~n6678 & ~n6693 ;
  assign n6703 = n6702 ^ n6694 ;
  assign n6743 = ~n3248 & ~n3850 ;
  assign n6742 = ~n2935 & n3807 ;
  assign n6744 = n6743 ^ n6742 ;
  assign n6736 = n3437 ^ n2935 ;
  assign n6739 = n3518 & n6736 ;
  assign n6733 = ~n61 & ~n3022 ;
  assign n6740 = n6739 ^ n6733 ;
  assign n6741 = x31 & n6740 ;
  assign n6745 = n6744 ^ n6741 ;
  assign n6710 = n5732 ^ n508 ;
  assign n6709 = n6325 ^ n4710 ;
  assign n6711 = n6710 ^ n6709 ;
  assign n4968 = n1189 ^ n382 ;
  assign n4969 = n4968 ^ n610 ;
  assign n4970 = n4969 ^ n1008 ;
  assign n4967 = n2993 ^ n457 ;
  assign n4971 = n4970 ^ n4967 ;
  assign n6712 = n6711 ^ n4971 ;
  assign n6706 = n3069 ^ n905 ;
  assign n6705 = n1139 ^ n622 ;
  assign n6707 = n6706 ^ n6705 ;
  assign n6704 = n5638 ^ n3736 ;
  assign n6708 = n6707 ^ n6704 ;
  assign n6713 = n6712 ^ n6708 ;
  assign n6714 = n6713 ^ n1320 ;
  assign n6726 = n795 ^ n118 ;
  assign n6727 = n6726 ^ n180 ;
  assign n6724 = n5573 ^ n2445 ;
  assign n6723 = n3645 ^ n557 ;
  assign n6725 = n6724 ^ n6723 ;
  assign n6728 = n6727 ^ n6725 ;
  assign n6721 = n2603 ^ n1376 ;
  assign n6722 = n6721 ^ n1210 ;
  assign n6729 = n6728 ^ n6722 ;
  assign n6717 = n3295 ^ n719 ;
  assign n6716 = n1362 ^ n234 ;
  assign n6718 = n6717 ^ n6716 ;
  assign n6719 = n6718 ^ n2133 ;
  assign n6715 = n3414 ^ n2376 ;
  assign n6720 = n6719 ^ n6715 ;
  assign n6730 = n6729 ^ n6720 ;
  assign n6731 = n6730 ^ n5531 ;
  assign n6732 = ~n6714 & ~n6731 ;
  assign n6746 = n6745 ^ n6732 ;
  assign n6801 = n2693 ^ n419 ;
  assign n6800 = n1981 ^ n974 ;
  assign n6802 = n6801 ^ n6800 ;
  assign n6803 = n6802 ^ n2875 ;
  assign n6796 = n2905 ^ n171 ;
  assign n6797 = n6796 ^ n507 ;
  assign n6793 = n546 ^ n214 ;
  assign n6794 = n6793 ^ n296 ;
  assign n6791 = n743 ^ n517 ;
  assign n6792 = n6791 ^ n575 ;
  assign n6795 = n6794 ^ n6792 ;
  assign n6798 = n6797 ^ n6795 ;
  assign n6799 = n6798 ^ n606 ;
  assign n6804 = n6803 ^ n6799 ;
  assign n6788 = n1753 ^ n584 ;
  assign n6787 = n770 ^ n522 ;
  assign n6789 = n6788 ^ n6787 ;
  assign n6785 = n4777 ^ n3647 ;
  assign n6783 = n542 ^ n339 ;
  assign n6784 = n6783 ^ n3756 ;
  assign n6786 = n6785 ^ n6784 ;
  assign n6790 = n6789 ^ n6786 ;
  assign n6805 = n6804 ^ n6790 ;
  assign n6777 = n514 ^ n378 ;
  assign n6778 = n6777 ^ n437 ;
  assign n6775 = n3140 ^ n803 ;
  assign n6776 = n6775 ^ n1008 ;
  assign n6779 = n6778 ^ n6776 ;
  assign n6774 = n1915 ^ n1397 ;
  assign n6780 = n6779 ^ n6774 ;
  assign n6771 = n5539 ^ n4710 ;
  assign n3770 = n825 ^ n385 ;
  assign n6770 = n6682 ^ n3770 ;
  assign n6772 = n6771 ^ n6770 ;
  assign n6773 = n6772 ^ n3383 ;
  assign n6781 = n6780 ^ n6773 ;
  assign n4944 = n2969 ^ n230 ;
  assign n6769 = n5735 ^ n4944 ;
  assign n6782 = n6781 ^ n6769 ;
  assign n6806 = n6805 ^ n6782 ;
  assign n6807 = ~n5598 & ~n6806 ;
  assign n6747 = n3434 ^ n3199 ;
  assign n6748 = n6747 ^ n3435 ;
  assign n6749 = n6748 ^ n3434 ;
  assign n6750 = n6749 ^ n6733 ;
  assign n6751 = n6750 ^ n3518 ;
  assign n6752 = n6751 ^ n6750 ;
  assign n6753 = n6749 ^ n3248 ;
  assign n6755 = n6753 ^ n3022 ;
  assign n6754 = n6753 ^ n3055 ;
  assign n6756 = n6755 ^ n6754 ;
  assign n6759 = x30 & n6756 ;
  assign n6760 = n6759 ^ n6755 ;
  assign n6761 = ~n3518 & ~n6760 ;
  assign n6762 = n6761 ^ n6753 ;
  assign n6763 = n6762 ^ n6733 ;
  assign n6764 = n6763 ^ n6750 ;
  assign n6765 = ~n6752 & ~n6764 ;
  assign n6766 = n6765 ^ n6750 ;
  assign n6767 = ~x31 & ~n6766 ;
  assign n6768 = n6767 ^ n6762 ;
  assign n6808 = n6807 ^ n6768 ;
  assign n6856 = x30 & ~n3055 ;
  assign n6857 = n6856 ^ n3022 ;
  assign n6858 = ~n3518 & ~n6857 ;
  assign n6839 = n3434 ^ n3198 ;
  assign n6840 = n6839 ^ n3022 ;
  assign n6842 = n6840 ^ n3055 ;
  assign n6841 = n6840 ^ n3196 ;
  assign n6843 = n6842 ^ n6841 ;
  assign n6846 = x30 & n6843 ;
  assign n6847 = n6846 ^ n6842 ;
  assign n6848 = ~n3518 & ~n6847 ;
  assign n6849 = n6848 ^ n6840 ;
  assign n6850 = n6849 ^ n3022 ;
  assign n6859 = n6858 ^ n6850 ;
  assign n6860 = ~x31 & ~n6859 ;
  assign n6861 = n6860 ^ n6849 ;
  assign n6831 = n2868 ^ n269 ;
  assign n6832 = n6831 ^ n395 ;
  assign n6830 = n615 ^ n478 ;
  assign n6833 = n6832 ^ n6830 ;
  assign n6834 = n6833 ^ n738 ;
  assign n6835 = n6834 ^ n1614 ;
  assign n4037 = n602 ^ n440 ;
  assign n4036 = n465 ^ n389 ;
  assign n4038 = n4037 ^ n4036 ;
  assign n6827 = n4038 ^ n2344 ;
  assign n6825 = n571 ^ n464 ;
  assign n3583 = n1925 ^ n241 ;
  assign n6826 = n6825 ^ n3583 ;
  assign n6828 = n6827 ^ n6826 ;
  assign n6822 = n2905 ^ n1719 ;
  assign n6821 = n3166 ^ n437 ;
  assign n6823 = n6822 ^ n6821 ;
  assign n6820 = n1220 ^ n658 ;
  assign n6824 = n6823 ^ n6820 ;
  assign n6829 = n6828 ^ n6824 ;
  assign n6836 = n6835 ^ n6829 ;
  assign n6816 = n3366 ^ n778 ;
  assign n6815 = n802 ^ n570 ;
  assign n6817 = n6816 ^ n6815 ;
  assign n6813 = n1048 ^ n831 ;
  assign n6812 = n490 ^ n184 ;
  assign n6814 = n6813 ^ n6812 ;
  assign n6818 = n6817 ^ n6814 ;
  assign n6809 = n2205 ^ n520 ;
  assign n6810 = n6809 ^ n1898 ;
  assign n3897 = n1179 ^ n562 ;
  assign n6811 = n6810 ^ n3897 ;
  assign n6819 = n6818 ^ n6811 ;
  assign n6837 = n6836 ^ n6819 ;
  assign n6838 = n2790 & ~n6837 ;
  assign n6862 = n6861 ^ n6838 ;
  assign n6900 = n1087 ^ n336 ;
  assign n6901 = n6900 ^ n1036 ;
  assign n6902 = n6901 ^ n2949 ;
  assign n6903 = n6902 ^ n6825 ;
  assign n6896 = n3296 ^ n1300 ;
  assign n6895 = n1106 ^ n470 ;
  assign n6897 = n6896 ^ n6895 ;
  assign n6893 = n1624 ^ n385 ;
  assign n6894 = n6893 ^ n2796 ;
  assign n6898 = n6897 ^ n6894 ;
  assign n6891 = n4181 ^ n3200 ;
  assign n6892 = n6891 ^ n904 ;
  assign n6899 = n6898 ^ n6892 ;
  assign n6904 = n6903 ^ n6899 ;
  assign n6888 = n2358 ^ n774 ;
  assign n6889 = n6888 ^ n1607 ;
  assign n6885 = n510 ^ n322 ;
  assign n6886 = n6885 ^ n528 ;
  assign n6887 = n6886 ^ n2162 ;
  assign n6890 = n6889 ^ n6887 ;
  assign n6905 = n6904 ^ n6890 ;
  assign n3773 = n2403 ^ n256 ;
  assign n6917 = n3773 ^ n272 ;
  assign n6918 = n6917 ^ n640 ;
  assign n3603 = n1498 ^ n567 ;
  assign n6915 = n3603 ^ n378 ;
  assign n6916 = n6915 ^ n1066 ;
  assign n6919 = n6918 ^ n6916 ;
  assign n6920 = n6919 ^ n3192 ;
  assign n6911 = n1823 ^ n886 ;
  assign n4111 = n618 ^ n317 ;
  assign n6910 = n4111 ^ n2316 ;
  assign n6912 = n6911 ^ n6910 ;
  assign n6913 = n6912 ^ n2335 ;
  assign n6907 = n3317 ^ n240 ;
  assign n6908 = n6907 ^ n589 ;
  assign n6906 = n818 ^ n798 ;
  assign n6909 = n6908 ^ n6906 ;
  assign n6914 = n6913 ^ n6909 ;
  assign n6921 = n6920 ^ n6914 ;
  assign n6922 = n6921 ^ n2131 ;
  assign n6923 = ~n6905 & ~n6922 ;
  assign n6877 = x30 & ~n3196 ;
  assign n6878 = n6877 ^ n3055 ;
  assign n6879 = ~n3518 & ~n6878 ;
  assign n6880 = n6879 ^ n3055 ;
  assign n6863 = n3433 ^ n3197 ;
  assign n6864 = n6863 ^ n3055 ;
  assign n6881 = n6880 ^ n6864 ;
  assign n6866 = n6864 ^ n3124 ;
  assign n6865 = n6864 ^ n3196 ;
  assign n6867 = n6866 ^ n6865 ;
  assign n6870 = ~x30 & n6867 ;
  assign n6871 = n6870 ^ n6866 ;
  assign n6872 = ~n3518 & ~n6871 ;
  assign n6882 = n6881 ^ n6872 ;
  assign n6883 = x31 & ~n6882 ;
  assign n6884 = n6883 ^ n6880 ;
  assign n6924 = n6923 ^ n6884 ;
  assign n6956 = ~n3431 & ~n3801 ;
  assign n6957 = n6956 ^ n3196 ;
  assign n6958 = n3518 & ~n6957 ;
  assign n6959 = n6958 ^ n3801 ;
  assign n6951 = n3124 & ~n3850 ;
  assign n6960 = n6959 ^ n6951 ;
  assign n6950 = ~n3429 & n22543 ;
  assign n6961 = n6960 ^ n6950 ;
  assign n4046 = n2082 ^ n585 ;
  assign n4047 = n4046 ^ n1374 ;
  assign n4045 = n2032 ^ n1542 ;
  assign n4048 = n4047 ^ n4045 ;
  assign n4043 = n514 ^ n150 ;
  assign n4042 = n753 ^ n454 ;
  assign n4044 = n4043 ^ n4042 ;
  assign n4049 = n4048 ^ n4044 ;
  assign n4050 = n4049 ^ n1063 ;
  assign n4039 = n4038 ^ n655 ;
  assign n4040 = n4039 ^ n4035 ;
  assign n4032 = n762 ^ n178 ;
  assign n4033 = n4032 ^ n399 ;
  assign n4041 = n4040 ^ n4033 ;
  assign n4051 = n4050 ^ n4041 ;
  assign n6925 = n4051 ^ n1401 ;
  assign n6942 = n6783 ^ n919 ;
  assign n6941 = n2432 ^ n1735 ;
  assign n6943 = n6942 ^ n6941 ;
  assign n6938 = n896 ^ n248 ;
  assign n6939 = n6938 ^ n609 ;
  assign n6937 = n908 ^ n744 ;
  assign n6940 = n6939 ^ n6937 ;
  assign n6944 = n6943 ^ n6940 ;
  assign n6935 = n701 ^ n251 ;
  assign n6936 = n6935 ^ n675 ;
  assign n6945 = n6944 ^ n6936 ;
  assign n6931 = n2310 ^ n357 ;
  assign n6932 = n6931 ^ n798 ;
  assign n6929 = n2358 ^ n347 ;
  assign n6930 = n6929 ^ n1001 ;
  assign n6933 = n6932 ^ n6930 ;
  assign n6926 = n956 ^ n256 ;
  assign n6927 = n6926 ^ n1298 ;
  assign n6928 = n6927 ^ n2623 ;
  assign n6934 = n6933 ^ n6928 ;
  assign n6946 = n6945 ^ n6934 ;
  assign n6947 = n6946 ^ n3301 ;
  assign n4976 = n1838 ^ n1106 ;
  assign n4975 = n950 ^ n556 ;
  assign n4977 = n4976 ^ n4975 ;
  assign n4973 = n2445 ^ n390 ;
  assign n4974 = n4973 ^ n767 ;
  assign n4978 = n4977 ^ n4974 ;
  assign n4966 = n917 ^ n747 ;
  assign n4972 = n4971 ^ n4966 ;
  assign n4979 = n4978 ^ n4972 ;
  assign n4964 = n3234 ^ n2080 ;
  assign n4960 = n1360 ^ n826 ;
  assign n4961 = n4960 ^ n570 ;
  assign n4962 = n4961 ^ n1604 ;
  assign n4211 = n2519 ^ n182 ;
  assign n4963 = n4962 ^ n4211 ;
  assign n4965 = n4964 ^ n4963 ;
  assign n4980 = n4979 ^ n4965 ;
  assign n6948 = n6947 ^ n4980 ;
  assign n6949 = ~n6925 & ~n6948 ;
  assign n6963 = n6961 ^ n6949 ;
  assign n6962 = n6949 & n6961 ;
  assign n6964 = n6963 ^ n6962 ;
  assign n6965 = n6964 ^ n6884 ;
  assign n6966 = n6924 & n6965 ;
  assign n6967 = n6966 ^ n6884 ;
  assign n6968 = n6967 ^ n6861 ;
  assign n6969 = ~n6862 & ~n6968 ;
  assign n6970 = n6969 ^ n6861 ;
  assign n6971 = n6970 ^ n6768 ;
  assign n6972 = n6808 & n6971 ;
  assign n6973 = n6972 ^ n6970 ;
  assign n6974 = n6973 ^ n6745 ;
  assign n6975 = ~n6746 & n6974 ;
  assign n6976 = n6975 ^ n6745 ;
  assign n6977 = n6976 ^ n6702 ;
  assign n6978 = ~n6703 & n6977 ;
  assign n6979 = n6978 ^ n6702 ;
  assign n6980 = n6979 ^ n6659 ;
  assign n6981 = n6662 & n6980 ;
  assign n6660 = n6659 ^ n6650 ;
  assign n6982 = n6981 ^ n6660 ;
  assign n6983 = n6651 & ~n6982 ;
  assign n6984 = n6983 ^ n6650 ;
  assign n6985 = n6984 ^ n6629 ;
  assign n6986 = ~n6640 & n6985 ;
  assign n6987 = n6986 ^ n6629 ;
  assign n6988 = n6987 ^ n6620 ;
  assign n6989 = ~n6621 & ~n6988 ;
  assign n6990 = n6989 ^ n6620 ;
  assign n6991 = n6990 ^ n6609 ;
  assign n6992 = n6611 & n6991 ;
  assign n6993 = n6992 ^ n6990 ;
  assign n6994 = n6993 ^ n6590 ;
  assign n6995 = n6598 & n6994 ;
  assign n6996 = n6995 ^ n6590 ;
  assign n6588 = n6479 ^ n6469 ;
  assign n6997 = n6996 ^ n6588 ;
  assign n7007 = ~n1541 & n4651 ;
  assign n7005 = ~n40 & ~n1819 ;
  assign n7003 = n6588 ^ x23 ;
  assign n5239 = x23 ^ x22 ;
  assign n7000 = ~n4985 & ~n5239 ;
  assign n7001 = n7000 ^ n4986 ;
  assign n7002 = n35 & n7001 ;
  assign n7004 = n7003 ^ n7002 ;
  assign n7006 = n7005 ^ n7004 ;
  assign n7008 = n7007 ^ n7006 ;
  assign n7009 = n6997 & ~n7008 ;
  assign n7010 = n7009 ^ n6996 ;
  assign n7011 = n7010 ^ n6579 ;
  assign n7012 = ~n6587 & ~n7011 ;
  assign n7013 = n7012 ^ n6579 ;
  assign n7014 = n7013 ^ n6569 ;
  assign n7015 = n6577 & ~n7014 ;
  assign n7016 = n7015 ^ n6569 ;
  assign n7017 = n7016 ^ n6559 ;
  assign n7018 = n6565 & n7017 ;
  assign n6566 = n6559 ^ n6554 ;
  assign n7019 = n7018 ^ n6566 ;
  assign n7020 = ~n6555 & n7019 ;
  assign n7021 = n7020 ^ n6554 ;
  assign n7023 = n7022 ^ n7021 ;
  assign n7140 = x9 ^ x8 ;
  assign n7149 = x11 & n7140 ;
  assign n7138 = x8 & x9 ;
  assign n7139 = n7138 ^ x10 ;
  assign n20239 = n7149 ^ n7139 ;
  assign n7141 = x10 & n7140 ;
  assign n7142 = n7141 ^ n7139 ;
  assign n20240 = n20239 ^ n7142 ;
  assign n7157 = ~n3509 & n20240 ;
  assign n20254 = x10 ^ x9 ;
  assign n20255 = ~n7140 & ~n20254 ;
  assign n20257 = n20255 ^ x11 ;
  assign n7146 = x10 & n7138 ;
  assign n7145 = ~x11 & ~n20255 ;
  assign n7147 = n7146 ^ n7145 ;
  assign n7148 = ~n20257 ^ n7147 ;
  assign n7158 = n7157 ^ n7148 ;
  assign n7159 = ~n368 & n7158 ;
  assign n7160 = n7159 ^ x11 ;
  assign n7059 = ~n4359 & n6163 ;
  assign n7056 = ~n856 & n6148 ;
  assign n7054 = ~n1248 & n20437 ;
  assign n7052 = n7010 ^ n6587 ;
  assign n7053 = n7052 ^ x17 ;
  assign n7055 = n7054 ^ n7053 ;
  assign n7057 = n7056 ^ n7055 ;
  assign n7051 = ~n1119 & n6143 ;
  assign n7058 = n7057 ^ n7051 ;
  assign n7060 = n7059 ^ n7058 ;
  assign n7069 = n4475 & n5221 ;
  assign n7064 = n7008 ^ n6996 ;
  assign n7065 = n7064 ^ x20 ;
  assign n7063 = ~n1345 & n5220 ;
  assign n7066 = n7065 ^ n7063 ;
  assign n7062 = ~n1751 & n13433 ;
  assign n7067 = n7066 ^ n7062 ;
  assign n7061 = ~n1450 & n5426 ;
  assign n7068 = n7067 ^ n7061 ;
  assign n7070 = n7069 ^ n7068 ;
  assign n7079 = ~n4495 & n5221 ;
  assign n7076 = ~n1751 & n5426 ;
  assign n7074 = ~n1670 & n13433 ;
  assign n7072 = n6993 ^ n6598 ;
  assign n7073 = n7072 ^ x20 ;
  assign n7075 = n7074 ^ n7073 ;
  assign n7077 = n7076 ^ n7075 ;
  assign n7071 = ~n1450 & n5220 ;
  assign n7078 = n7077 ^ n7071 ;
  assign n7080 = n7079 ^ n7078 ;
  assign n7089 = n6990 ^ n6611 ;
  assign n7085 = n4656 & ~n4892 ;
  assign n7084 = ~n1897 & n4651 ;
  assign n7086 = n7085 ^ n7084 ;
  assign n7087 = n7086 ^ x23 ;
  assign n7082 = ~n40 & ~n1972 ;
  assign n7081 = ~n1541 & n4655 ;
  assign n7083 = n7082 ^ n7081 ;
  assign n7088 = n7087 ^ n7083 ;
  assign n7090 = n7089 ^ n7088 ;
  assign n7099 = n6987 ^ n6621 ;
  assign n7124 = n7099 ^ n7089 ;
  assign n7097 = ~n4435 & n5480 ;
  assign n7095 = ~n2288 & n4600 ;
  assign n7092 = ~n2199 & ~n4434 ;
  assign n7091 = ~n2371 & n20603 ;
  assign n7093 = n7092 ^ n7091 ;
  assign n7094 = n7093 ^ x26 ;
  assign n7096 = n7095 ^ n7094 ;
  assign n7098 = n7097 ^ n7096 ;
  assign n7100 = n7099 ^ n7098 ;
  assign n7110 = ~n4435 & n6449 ;
  assign n7108 = ~n2467 & n20603 ;
  assign n7105 = ~n2288 & ~n4434 ;
  assign n7104 = ~n2371 & n4600 ;
  assign n7106 = n7105 ^ n7104 ;
  assign n7107 = n7106 ^ x26 ;
  assign n7109 = n7108 ^ n7107 ;
  assign n7111 = n7110 ^ n7109 ;
  assign n7121 = n7111 ^ n7099 ;
  assign n7116 = ~n2589 & n3985 ;
  assign n7112 = n7111 ^ x29 ;
  assign n7103 = ~n2552 & n4369 ;
  assign n7113 = n7112 ^ n7103 ;
  assign n7102 = ~n2657 & n3837 ;
  assign n7114 = n7113 ^ n7102 ;
  assign n7101 = n3983 & n6212 ;
  assign n7115 = n7114 ^ n7101 ;
  assign n7117 = n7116 ^ n7115 ;
  assign n7118 = n6984 ^ n6640 ;
  assign n7119 = n7118 ^ n7111 ;
  assign n7120 = n7117 & n7119 ;
  assign n7122 = n7121 ^ n7120 ;
  assign n7123 = n7100 & n7122 ;
  assign n7125 = n7124 ^ n7123 ;
  assign n7126 = ~n7090 & ~n7125 ;
  assign n7127 = n7126 ^ n7089 ;
  assign n7128 = n7127 ^ n7072 ;
  assign n7129 = n7080 & ~n7128 ;
  assign n7130 = n7129 ^ n7072 ;
  assign n7131 = n7130 ^ n7064 ;
  assign n7132 = n7070 & n7131 ;
  assign n7133 = n7132 ^ n7064 ;
  assign n7134 = n7133 ^ n7052 ;
  assign n7135 = ~n7060 & ~n7134 ;
  assign n7136 = n7135 ^ n7052 ;
  assign n7030 = ~n540 & ~n6547 ;
  assign n7029 = ~n408 & ~n6529 ;
  assign n7031 = n7030 ^ n7029 ;
  assign n7026 = ~x13 & ~n3839 ;
  assign n7027 = n7026 ^ n3505 ;
  assign n7028 = n6391 & ~n7027 ;
  assign n7032 = n7031 ^ n7028 ;
  assign n7033 = x14 & n7032 ;
  assign n7035 = ~x14 & n6528 ;
  assign n7040 = ~n3505 & n7035 ;
  assign n7034 = n7031 ^ x14 ;
  assign n7041 = n7040 ^ n7034 ;
  assign n7042 = ~n7033 & ~n7041 ;
  assign n7046 = n6535 ^ n6403 ;
  assign n7047 = n7046 ^ n6534 ;
  assign n7048 = n3840 & n7047 ;
  assign n7049 = n7042 & n7048 ;
  assign n7043 = n7013 ^ n6577 ;
  assign n7044 = n7043 ^ n7033 ;
  assign n7045 = n7044 ^ n7042 ;
  assign n7050 = n7049 ^ n7045 ;
  assign n7137 = n7136 ^ n7050 ;
  assign n7161 = n7160 ^ n7137 ;
  assign n7184 = n7133 ^ n7060 ;
  assign n7281 = n7184 ^ n7160 ;
  assign n7168 = ~n698 & ~n6547 ;
  assign n7167 = ~n540 & ~n6529 ;
  assign n7169 = n7168 ^ n7167 ;
  assign n7164 = ~x13 & ~n3811 ;
  assign n7165 = n7164 ^ n408 ;
  assign n7166 = n6391 & ~n7165 ;
  assign n7170 = n7169 ^ n7166 ;
  assign n7171 = x14 & n7170 ;
  assign n7177 = ~n408 & n7035 ;
  assign n7172 = n7169 ^ x14 ;
  assign n7178 = n7177 ^ n7172 ;
  assign n7179 = ~n7171 & ~n7178 ;
  assign n7181 = n3812 & n7047 ;
  assign n7182 = n7179 & n7181 ;
  assign n7180 = n7179 ^ n7171 ;
  assign n7183 = n7182 ^ n7180 ;
  assign n7185 = n7184 ^ n7183 ;
  assign n7194 = ~n4336 & n6163 ;
  assign n7192 = ~n1248 & n6143 ;
  assign n7189 = ~n1119 & n6148 ;
  assign n7188 = ~n990 & n20437 ;
  assign n7190 = n7189 ^ n7188 ;
  assign n7191 = n7190 ^ x17 ;
  assign n7193 = n7192 ^ n7191 ;
  assign n7195 = n7194 ^ n7193 ;
  assign n7186 = n7130 ^ n7070 ;
  assign n7196 = n7195 ^ n7186 ;
  assign n7205 = n4580 & n6163 ;
  assign n7202 = ~n1248 & n6148 ;
  assign n7200 = ~n1345 & n20437 ;
  assign n7198 = n7127 ^ n7080 ;
  assign n7199 = n7198 ^ x17 ;
  assign n7201 = n7200 ^ n7199 ;
  assign n7203 = n7202 ^ n7201 ;
  assign n7197 = ~n990 & n6143 ;
  assign n7204 = n7203 ^ n7197 ;
  assign n7206 = n7205 ^ n7204 ;
  assign n7216 = n4690 & n5221 ;
  assign n7214 = ~n1670 & n5426 ;
  assign n7211 = ~n1819 & n13433 ;
  assign n7210 = ~n1751 & n5220 ;
  assign n7212 = n7211 ^ n7210 ;
  assign n7213 = n7212 ^ x20 ;
  assign n7215 = n7214 ^ n7213 ;
  assign n7217 = n7216 ^ n7215 ;
  assign n7209 = n7125 ^ n7088 ;
  assign n7218 = n7217 ^ n7209 ;
  assign n7267 = ~n2095 & n4651 ;
  assign n7240 = n7118 ^ n7117 ;
  assign n7226 = ~n4435 & n5696 ;
  assign n7224 = ~n2552 & n20603 ;
  assign n7221 = ~n2467 & n4600 ;
  assign n7220 = ~n2371 & ~n4434 ;
  assign n7222 = n7221 ^ n7220 ;
  assign n7223 = n7222 ^ x26 ;
  assign n7225 = n7224 ^ n7223 ;
  assign n7227 = n7226 ^ n7225 ;
  assign n7219 = n6982 ^ n6641 ;
  assign n7228 = n7227 ^ n7219 ;
  assign n7236 = ~n2657 & n3985 ;
  assign n7232 = n7227 ^ x29 ;
  assign n7231 = ~n2712 & n3837 ;
  assign n7233 = n7232 ^ n7231 ;
  assign n7230 = ~n2589 & n4369 ;
  assign n7234 = n7233 ^ n7230 ;
  assign n6079 = n6078 ^ n2589 ;
  assign n7229 = n3983 & n6079 ;
  assign n7235 = n7234 ^ n7229 ;
  assign n7237 = n7236 ^ n7235 ;
  assign n7238 = n7228 & n7237 ;
  assign n7239 = n7238 ^ n7227 ;
  assign n7241 = n7240 ^ n7239 ;
  assign n7251 = ~n2199 & n4651 ;
  assign n7249 = ~n40 & ~n2095 ;
  assign n7247 = n7239 ^ x23 ;
  assign n7244 = ~n4884 & n5239 ;
  assign n7245 = n7244 ^ n1897 ;
  assign n7246 = n35 & ~n7245 ;
  assign n7248 = n7247 ^ n7246 ;
  assign n7250 = n7249 ^ n7248 ;
  assign n7252 = n7251 ^ n7250 ;
  assign n7253 = n7241 & ~n7252 ;
  assign n7254 = n7253 ^ n7240 ;
  assign n7264 = n7254 ^ x23 ;
  assign n7261 = n5239 & n5286 ;
  assign n7262 = n7261 ^ n1972 ;
  assign n7263 = n35 & ~n7262 ;
  assign n7265 = n7264 ^ n7263 ;
  assign n7256 = ~n40 & ~n1897 ;
  assign n7266 = n7265 ^ n7256 ;
  assign n7268 = n7267 ^ n7266 ;
  assign n7269 = n7122 ^ n7098 ;
  assign n7270 = n7269 ^ n7254 ;
  assign n7271 = n7268 & n7270 ;
  assign n7255 = n7254 ^ n7209 ;
  assign n7272 = n7271 ^ n7255 ;
  assign n7273 = ~n7218 & n7272 ;
  assign n7274 = n7273 ^ n7217 ;
  assign n7275 = n7274 ^ n7198 ;
  assign n7276 = ~n7206 & ~n7275 ;
  assign n7207 = n7198 ^ n7186 ;
  assign n7277 = n7276 ^ n7207 ;
  assign n7278 = n7196 & ~n7277 ;
  assign n7187 = n7186 ^ n7183 ;
  assign n7279 = n7278 ^ n7187 ;
  assign n7280 = n7185 & n7279 ;
  assign n7282 = n7281 ^ n7280 ;
  assign n7283 = ~n7161 & ~n7282 ;
  assign n7284 = n7283 ^ n7160 ;
  assign n7285 = n7136 ^ n7043 ;
  assign n7286 = ~n7050 & n7285 ;
  assign n7287 = n7286 ^ n7136 ;
  assign n7288 = n7287 ^ n7284 ;
  assign n7289 = n7016 ^ n6565 ;
  assign n7290 = n7289 ^ n7284 ;
  assign n7291 = n7288 & ~n7290 ;
  assign n7292 = ~n7284 & n7291 ;
  assign n7293 = n7019 ^ n6527 ;
  assign n7294 = n7293 ^ n7291 ;
  assign n7302 = n3515 & n20240 ;
  assign n7298 = n7279 ^ n7184 ;
  assign n7299 = n7298 ^ x11 ;
  assign n7297 = ~n368 & n7142 ;
  assign n7300 = n7299 ^ n7297 ;
  assign n7296 = ~n3505 & n7148 ;
  assign n7301 = n7300 ^ n7296 ;
  assign n7303 = n7302 ^ n7301 ;
  assign n7319 = n7274 ^ n7206 ;
  assign n7306 = ~n856 & ~n6529 ;
  assign n7305 = ~n1119 & ~n6547 ;
  assign n7307 = n7306 ^ n7305 ;
  assign n7318 = n7307 ^ x14 ;
  assign n7320 = n7319 ^ n7318 ;
  assign n7310 = x14 ^ x13 ;
  assign n7311 = n7310 ^ n698 ;
  assign n7308 = n7307 ^ n698 ;
  assign n7312 = n7311 ^ n7308 ;
  assign n7315 = n3495 & n7312 ;
  assign n7316 = n7315 ^ n7308 ;
  assign n7317 = n6391 & ~n7316 ;
  assign n7321 = n7320 ^ n7317 ;
  assign n7331 = n4986 & n5221 ;
  assign n7328 = ~n1541 & n13433 ;
  assign n7326 = ~n1819 & n5426 ;
  assign n7324 = n7269 ^ n7268 ;
  assign n7325 = n7324 ^ x20 ;
  assign n7327 = n7326 ^ n7325 ;
  assign n7329 = n7328 ^ n7327 ;
  assign n7323 = ~n1670 & n5220 ;
  assign n7330 = n7329 ^ n7323 ;
  assign n7332 = n7331 ^ n7330 ;
  assign n7341 = ~n5154 & n5221 ;
  assign n7338 = ~n1541 & n5426 ;
  assign n7336 = ~n1819 & n5220 ;
  assign n7334 = n7252 ^ n7240 ;
  assign n7335 = n7334 ^ x20 ;
  assign n7337 = n7336 ^ n7335 ;
  assign n7339 = n7338 ^ n7337 ;
  assign n7333 = ~n1972 & n13433 ;
  assign n7340 = n7339 ^ n7333 ;
  assign n7342 = n7341 ^ n7340 ;
  assign n7351 = ~n2288 & n4651 ;
  assign n7348 = ~n40 & ~n2199 ;
  assign n7346 = n4656 & n5760 ;
  assign n7344 = n7237 ^ n7219 ;
  assign n7345 = n7344 ^ x23 ;
  assign n7347 = n7346 ^ n7345 ;
  assign n7349 = n7348 ^ n7347 ;
  assign n7343 = ~n2095 & n4655 ;
  assign n7350 = n7349 ^ n7343 ;
  assign n7352 = n7351 ^ n7350 ;
  assign n7493 = n6979 ^ n6662 ;
  assign n7363 = ~n2748 & n3985 ;
  assign n7360 = ~n2839 & n3837 ;
  assign n7358 = ~n3324 & n4369 ;
  assign n7356 = n6973 ^ n6746 ;
  assign n7357 = n7356 ^ x29 ;
  assign n7359 = n7358 ^ n7357 ;
  assign n7361 = n7360 ^ n7359 ;
  assign n7354 = n6643 ^ n3324 ;
  assign n7355 = n3983 & n7354 ;
  assign n7362 = n7361 ^ n7355 ;
  assign n7364 = n7363 ^ n7362 ;
  assign n7374 = ~n3248 & n3837 ;
  assign n7369 = n6967 ^ n6862 ;
  assign n7370 = n7369 ^ x29 ;
  assign n7368 = n3983 & ~n6695 ;
  assign n7371 = n7370 ^ n7368 ;
  assign n7367 = ~n2935 & n3985 ;
  assign n7372 = n7371 ^ n7367 ;
  assign n7366 = ~n2839 & n4369 ;
  assign n7373 = n7372 ^ n7366 ;
  assign n7375 = n7374 ^ n7373 ;
  assign n7384 = n6964 ^ n6924 ;
  assign n7379 = ~n3022 & n3837 ;
  assign n7378 = ~n2935 & n4369 ;
  assign n7380 = n7379 ^ n7378 ;
  assign n7381 = n7380 ^ x29 ;
  assign n7377 = n3983 & n6736 ;
  assign n7382 = n7381 ^ n7377 ;
  assign n7376 = ~n3248 & n3985 ;
  assign n7383 = n7382 ^ n7376 ;
  assign n7385 = n7384 ^ n7383 ;
  assign n7396 = ~n3055 & n3837 ;
  assign n7394 = ~n3022 & n3985 ;
  assign n7390 = n5065 & ~n6749 ;
  assign n7391 = n7390 ^ n3248 ;
  assign n7392 = n3833 & ~n7391 ;
  assign n7393 = n7392 ^ x29 ;
  assign n7395 = n7394 ^ n7393 ;
  assign n7397 = n7396 ^ n7395 ;
  assign n7411 = ~n3196 & n3985 ;
  assign n7410 = ~n3124 & n3837 ;
  assign n7412 = n7411 ^ n7410 ;
  assign n7408 = n3983 & ~n6863 ;
  assign n7407 = ~n3055 & n3833 ;
  assign n7409 = n7408 ^ n7407 ;
  assign n7413 = n7412 ^ n7409 ;
  assign n7423 = ~n3429 & n3837 ;
  assign n7422 = ~n3124 & n3985 ;
  assign n7424 = n7423 ^ n7422 ;
  assign n7419 = n3431 & n5065 ;
  assign n7420 = n7419 ^ n3196 ;
  assign n7421 = n3833 & ~n7420 ;
  assign n7425 = n7424 ^ n7421 ;
  assign n7426 = ~n3124 & n3833 ;
  assign n7427 = ~n3429 & n3835 ;
  assign n7428 = ~n7426 & n7427 ;
  assign n7429 = n7428 ^ n7426 ;
  assign n7430 = ~n7425 & ~n7429 ;
  assign n7433 = ~x30 & ~n3429 ;
  assign n7436 = ~n7430 & ~n7433 ;
  assign n7437 = x29 & n7436 ;
  assign n7438 = n7437 ^ x29 ;
  assign n7414 = ~n60 & ~n3429 ;
  assign n7439 = n7438 ^ n7414 ;
  assign n7440 = ~n7413 & n7439 ;
  assign n7441 = n7440 ^ n7414 ;
  assign n7402 = ~n3022 & n4369 ;
  assign n7401 = ~n3196 & n3837 ;
  assign n7403 = n7402 ^ n7401 ;
  assign n7404 = n7403 ^ x29 ;
  assign n7400 = n3983 & n6840 ;
  assign n7405 = n7404 ^ n7400 ;
  assign n7399 = ~n3055 & n3985 ;
  assign n7406 = n7405 ^ n7399 ;
  assign n7442 = n7441 ^ n7406 ;
  assign n7444 = ~n3124 & n3518 ;
  assign n7443 = ~n3429 & ~n3801 ;
  assign n7445 = n7444 ^ n7443 ;
  assign n7446 = n7445 ^ n7406 ;
  assign n7447 = n7442 & ~n7446 ;
  assign n7448 = n7447 ^ n7441 ;
  assign n7453 = n7397 & n7448 ;
  assign n7398 = n7397 ^ n6962 ;
  assign n7449 = n7448 ^ n7397 ;
  assign n7450 = ~n7398 & ~n7449 ;
  assign n7451 = n7450 ^ n6962 ;
  assign n7454 = n7453 ^ n7451 ;
  assign n7452 = n7451 ^ n7383 ;
  assign n7457 = n7452 ^ n6964 ;
  assign n7458 = n7457 ^ n7452 ;
  assign n7459 = ~n7454 & ~n7458 ;
  assign n7460 = n7459 ^ n7452 ;
  assign n7461 = ~n7385 & ~n7460 ;
  assign n7462 = n7461 ^ n7383 ;
  assign n7463 = n7462 ^ n7369 ;
  assign n7464 = n7375 & n7463 ;
  assign n7465 = n7464 ^ n7369 ;
  assign n7365 = n6970 ^ n6808 ;
  assign n7466 = n7465 ^ n7365 ;
  assign n7474 = ~n2839 & n3985 ;
  assign n7470 = n7365 ^ x29 ;
  assign n7469 = ~n2748 & n4369 ;
  assign n7471 = n7470 ^ n7469 ;
  assign n7468 = ~n2935 & n3837 ;
  assign n7472 = n7471 ^ n7468 ;
  assign n7467 = n3983 & ~n6302 ;
  assign n7473 = n7472 ^ n7467 ;
  assign n7475 = n7474 ^ n7473 ;
  assign n7476 = ~n7466 & n7475 ;
  assign n7477 = n7476 ^ n7465 ;
  assign n7478 = n7477 ^ n7356 ;
  assign n7479 = ~n7364 & ~n7478 ;
  assign n7480 = n7479 ^ n7356 ;
  assign n7353 = n6976 ^ n6703 ;
  assign n7481 = n7480 ^ n7353 ;
  assign n7489 = ~n3324 & n3985 ;
  assign n7485 = n7353 ^ x29 ;
  assign n7484 = ~n2748 & n3837 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7483 = ~n2712 & n4369 ;
  assign n7487 = n7486 ^ n7483 ;
  assign n7482 = n3983 & n6623 ;
  assign n7488 = n7487 ^ n7482 ;
  assign n7490 = n7489 ^ n7488 ;
  assign n7491 = n7481 & n7490 ;
  assign n7492 = n7491 ^ n7480 ;
  assign n7494 = n7493 ^ n7492 ;
  assign n7502 = ~n4435 & n6008 ;
  assign n7498 = n7493 ^ x26 ;
  assign n7497 = ~n2552 & n4600 ;
  assign n7499 = n7498 ^ n7497 ;
  assign n7496 = ~n2589 & n20603 ;
  assign n7500 = n7499 ^ n7496 ;
  assign n7495 = ~n2467 & ~n4434 ;
  assign n7501 = n7500 ^ n7495 ;
  assign n7503 = n7502 ^ n7501 ;
  assign n7504 = ~n7494 & n7503 ;
  assign n7505 = n7504 ^ n7493 ;
  assign n7506 = n7505 ^ n7344 ;
  assign n7507 = n7352 & n7506 ;
  assign n7508 = n7507 ^ n7344 ;
  assign n7509 = n7508 ^ n7334 ;
  assign n7510 = n7342 & n7509 ;
  assign n7511 = n7510 ^ n7334 ;
  assign n7512 = n7511 ^ n7324 ;
  assign n7513 = n7332 & n7512 ;
  assign n7514 = n7513 ^ n7324 ;
  assign n7322 = n7272 ^ n7217 ;
  assign n7515 = n7514 ^ n7322 ;
  assign n7523 = n4307 & n6163 ;
  assign n7519 = n7322 ^ x17 ;
  assign n7518 = ~n1450 & n20437 ;
  assign n7520 = n7519 ^ n7518 ;
  assign n7517 = ~n990 & n6148 ;
  assign n7521 = n7520 ^ n7517 ;
  assign n7516 = ~n1345 & n6143 ;
  assign n7522 = n7521 ^ n7516 ;
  assign n7524 = n7523 ^ n7522 ;
  assign n7525 = ~n7515 & n7524 ;
  assign n7526 = n7525 ^ n7514 ;
  assign n7527 = n7526 ^ n7319 ;
  assign n7528 = ~n7321 & ~n7527 ;
  assign n7529 = n7528 ^ n7319 ;
  assign n7304 = n7277 ^ n7195 ;
  assign n7530 = n7529 ^ n7304 ;
  assign n7538 = ~n698 & ~n6529 ;
  assign n7537 = ~n856 & ~n6547 ;
  assign n7539 = n7538 ^ n7537 ;
  assign n7534 = ~x13 & ~n3955 ;
  assign n7535 = n7534 ^ n540 ;
  assign n7536 = n6391 & ~n7535 ;
  assign n7540 = n7539 ^ n7536 ;
  assign n7541 = x14 & n7540 ;
  assign n7547 = ~n540 & n7035 ;
  assign n7542 = n7539 ^ x14 ;
  assign n7548 = n7547 ^ n7542 ;
  assign n7549 = ~n7541 & ~n7548 ;
  assign n7552 = n3968 & n7047 ;
  assign n7553 = n7549 & n7552 ;
  assign n7550 = n7541 ^ n7304 ;
  assign n7551 = n7550 ^ n7549 ;
  assign n7554 = n7553 ^ n7551 ;
  assign n7555 = n7530 & ~n7554 ;
  assign n7556 = n7555 ^ n7529 ;
  assign n7557 = n7556 ^ n7298 ;
  assign n7558 = n7303 & ~n7557 ;
  assign n7559 = n7558 ^ n7298 ;
  assign n7295 = n7282 ^ n7137 ;
  assign n7560 = n7559 ^ n7295 ;
  assign n11827 = ~n3505 & n7142 ;
  assign n11825 = ~n408 & n7148 ;
  assign n11822 = ~n3513 & n20240 ;
  assign n11821 = ~n368 & n7140 ;
  assign n11823 = n11822 ^ n11821 ;
  assign n11824 = n11823 ^ x11 ;
  assign n11826 = n11825 ^ n11824 ;
  assign n11828 = n11827 ^ n11826 ;
  assign n11820 = n7554 ^ n7529 ;
  assign n11829 = n11828 ^ n11820 ;
  assign n8137 = x6 ^ x5 ;
  assign n8145 = x8 & n8137 ;
  assign n8146 = n8145 ^ n8137 ;
  assign n8147 = n8146 ^ x7 ;
  assign n8138 = x7 & n8137 ;
  assign n8148 = n8147 ^ n8138 ;
  assign n8149 = n8148 ^ n8145 ;
  assign n8150 = n8149 ^ n8147 ;
  assign n8166 = n3515 & n8150 ;
  assign n8133 = x5 & x6 ;
  assign n8136 = n8133 ^ x7 ;
  assign n8139 = n8138 ^ n8136 ;
  assign n19031 = n8139 ^ n8137 ;
  assign n8143 = x8 & n19031 ;
  assign n8134 = x7 & n8133 ;
  assign n8135 = n8134 ^ x8 ;
  assign n8144 = n8143 ^ n8135 ;
  assign n8164 = ~n3505 & n8144 ;
  assign n8162 = ~n368 & n8139 ;
  assign n8126 = n3812 & n20240 ;
  assign n8124 = ~n698 & n7148 ;
  assign n8121 = ~n540 & n7142 ;
  assign n7150 = n7149 ^ n7140 ;
  assign n7151 = n7150 ^ n7141 ;
  assign n8120 = ~n408 & n7151 ;
  assign n8122 = n8121 ^ n8120 ;
  assign n8123 = n8122 ^ x11 ;
  assign n8125 = n8124 ^ n8123 ;
  assign n8127 = n8126 ^ n8125 ;
  assign n7602 = ~n4495 & n6163 ;
  assign n7599 = ~n1751 & n6143 ;
  assign n7597 = ~n1450 & n6148 ;
  assign n7595 = n7508 ^ n7342 ;
  assign n7596 = n7595 ^ x17 ;
  assign n7598 = n7597 ^ n7596 ;
  assign n7600 = n7599 ^ n7598 ;
  assign n7594 = ~n1670 & n20437 ;
  assign n7601 = n7600 ^ n7594 ;
  assign n7603 = n7602 ^ n7601 ;
  assign n7612 = ~n4892 & n5221 ;
  assign n7609 = ~n1972 & n5426 ;
  assign n7607 = ~n1897 & n13433 ;
  assign n7605 = n7505 ^ n7352 ;
  assign n7606 = n7605 ^ x20 ;
  assign n7608 = n7607 ^ n7606 ;
  assign n7610 = n7609 ^ n7608 ;
  assign n7604 = ~n1541 & n5220 ;
  assign n7611 = n7610 ^ n7604 ;
  assign n7613 = n7612 ^ n7611 ;
  assign n7622 = ~n2371 & n4651 ;
  assign n7617 = n7503 ^ n7492 ;
  assign n7618 = n7617 ^ x23 ;
  assign n7616 = n4656 & n5480 ;
  assign n7619 = n7618 ^ n7616 ;
  assign n7615 = ~n40 & ~n2288 ;
  assign n7620 = n7619 ^ n7615 ;
  assign n7614 = ~n2199 & n4655 ;
  assign n7621 = n7620 ^ n7614 ;
  assign n7623 = n7622 ^ n7621 ;
  assign n7633 = ~n4435 & n6079 ;
  assign n7630 = ~n2657 & n4600 ;
  assign n7628 = ~n2712 & n20603 ;
  assign n7626 = n7477 ^ n7364 ;
  assign n7627 = n7626 ^ x26 ;
  assign n7629 = n7628 ^ n7627 ;
  assign n7631 = n7630 ^ n7629 ;
  assign n7625 = ~n2589 & ~n4434 ;
  assign n7632 = n7631 ^ n7625 ;
  assign n7634 = n7633 ^ n7632 ;
  assign n7644 = ~n4435 & n6623 ;
  assign n7641 = ~n2712 & ~n4434 ;
  assign n7639 = ~n3324 & n4600 ;
  assign n7637 = n7462 ^ n7375 ;
  assign n7638 = n7637 ^ x26 ;
  assign n7640 = n7639 ^ n7638 ;
  assign n7642 = n7641 ^ n7640 ;
  assign n7636 = ~n2748 & n20603 ;
  assign n7643 = n7642 ^ n7636 ;
  assign n7645 = n7644 ^ n7643 ;
  assign n7656 = ~n4435 & n7354 ;
  assign n7653 = ~n2839 & n20603 ;
  assign n7651 = ~n2748 & n4600 ;
  assign n7648 = n7452 ^ n6924 ;
  assign n7647 = ~n6964 & n7454 ;
  assign n7649 = n7648 ^ n7647 ;
  assign n7650 = n7649 ^ x26 ;
  assign n7652 = n7651 ^ n7650 ;
  assign n7654 = n7653 ^ n7652 ;
  assign n7646 = ~n3324 & ~n4434 ;
  assign n7655 = n7654 ^ n7646 ;
  assign n7657 = n7656 ^ n7655 ;
  assign n7749 = n7446 ^ n7441 ;
  assign n7729 = ~n4435 & n6753 ;
  assign n7727 = ~n3055 & n20603 ;
  assign n7724 = ~n3022 & n4600 ;
  assign n7723 = ~n3248 & ~n4434 ;
  assign n7725 = n7724 ^ n7723 ;
  assign n7726 = n7725 ^ x26 ;
  assign n7728 = n7727 ^ n7726 ;
  assign n7730 = n7729 ^ n7728 ;
  assign n7674 = ~n4435 & n6840 ;
  assign n7672 = ~n3022 & ~n4434 ;
  assign n7669 = ~n3196 & n20603 ;
  assign n7668 = ~n3055 & n4600 ;
  assign n7670 = n7669 ^ n7668 ;
  assign n7671 = n7670 ^ x26 ;
  assign n7673 = n7672 ^ n7671 ;
  assign n7675 = n7674 ^ n7673 ;
  assign n7666 = ~n3429 & n3832 ;
  assign n7667 = n7666 ^ n7426 ;
  assign n7676 = n7675 ^ n7667 ;
  assign n7677 = ~n3429 & n3833 ;
  assign n7678 = n4600 ^ n96 ;
  assign n7679 = n96 & ~n3124 ;
  assign n7680 = x26 & ~n7679 ;
  assign n7681 = n7678 & n7680 ;
  assign n7682 = ~n3429 & n7681 ;
  assign n7683 = n7682 ^ n7680 ;
  assign n7694 = n96 & ~n3196 ;
  assign n7701 = n285 & ~n3124 ;
  assign n7702 = n7694 & n7701 ;
  assign n7703 = n7702 ^ n7694 ;
  assign n7695 = ~n20603 ^ n7694 ;
  assign n7704 = n7703 ^ n7695 ;
  assign n7705 = n3429 & ~n7704 ;
  assign n7706 = n7705 ^ n7695 ;
  assign n7688 = n3196 & n3429 ;
  assign n7691 = ~n4435 & n7688 ;
  assign n7692 = n7691 ^ n4600 ;
  assign n7693 = ~n3124 & n7692 ;
  assign n7707 = n7706 ^ n7693 ;
  assign n7708 = n7683 & n7707 ;
  assign n7709 = ~n7677 & ~n7708 ;
  assign n7716 = ~n4435 & n6864 ;
  assign n7714 = ~n3124 & n20603 ;
  assign n7711 = ~n3196 & n4600 ;
  assign n7710 = ~n3055 & ~n4434 ;
  assign n7712 = n7711 ^ n7710 ;
  assign n7713 = n7712 ^ x26 ;
  assign n7715 = n7714 ^ n7713 ;
  assign n7717 = n7716 ^ n7715 ;
  assign n7718 = n7709 & n7717 ;
  assign n7719 = n7718 ^ n7717 ;
  assign n7720 = n7719 ^ n7667 ;
  assign n7721 = n7676 & ~n7720 ;
  assign n7722 = n7721 ^ n7675 ;
  assign n7731 = n7730 ^ n7722 ;
  assign n7733 = n7730 ^ n7425 ;
  assign n7732 = x29 & n7429 ;
  assign n7734 = n7733 ^ n7732 ;
  assign n7735 = n7731 & n7734 ;
  assign n7736 = n7735 ^ n7730 ;
  assign n7664 = n7414 ^ n7413 ;
  assign n7661 = n7433 ^ n7414 ;
  assign n7662 = n7661 ^ n7430 ;
  assign n7663 = x29 & ~n7662 ;
  assign n7665 = n7664 ^ n7663 ;
  assign n7737 = n7736 ^ n7665 ;
  assign n7745 = ~n4435 & n6736 ;
  assign n7741 = n7665 ^ x26 ;
  assign n7740 = ~n3022 & n20603 ;
  assign n7742 = n7741 ^ n7740 ;
  assign n7739 = ~n3248 & n4600 ;
  assign n7743 = n7742 ^ n7739 ;
  assign n7738 = ~n2935 & ~n4434 ;
  assign n7744 = n7743 ^ n7738 ;
  assign n7746 = n7745 ^ n7744 ;
  assign n7747 = n7737 & ~n7746 ;
  assign n7748 = n7747 ^ n7736 ;
  assign n7750 = n7749 ^ n7748 ;
  assign n7758 = ~n4435 & ~n6695 ;
  assign n7754 = n7749 ^ x26 ;
  assign n7753 = ~n3248 & n20603 ;
  assign n7755 = n7754 ^ n7753 ;
  assign n7752 = ~n2935 & n4600 ;
  assign n7756 = n7755 ^ n7752 ;
  assign n7751 = ~n2839 & ~n4434 ;
  assign n7757 = n7756 ^ n7751 ;
  assign n7759 = n7758 ^ n7757 ;
  assign n7760 = n7750 & n7759 ;
  assign n7761 = n7760 ^ n7749 ;
  assign n7658 = n7397 ^ n6961 ;
  assign n7659 = n7658 ^ n6949 ;
  assign n7660 = n7659 ^ n7448 ;
  assign n7762 = n7761 ^ n7660 ;
  assign n7770 = ~n4435 & ~n6302 ;
  assign n7766 = n7660 ^ x26 ;
  assign n7765 = ~n2748 & ~n4434 ;
  assign n7767 = n7766 ^ n7765 ;
  assign n7764 = ~n2935 & n20603 ;
  assign n7768 = n7767 ^ n7764 ;
  assign n7763 = ~n2839 & n4600 ;
  assign n7769 = n7768 ^ n7763 ;
  assign n7771 = n7770 ^ n7769 ;
  assign n7772 = n7762 & ~n7771 ;
  assign n7773 = n7772 ^ n7761 ;
  assign n7774 = n7773 ^ n7649 ;
  assign n7775 = ~n7657 & ~n7774 ;
  assign n7776 = n7775 ^ n7649 ;
  assign n7777 = n7776 ^ n7637 ;
  assign n7778 = n7645 & ~n7777 ;
  assign n7779 = n7778 ^ n7637 ;
  assign n7635 = n7475 ^ n7465 ;
  assign n7780 = n7779 ^ n7635 ;
  assign n7788 = ~n4435 & n6229 ;
  assign n7784 = n7635 ^ x26 ;
  assign n7783 = ~n2712 & n4600 ;
  assign n7785 = n7784 ^ n7783 ;
  assign n7782 = ~n2657 & ~n4434 ;
  assign n7786 = n7785 ^ n7782 ;
  assign n7781 = ~n3324 & n20603 ;
  assign n7787 = n7786 ^ n7781 ;
  assign n7789 = n7788 ^ n7787 ;
  assign n7790 = ~n7780 & n7789 ;
  assign n7791 = n7790 ^ n7779 ;
  assign n7792 = n7791 ^ n7626 ;
  assign n7793 = ~n7634 & ~n7792 ;
  assign n7794 = n7793 ^ n7626 ;
  assign n7624 = n7490 ^ n7480 ;
  assign n7795 = n7794 ^ n7624 ;
  assign n7803 = ~n4435 & n6212 ;
  assign n7799 = n7624 ^ x26 ;
  assign n7798 = ~n2589 & n4600 ;
  assign n7800 = n7799 ^ n7798 ;
  assign n7797 = ~n2657 & n20603 ;
  assign n7801 = n7800 ^ n7797 ;
  assign n7796 = ~n2552 & ~n4434 ;
  assign n7802 = n7801 ^ n7796 ;
  assign n7804 = n7803 ^ n7802 ;
  assign n7805 = ~n7795 & ~n7804 ;
  assign n7806 = n7805 ^ n7794 ;
  assign n7807 = n7806 ^ n7617 ;
  assign n7808 = ~n7623 & n7807 ;
  assign n7809 = n7808 ^ n7617 ;
  assign n7810 = n7809 ^ n7605 ;
  assign n7811 = n7613 & ~n7810 ;
  assign n7812 = n7811 ^ n7605 ;
  assign n7813 = n7812 ^ n7595 ;
  assign n7814 = n7603 & n7813 ;
  assign n7815 = n7814 ^ n7595 ;
  assign n7592 = n4475 & n6163 ;
  assign n7589 = ~n1751 & n20437 ;
  assign n7587 = ~n1345 & n6148 ;
  assign n7585 = n7511 ^ n7332 ;
  assign n7586 = n7585 ^ x17 ;
  assign n7588 = n7587 ^ n7586 ;
  assign n7590 = n7589 ^ n7588 ;
  assign n7584 = ~n1450 & n6143 ;
  assign n7591 = n7590 ^ n7584 ;
  assign n7593 = n7592 ^ n7591 ;
  assign n7816 = n7815 ^ n7593 ;
  assign n7565 = ~n1248 & ~n6529 ;
  assign n7564 = ~n990 & ~n6547 ;
  assign n7566 = n7565 ^ n7564 ;
  assign n7567 = ~n4336 & ~n7566 ;
  assign n7568 = n7567 ^ n1119 ;
  assign n7569 = x13 & ~n7568 ;
  assign n7570 = n7569 ^ n1119 ;
  assign n7571 = n6391 & ~n7570 ;
  assign n7572 = n7571 ^ n7566 ;
  assign n7573 = ~x14 & n7572 ;
  assign n7817 = n7816 ^ n7573 ;
  assign n7575 = x14 & n7047 ;
  assign n7580 = ~n1119 & n7575 ;
  assign n7574 = n7566 ^ x14 ;
  assign n7581 = n7580 ^ n7574 ;
  assign n7582 = ~n7573 & n7581 ;
  assign n7818 = n7817 ^ n7582 ;
  assign n7561 = ~n4336 & n6528 ;
  assign n7583 = n7561 & n7582 ;
  assign n7819 = n7818 ^ n7583 ;
  assign n7856 = n4690 & n6163 ;
  assign n7853 = ~n1751 & n6148 ;
  assign n7851 = ~n1819 & n20437 ;
  assign n7849 = n7809 ^ n7613 ;
  assign n7850 = n7849 ^ x17 ;
  assign n7852 = n7851 ^ n7850 ;
  assign n7854 = n7853 ^ n7852 ;
  assign n7848 = ~n1670 & n6143 ;
  assign n7855 = n7854 ^ n7848 ;
  assign n7857 = n7856 ^ n7855 ;
  assign n7866 = n5221 & ~n5287 ;
  assign n7863 = ~n1972 & n5220 ;
  assign n7861 = ~n2095 & n13433 ;
  assign n7859 = n7806 ^ n7623 ;
  assign n7860 = n7859 ^ x20 ;
  assign n7862 = n7861 ^ n7860 ;
  assign n7864 = n7863 ^ n7862 ;
  assign n7858 = ~n1897 & n5426 ;
  assign n7865 = n7864 ^ n7858 ;
  assign n7867 = n7866 ^ n7865 ;
  assign n7877 = ~n2371 & n4655 ;
  assign n7874 = ~n40 & ~n2467 ;
  assign n7872 = n4656 & n5696 ;
  assign n7870 = n7791 ^ n7634 ;
  assign n7871 = n7870 ^ x23 ;
  assign n7873 = n7872 ^ n7871 ;
  assign n7875 = n7874 ^ n7873 ;
  assign n7869 = ~n2552 & n4651 ;
  assign n7876 = n7875 ^ n7869 ;
  assign n7878 = n7877 ^ n7876 ;
  assign n7888 = ~n2657 & n4651 ;
  assign n7885 = ~n40 & ~n2589 ;
  assign n7883 = n4656 & n6212 ;
  assign n7881 = n7776 ^ n7645 ;
  assign n7882 = n7881 ^ x23 ;
  assign n7884 = n7883 ^ n7882 ;
  assign n7886 = n7885 ^ n7884 ;
  assign n7880 = ~n2552 & n4655 ;
  assign n7887 = n7886 ^ n7880 ;
  assign n7889 = n7888 ^ n7887 ;
  assign n8016 = n7771 ^ n7761 ;
  assign n7991 = n7746 ^ n7736 ;
  assign n7898 = n4656 & ~n6695 ;
  assign n7897 = ~n40 & ~n2935 ;
  assign n7899 = n7898 ^ n7897 ;
  assign n7900 = n7899 ^ x23 ;
  assign n7895 = ~n3248 & n4651 ;
  assign n7894 = ~n2839 & n4655 ;
  assign n7896 = n7895 ^ n7894 ;
  assign n7901 = n7900 ^ n7896 ;
  assign n7893 = n7719 ^ n7676 ;
  assign n7902 = n7901 ^ n7893 ;
  assign n7909 = n4656 & n6736 ;
  assign n7908 = ~n40 & ~n3248 ;
  assign n7910 = n7909 ^ n7908 ;
  assign n7911 = n7910 ^ x23 ;
  assign n7906 = ~n3022 & n4651 ;
  assign n7905 = ~n2935 & n4655 ;
  assign n7907 = n7906 ^ n7905 ;
  assign n7912 = n7911 ^ n7907 ;
  assign n7903 = n7708 ^ n7677 ;
  assign n7904 = n7903 ^ n7717 ;
  assign n7913 = n7912 ^ n7904 ;
  assign n7684 = n7683 ^ x26 ;
  assign n7923 = n7707 ^ n7684 ;
  assign n7918 = n4656 & n6753 ;
  assign n7917 = ~n40 & ~n3022 ;
  assign n7919 = n7918 ^ n7917 ;
  assign n7920 = n7919 ^ x23 ;
  assign n7915 = ~n3248 & n4655 ;
  assign n7914 = ~n3055 & n4651 ;
  assign n7916 = n7915 ^ n7914 ;
  assign n7921 = n7920 ^ n7916 ;
  assign n7924 = n7923 ^ n7921 ;
  assign n7932 = n4656 & n6840 ;
  assign n7931 = ~n40 & ~n3055 ;
  assign n7933 = n7932 ^ n7931 ;
  assign n7934 = n7933 ^ x23 ;
  assign n7929 = ~n3022 & n4655 ;
  assign n7928 = ~n3196 & n4651 ;
  assign n7930 = n7929 ^ n7928 ;
  assign n7935 = n7934 ^ n7930 ;
  assign n7925 = n133 ^ n89 ;
  assign n7926 = ~n3429 & ~n7925 ;
  assign n7927 = n7926 ^ n7679 ;
  assign n7936 = n7935 ^ n7927 ;
  assign n7937 = n96 & ~n3429 ;
  assign n7938 = n35 & ~n3124 ;
  assign n7939 = x23 & ~n7938 ;
  assign n7940 = ~n42 & n7939 ;
  assign n7941 = ~n3429 & n7940 ;
  assign n7942 = n7941 ^ n7939 ;
  assign n7953 = ~n3429 & n4651 ;
  assign n7952 = n35 & ~n3196 ;
  assign n7954 = n7953 ^ n7952 ;
  assign n7949 = n3429 & n4656 ;
  assign n7950 = n7949 ^ n40 ;
  assign n7951 = ~n3124 & ~n7950 ;
  assign n7955 = n7954 ^ n7951 ;
  assign n7956 = n7942 & ~n7955 ;
  assign n7957 = ~n7937 & ~n7956 ;
  assign n7962 = n4656 & n6864 ;
  assign n7961 = ~n40 & ~n3196 ;
  assign n7963 = n7962 ^ n7961 ;
  assign n7964 = n7963 ^ x23 ;
  assign n7959 = ~n3124 & n4651 ;
  assign n7958 = ~n3055 & n4655 ;
  assign n7960 = n7959 ^ n7958 ;
  assign n7965 = n7964 ^ n7960 ;
  assign n7966 = n7957 & n7965 ;
  assign n7967 = n7966 ^ n7965 ;
  assign n7968 = n7967 ^ n7927 ;
  assign n7969 = n7936 & ~n7968 ;
  assign n7970 = n7969 ^ n7935 ;
  assign n7971 = n7970 ^ n7921 ;
  assign n7972 = ~n7924 & n7971 ;
  assign n7922 = n7921 ^ n7904 ;
  assign n7973 = n7972 ^ n7922 ;
  assign n7974 = n7913 & ~n7973 ;
  assign n7975 = n7974 ^ n7912 ;
  assign n7976 = n7975 ^ n7901 ;
  assign n7977 = n7902 & n7976 ;
  assign n7978 = n7977 ^ n7901 ;
  assign n7892 = n7734 ^ n7722 ;
  assign n7979 = n7978 ^ n7892 ;
  assign n7987 = ~n2935 & n4651 ;
  assign n7983 = n7892 ^ x23 ;
  assign n7982 = n4656 & ~n6302 ;
  assign n7984 = n7983 ^ n7982 ;
  assign n7981 = ~n40 & ~n2839 ;
  assign n7985 = n7984 ^ n7981 ;
  assign n7980 = ~n2748 & n4655 ;
  assign n7986 = n7985 ^ n7980 ;
  assign n7988 = n7987 ^ n7986 ;
  assign n7989 = n7979 & ~n7988 ;
  assign n7990 = n7989 ^ n7978 ;
  assign n7992 = n7991 ^ n7990 ;
  assign n8000 = ~n3324 & n4655 ;
  assign n7996 = n7991 ^ x23 ;
  assign n7995 = n4656 & n7354 ;
  assign n7997 = n7996 ^ n7995 ;
  assign n7994 = ~n2839 & n4651 ;
  assign n7998 = n7997 ^ n7994 ;
  assign n7993 = ~n40 & ~n2748 ;
  assign n7999 = n7998 ^ n7993 ;
  assign n8001 = n8000 ^ n7999 ;
  assign n8002 = n7992 & n8001 ;
  assign n8003 = n8002 ^ n7991 ;
  assign n7891 = n7759 ^ n7748 ;
  assign n8004 = n8003 ^ n7891 ;
  assign n8012 = ~n2712 & n4655 ;
  assign n8008 = n7891 ^ x23 ;
  assign n8007 = n4656 & n6623 ;
  assign n8009 = n8008 ^ n8007 ;
  assign n8006 = ~n40 & ~n3324 ;
  assign n8010 = n8009 ^ n8006 ;
  assign n8005 = ~n2748 & n4651 ;
  assign n8011 = n8010 ^ n8005 ;
  assign n8013 = n8012 ^ n8011 ;
  assign n8014 = n8004 & ~n8013 ;
  assign n8015 = n8014 ^ n8003 ;
  assign n8017 = n8016 ^ n8015 ;
  assign n8025 = ~n2657 & n4655 ;
  assign n8021 = n8016 ^ x23 ;
  assign n8020 = n4656 & n6229 ;
  assign n8022 = n8021 ^ n8020 ;
  assign n8019 = ~n40 & ~n2712 ;
  assign n8023 = n8022 ^ n8019 ;
  assign n8018 = ~n3324 & n4651 ;
  assign n8024 = n8023 ^ n8018 ;
  assign n8026 = n8025 ^ n8024 ;
  assign n8027 = n8017 & n8026 ;
  assign n8028 = n8027 ^ n8016 ;
  assign n7890 = n7773 ^ n7657 ;
  assign n8029 = n8028 ^ n7890 ;
  assign n8037 = ~n2589 & n4655 ;
  assign n8033 = n7890 ^ x23 ;
  assign n8032 = n4656 & n6079 ;
  assign n8034 = n8033 ^ n8032 ;
  assign n8031 = ~n40 & ~n2657 ;
  assign n8035 = n8034 ^ n8031 ;
  assign n8030 = ~n2712 & n4651 ;
  assign n8036 = n8035 ^ n8030 ;
  assign n8038 = n8037 ^ n8036 ;
  assign n8039 = ~n8029 & n8038 ;
  assign n8040 = n8039 ^ n8028 ;
  assign n8041 = n8040 ^ n7881 ;
  assign n8042 = ~n7889 & ~n8041 ;
  assign n8043 = n8042 ^ n7881 ;
  assign n7879 = n7789 ^ n7779 ;
  assign n8044 = n8043 ^ n7879 ;
  assign n8052 = ~n2589 & n4651 ;
  assign n8048 = n7879 ^ x23 ;
  assign n8047 = n4656 & n6008 ;
  assign n8049 = n8048 ^ n8047 ;
  assign n8046 = ~n40 & ~n2552 ;
  assign n8050 = n8049 ^ n8046 ;
  assign n8045 = ~n2467 & n4655 ;
  assign n8051 = n8050 ^ n8045 ;
  assign n8053 = n8052 ^ n8051 ;
  assign n8054 = n8044 & n8053 ;
  assign n8055 = n8054 ^ n8043 ;
  assign n8056 = n8055 ^ n7870 ;
  assign n8057 = ~n7878 & n8056 ;
  assign n8058 = n8057 ^ n7870 ;
  assign n7868 = n7804 ^ n7794 ;
  assign n8059 = n8058 ^ n7868 ;
  assign n8067 = ~n2288 & n4655 ;
  assign n8063 = n7868 ^ x23 ;
  assign n8062 = n4656 & n6449 ;
  assign n8064 = n8063 ^ n8062 ;
  assign n8061 = ~n40 & ~n2371 ;
  assign n8065 = n8064 ^ n8061 ;
  assign n8060 = ~n2467 & n4651 ;
  assign n8066 = n8065 ^ n8060 ;
  assign n8068 = n8067 ^ n8066 ;
  assign n8069 = n8059 & n8068 ;
  assign n8070 = n8069 ^ n8058 ;
  assign n8071 = n8070 ^ n7859 ;
  assign n8072 = n7867 & ~n8071 ;
  assign n8073 = n8072 ^ n7859 ;
  assign n8074 = n8073 ^ n7849 ;
  assign n8075 = ~n7857 & ~n8074 ;
  assign n8076 = n8075 ^ n7849 ;
  assign n7847 = n7812 ^ n7603 ;
  assign n8077 = n8076 ^ n7847 ;
  assign n8085 = ~n1345 & ~n6547 ;
  assign n8084 = ~n990 & ~n6529 ;
  assign n8086 = n8085 ^ n8084 ;
  assign n8081 = x13 & ~n4333 ;
  assign n8082 = n8081 ^ n1248 ;
  assign n8083 = n6391 & ~n8082 ;
  assign n8087 = n8086 ^ n8083 ;
  assign n8088 = ~x14 & n8087 ;
  assign n8098 = n8088 ^ n7847 ;
  assign n8094 = ~n1248 & n7575 ;
  assign n8089 = n8086 ^ x14 ;
  assign n8095 = n8094 ^ n8089 ;
  assign n8096 = ~n8088 & n8095 ;
  assign n8099 = n8098 ^ n8096 ;
  assign n8078 = n4580 & n6528 ;
  assign n8097 = n8078 & n8096 ;
  assign n8100 = n8099 ^ n8097 ;
  assign n8101 = ~n8077 & ~n8100 ;
  assign n8102 = n8101 ^ n8076 ;
  assign n7840 = n7524 ^ n7514 ;
  assign n7841 = n7840 ^ x14 ;
  assign n7838 = n7047 ^ n6537 ;
  assign n7825 = ~n1248 & ~n6547 ;
  assign n7824 = ~n1119 & ~n6529 ;
  assign n7826 = n7825 ^ n7824 ;
  assign n7839 = n7838 ^ n7826 ;
  assign n7842 = n7841 ^ n7839 ;
  assign n7831 = ~n856 & n7826 ;
  assign n7832 = x14 & n7831 ;
  assign n7833 = n7832 ^ x14 ;
  assign n7834 = n7833 ^ x13 ;
  assign n7835 = ~n3493 & n7834 ;
  assign n7836 = n7835 ^ n856 ;
  assign n7837 = n6391 & ~n7836 ;
  assign n7843 = n7842 ^ n7837 ;
  assign n7820 = n7815 ^ n7585 ;
  assign n7821 = ~n7593 & n7820 ;
  assign n7822 = n7821 ^ n7815 ;
  assign n7844 = n7843 ^ n7822 ;
  assign n7845 = n7844 ^ n7816 ;
  assign n7846 = n7845 ^ n7844 ;
  assign n8103 = n8102 ^ n7846 ;
  assign n8104 = n7819 & ~n8103 ;
  assign n8105 = n8104 ^ n7845 ;
  assign n8160 = n8127 ^ n8105 ;
  assign n8161 = n8160 ^ x8 ;
  assign n8163 = n8162 ^ n8161 ;
  assign n8165 = n8164 ^ n8163 ;
  assign n8167 = n8166 ^ n8165 ;
  assign n8177 = ~n3930 & n20240 ;
  assign n8174 = ~n1119 & n7148 ;
  assign n8172 = ~n698 & n7151 ;
  assign n8170 = n8100 ^ n8076 ;
  assign n8171 = n8170 ^ x11 ;
  assign n8173 = n8172 ^ n8171 ;
  assign n8175 = n8174 ^ n8173 ;
  assign n8169 = ~n856 & n7142 ;
  assign n8176 = n8175 ^ n8169 ;
  assign n8178 = n8177 ^ n8176 ;
  assign n8186 = ~n1450 & ~n6547 ;
  assign n8185 = ~n1345 & ~n6529 ;
  assign n8187 = n8186 ^ n8185 ;
  assign n8182 = x13 & ~n3486 ;
  assign n8183 = n8182 ^ n990 ;
  assign n8184 = n6391 & ~n8183 ;
  assign n8188 = n8187 ^ n8184 ;
  assign n8189 = ~x14 & n8188 ;
  assign n8195 = ~n990 & n7575 ;
  assign n8190 = n8187 ^ x14 ;
  assign n8196 = n8195 ^ n8190 ;
  assign n8197 = ~n8189 & n8196 ;
  assign n8201 = n4307 & n6528 ;
  assign n8202 = n8197 & n8201 ;
  assign n8198 = n8073 ^ n7857 ;
  assign n8199 = n8198 ^ n8189 ;
  assign n8200 = n8199 ^ n8197 ;
  assign n8203 = n8202 ^ n8200 ;
  assign n8212 = n4986 & n6163 ;
  assign n8209 = ~n1541 & n20437 ;
  assign n8207 = ~n1819 & n6143 ;
  assign n8205 = n8070 ^ n7867 ;
  assign n8206 = n8205 ^ x17 ;
  assign n8208 = n8207 ^ n8206 ;
  assign n8210 = n8209 ^ n8208 ;
  assign n8204 = ~n1670 & n6148 ;
  assign n8211 = n8210 ^ n8204 ;
  assign n8213 = n8212 ^ n8211 ;
  assign n8223 = n5221 & n5760 ;
  assign n8220 = ~n2199 & n5426 ;
  assign n8218 = ~n2095 & n5220 ;
  assign n8216 = n8055 ^ n7878 ;
  assign n8217 = n8216 ^ x20 ;
  assign n8219 = n8218 ^ n8217 ;
  assign n8221 = n8220 ^ n8219 ;
  assign n8215 = ~n2288 & n13433 ;
  assign n8222 = n8221 ^ n8215 ;
  assign n8224 = n8223 ^ n8222 ;
  assign n8234 = n5221 & n6449 ;
  assign n8231 = ~n2288 & n5220 ;
  assign n8229 = ~n2467 & n13433 ;
  assign n8227 = n8040 ^ n7889 ;
  assign n8228 = n8227 ^ x20 ;
  assign n8230 = n8229 ^ n8228 ;
  assign n8232 = n8231 ^ n8230 ;
  assign n8226 = ~n2371 & n5426 ;
  assign n8233 = n8232 ^ n8226 ;
  assign n8235 = n8234 ^ n8233 ;
  assign n8412 = n8038 ^ n8028 ;
  assign n8243 = n5221 & n6008 ;
  assign n8241 = ~n2589 & n13433 ;
  assign n8238 = ~n2467 & n5220 ;
  assign n8237 = ~n2552 & n5426 ;
  assign n8239 = n8238 ^ n8237 ;
  assign n8240 = n8239 ^ x20 ;
  assign n8242 = n8241 ^ n8240 ;
  assign n8244 = n8243 ^ n8242 ;
  assign n8236 = n8026 ^ n8015 ;
  assign n8245 = n8244 ^ n8236 ;
  assign n8396 = n8013 ^ n8003 ;
  assign n8408 = n8396 ^ n8244 ;
  assign n8383 = n8001 ^ n7990 ;
  assign n8358 = n7975 ^ n7902 ;
  assign n8255 = n5221 & ~n6302 ;
  assign n8253 = ~n2748 & n5220 ;
  assign n8250 = ~n2935 & n13433 ;
  assign n8249 = ~n2839 & n5426 ;
  assign n8251 = n8250 ^ n8249 ;
  assign n8252 = n8251 ^ x20 ;
  assign n8254 = n8253 ^ n8252 ;
  assign n8256 = n8255 ^ n8254 ;
  assign n8248 = n7970 ^ n7924 ;
  assign n8257 = n8256 ^ n8248 ;
  assign n8265 = n5221 & ~n6695 ;
  assign n8263 = ~n3248 & n13433 ;
  assign n8260 = ~n2935 & n5426 ;
  assign n8259 = ~n2839 & n5220 ;
  assign n8261 = n8260 ^ n8259 ;
  assign n8262 = n8261 ^ x20 ;
  assign n8264 = n8263 ^ n8262 ;
  assign n8266 = n8265 ^ n8264 ;
  assign n8258 = n7967 ^ n7936 ;
  assign n8267 = n8266 ^ n8258 ;
  assign n8276 = n5221 & n6736 ;
  assign n8274 = ~n2935 & n5220 ;
  assign n8271 = ~n3022 & n13433 ;
  assign n8270 = ~n3248 & n5426 ;
  assign n8272 = n8271 ^ n8270 ;
  assign n8273 = n8272 ^ x20 ;
  assign n8275 = n8274 ^ n8273 ;
  assign n8277 = n8276 ^ n8275 ;
  assign n8268 = n7956 ^ n7937 ;
  assign n8269 = n8268 ^ n7965 ;
  assign n8278 = n8277 ^ n8269 ;
  assign n8286 = n5221 & n6753 ;
  assign n8284 = ~n3055 & n13433 ;
  assign n8281 = ~n3022 & n5426 ;
  assign n8280 = ~n3248 & n5220 ;
  assign n8282 = n8281 ^ n8280 ;
  assign n8283 = n8282 ^ x20 ;
  assign n8285 = n8284 ^ n8283 ;
  assign n8287 = n8286 ^ n8285 ;
  assign n7943 = n7942 ^ x23 ;
  assign n8279 = n7955 ^ n7943 ;
  assign n8288 = n8287 ^ n8279 ;
  assign n8298 = n5221 & n6840 ;
  assign n8296 = ~n3022 & n5220 ;
  assign n8293 = ~n3196 & n13433 ;
  assign n8292 = ~n3055 & n5426 ;
  assign n8294 = n8293 ^ n8292 ;
  assign n8295 = n8294 ^ x20 ;
  assign n8297 = n8296 ^ n8295 ;
  assign n8299 = n8298 ^ n8297 ;
  assign n8289 = n37 ^ x22 ;
  assign n8290 = ~n3429 & ~n8289 ;
  assign n8291 = n8290 ^ n7938 ;
  assign n8300 = n8299 ^ n8291 ;
  assign n8301 = n35 & ~n3429 ;
  assign n8302 = ~n3196 & n5215 ;
  assign n8309 = ~n3124 & n5224 ;
  assign n8310 = n8302 & n8309 ;
  assign n8311 = n8310 ^ n8302 ;
  assign n8303 = n13433 ^ n8302 ;
  assign n8312 = n8311 ^ n8303 ;
  assign n8313 = n3429 & n8312 ;
  assign n8314 = n8313 ^ n8303 ;
  assign n8315 = x20 & ~n8314 ;
  assign n8316 = n5426 ^ n5215 ;
  assign n8317 = ~n3430 & n8316 ;
  assign n8318 = n8315 & n8317 ;
  assign n8319 = n8318 ^ n8315 ;
  assign n8320 = ~n8301 & ~n8319 ;
  assign n8327 = n5221 & n6864 ;
  assign n8325 = ~n3196 & n5426 ;
  assign n8322 = ~n3124 & n13433 ;
  assign n8321 = ~n3055 & n5220 ;
  assign n8323 = n8322 ^ n8321 ;
  assign n8324 = n8323 ^ x20 ;
  assign n8326 = n8325 ^ n8324 ;
  assign n8328 = n8327 ^ n8326 ;
  assign n8329 = n8320 & n8328 ;
  assign n8330 = n8329 ^ n8328 ;
  assign n8331 = n8330 ^ n8291 ;
  assign n8332 = n8300 & ~n8331 ;
  assign n8333 = n8332 ^ n8299 ;
  assign n8334 = n8333 ^ n8287 ;
  assign n8335 = n8288 & n8334 ;
  assign n8336 = n8335 ^ n8287 ;
  assign n8337 = n8336 ^ n8277 ;
  assign n8338 = n8278 & n8337 ;
  assign n8339 = n8338 ^ n8277 ;
  assign n8340 = n8339 ^ n8266 ;
  assign n8341 = n8267 & n8340 ;
  assign n8342 = n8341 ^ n8266 ;
  assign n8343 = n8342 ^ n8256 ;
  assign n8344 = ~n8257 & n8343 ;
  assign n8345 = n8344 ^ n8256 ;
  assign n8247 = n7973 ^ n7912 ;
  assign n8346 = n8345 ^ n8247 ;
  assign n8354 = n5221 & n7354 ;
  assign n8350 = n8247 ^ x20 ;
  assign n8349 = ~n2748 & n5426 ;
  assign n8351 = n8350 ^ n8349 ;
  assign n8348 = ~n2839 & n13433 ;
  assign n8352 = n8351 ^ n8348 ;
  assign n8347 = ~n3324 & n5220 ;
  assign n8353 = n8352 ^ n8347 ;
  assign n8355 = n8354 ^ n8353 ;
  assign n8356 = n8346 & ~n8355 ;
  assign n8357 = n8356 ^ n8345 ;
  assign n8359 = n8358 ^ n8357 ;
  assign n8367 = n5221 & n6623 ;
  assign n8363 = n8358 ^ x20 ;
  assign n8362 = ~n2748 & n13433 ;
  assign n8364 = n8363 ^ n8362 ;
  assign n8361 = ~n3324 & n5426 ;
  assign n8365 = n8364 ^ n8361 ;
  assign n8360 = ~n2712 & n5220 ;
  assign n8366 = n8365 ^ n8360 ;
  assign n8368 = n8367 ^ n8366 ;
  assign n8369 = n8359 & n8368 ;
  assign n8370 = n8369 ^ n8358 ;
  assign n8246 = n7988 ^ n7978 ;
  assign n8371 = n8370 ^ n8246 ;
  assign n8379 = n5221 & n6229 ;
  assign n8375 = n8246 ^ x20 ;
  assign n8374 = ~n3324 & n13433 ;
  assign n8376 = n8375 ^ n8374 ;
  assign n8373 = ~n2712 & n5426 ;
  assign n8377 = n8376 ^ n8373 ;
  assign n8372 = ~n2657 & n5220 ;
  assign n8378 = n8377 ^ n8372 ;
  assign n8380 = n8379 ^ n8378 ;
  assign n8381 = n8371 & ~n8380 ;
  assign n8382 = n8381 ^ n8370 ;
  assign n8384 = n8383 ^ n8382 ;
  assign n8392 = n5221 & n6079 ;
  assign n8388 = n8383 ^ x20 ;
  assign n8387 = ~n2712 & n13433 ;
  assign n8389 = n8388 ^ n8387 ;
  assign n8386 = ~n2657 & n5426 ;
  assign n8390 = n8389 ^ n8386 ;
  assign n8385 = ~n2589 & n5220 ;
  assign n8391 = n8390 ^ n8385 ;
  assign n8393 = n8392 ^ n8391 ;
  assign n8394 = n8384 & n8393 ;
  assign n8395 = n8394 ^ n8383 ;
  assign n8397 = n8396 ^ n8395 ;
  assign n8405 = n5221 & n6212 ;
  assign n8401 = n8396 ^ x20 ;
  assign n8400 = ~n2589 & n5426 ;
  assign n8402 = n8401 ^ n8400 ;
  assign n8399 = ~n2657 & n13433 ;
  assign n8403 = n8402 ^ n8399 ;
  assign n8398 = ~n2552 & n5220 ;
  assign n8404 = n8403 ^ n8398 ;
  assign n8406 = n8405 ^ n8404 ;
  assign n8407 = n8397 & n8406 ;
  assign n8409 = n8408 ^ n8407 ;
  assign n8410 = n8245 & n8409 ;
  assign n8411 = n8410 ^ n8244 ;
  assign n8413 = n8412 ^ n8411 ;
  assign n8421 = n5221 & n5696 ;
  assign n8417 = n8412 ^ x20 ;
  assign n8416 = ~n2467 & n5426 ;
  assign n8418 = n8417 ^ n8416 ;
  assign n8415 = ~n2552 & n13433 ;
  assign n8419 = n8418 ^ n8415 ;
  assign n8414 = ~n2371 & n5220 ;
  assign n8420 = n8419 ^ n8414 ;
  assign n8422 = n8421 ^ n8420 ;
  assign n8423 = ~n8413 & ~n8422 ;
  assign n8424 = n8423 ^ n8412 ;
  assign n8425 = n8424 ^ n8227 ;
  assign n8426 = ~n8235 & n8425 ;
  assign n8427 = n8426 ^ n8227 ;
  assign n8225 = n8053 ^ n8043 ;
  assign n8428 = n8427 ^ n8225 ;
  assign n8436 = n5221 & n5480 ;
  assign n8432 = n8225 ^ x20 ;
  assign n8431 = ~n2288 & n5426 ;
  assign n8433 = n8432 ^ n8431 ;
  assign n8430 = ~n2371 & n13433 ;
  assign n8434 = n8433 ^ n8430 ;
  assign n8429 = ~n2199 & n5220 ;
  assign n8435 = n8434 ^ n8429 ;
  assign n8437 = n8436 ^ n8435 ;
  assign n8438 = ~n8428 & ~n8437 ;
  assign n8439 = n8438 ^ n8427 ;
  assign n8440 = n8439 ^ n8216 ;
  assign n8441 = n8224 & ~n8440 ;
  assign n8442 = n8441 ^ n8216 ;
  assign n8214 = n8068 ^ n8058 ;
  assign n8443 = n8442 ^ n8214 ;
  assign n8452 = ~n2095 & n5426 ;
  assign n8450 = ~n2199 & n13433 ;
  assign n8449 = n8214 ^ x20 ;
  assign n8451 = n8450 ^ n8449 ;
  assign n8453 = n8452 ^ n8451 ;
  assign n8444 = n5824 ^ n5224 ;
  assign n8445 = n8444 ^ n5824 ;
  assign n8446 = ~n4884 & ~n8445 ;
  assign n8447 = n8446 ^ n5824 ;
  assign n8448 = n5215 & n8447 ;
  assign n8454 = n8453 ^ n8448 ;
  assign n8455 = n8443 & ~n8454 ;
  assign n8456 = n8455 ^ n8442 ;
  assign n8457 = n8456 ^ n8205 ;
  assign n8458 = ~n8213 & ~n8457 ;
  assign n8459 = n8458 ^ n8205 ;
  assign n8460 = n8459 ^ n8198 ;
  assign n8461 = ~n8203 & n8460 ;
  assign n8462 = n8461 ^ n8198 ;
  assign n8463 = n8462 ^ n8170 ;
  assign n8464 = ~n8178 & n8463 ;
  assign n8465 = n8464 ^ n8170 ;
  assign n8168 = n8102 ^ n7819 ;
  assign n8466 = n8465 ^ n8168 ;
  assign n8474 = n3968 & n20240 ;
  assign n8470 = n8168 ^ x11 ;
  assign n8469 = ~n856 & n7148 ;
  assign n8471 = n8470 ^ n8469 ;
  assign n8468 = ~n540 & n7151 ;
  assign n8472 = n8471 ^ n8468 ;
  assign n8467 = ~n698 & n7142 ;
  assign n8473 = n8472 ^ n8467 ;
  assign n8475 = n8474 ^ n8473 ;
  assign n8476 = n8466 & n8475 ;
  assign n8477 = n8476 ^ n8465 ;
  assign n8478 = n8477 ^ n8160 ;
  assign n8479 = ~n8167 & n8478 ;
  assign n8480 = n8479 ^ n8160 ;
  assign n8155 = ~n3509 & n8150 ;
  assign n8156 = n8155 ^ n8144 ;
  assign n8157 = ~n368 & n8156 ;
  assign n8158 = n8157 ^ x8 ;
  assign n8116 = n7840 ^ n7822 ;
  assign n8117 = ~n7843 & ~n8116 ;
  assign n8118 = n8117 ^ n7840 ;
  assign n8114 = n3840 & n20240 ;
  assign n8111 = ~n3505 & n7151 ;
  assign n8109 = ~n408 & n7142 ;
  assign n8107 = n7526 ^ n7321 ;
  assign n8108 = n8107 ^ x11 ;
  assign n8110 = n8109 ^ n8108 ;
  assign n8112 = n8111 ^ n8110 ;
  assign n8106 = ~n540 & n7148 ;
  assign n8113 = n8112 ^ n8106 ;
  assign n8115 = n8114 ^ n8113 ;
  assign n8119 = n8118 ^ n8115 ;
  assign n8129 = n8119 ^ n7844 ;
  assign n8128 = n8127 ^ n8119 ;
  assign n8130 = n8129 ^ n8128 ;
  assign n8131 = ~n8105 & ~n8130 ;
  assign n8132 = n8131 ^ n8129 ;
  assign n8159 = n8158 ^ n8132 ;
  assign n8481 = n8480 ^ n8159 ;
  assign n8512 = ~n4892 & n6163 ;
  assign n8509 = ~n1541 & n6148 ;
  assign n8507 = ~n1972 & n6143 ;
  assign n8505 = n8439 ^ n8224 ;
  assign n8506 = n8505 ^ x17 ;
  assign n8508 = n8507 ^ n8506 ;
  assign n8510 = n8509 ^ n8508 ;
  assign n8504 = ~n1897 & n20437 ;
  assign n8511 = n8510 ^ n8504 ;
  assign n8513 = n8512 ^ n8511 ;
  assign n8523 = n5824 & n6163 ;
  assign n8520 = ~n2199 & n20437 ;
  assign n8518 = ~n2095 & n6143 ;
  assign n8516 = n8424 ^ n8235 ;
  assign n8517 = n8516 ^ x17 ;
  assign n8519 = n8518 ^ n8517 ;
  assign n8521 = n8520 ^ n8519 ;
  assign n8515 = ~n1897 & n6148 ;
  assign n8522 = n8521 ^ n8515 ;
  assign n8524 = n8523 ^ n8522 ;
  assign n8748 = n8409 ^ n8236 ;
  assign n8536 = n6163 & n6212 ;
  assign n8533 = ~n2657 & n20437 ;
  assign n8531 = ~n2552 & n6148 ;
  assign n8529 = n8368 ^ n8357 ;
  assign n8530 = n8529 ^ x17 ;
  assign n8532 = n8531 ^ n8530 ;
  assign n8534 = n8533 ^ n8532 ;
  assign n8528 = ~n2589 & n6143 ;
  assign n8535 = n8534 ^ n8528 ;
  assign n8537 = n8536 ^ n8535 ;
  assign n8679 = n8342 ^ n8257 ;
  assign n8654 = n8336 ^ n8278 ;
  assign n8548 = n6163 & ~n6695 ;
  assign n8546 = ~n3248 & n20437 ;
  assign n8543 = ~n2935 & n6143 ;
  assign n8542 = ~n2839 & n6148 ;
  assign n8544 = n8543 ^ n8542 ;
  assign n8545 = n8544 ^ x17 ;
  assign n8547 = n8546 ^ n8545 ;
  assign n8549 = n8548 ^ n8547 ;
  assign n8541 = n8330 ^ n8300 ;
  assign n8550 = n8549 ^ n8541 ;
  assign n8559 = n6163 & n6736 ;
  assign n8557 = ~n3248 & n6143 ;
  assign n8554 = ~n3022 & n20437 ;
  assign n8553 = ~n2935 & n6148 ;
  assign n8555 = n8554 ^ n8553 ;
  assign n8556 = n8555 ^ x17 ;
  assign n8558 = n8557 ^ n8556 ;
  assign n8560 = n8559 ^ n8558 ;
  assign n8551 = n8319 ^ n8301 ;
  assign n8552 = n8551 ^ n8328 ;
  assign n8561 = n8560 ^ n8552 ;
  assign n8615 = n6163 & n6753 ;
  assign n8613 = ~n3022 & n6143 ;
  assign n8610 = ~n3248 & n6148 ;
  assign n8609 = ~n3055 & n20437 ;
  assign n8611 = n8610 ^ n8609 ;
  assign n8612 = n8611 ^ x17 ;
  assign n8614 = n8613 ^ n8612 ;
  assign n8616 = n8615 ^ n8614 ;
  assign n8572 = n6163 & n6840 ;
  assign n8570 = ~n3055 & n6143 ;
  assign n8567 = ~n3022 & n6148 ;
  assign n8566 = ~n3196 & n20437 ;
  assign n8568 = n8567 ^ n8566 ;
  assign n8569 = n8568 ^ x17 ;
  assign n8571 = n8570 ^ n8569 ;
  assign n8573 = n8572 ^ n8571 ;
  assign n8563 = n5213 ^ x19 ;
  assign n8564 = ~n3429 & n8563 ;
  assign n8562 = ~n3124 & n5215 ;
  assign n8565 = n8564 ^ n8562 ;
  assign n8574 = n8573 ^ n8565 ;
  assign n8575 = ~n3429 & n5215 ;
  assign n8576 = ~n3124 & n6141 ;
  assign n8577 = x17 & ~n8576 ;
  assign n8578 = n6154 & n8577 ;
  assign n8579 = ~n3429 & n8578 ;
  assign n8580 = n8579 ^ n8577 ;
  assign n8591 = ~n3429 & n20437 ;
  assign n8588 = n3429 & n6163 ;
  assign n8589 = n8588 ^ n6143 ;
  assign n8590 = ~n3124 & n8589 ;
  assign n8592 = n8591 ^ n8590 ;
  assign n8583 = ~n3196 & n6141 ;
  assign n8593 = n8592 ^ n8583 ;
  assign n8594 = n8580 & ~n8593 ;
  assign n8595 = ~n8575 & ~n8594 ;
  assign n8602 = n6163 & n6864 ;
  assign n8600 = ~n3124 & n20437 ;
  assign n8597 = ~n3196 & n6143 ;
  assign n8596 = ~n3055 & n6148 ;
  assign n8598 = n8597 ^ n8596 ;
  assign n8599 = n8598 ^ x17 ;
  assign n8601 = n8600 ^ n8599 ;
  assign n8603 = n8602 ^ n8601 ;
  assign n8604 = n8595 & n8603 ;
  assign n8605 = n8604 ^ n8603 ;
  assign n8606 = n8605 ^ n8565 ;
  assign n8607 = n8574 & ~n8606 ;
  assign n8608 = n8607 ^ n8573 ;
  assign n8617 = n8616 ^ n8608 ;
  assign n8630 = n8616 ^ n8314 ;
  assign n8619 = n5226 ^ x19 ;
  assign n8618 = ~x19 & ~n5214 ;
  assign n8620 = n8619 ^ n8618 ;
  assign n8631 = n8630 ^ n8620 ;
  assign n8627 = n5221 & n7688 ;
  assign n8628 = n8627 ^ n5426 ;
  assign n8629 = ~n3124 & n8628 ;
  assign n8632 = n8631 ^ n8629 ;
  assign n8621 = n3429 & ~n8562 ;
  assign n8622 = ~n8620 & n8621 ;
  assign n8633 = n8632 ^ n8622 ;
  assign n8634 = n8617 & ~n8633 ;
  assign n8635 = n8634 ^ n8616 ;
  assign n8636 = n8635 ^ n8560 ;
  assign n8637 = n8561 & n8636 ;
  assign n8638 = n8637 ^ n8560 ;
  assign n8639 = n8638 ^ n8549 ;
  assign n8640 = n8550 & n8639 ;
  assign n8641 = n8640 ^ n8549 ;
  assign n8540 = n8333 ^ n8288 ;
  assign n8642 = n8641 ^ n8540 ;
  assign n8650 = n6163 & ~n6302 ;
  assign n8646 = n8540 ^ x17 ;
  assign n8645 = ~n2748 & n6148 ;
  assign n8647 = n8646 ^ n8645 ;
  assign n8644 = ~n2839 & n6143 ;
  assign n8648 = n8647 ^ n8644 ;
  assign n8643 = ~n2935 & n20437 ;
  assign n8649 = n8648 ^ n8643 ;
  assign n8651 = n8650 ^ n8649 ;
  assign n8652 = n8642 & ~n8651 ;
  assign n8653 = n8652 ^ n8641 ;
  assign n8655 = n8654 ^ n8653 ;
  assign n8663 = n6163 & n7354 ;
  assign n8659 = n8654 ^ x17 ;
  assign n8658 = ~n3324 & n6148 ;
  assign n8660 = n8659 ^ n8658 ;
  assign n8657 = ~n2839 & n20437 ;
  assign n8661 = n8660 ^ n8657 ;
  assign n8656 = ~n2748 & n6143 ;
  assign n8662 = n8661 ^ n8656 ;
  assign n8664 = n8663 ^ n8662 ;
  assign n8665 = n8655 & n8664 ;
  assign n8666 = n8665 ^ n8654 ;
  assign n8539 = n8339 ^ n8267 ;
  assign n8667 = n8666 ^ n8539 ;
  assign n8675 = n6163 & n6623 ;
  assign n8671 = n8539 ^ x17 ;
  assign n8670 = ~n3324 & n6143 ;
  assign n8672 = n8671 ^ n8670 ;
  assign n8669 = ~n2712 & n6148 ;
  assign n8673 = n8672 ^ n8669 ;
  assign n8668 = ~n2748 & n20437 ;
  assign n8674 = n8673 ^ n8668 ;
  assign n8676 = n8675 ^ n8674 ;
  assign n8677 = n8667 & ~n8676 ;
  assign n8678 = n8677 ^ n8666 ;
  assign n8680 = n8679 ^ n8678 ;
  assign n8688 = n6163 & n6229 ;
  assign n8684 = n8679 ^ x17 ;
  assign n8683 = ~n3324 & n20437 ;
  assign n8685 = n8684 ^ n8683 ;
  assign n8682 = ~n2657 & n6148 ;
  assign n8686 = n8685 ^ n8682 ;
  assign n8681 = ~n2712 & n6143 ;
  assign n8687 = n8686 ^ n8681 ;
  assign n8689 = n8688 ^ n8687 ;
  assign n8690 = ~n8680 & ~n8689 ;
  assign n8691 = n8690 ^ n8679 ;
  assign n8538 = n8355 ^ n8345 ;
  assign n8692 = n8691 ^ n8538 ;
  assign n8700 = n6079 & n6163 ;
  assign n8696 = n8538 ^ x17 ;
  assign n8695 = ~n2712 & n20437 ;
  assign n8697 = n8696 ^ n8695 ;
  assign n8694 = ~n2589 & n6148 ;
  assign n8698 = n8697 ^ n8694 ;
  assign n8693 = ~n2657 & n6143 ;
  assign n8699 = n8698 ^ n8693 ;
  assign n8701 = n8700 ^ n8699 ;
  assign n8702 = ~n8692 & ~n8701 ;
  assign n8703 = n8702 ^ n8691 ;
  assign n8704 = n8703 ^ n8529 ;
  assign n8705 = n8537 & ~n8704 ;
  assign n8706 = n8705 ^ n8529 ;
  assign n8527 = n8380 ^ n8370 ;
  assign n8707 = n8706 ^ n8527 ;
  assign n8715 = n6008 & n6163 ;
  assign n8711 = n8527 ^ x17 ;
  assign n8710 = ~n2467 & n6148 ;
  assign n8712 = n8711 ^ n8710 ;
  assign n8709 = ~n2589 & n20437 ;
  assign n8713 = n8712 ^ n8709 ;
  assign n8708 = ~n2552 & n6143 ;
  assign n8714 = n8713 ^ n8708 ;
  assign n8716 = n8715 ^ n8714 ;
  assign n8717 = n8707 & ~n8716 ;
  assign n8718 = n8717 ^ n8706 ;
  assign n8526 = n8393 ^ n8382 ;
  assign n8720 = n8718 ^ n8526 ;
  assign n8719 = ~n8526 & ~n8718 ;
  assign n8721 = n8720 ^ n8719 ;
  assign n8727 = n5696 & n6163 ;
  assign n8724 = ~n2552 & n20437 ;
  assign n8723 = ~n2371 & n6148 ;
  assign n8725 = n8724 ^ n8723 ;
  assign n8722 = ~n2467 & n6143 ;
  assign n8726 = n8725 ^ n8722 ;
  assign n8728 = n8727 ^ n8726 ;
  assign n8729 = n8728 ^ x17 ;
  assign n8738 = n8406 ^ n8395 ;
  assign n8735 = n6163 & n6449 ;
  assign n8732 = ~n2288 & n6148 ;
  assign n8731 = ~n2371 & n6143 ;
  assign n8733 = n8732 ^ n8731 ;
  assign n8730 = ~n2467 & n20437 ;
  assign n8734 = n8733 ^ n8730 ;
  assign n8736 = n8735 ^ n8734 ;
  assign n8737 = n8736 ^ n8728 ;
  assign n8739 = n8738 ^ n8737 ;
  assign n8740 = ~n8729 & n8739 ;
  assign n8741 = n8721 & n8740 ;
  assign n8742 = n8738 ^ n8719 ;
  assign n8743 = n8736 ^ x17 ;
  assign n8744 = n8743 ^ n8719 ;
  assign n8745 = ~n8742 & ~n8744 ;
  assign n8746 = n8745 ^ n8719 ;
  assign n8747 = ~n8741 & ~n8746 ;
  assign n8749 = n8748 ^ n8747 ;
  assign n8757 = n5480 & n6163 ;
  assign n8753 = n8748 ^ x17 ;
  assign n8752 = ~n2199 & n6148 ;
  assign n8754 = n8753 ^ n8752 ;
  assign n8751 = ~n2288 & n6143 ;
  assign n8755 = n8754 ^ n8751 ;
  assign n8750 = ~n2371 & n20437 ;
  assign n8756 = n8755 ^ n8750 ;
  assign n8758 = n8757 ^ n8756 ;
  assign n8759 = n8749 & n8758 ;
  assign n8760 = n8759 ^ n8748 ;
  assign n8525 = n8422 ^ n8411 ;
  assign n8761 = n8760 ^ n8525 ;
  assign n8769 = n5760 & n6163 ;
  assign n8765 = n8525 ^ x17 ;
  assign n8764 = ~n2095 & n6148 ;
  assign n8766 = n8765 ^ n8764 ;
  assign n8763 = ~n2288 & n20437 ;
  assign n8767 = n8766 ^ n8763 ;
  assign n8762 = ~n2199 & n6143 ;
  assign n8768 = n8767 ^ n8762 ;
  assign n8770 = n8769 ^ n8768 ;
  assign n8771 = ~n8761 & n8770 ;
  assign n8772 = n8771 ^ n8760 ;
  assign n8773 = n8772 ^ n8516 ;
  assign n8774 = n8524 & n8773 ;
  assign n8775 = n8774 ^ n8516 ;
  assign n8514 = n8437 ^ n8427 ;
  assign n8776 = n8775 ^ n8514 ;
  assign n8784 = ~n5287 & n6163 ;
  assign n8780 = n8514 ^ x17 ;
  assign n8779 = ~n2095 & n20437 ;
  assign n8781 = n8780 ^ n8779 ;
  assign n8778 = ~n1972 & n6148 ;
  assign n8782 = n8781 ^ n8778 ;
  assign n8777 = ~n1897 & n6143 ;
  assign n8783 = n8782 ^ n8777 ;
  assign n8785 = n8784 ^ n8783 ;
  assign n8786 = ~n8776 & n8785 ;
  assign n8787 = n8786 ^ n8775 ;
  assign n8788 = n8787 ^ n8505 ;
  assign n8789 = ~n8513 & ~n8788 ;
  assign n8790 = n8789 ^ n8505 ;
  assign n8503 = n8454 ^ n8442 ;
  assign n8791 = n8790 ^ n8503 ;
  assign n8799 = ~n5154 & n6163 ;
  assign n8795 = n8503 ^ x17 ;
  assign n8794 = ~n1819 & n6148 ;
  assign n8796 = n8795 ^ n8794 ;
  assign n8793 = ~n1541 & n6143 ;
  assign n8797 = n8796 ^ n8793 ;
  assign n8792 = ~n1972 & n20437 ;
  assign n8798 = n8797 ^ n8792 ;
  assign n8800 = n8799 ^ n8798 ;
  assign n8801 = ~n8791 & ~n8800 ;
  assign n8802 = n8801 ^ n8790 ;
  assign n8500 = n8456 ^ n8213 ;
  assign n8490 = ~n1450 & ~n6529 ;
  assign n8489 = ~n1751 & ~n6547 ;
  assign n8491 = n8490 ^ n8489 ;
  assign n8499 = n8491 ^ x14 ;
  assign n8501 = n8500 ^ n8499 ;
  assign n8492 = n8491 ^ n1345 ;
  assign n8487 = n7310 ^ n1345 ;
  assign n8493 = n8492 ^ n8487 ;
  assign n8496 = n3483 & n8493 ;
  assign n8497 = n8496 ^ n8487 ;
  assign n8498 = n6391 & ~n8497 ;
  assign n8502 = n8501 ^ n8498 ;
  assign n8848 = n8802 ^ n8502 ;
  assign n8824 = ~n1248 & n7142 ;
  assign n8823 = ~n990 & n7148 ;
  assign n8825 = n8824 ^ n8823 ;
  assign n8826 = n8825 ^ n7149 ;
  assign n8827 = n8826 ^ x11 ;
  assign n8828 = n8825 ^ x11 ;
  assign n8835 = n4335 & n8828 ;
  assign n8829 = n8828 ^ n7150 ;
  assign n8836 = n8835 ^ n8829 ;
  assign n8830 = n8829 ^ n1119 ;
  assign n8831 = n8830 ^ x10 ;
  assign n8832 = n8831 ^ n8828 ;
  assign n8839 = n8832 ^ n8830 ;
  assign n8840 = n4335 & n8839 ;
  assign n8841 = n8840 ^ n8830 ;
  assign n8842 = ~n8829 & ~n8841 ;
  assign n8843 = ~n8836 & n8842 ;
  assign n8844 = n8843 ^ n8840 ;
  assign n8845 = n8844 ^ n7150 ;
  assign n8846 = n8845 ^ n8830 ;
  assign n8847 = ~n8827 & n8846 ;
  assign n8849 = n8848 ^ n8847 ;
  assign n9396 = n8800 ^ n8790 ;
  assign n8872 = n8787 ^ n8513 ;
  assign n8851 = ~n1670 & ~n6529 ;
  assign n8850 = ~n1819 & ~n6547 ;
  assign n8852 = n8851 ^ n8850 ;
  assign n8853 = n8852 ^ n6537 ;
  assign n8854 = n8853 ^ x14 ;
  assign n8863 = n8852 ^ x14 ;
  assign n8866 = ~x13 & ~n4492 ;
  assign n8867 = n8866 ^ n1751 ;
  assign n8868 = ~n8863 & n8867 ;
  assign n8869 = n8868 ^ n1751 ;
  assign n8855 = n6404 ^ x13 ;
  assign n8856 = n8855 ^ n6547 ;
  assign n8857 = n4690 ^ n4492 ;
  assign n8860 = ~n6539 & ~n8857 ;
  assign n8861 = n8860 ^ n4690 ;
  assign n8862 = n8856 & n8861 ;
  assign n8870 = n8869 ^ n8862 ;
  assign n8871 = ~n8854 & ~n8870 ;
  assign n8873 = n8872 ^ n8871 ;
  assign n8893 = n8785 ^ n8775 ;
  assign n8880 = ~n1819 & ~n6529 ;
  assign n8879 = ~n1541 & ~n6547 ;
  assign n8881 = n8880 ^ n8879 ;
  assign n8876 = x13 & ~n4985 ;
  assign n8877 = n8876 ^ n1670 ;
  assign n8878 = n6391 & ~n8877 ;
  assign n8882 = n8881 ^ n8878 ;
  assign n8883 = ~x14 & n8882 ;
  assign n8886 = n4986 ^ x13 ;
  assign n8887 = n8886 ^ n4986 ;
  assign n8888 = ~n4985 & n8887 ;
  assign n8889 = n8888 ^ n4986 ;
  assign n8890 = n6537 & n8889 ;
  assign n8884 = n8881 ^ x14 ;
  assign n8891 = n8890 ^ n8884 ;
  assign n8892 = ~n8883 & ~n8891 ;
  assign n8894 = n8893 ^ n8892 ;
  assign n8902 = ~n1897 & ~n6547 ;
  assign n8901 = ~n1972 & ~n6529 ;
  assign n8903 = n8902 ^ n8901 ;
  assign n8898 = ~x13 & n4891 ;
  assign n8899 = n8898 ^ n1541 ;
  assign n8900 = n6391 & ~n8899 ;
  assign n8904 = n8903 ^ n8900 ;
  assign n8905 = x14 & n8904 ;
  assign n8911 = ~n1541 & n7035 ;
  assign n8906 = n8903 ^ x14 ;
  assign n8912 = n8911 ^ n8906 ;
  assign n8913 = ~n8905 & ~n8912 ;
  assign n8917 = ~n4892 & n7047 ;
  assign n8918 = n8913 & n8917 ;
  assign n8914 = n8770 ^ n8760 ;
  assign n8915 = n8914 ^ n8905 ;
  assign n8916 = n8915 ^ n8913 ;
  assign n8919 = n8918 ^ n8916 ;
  assign n9357 = n8758 ^ n8747 ;
  assign n8930 = ~n2199 & ~n6529 ;
  assign n8929 = ~n2288 & ~n6547 ;
  assign n8931 = n8930 ^ n8929 ;
  assign n8926 = x13 & ~n5759 ;
  assign n8927 = n8926 ^ n2095 ;
  assign n8928 = n6391 & ~n8927 ;
  assign n8932 = n8931 ^ n8928 ;
  assign n8933 = ~x14 & n8932 ;
  assign n8939 = ~n2095 & n7575 ;
  assign n8934 = n8931 ^ x14 ;
  assign n8940 = n8939 ^ n8934 ;
  assign n8941 = ~n8933 & n8940 ;
  assign n8945 = n5760 & n6528 ;
  assign n8946 = n8941 & n8945 ;
  assign n8942 = n8729 ^ n8720 ;
  assign n8943 = n8942 ^ n8933 ;
  assign n8944 = n8943 ^ n8941 ;
  assign n8947 = n8946 ^ n8944 ;
  assign n8955 = ~n2288 & ~n6529 ;
  assign n8954 = ~n2371 & ~n6547 ;
  assign n8956 = n8955 ^ n8954 ;
  assign n8951 = x13 & ~n5479 ;
  assign n8952 = n8951 ^ n2199 ;
  assign n8953 = n6391 & ~n8952 ;
  assign n8957 = n8956 ^ n8953 ;
  assign n8958 = ~x14 & n8957 ;
  assign n8964 = ~n2199 & n7575 ;
  assign n8959 = n8956 ^ x14 ;
  assign n8965 = n8964 ^ n8959 ;
  assign n8966 = ~n8958 & n8965 ;
  assign n8970 = n5480 & n6528 ;
  assign n8971 = n8966 & n8970 ;
  assign n8967 = n8716 ^ n8706 ;
  assign n8968 = n8967 ^ n8958 ;
  assign n8969 = n8968 ^ n8966 ;
  assign n8972 = n8971 ^ n8969 ;
  assign n9303 = n8703 ^ n8537 ;
  assign n8977 = ~n2552 & ~n6529 ;
  assign n8976 = ~n2589 & ~n6547 ;
  assign n8978 = n8977 ^ n8976 ;
  assign n8987 = n8978 ^ x14 ;
  assign n8986 = n8689 ^ n8678 ;
  assign n8988 = n8987 ^ n8986 ;
  assign n8979 = n8978 ^ n2467 ;
  assign n8974 = n7310 ^ n2467 ;
  assign n8980 = n8979 ^ n8974 ;
  assign n8983 = n6007 & n8980 ;
  assign n8984 = n8983 ^ n8974 ;
  assign n8985 = n6391 & ~n8984 ;
  assign n8989 = n8988 ^ n8985 ;
  assign n8997 = ~n2589 & ~n6529 ;
  assign n8996 = ~n2657 & ~n6547 ;
  assign n8998 = n8997 ^ n8996 ;
  assign n8993 = ~x13 & ~n6211 ;
  assign n8994 = n8993 ^ n2552 ;
  assign n8995 = n6391 & ~n8994 ;
  assign n8999 = n8998 ^ n8995 ;
  assign n9000 = x14 & n8999 ;
  assign n9006 = ~n2552 & n7035 ;
  assign n9001 = n8998 ^ x14 ;
  assign n9007 = n9006 ^ n9001 ;
  assign n9008 = ~n9000 & ~n9007 ;
  assign n9012 = n6212 & n7047 ;
  assign n9013 = n9008 & n9012 ;
  assign n9009 = n8676 ^ n8666 ;
  assign n9010 = n9009 ^ n9000 ;
  assign n9011 = n9010 ^ n9008 ;
  assign n9014 = n9013 ^ n9011 ;
  assign n9021 = ~n2712 & ~n6547 ;
  assign n9020 = ~n2657 & ~n6529 ;
  assign n9022 = n9021 ^ n9020 ;
  assign n9017 = x13 & ~n6078 ;
  assign n9018 = n9017 ^ n2589 ;
  assign n9019 = n6391 & ~n9018 ;
  assign n9023 = n9022 ^ n9019 ;
  assign n9024 = ~x14 & n9023 ;
  assign n9030 = ~n2589 & n7575 ;
  assign n9025 = n9022 ^ x14 ;
  assign n9031 = n9030 ^ n9025 ;
  assign n9032 = ~n9024 & n9031 ;
  assign n9036 = n6079 & n6528 ;
  assign n9037 = n9032 & n9036 ;
  assign n9033 = n8664 ^ n8653 ;
  assign n9034 = n9033 ^ n9024 ;
  assign n9035 = n9034 ^ n9032 ;
  assign n9038 = n9037 ^ n9035 ;
  assign n9040 = ~n3324 & ~n6547 ;
  assign n9039 = ~n2712 & ~n6529 ;
  assign n9041 = n9040 ^ n9039 ;
  assign n9054 = n9041 ^ x14 ;
  assign n9053 = n8651 ^ n8641 ;
  assign n9055 = n9054 ^ n9053 ;
  assign n17173 = n6539 ^ x13 ;
  assign n9042 = n9041 ^ n7310 ;
  assign n9044 = n17173 ^ n9042 ;
  assign n9045 = n7310 ^ n2657 ;
  assign n9046 = n9045 ^ n9041 ;
  assign n9047 = n17173 ^ n9046 ;
  assign n9048 = ~n9044 & n9047 ;
  assign n9049 = n17173 ^ n9048 ;
  assign n9050 = n6228 & ~n9049 ;
  assign n9051 = n9050 ^ n9045 ;
  assign n9052 = n6391 & ~n9051 ;
  assign n9056 = n9055 ^ n9052 ;
  assign n9260 = n8638 ^ n8550 ;
  assign n9059 = ~n2748 & ~n6529 ;
  assign n9058 = ~n2839 & ~n6547 ;
  assign n9060 = n9059 ^ n9058 ;
  assign n9061 = n9060 ^ n6537 ;
  assign n9062 = n9061 ^ x14 ;
  assign n9075 = x13 & ~n7354 ;
  assign n9074 = ~n3324 & n8856 ;
  assign n9076 = n9075 ^ n9074 ;
  assign n9077 = ~n6539 & n9076 ;
  assign n9063 = n9060 ^ x14 ;
  assign n9070 = ~x13 & ~n6643 ;
  assign n9071 = n9070 ^ n3324 ;
  assign n9072 = ~n9063 & n9071 ;
  assign n9067 = n8856 ^ n6643 ;
  assign n9073 = n9072 ^ n9067 ;
  assign n9078 = n9077 ^ n9073 ;
  assign n9079 = ~n9062 & n9078 ;
  assign n9057 = n8635 ^ n8561 ;
  assign n9080 = n9079 ^ n9057 ;
  assign n9104 = n8633 ^ n8608 ;
  assign n9088 = ~n2935 & ~n6547 ;
  assign n9087 = ~n2839 & ~n6529 ;
  assign n9089 = n9088 ^ n9087 ;
  assign n9084 = ~x13 & n6301 ;
  assign n9085 = n9084 ^ n2748 ;
  assign n9086 = n6391 & ~n9085 ;
  assign n9090 = n9089 ^ n9086 ;
  assign n9091 = x14 & n9090 ;
  assign n9097 = ~n2748 & n7035 ;
  assign n9092 = n9089 ^ x14 ;
  assign n9098 = n9097 ^ n9092 ;
  assign n9099 = ~n9091 & ~n9098 ;
  assign n9101 = ~n6302 & n7047 ;
  assign n9102 = n9099 & n9101 ;
  assign n9100 = n9099 ^ n9091 ;
  assign n9103 = n9102 ^ n9100 ;
  assign n9105 = n9104 ^ n9103 ;
  assign n9109 = ~n3248 & ~n6547 ;
  assign n9108 = ~n2935 & ~n6529 ;
  assign n9110 = n9109 ^ n9108 ;
  assign n9115 = ~x14 & ~n2839 ;
  assign n9111 = n7310 ^ n2839 ;
  assign n9116 = n9115 ^ n9111 ;
  assign n9117 = ~n3439 & ~n9116 ;
  assign n9118 = n9117 ^ n9111 ;
  assign n9119 = n6391 & ~n9118 ;
  assign n9120 = ~n9110 & ~n9119 ;
  assign n9121 = n9120 ^ x14 ;
  assign n9107 = n3440 & n6537 ;
  assign n9122 = n9121 ^ n9107 ;
  assign n9106 = n8605 ^ n8574 ;
  assign n9123 = n9122 ^ n9106 ;
  assign n9147 = n8594 ^ n8575 ;
  assign n9148 = n9147 ^ n8603 ;
  assign n9131 = ~n3022 & ~n6547 ;
  assign n9130 = ~n3248 & ~n6529 ;
  assign n9132 = n9131 ^ n9130 ;
  assign n9127 = x13 & ~n3437 ;
  assign n9128 = n9127 ^ n2935 ;
  assign n9129 = n6391 & ~n9128 ;
  assign n9133 = n9132 ^ n9129 ;
  assign n9134 = ~x14 & n9133 ;
  assign n9140 = ~n2935 & n7575 ;
  assign n9135 = n9132 ^ x14 ;
  assign n9141 = n9140 ^ n9135 ;
  assign n9142 = ~n9134 & n9141 ;
  assign n9144 = n6528 & n6736 ;
  assign n9145 = n9142 & n9144 ;
  assign n9143 = n9142 ^ n9134 ;
  assign n9146 = n9145 ^ n9143 ;
  assign n9149 = n9148 ^ n9146 ;
  assign n8581 = n8580 ^ x17 ;
  assign n9172 = n8593 ^ n8581 ;
  assign n9156 = ~n3022 & ~n6529 ;
  assign n9155 = ~n3055 & ~n6547 ;
  assign n9157 = n9156 ^ n9155 ;
  assign n9152 = x13 & ~n6749 ;
  assign n9153 = n9152 ^ n3248 ;
  assign n9154 = n6391 & ~n9153 ;
  assign n9158 = n9157 ^ n9154 ;
  assign n9159 = ~x14 & n9158 ;
  assign n9165 = ~n3248 & n7575 ;
  assign n9160 = n9157 ^ x14 ;
  assign n9166 = n9165 ^ n9160 ;
  assign n9167 = ~n9159 & n9166 ;
  assign n9169 = n6528 & n6753 ;
  assign n9170 = n9167 & n9169 ;
  assign n9168 = n9167 ^ n9159 ;
  assign n9171 = n9170 ^ n9168 ;
  assign n9173 = n9172 ^ n9171 ;
  assign n9183 = ~n3196 & ~n6529 ;
  assign n9182 = ~n3124 & ~n6547 ;
  assign n9184 = n9183 ^ n9182 ;
  assign n9179 = ~x13 & ~n6863 ;
  assign n9180 = n9179 ^ n3055 ;
  assign n9181 = n6391 & ~n9180 ;
  assign n9185 = n9184 ^ n9181 ;
  assign n9186 = x14 & n9185 ;
  assign n9192 = ~n3055 & n7035 ;
  assign n9187 = n9184 ^ x14 ;
  assign n9193 = n9192 ^ n9187 ;
  assign n9194 = ~n9186 & ~n9193 ;
  assign n9196 = n6864 & n7047 ;
  assign n9197 = n9194 & n9196 ;
  assign n9195 = n9194 ^ n9186 ;
  assign n9198 = n9197 ^ n9195 ;
  assign n9199 = ~n3429 & n6141 ;
  assign n9200 = n6391 ^ n3429 ;
  assign n9202 = ~n3124 & n6391 ;
  assign n9201 = n6532 ^ n3429 ;
  assign n9203 = n9202 ^ n9201 ;
  assign n9204 = n9203 ^ n3429 ;
  assign n9205 = ~n9200 & n9204 ;
  assign n9206 = n9205 ^ n3429 ;
  assign n9207 = x14 & ~n9206 ;
  assign n9208 = n9207 ^ x14 ;
  assign n9215 = ~n3429 & ~n6547 ;
  assign n9214 = ~n3124 & ~n6529 ;
  assign n9216 = n9215 ^ n9214 ;
  assign n9211 = n3431 & n7310 ;
  assign n9212 = n9211 ^ n3196 ;
  assign n9213 = n6391 & ~n9212 ;
  assign n9217 = n9216 ^ n9213 ;
  assign n9218 = n9208 & ~n9217 ;
  assign n9219 = ~n9199 & ~n9218 ;
  assign n9220 = ~n9198 & n9219 ;
  assign n9221 = n9220 ^ n9198 ;
  assign n6140 = n6139 ^ x16 ;
  assign n9174 = ~n3429 & n6140 ;
  assign n9175 = n9174 ^ n8576 ;
  assign n9222 = n9221 ^ n9175 ;
  assign n9237 = ~n3022 & n6391 ;
  assign n9233 = ~n3196 & ~n6547 ;
  assign n9232 = ~n3055 & ~n6529 ;
  assign n9234 = n9233 ^ n9232 ;
  assign n9239 = n6839 & ~n9234 ;
  assign n9240 = n9237 & n9239 ;
  assign n9241 = x14 & ~n9240 ;
  assign n9227 = ~x14 & ~n3022 ;
  assign n9223 = n7310 ^ n3022 ;
  assign n9228 = n9227 ^ n9223 ;
  assign n9229 = n6839 & ~n9228 ;
  assign n9230 = n9229 ^ n9223 ;
  assign n9231 = n6391 & ~n9230 ;
  assign n9235 = n9234 ^ n9231 ;
  assign n9236 = n9235 ^ n9221 ;
  assign n9242 = n9241 ^ n9236 ;
  assign n9243 = ~n9222 & ~n9242 ;
  assign n9244 = n9243 ^ n9221 ;
  assign n9245 = n9244 ^ n9171 ;
  assign n9246 = n9173 & n9245 ;
  assign n9247 = n9246 ^ n9172 ;
  assign n9248 = n9247 ^ n9146 ;
  assign n9249 = n9149 & n9248 ;
  assign n9250 = n9249 ^ n9146 ;
  assign n9251 = n9250 ^ n9122 ;
  assign n9252 = ~n9123 & ~n9251 ;
  assign n9253 = n9252 ^ n9122 ;
  assign n9254 = n9253 ^ n9103 ;
  assign n9255 = n9105 & n9254 ;
  assign n9256 = n9255 ^ n9103 ;
  assign n9257 = n9256 ^ n9057 ;
  assign n9258 = ~n9080 & ~n9257 ;
  assign n9259 = n9258 ^ n9057 ;
  assign n9261 = n9260 ^ n9259 ;
  assign n9270 = n9260 ^ x14 ;
  assign n9269 = ~n3324 & ~n6529 ;
  assign n9271 = n9270 ^ n9269 ;
  assign n9268 = ~n2748 & ~n6547 ;
  assign n9272 = n9271 ^ n9268 ;
  assign n9262 = n6623 ^ n2712 ;
  assign n9265 = n7310 & ~n9262 ;
  assign n9266 = n9265 ^ n2712 ;
  assign n9267 = n6391 & ~n9266 ;
  assign n9273 = n9272 ^ n9267 ;
  assign n9274 = n9261 & n9273 ;
  assign n9275 = n9274 ^ n9260 ;
  assign n9276 = n9275 ^ n9053 ;
  assign n9277 = n9056 & n9276 ;
  assign n9278 = n9277 ^ n9053 ;
  assign n9279 = n9278 ^ n9033 ;
  assign n9280 = n9038 & n9279 ;
  assign n9281 = n9280 ^ n9033 ;
  assign n9282 = n9281 ^ n9009 ;
  assign n9283 = ~n9014 & n9282 ;
  assign n9284 = n9283 ^ n9009 ;
  assign n9285 = n9284 ^ n8986 ;
  assign n9286 = ~n8989 & ~n9285 ;
  assign n9287 = n9286 ^ n8986 ;
  assign n8973 = n8701 ^ n8691 ;
  assign n9288 = n9287 ^ n8973 ;
  assign n9297 = n8973 ^ x14 ;
  assign n9296 = ~n2552 & ~n6547 ;
  assign n9298 = n9297 ^ n9296 ;
  assign n9295 = ~n2467 & ~n6529 ;
  assign n9299 = n9298 ^ n9295 ;
  assign n9292 = ~n5695 & ~n7310 ;
  assign n9293 = n9292 ^ n5696 ;
  assign n9294 = n6391 & n9293 ;
  assign n9300 = n9299 ^ n9294 ;
  assign n9301 = n9288 & n9300 ;
  assign n9302 = n9301 ^ n9287 ;
  assign n9304 = n9303 ^ n9302 ;
  assign n9306 = n2288 ^ x14 ;
  assign n9307 = n9306 ^ x13 ;
  assign n9308 = n9307 ^ x14 ;
  assign n9311 = ~n5814 & ~n9308 ;
  assign n9312 = n9311 ^ x14 ;
  assign n9313 = n6391 & n9312 ;
  assign n9314 = n9313 ^ x14 ;
  assign n9324 = n9314 ^ n9303 ;
  assign n9318 = ~n2467 & ~n6547 ;
  assign n9317 = ~n2371 & ~n6529 ;
  assign n9319 = n9318 ^ n9317 ;
  assign n9320 = ~x14 & ~n2288 ;
  assign n9321 = n5814 & n6391 ;
  assign n9322 = n9320 & n9321 ;
  assign n9323 = ~n9319 & ~n9322 ;
  assign n9325 = n9324 ^ n9323 ;
  assign n9305 = n5479 ^ n3331 ;
  assign n9315 = x14 & ~n9314 ;
  assign n9316 = ~n9305 & n9315 ;
  assign n9326 = n9325 ^ n9316 ;
  assign n9327 = n9304 & n9326 ;
  assign n9328 = n9327 ^ n9303 ;
  assign n9329 = n9328 ^ n8967 ;
  assign n9330 = n8972 & ~n9329 ;
  assign n9331 = n9330 ^ n8967 ;
  assign n9332 = n9331 ^ n8942 ;
  assign n9333 = n8947 & n9332 ;
  assign n9334 = n9333 ^ n8942 ;
  assign n8920 = n8729 ^ n8718 ;
  assign n8921 = n8729 ^ n8526 ;
  assign n8922 = n8920 & n8921 ;
  assign n8923 = n8922 ^ n8739 ;
  assign n9335 = n9334 ^ n8923 ;
  assign n9352 = x14 & n5285 ;
  assign n9353 = n6391 & n9352 ;
  assign n9347 = ~n2095 & ~n6529 ;
  assign n9346 = ~n2199 & ~n6547 ;
  assign n9348 = n9347 ^ n9346 ;
  assign n9345 = n8923 ^ x14 ;
  assign n9349 = n9348 ^ n9345 ;
  assign n9340 = ~x14 & ~n1897 ;
  assign n9336 = n7310 ^ n1897 ;
  assign n9341 = n9340 ^ n9336 ;
  assign n9342 = n4884 & ~n9341 ;
  assign n9343 = n9342 ^ n9336 ;
  assign n9344 = n6391 & ~n9343 ;
  assign n9350 = n9349 ^ n9344 ;
  assign n9354 = n9353 ^ n9350 ;
  assign n9355 = n9335 & ~n9354 ;
  assign n9356 = n9355 ^ n9334 ;
  assign n9358 = n9357 ^ n9356 ;
  assign n9366 = n9357 ^ x14 ;
  assign n9365 = ~n2095 & ~n6547 ;
  assign n9367 = n9366 ^ n9365 ;
  assign n9364 = ~n1897 & ~n6529 ;
  assign n9368 = n9367 ^ n9364 ;
  assign n9361 = n5286 & ~n7310 ;
  assign n9362 = n9361 ^ n5287 ;
  assign n9363 = n6391 & ~n9362 ;
  assign n9369 = n9368 ^ n9363 ;
  assign n9370 = n9358 & n9369 ;
  assign n9371 = n9370 ^ n9357 ;
  assign n9372 = n9371 ^ n8914 ;
  assign n9373 = n8919 & ~n9372 ;
  assign n9374 = n9373 ^ n8914 ;
  assign n8895 = n8772 ^ n8524 ;
  assign n9375 = n9374 ^ n8895 ;
  assign n9385 = ~n1972 & ~n6547 ;
  assign n9383 = ~n1541 & ~n6529 ;
  assign n9382 = n8895 ^ x14 ;
  assign n9384 = n9383 ^ n9382 ;
  assign n9386 = n9385 ^ n9384 ;
  assign n9379 = n4488 & ~n7310 ;
  assign n9380 = n9379 ^ n5154 ;
  assign n9381 = n6391 & ~n9380 ;
  assign n9387 = n9386 ^ n9381 ;
  assign n9388 = ~n9375 & ~n9387 ;
  assign n9389 = n9388 ^ n9374 ;
  assign n9390 = n9389 ^ n8893 ;
  assign n9391 = n8894 & n9390 ;
  assign n9392 = n9391 ^ n8893 ;
  assign n9393 = n9392 ^ n8872 ;
  assign n9394 = n8873 & n9393 ;
  assign n9395 = n9394 ^ n8872 ;
  assign n9397 = n9396 ^ n9395 ;
  assign n9416 = n9396 ^ x14 ;
  assign n9401 = ~n1670 & ~n6547 ;
  assign n9400 = ~n1751 & ~n6529 ;
  assign n9402 = n9401 ^ n9400 ;
  assign n9417 = n9416 ^ n9402 ;
  assign n9413 = n1450 ^ x14 ;
  assign n9414 = n9413 ^ x13 ;
  assign n9415 = n6391 & ~n9414 ;
  assign n9418 = n9417 ^ n9415 ;
  assign n9407 = ~x14 & n9402 ;
  assign n9408 = ~n1450 & n9407 ;
  assign n9409 = n9408 ^ n1450 ;
  assign n9398 = n7310 ^ n1450 ;
  assign n9410 = n9409 ^ n9398 ;
  assign n9411 = n6391 & n9410 ;
  assign n9412 = ~n4494 & n9411 ;
  assign n9419 = n9418 ^ n9412 ;
  assign n9420 = n9397 & ~n9419 ;
  assign n9421 = n9420 ^ n9396 ;
  assign n9422 = n9421 ^ n8848 ;
  assign n9423 = ~n8849 & ~n9422 ;
  assign n9424 = n9423 ^ n8848 ;
  assign n8821 = ~n540 & n8139 ;
  assign n8814 = ~n4359 & n20240 ;
  assign n8811 = ~n856 & n7151 ;
  assign n8809 = ~n1248 & n7148 ;
  assign n8807 = n8459 ^ n8203 ;
  assign n8808 = n8807 ^ x11 ;
  assign n8810 = n8809 ^ n8808 ;
  assign n8812 = n8811 ^ n8810 ;
  assign n8806 = ~n1119 & n7142 ;
  assign n8813 = n8812 ^ n8806 ;
  assign n8815 = n8814 ^ n8813 ;
  assign n8803 = n8802 ^ n8500 ;
  assign n8804 = ~n8502 & n8803 ;
  assign n8805 = n8804 ^ n8500 ;
  assign n8816 = n8815 ^ n8805 ;
  assign n8817 = n8816 ^ x8 ;
  assign n8486 = ~n698 & n8144 ;
  assign n8818 = n8817 ^ n8486 ;
  assign n8484 = n8148 ^ x7 ;
  assign n8485 = ~n408 & n8484 ;
  assign n8819 = n8818 ^ n8485 ;
  assign n8482 = n3812 & n8150 ;
  assign n8820 = n8819 ^ n8482 ;
  assign n8822 = n8821 ^ n8820 ;
  assign n9425 = n9424 ^ n8822 ;
  assign n9434 = ~n698 & n8139 ;
  assign n9429 = n9421 ^ n8849 ;
  assign n9430 = n9429 ^ x8 ;
  assign n9428 = ~n856 & n8144 ;
  assign n9431 = n9430 ^ n9428 ;
  assign n9427 = ~n540 & n8484 ;
  assign n9432 = n9431 ^ n9427 ;
  assign n9426 = n3968 & n8150 ;
  assign n9433 = n9432 ^ n9426 ;
  assign n9435 = n9434 ^ n9433 ;
  assign n9444 = n4580 & n20240 ;
  assign n9441 = ~n990 & n7142 ;
  assign n9439 = ~n1345 & n7148 ;
  assign n9437 = n9419 ^ n9395 ;
  assign n9438 = n9437 ^ x11 ;
  assign n9440 = n9439 ^ n9438 ;
  assign n9442 = n9441 ^ n9440 ;
  assign n9436 = ~n1248 & n7151 ;
  assign n9443 = n9442 ^ n9436 ;
  assign n9445 = n9444 ^ n9443 ;
  assign n9454 = n4307 & n20240 ;
  assign n9451 = ~n990 & n7151 ;
  assign n9449 = ~n1345 & n7142 ;
  assign n9447 = n9392 ^ n8873 ;
  assign n9448 = n9447 ^ x11 ;
  assign n9450 = n9449 ^ n9448 ;
  assign n9452 = n9451 ^ n9450 ;
  assign n9446 = ~n1450 & n7148 ;
  assign n9453 = n9452 ^ n9446 ;
  assign n9455 = n9454 ^ n9453 ;
  assign n9465 = ~n4495 & n20240 ;
  assign n9462 = ~n1751 & n7142 ;
  assign n9460 = ~n1450 & n7151 ;
  assign n9458 = n9387 ^ n9374 ;
  assign n9459 = n9458 ^ x11 ;
  assign n9461 = n9460 ^ n9459 ;
  assign n9463 = n9462 ^ n9461 ;
  assign n9457 = ~n1670 & n7148 ;
  assign n9464 = n9463 ^ n9457 ;
  assign n9466 = n9465 ^ n9464 ;
  assign n9856 = n9371 ^ n8919 ;
  assign n9476 = ~n5154 & n20240 ;
  assign n9473 = ~n1541 & n7142 ;
  assign n9471 = ~n1819 & n7151 ;
  assign n9469 = n9354 ^ n9334 ;
  assign n9470 = n9469 ^ x11 ;
  assign n9472 = n9471 ^ n9470 ;
  assign n9474 = n9473 ^ n9472 ;
  assign n9468 = ~n1972 & n7148 ;
  assign n9475 = n9474 ^ n9468 ;
  assign n9477 = n9476 ^ n9475 ;
  assign n9486 = ~n4892 & n20240 ;
  assign n9483 = ~n1541 & n7151 ;
  assign n9481 = ~n1972 & n7142 ;
  assign n9479 = n9331 ^ n8947 ;
  assign n9480 = n9479 ^ x11 ;
  assign n9482 = n9481 ^ n9480 ;
  assign n9484 = n9483 ^ n9482 ;
  assign n9478 = ~n1897 & n7148 ;
  assign n9485 = n9484 ^ n9478 ;
  assign n9487 = n9486 ^ n9485 ;
  assign n9496 = ~n5287 & n20240 ;
  assign n9493 = ~n2095 & n7148 ;
  assign n9491 = ~n1897 & n7142 ;
  assign n9489 = n9328 ^ n8972 ;
  assign n9490 = n9489 ^ x11 ;
  assign n9492 = n9491 ^ n9490 ;
  assign n9494 = n9493 ^ n9492 ;
  assign n9488 = ~n1972 & n7151 ;
  assign n9495 = n9494 ^ n9488 ;
  assign n9497 = n9496 ^ n9495 ;
  assign n9509 = ~n2199 & n7142 ;
  assign n9507 = ~n2288 & n7148 ;
  assign n9505 = n9300 ^ n9287 ;
  assign n9506 = n9505 ^ x11 ;
  assign n9508 = n9507 ^ n9506 ;
  assign n9510 = n9509 ^ n9508 ;
  assign n9499 = x11 ^ x10 ;
  assign n9502 = ~n5759 & ~n9499 ;
  assign n9503 = n9502 ^ n5760 ;
  assign n9504 = n7140 & n9503 ;
  assign n9511 = n9510 ^ n9504 ;
  assign n9519 = n5480 & n20240 ;
  assign n9517 = ~n2288 & n7142 ;
  assign n9514 = ~n2199 & n7151 ;
  assign n9513 = ~n2371 & n7148 ;
  assign n9515 = n9514 ^ n9513 ;
  assign n9516 = n9515 ^ x11 ;
  assign n9518 = n9517 ^ n9516 ;
  assign n9520 = n9519 ^ n9518 ;
  assign n9512 = n9284 ^ n8989 ;
  assign n9521 = n9520 ^ n9512 ;
  assign n9529 = n9281 ^ n9014 ;
  assign n9527 = n6449 & n20240 ;
  assign n9524 = ~n2288 & n7151 ;
  assign n9523 = ~n2371 & n7142 ;
  assign n9525 = n9524 ^ n9523 ;
  assign n9522 = ~n2467 & n7148 ;
  assign n9526 = n9525 ^ n9522 ;
  assign n9528 = n9527 ^ n9526 ;
  assign n9530 = n9529 ^ n9528 ;
  assign n9791 = n5696 & n20240 ;
  assign n9788 = ~n2552 & n7148 ;
  assign n9787 = ~n2371 & n7151 ;
  assign n9789 = n9788 ^ n9787 ;
  assign n9786 = ~n2467 & n7142 ;
  assign n9790 = n9789 ^ n9786 ;
  assign n9792 = n9791 ^ n9790 ;
  assign n9805 = n9792 ^ n9528 ;
  assign n9772 = n9275 ^ n9056 ;
  assign n9539 = n6212 & n20240 ;
  assign n9537 = ~n2589 & n7142 ;
  assign n9534 = ~n2552 & n7151 ;
  assign n9533 = ~n2657 & n7148 ;
  assign n9535 = n9534 ^ n9533 ;
  assign n9536 = n9535 ^ x11 ;
  assign n9538 = n9537 ^ n9536 ;
  assign n9540 = n9539 ^ n9538 ;
  assign n9532 = n9273 ^ n9259 ;
  assign n9541 = n9540 ^ n9532 ;
  assign n9756 = n9256 ^ n9080 ;
  assign n9768 = n9756 ^ n9540 ;
  assign n9741 = n9253 ^ n9105 ;
  assign n9701 = ~n6302 & n20240 ;
  assign n9699 = ~n2839 & n7142 ;
  assign n9696 = ~n2748 & n7151 ;
  assign n9695 = ~n2935 & n7148 ;
  assign n9697 = n9696 ^ n9695 ;
  assign n9698 = n9697 ^ x11 ;
  assign n9700 = n9699 ^ n9698 ;
  assign n9702 = n9701 ^ n9700 ;
  assign n9550 = ~n6695 & n20240 ;
  assign n9548 = ~n3248 & n7148 ;
  assign n9545 = ~n2935 & n7142 ;
  assign n9544 = ~n2839 & n7151 ;
  assign n9546 = n9545 ^ n9544 ;
  assign n9547 = n9546 ^ x11 ;
  assign n9549 = n9548 ^ n9547 ;
  assign n9551 = n9550 ^ n9549 ;
  assign n9543 = n9242 ^ n9175 ;
  assign n9552 = n9551 ^ n9543 ;
  assign n9562 = n6736 & n20240 ;
  assign n9559 = ~n2935 & n7151 ;
  assign n9557 = ~n3022 & n7148 ;
  assign n9554 = n9218 ^ n9199 ;
  assign n9555 = n9554 ^ n9198 ;
  assign n9556 = n9555 ^ x11 ;
  assign n9558 = n9557 ^ n9556 ;
  assign n9560 = n9559 ^ n9558 ;
  assign n9553 = ~n3248 & n7142 ;
  assign n9561 = n9560 ^ n9553 ;
  assign n9563 = n9562 ^ n9561 ;
  assign n9571 = n6753 & n20240 ;
  assign n9569 = ~n3022 & n7142 ;
  assign n9566 = ~n3248 & n7151 ;
  assign n9565 = ~n3055 & n7148 ;
  assign n9567 = n9566 ^ n9565 ;
  assign n9568 = n9567 ^ x11 ;
  assign n9570 = n9569 ^ n9568 ;
  assign n9572 = n9571 ^ n9570 ;
  assign n9564 = n9217 ^ n9207 ;
  assign n9573 = n9572 ^ n9564 ;
  assign n9606 = n6864 & n20240 ;
  assign n9603 = ~n3196 & n7142 ;
  assign n9602 = ~n3124 & n7148 ;
  assign n9604 = n9603 ^ n9602 ;
  assign n9601 = ~n3055 & n7151 ;
  assign n9605 = n9604 ^ n9601 ;
  assign n9607 = n9606 ^ n9605 ;
  assign n9583 = x11 & ~n20255 ;
  assign n9584 = ~n3124 & n7140 ;
  assign n9585 = n3429 & ~n9584 ;
  assign n9586 = n9583 & n9585 ;
  assign n9587 = n9586 ^ n9583 ;
  assign n9588 = n9587 ^ x11 ;
  assign n9597 = ~n3429 & n7148 ;
  assign n9596 = ~n3196 & n7140 ;
  assign n9598 = n9597 ^ n9596 ;
  assign n9593 = n3429 & n20240 ;
  assign n9594 = n9593 ^ n7142 ;
  assign n9595 = ~n3124 & n9594 ;
  assign n9599 = n9598 ^ n9595 ;
  assign n9600 = n9588 & ~n9599 ;
  assign n9608 = n9607 ^ n9600 ;
  assign n9611 = n9608 ^ x11 ;
  assign n9612 = n9611 ^ n3429 ;
  assign n9672 = n9612 ^ x12 ;
  assign n9673 = n9672 ^ x11 ;
  assign n9674 = n9673 ^ n9607 ;
  assign n9676 = n9674 ^ n9672 ;
  assign n9626 = n9607 & ~n9608 ;
  assign n9627 = n9626 ^ n9611 ;
  assign n9616 = n9608 ^ x12 ;
  assign n9628 = n9627 ^ n9616 ;
  assign n9629 = n9628 ^ n9600 ;
  assign n9630 = n9616 ^ n3429 ;
  assign n9631 = n9630 ^ n9600 ;
  assign n9632 = n9629 & ~n9631 ;
  assign n9615 = n9612 ^ x11 ;
  assign n9617 = n9616 ^ n9615 ;
  assign n9633 = n9617 ^ n9612 ;
  assign n9619 = n9617 ^ n9600 ;
  assign n9634 = n9633 ^ n9619 ;
  assign n9635 = n9617 ^ n9611 ;
  assign n9636 = n9635 ^ n9619 ;
  assign n9637 = n9634 & n9636 ;
  assign n9638 = n9632 & n9637 ;
  assign n9639 = n9638 ^ n9626 ;
  assign n9640 = n9639 ^ n3429 ;
  assign n9620 = n9619 ^ n9615 ;
  assign n9669 = n9640 ^ n9620 ;
  assign n9670 = n9669 ^ n9619 ;
  assign n9613 = n9612 ^ n9608 ;
  assign n9645 = n9613 ^ x12 ;
  assign n9671 = n9670 ^ n9645 ;
  assign n9677 = n9676 ^ n9671 ;
  assign n9678 = n9677 ^ n9600 ;
  assign n9679 = n9678 ^ n9674 ;
  assign n9580 = n6840 & n20240 ;
  assign n9578 = ~n3055 & n7142 ;
  assign n9575 = ~n3022 & n7151 ;
  assign n9574 = ~n3196 & n7148 ;
  assign n9576 = n9575 ^ n9574 ;
  assign n9577 = n9576 ^ x11 ;
  assign n9579 = n9578 ^ n9577 ;
  assign n9581 = n9580 ^ n9579 ;
  assign n9680 = n9679 ^ n9581 ;
  assign n9682 = n9581 ^ n9202 ;
  assign n9681 = ~n3429 & ~n6531 ;
  assign n9683 = n9682 ^ n9681 ;
  assign n9684 = n9680 & ~n9683 ;
  assign n9685 = n9684 ^ n9679 ;
  assign n9686 = n9685 ^ n9572 ;
  assign n9687 = n9573 & n9686 ;
  assign n9688 = n9687 ^ n9572 ;
  assign n9689 = n9688 ^ n9555 ;
  assign n9690 = ~n9563 & ~n9689 ;
  assign n9691 = n9690 ^ n9555 ;
  assign n9692 = n9691 ^ n9551 ;
  assign n9693 = ~n9552 & ~n9692 ;
  assign n9694 = n9693 ^ n9551 ;
  assign n9703 = n9702 ^ n9694 ;
  assign n9704 = n9694 ^ n9173 ;
  assign n9705 = n9704 ^ n9244 ;
  assign n9706 = n9703 & n9705 ;
  assign n9707 = n9706 ^ n9702 ;
  assign n9542 = n9247 ^ n9149 ;
  assign n9709 = n9707 ^ n9542 ;
  assign n9708 = n9542 & n9707 ;
  assign n9710 = n9709 ^ n9708 ;
  assign n9716 = n7354 & n20240 ;
  assign n9713 = ~n2748 & n7142 ;
  assign n9712 = ~n3324 & n7151 ;
  assign n9714 = n9713 ^ n9712 ;
  assign n9711 = ~n2839 & n7148 ;
  assign n9715 = n9714 ^ n9711 ;
  assign n9717 = n9716 ^ n9715 ;
  assign n9718 = n9717 ^ x11 ;
  assign n9731 = n9250 ^ n9123 ;
  assign n9727 = ~n2748 & n7148 ;
  assign n9726 = ~n3324 & n7142 ;
  assign n9728 = n9727 ^ n9726 ;
  assign n9723 = ~n9262 & n9499 ;
  assign n9724 = n9723 ^ n2712 ;
  assign n9725 = n7140 & ~n9724 ;
  assign n9729 = n9728 ^ n9725 ;
  assign n9730 = n9729 ^ n9717 ;
  assign n9732 = n9731 ^ n9730 ;
  assign n9733 = n9718 & n9732 ;
  assign n9734 = n9710 & n9733 ;
  assign n9735 = n9731 ^ n9708 ;
  assign n9736 = n9729 ^ x11 ;
  assign n9737 = n9736 ^ n9708 ;
  assign n9738 = ~n9735 & n9737 ;
  assign n9739 = n9738 ^ n9708 ;
  assign n9740 = ~n9734 & ~n9739 ;
  assign n9742 = n9741 ^ n9740 ;
  assign n9751 = ~n3324 & n7148 ;
  assign n9749 = ~n2712 & n7142 ;
  assign n9748 = n9741 ^ x11 ;
  assign n9750 = n9749 ^ n9748 ;
  assign n9752 = n9751 ^ n9750 ;
  assign n9745 = ~n6228 & ~n9499 ;
  assign n9746 = n9745 ^ n6229 ;
  assign n9747 = n7140 & n9746 ;
  assign n9753 = n9752 ^ n9747 ;
  assign n9754 = n9742 & ~n9753 ;
  assign n9755 = n9754 ^ n9741 ;
  assign n9757 = n9756 ^ n9755 ;
  assign n9765 = n6079 & n20240 ;
  assign n9761 = n9756 ^ x11 ;
  assign n9760 = ~n2589 & n7151 ;
  assign n9762 = n9761 ^ n9760 ;
  assign n9759 = ~n2657 & n7142 ;
  assign n9763 = n9762 ^ n9759 ;
  assign n9758 = ~n2712 & n7148 ;
  assign n9764 = n9763 ^ n9758 ;
  assign n9766 = n9765 ^ n9764 ;
  assign n9767 = ~n9757 & n9766 ;
  assign n9769 = n9768 ^ n9767 ;
  assign n9770 = n9541 & n9769 ;
  assign n9771 = n9770 ^ n9540 ;
  assign n9773 = n9772 ^ n9771 ;
  assign n9781 = n6008 & n20240 ;
  assign n9777 = n9772 ^ x11 ;
  assign n9776 = ~n2467 & n7151 ;
  assign n9778 = n9777 ^ n9776 ;
  assign n9775 = ~n2589 & n7148 ;
  assign n9779 = n9778 ^ n9775 ;
  assign n9774 = ~n2552 & n7142 ;
  assign n9780 = n9779 ^ n9774 ;
  assign n9782 = n9781 ^ n9780 ;
  assign n9783 = n9773 & n9782 ;
  assign n9784 = n9783 ^ n9772 ;
  assign n9531 = n9278 ^ n9038 ;
  assign n9785 = n9784 ^ n9531 ;
  assign n9806 = n9805 ^ n9785 ;
  assign n9807 = n9806 ^ n9805 ;
  assign n9808 = n9792 ^ n9784 ;
  assign n9811 = ~n9807 & n9808 ;
  assign n9812 = n9811 ^ n9805 ;
  assign n9813 = ~n9530 & ~n9812 ;
  assign n9800 = n9784 ^ n9529 ;
  assign n9793 = n9792 ^ x11 ;
  assign n9794 = n9793 ^ n9792 ;
  assign n9795 = n9792 ^ n9531 ;
  assign n9796 = n9795 ^ n9792 ;
  assign n9797 = n9794 & n9796 ;
  assign n9798 = n9797 ^ n9792 ;
  assign n9799 = n9785 & n9798 ;
  assign n9801 = n9800 ^ n9799 ;
  assign n9802 = n9530 & ~n9801 ;
  assign n9815 = n9813 ^ n9802 ;
  assign n9816 = ~x11 & n9815 ;
  assign n9803 = n9802 ^ n9529 ;
  assign n9804 = n9803 ^ n9512 ;
  assign n9817 = n9816 ^ n9804 ;
  assign n9818 = ~n9521 & ~n9817 ;
  assign n9819 = n9818 ^ n9520 ;
  assign n9820 = n9819 ^ n9505 ;
  assign n9821 = n9511 & n9820 ;
  assign n9822 = n9821 ^ n9505 ;
  assign n9498 = n9326 ^ n9302 ;
  assign n9823 = n9822 ^ n9498 ;
  assign n9831 = n5824 & n20240 ;
  assign n9827 = n9498 ^ x11 ;
  assign n9826 = ~n2095 & n7142 ;
  assign n9828 = n9827 ^ n9826 ;
  assign n9825 = ~n2199 & n7148 ;
  assign n9829 = n9828 ^ n9825 ;
  assign n9824 = ~n1897 & n7151 ;
  assign n9830 = n9829 ^ n9824 ;
  assign n9832 = n9831 ^ n9830 ;
  assign n9833 = ~n9823 & n9832 ;
  assign n9834 = n9833 ^ n9822 ;
  assign n9835 = n9834 ^ n9489 ;
  assign n9836 = ~n9497 & ~n9835 ;
  assign n9837 = n9836 ^ n9489 ;
  assign n9838 = n9837 ^ n9479 ;
  assign n9839 = n9487 & ~n9838 ;
  assign n9840 = n9839 ^ n9479 ;
  assign n9841 = n9840 ^ n9469 ;
  assign n9842 = n9477 & n9841 ;
  assign n9843 = n9842 ^ n9469 ;
  assign n9467 = n9369 ^ n9356 ;
  assign n9844 = n9843 ^ n9467 ;
  assign n9852 = n4986 & n20240 ;
  assign n9848 = n9467 ^ x11 ;
  assign n9847 = ~n1819 & n7142 ;
  assign n9849 = n9848 ^ n9847 ;
  assign n9846 = ~n1541 & n7148 ;
  assign n9850 = n9849 ^ n9846 ;
  assign n9845 = ~n1670 & n7151 ;
  assign n9851 = n9850 ^ n9845 ;
  assign n9853 = n9852 ^ n9851 ;
  assign n9854 = n9844 & ~n9853 ;
  assign n9855 = n9854 ^ n9843 ;
  assign n9857 = n9856 ^ n9855 ;
  assign n9865 = n4690 & n20240 ;
  assign n9861 = n9856 ^ x11 ;
  assign n9860 = ~n1819 & n7148 ;
  assign n9862 = n9861 ^ n9860 ;
  assign n9859 = ~n1751 & n7151 ;
  assign n9863 = n9862 ^ n9859 ;
  assign n9858 = ~n1670 & n7142 ;
  assign n9864 = n9863 ^ n9858 ;
  assign n9866 = n9865 ^ n9864 ;
  assign n9867 = n9857 & n9866 ;
  assign n9868 = n9867 ^ n9856 ;
  assign n9869 = n9868 ^ n9458 ;
  assign n9870 = ~n9466 & ~n9869 ;
  assign n9871 = n9870 ^ n9458 ;
  assign n9456 = n9389 ^ n8894 ;
  assign n9872 = n9871 ^ n9456 ;
  assign n9880 = n4475 & n20240 ;
  assign n9876 = n9456 ^ x11 ;
  assign n9875 = ~n1345 & n7151 ;
  assign n9877 = n9876 ^ n9875 ;
  assign n9874 = ~n1751 & n7148 ;
  assign n9878 = n9877 ^ n9874 ;
  assign n9873 = ~n1450 & n7142 ;
  assign n9879 = n9878 ^ n9873 ;
  assign n9881 = n9880 ^ n9879 ;
  assign n9882 = n9872 & n9881 ;
  assign n9883 = n9882 ^ n9871 ;
  assign n9884 = n9883 ^ n9447 ;
  assign n9885 = ~n9455 & n9884 ;
  assign n9886 = n9885 ^ n9447 ;
  assign n9887 = n9886 ^ n9437 ;
  assign n9888 = n9445 & ~n9887 ;
  assign n9889 = n9888 ^ n9437 ;
  assign n9890 = n9889 ^ n9429 ;
  assign n9891 = n9435 & n9890 ;
  assign n9892 = n9891 ^ n9429 ;
  assign n9893 = n9425 & ~n9892 ;
  assign n9907 = n9886 ^ n9445 ;
  assign n9903 = ~n856 & n8139 ;
  assign n9902 = ~n1119 & n8144 ;
  assign n9904 = n9903 ^ n9902 ;
  assign n9905 = n9904 ^ x8 ;
  assign n9896 = x8 ^ x7 ;
  assign n9899 = n3495 & ~n9896 ;
  assign n9900 = n9899 ^ n3930 ;
  assign n9901 = n8137 & ~n9900 ;
  assign n9906 = n9905 ^ n9901 ;
  assign n9908 = n9907 ^ n9906 ;
  assign n9917 = ~n1119 & n8139 ;
  assign n9912 = n9883 ^ n9455 ;
  assign n9913 = n9912 ^ x8 ;
  assign n9911 = ~n1248 & n8144 ;
  assign n9914 = n9913 ^ n9911 ;
  assign n9910 = ~n856 & n8484 ;
  assign n9915 = n9914 ^ n9910 ;
  assign n9909 = ~n4359 & n8150 ;
  assign n9916 = n9915 ^ n9909 ;
  assign n9918 = n9917 ^ n9916 ;
  assign n9927 = ~n1248 & n8139 ;
  assign n9924 = ~n990 & n8144 ;
  assign n9922 = ~n1119 & n8484 ;
  assign n9920 = n9881 ^ n9871 ;
  assign n9921 = n9920 ^ x8 ;
  assign n9923 = n9922 ^ n9921 ;
  assign n9925 = n9924 ^ n9923 ;
  assign n9919 = ~n4336 & n8150 ;
  assign n9926 = n9925 ^ n9919 ;
  assign n9928 = n9927 ^ n9926 ;
  assign n9939 = ~n990 & n8139 ;
  assign n9937 = ~n1345 & n8144 ;
  assign n9930 = n1248 ^ x8 ;
  assign n9931 = n9930 ^ x7 ;
  assign n9932 = n9931 ^ n1248 ;
  assign n9933 = ~n4333 & n9932 ;
  assign n9934 = n9933 ^ n1248 ;
  assign n9935 = n8137 & ~n9934 ;
  assign n9936 = n9935 ^ x8 ;
  assign n9938 = n9937 ^ n9936 ;
  assign n9940 = n9939 ^ n9938 ;
  assign n9929 = n9868 ^ n9466 ;
  assign n9941 = n9940 ^ n9929 ;
  assign n9953 = ~n1670 & n8144 ;
  assign n9948 = n9840 ^ n9477 ;
  assign n9949 = n9948 ^ x8 ;
  assign n9947 = ~n1450 & n8484 ;
  assign n9950 = n9949 ^ n9947 ;
  assign n9946 = ~n1751 & n8139 ;
  assign n9951 = n9950 ^ n9946 ;
  assign n9945 = ~n4495 & n8150 ;
  assign n9952 = n9951 ^ n9945 ;
  assign n9954 = n9953 ^ n9952 ;
  assign n9963 = ~n1819 & n8144 ;
  assign n9958 = n9837 ^ n9487 ;
  assign n9959 = n9958 ^ x8 ;
  assign n9957 = ~n1670 & n8139 ;
  assign n9960 = n9959 ^ n9957 ;
  assign n9956 = ~n1751 & n8484 ;
  assign n9961 = n9960 ^ n9956 ;
  assign n9955 = n4690 & n8150 ;
  assign n9962 = n9961 ^ n9955 ;
  assign n9964 = n9963 ^ n9962 ;
  assign n9970 = ~n1819 & n8484 ;
  assign n9969 = ~n1541 & n8139 ;
  assign n9971 = n9970 ^ n9969 ;
  assign n9972 = n9971 ^ x8 ;
  assign n9968 = ~n5154 & n8150 ;
  assign n9973 = n9972 ^ n9968 ;
  assign n9967 = ~n1972 & n8144 ;
  assign n9974 = n9973 ^ n9967 ;
  assign n9966 = n9832 ^ n9822 ;
  assign n9975 = n9974 ^ n9966 ;
  assign n9987 = ~n2095 & n8144 ;
  assign n9985 = ~n1897 & n8139 ;
  assign n9982 = n9817 ^ n9520 ;
  assign n9983 = n9982 ^ x8 ;
  assign n9979 = n5286 & ~n9896 ;
  assign n9980 = n9979 ^ n5287 ;
  assign n9981 = n8137 & ~n9980 ;
  assign n9984 = n9983 ^ n9981 ;
  assign n9986 = n9985 ^ n9984 ;
  assign n9988 = n9987 ^ n9986 ;
  assign n10004 = ~n2199 & n8144 ;
  assign n9999 = n9805 ^ n9529 ;
  assign n9997 = n9793 ^ n9531 ;
  assign n9998 = ~n9785 & n9997 ;
  assign n10000 = n9999 ^ n9998 ;
  assign n10001 = n10000 ^ x8 ;
  assign n9994 = ~n4884 & n9896 ;
  assign n9995 = n9994 ^ n1897 ;
  assign n9996 = n8137 & ~n9995 ;
  assign n10002 = n10001 ^ n9996 ;
  assign n9989 = ~n2095 & n8139 ;
  assign n10003 = n10002 ^ n9989 ;
  assign n10005 = n10004 ^ n10003 ;
  assign n10230 = n9793 ^ n9785 ;
  assign n10014 = n9782 ^ n9771 ;
  assign n10012 = ~n2199 & n8484 ;
  assign n10010 = ~n2371 & n8144 ;
  assign n10007 = n5480 & n8150 ;
  assign n10006 = ~n2288 & n8139 ;
  assign n10008 = n10007 ^ n10006 ;
  assign n10009 = n10008 ^ x8 ;
  assign n10011 = n10010 ^ n10009 ;
  assign n10013 = n10012 ^ n10011 ;
  assign n10015 = n10014 ^ n10013 ;
  assign n10214 = n9769 ^ n9532 ;
  assign n10024 = ~n2467 & n8139 ;
  assign n10019 = n9766 ^ n9755 ;
  assign n10020 = n10019 ^ x8 ;
  assign n10018 = ~n2552 & n8144 ;
  assign n10021 = n10020 ^ n10018 ;
  assign n10017 = ~n2371 & n8484 ;
  assign n10022 = n10021 ^ n10017 ;
  assign n10016 = n5696 & n8150 ;
  assign n10023 = n10022 ^ n10016 ;
  assign n10025 = n10024 ^ n10023 ;
  assign n10030 = ~n2467 & n8484 ;
  assign n10029 = ~n2589 & n8144 ;
  assign n10031 = n10030 ^ n10029 ;
  assign n10032 = n10031 ^ x8 ;
  assign n10028 = n6008 & n8150 ;
  assign n10033 = n10032 ^ n10028 ;
  assign n10027 = ~n2552 & n8139 ;
  assign n10034 = n10033 ^ n10027 ;
  assign n10026 = n9753 ^ n9740 ;
  assign n10035 = n10034 ^ n10026 ;
  assign n10047 = ~n2589 & n8139 ;
  assign n10039 = n9718 ^ n9707 ;
  assign n10040 = n9718 ^ n9542 ;
  assign n10041 = n10039 & n10040 ;
  assign n10042 = n10041 ^ n9732 ;
  assign n10043 = n10042 ^ x8 ;
  assign n10038 = ~n2552 & n8484 ;
  assign n10044 = n10043 ^ n10038 ;
  assign n10037 = ~n2657 & n8144 ;
  assign n10045 = n10044 ^ n10037 ;
  assign n10036 = n6212 & n8150 ;
  assign n10046 = n10045 ^ n10036 ;
  assign n10048 = n10047 ^ n10046 ;
  assign n10060 = ~n2712 & n8139 ;
  assign n10054 = n9702 ^ n9173 ;
  assign n10053 = n9694 ^ n9244 ;
  assign n10055 = n10054 ^ n10053 ;
  assign n10056 = n10055 ^ x8 ;
  assign n10052 = ~n3324 & n8144 ;
  assign n10057 = n10056 ^ n10052 ;
  assign n10051 = ~n2657 & n8484 ;
  assign n10058 = n10057 ^ n10051 ;
  assign n10050 = n6229 & n8150 ;
  assign n10059 = n10058 ^ n10050 ;
  assign n10061 = n10060 ^ n10059 ;
  assign n10066 = ~n2748 & n8144 ;
  assign n10065 = ~n2712 & n8484 ;
  assign n10067 = n10066 ^ n10065 ;
  assign n10068 = n10067 ^ x8 ;
  assign n10064 = n6623 & n8150 ;
  assign n10069 = n10068 ^ n10064 ;
  assign n10063 = ~n3324 & n8139 ;
  assign n10070 = n10069 ^ n10063 ;
  assign n10062 = n9691 ^ n9552 ;
  assign n10071 = n10070 ^ n10062 ;
  assign n10080 = ~n2748 & n8139 ;
  assign n10077 = ~n2839 & n8144 ;
  assign n10075 = ~n3324 & n8484 ;
  assign n10073 = n9688 ^ n9563 ;
  assign n10074 = n10073 ^ x8 ;
  assign n10076 = n10075 ^ n10074 ;
  assign n10078 = n10077 ^ n10076 ;
  assign n10072 = n7354 & n8150 ;
  assign n10079 = n10078 ^ n10072 ;
  assign n10081 = n10080 ^ n10079 ;
  assign n10091 = ~n3248 & n8144 ;
  assign n10086 = n9683 ^ n9679 ;
  assign n10087 = n10086 ^ x8 ;
  assign n10085 = ~n2935 & n8139 ;
  assign n10088 = n10087 ^ n10085 ;
  assign n10084 = ~n2839 & n8484 ;
  assign n10089 = n10088 ^ n10084 ;
  assign n10083 = ~n6695 & n8150 ;
  assign n10090 = n10089 ^ n10083 ;
  assign n10092 = n10091 ^ n10090 ;
  assign n10104 = ~n3429 & n6391 ;
  assign n10098 = ~n3022 & n8144 ;
  assign n10097 = ~n2935 & n8484 ;
  assign n10099 = n10098 ^ n10097 ;
  assign n10100 = n10099 ^ x8 ;
  assign n10096 = n6736 & n8150 ;
  assign n10101 = n10100 ^ n10096 ;
  assign n10095 = ~n3248 & n8139 ;
  assign n10102 = n10101 ^ n10095 ;
  assign n10093 = n9600 ^ x11 ;
  assign n10094 = n10093 ^ n9607 ;
  assign n10103 = n10102 ^ n10094 ;
  assign n10105 = n10104 ^ n10103 ;
  assign n10110 = ~n3022 & n8139 ;
  assign n10109 = ~n3248 & n8484 ;
  assign n10111 = n10110 ^ n10109 ;
  assign n10112 = n10111 ^ x8 ;
  assign n10108 = n6753 & n8150 ;
  assign n10113 = n10112 ^ n10108 ;
  assign n10107 = ~n3055 & n8144 ;
  assign n10114 = n10113 ^ n10107 ;
  assign n10106 = n9599 ^ n9587 ;
  assign n10115 = n10114 ^ n10106 ;
  assign n10152 = ~n3022 & n8484 ;
  assign n10151 = ~n3196 & n8144 ;
  assign n10153 = n10152 ^ n10151 ;
  assign n10154 = n10153 ^ x8 ;
  assign n10150 = n6840 & n8150 ;
  assign n10155 = n10154 ^ n10150 ;
  assign n10149 = ~n3055 & n8139 ;
  assign n10156 = n10155 ^ n10149 ;
  assign n10120 = ~n3196 & n8139 ;
  assign n10119 = ~n3124 & n8144 ;
  assign n10121 = n10120 ^ n10119 ;
  assign n10117 = ~n6863 & n8150 ;
  assign n10116 = ~n3055 & n8137 ;
  assign n10118 = n10117 ^ n10116 ;
  assign n10122 = n10121 ^ n10118 ;
  assign n10123 = ~n3429 & n7140 ;
  assign n10124 = x8 & n10123 ;
  assign n10125 = ~n10122 & ~n10124 ;
  assign n10128 = ~n3124 & n8137 ;
  assign n10129 = ~n3429 & n19031 ;
  assign n10130 = x8 & ~n10129 ;
  assign n10131 = ~n10128 & n10130 ;
  assign n10142 = ~n3429 & n8144 ;
  assign n10141 = ~n3196 & n8137 ;
  assign n10143 = n10142 ^ n10141 ;
  assign n10138 = n3429 & n8150 ;
  assign n10139 = n10138 ^ n8139 ;
  assign n10140 = ~n3124 & n10139 ;
  assign n10144 = n10143 ^ n10140 ;
  assign n10145 = n10131 & ~n10144 ;
  assign n10126 = n10123 ^ n10122 ;
  assign n10127 = n10126 ^ n10124 ;
  assign n10146 = n10145 ^ n10127 ;
  assign n10147 = n10125 & ~n10146 ;
  assign n10148 = n10147 ^ n10127 ;
  assign n10157 = n10156 ^ n10148 ;
  assign n10159 = n10156 ^ n9584 ;
  assign n10158 = ~n3429 & n7139 ;
  assign n10160 = n10159 ^ n10158 ;
  assign n10161 = ~n10157 & n10160 ;
  assign n10162 = n10161 ^ n10156 ;
  assign n10163 = n10162 ^ n10114 ;
  assign n10164 = n10115 & n10163 ;
  assign n10165 = n10164 ^ n10114 ;
  assign n10166 = n10165 ^ n10102 ;
  assign n10167 = n10105 & n10166 ;
  assign n10168 = n10167 ^ n10102 ;
  assign n10169 = n10168 ^ n10086 ;
  assign n10170 = n10092 & n10169 ;
  assign n10171 = n10170 ^ n10086 ;
  assign n10082 = n9685 ^ n9573 ;
  assign n10172 = n10171 ^ n10082 ;
  assign n10180 = ~n2839 & n8139 ;
  assign n10176 = n10082 ^ x8 ;
  assign n10175 = ~n2748 & n8484 ;
  assign n10177 = n10176 ^ n10175 ;
  assign n10174 = ~n2935 & n8144 ;
  assign n10178 = n10177 ^ n10174 ;
  assign n10173 = ~n6302 & n8150 ;
  assign n10179 = n10178 ^ n10173 ;
  assign n10181 = n10180 ^ n10179 ;
  assign n10182 = n10172 & ~n10181 ;
  assign n10183 = n10182 ^ n10171 ;
  assign n10184 = n10183 ^ n10073 ;
  assign n10185 = ~n10081 & ~n10184 ;
  assign n10186 = n10185 ^ n10073 ;
  assign n10187 = n10186 ^ n10070 ;
  assign n10188 = n10071 & ~n10187 ;
  assign n10189 = n10188 ^ n10070 ;
  assign n10190 = n10189 ^ n10055 ;
  assign n10191 = ~n10061 & ~n10190 ;
  assign n10192 = n10191 ^ n10055 ;
  assign n10049 = n9718 ^ n9709 ;
  assign n10193 = n10192 ^ n10049 ;
  assign n10201 = ~n2657 & n8139 ;
  assign n10197 = n10049 ^ x8 ;
  assign n10196 = ~n2712 & n8144 ;
  assign n10198 = n10197 ^ n10196 ;
  assign n10195 = ~n2589 & n8484 ;
  assign n10199 = n10198 ^ n10195 ;
  assign n10194 = n6079 & n8150 ;
  assign n10200 = n10199 ^ n10194 ;
  assign n10202 = n10201 ^ n10200 ;
  assign n10203 = ~n10193 & ~n10202 ;
  assign n10204 = n10203 ^ n10192 ;
  assign n10205 = n10204 ^ n10042 ;
  assign n10206 = ~n10048 & n10205 ;
  assign n10207 = n10206 ^ n10042 ;
  assign n10208 = n10207 ^ n10034 ;
  assign n10209 = n10035 & ~n10208 ;
  assign n10210 = n10209 ^ n10034 ;
  assign n10211 = n10210 ^ n10019 ;
  assign n10212 = ~n10025 & ~n10211 ;
  assign n10213 = n10212 ^ n10019 ;
  assign n10215 = n10214 ^ n10213 ;
  assign n10223 = ~n2467 & n8144 ;
  assign n10219 = n10214 ^ x8 ;
  assign n10218 = n6449 & n8150 ;
  assign n10220 = n10219 ^ n10218 ;
  assign n10217 = ~n2371 & n8139 ;
  assign n10221 = n10220 ^ n10217 ;
  assign n10216 = ~n2288 & n8484 ;
  assign n10222 = n10221 ^ n10216 ;
  assign n10224 = n10223 ^ n10222 ;
  assign n10225 = ~n10215 & n10224 ;
  assign n10226 = n10225 ^ n10214 ;
  assign n10227 = n10226 ^ n10013 ;
  assign n10228 = n10015 & ~n10227 ;
  assign n10229 = n10228 ^ n10014 ;
  assign n10231 = n10230 ^ n10229 ;
  assign n10239 = ~n2199 & n8139 ;
  assign n10235 = n10230 ^ x8 ;
  assign n10234 = ~n2095 & n8484 ;
  assign n10236 = n10235 ^ n10234 ;
  assign n10233 = ~n2288 & n8144 ;
  assign n10237 = n10236 ^ n10233 ;
  assign n10232 = n5760 & n8150 ;
  assign n10238 = n10237 ^ n10232 ;
  assign n10240 = n10239 ^ n10238 ;
  assign n10241 = n10231 & n10240 ;
  assign n10242 = n10241 ^ n10230 ;
  assign n10243 = n10242 ^ n10000 ;
  assign n10244 = n10005 & ~n10243 ;
  assign n10245 = n10244 ^ n10242 ;
  assign n10246 = n10245 ^ n9982 ;
  assign n10247 = n9988 & n10246 ;
  assign n10248 = n10247 ^ n9982 ;
  assign n9976 = n9819 ^ n9511 ;
  assign n10249 = n10248 ^ n9976 ;
  assign n10257 = ~n1897 & n8144 ;
  assign n10253 = n9976 ^ x8 ;
  assign n10252 = ~n1972 & n8139 ;
  assign n10254 = n10253 ^ n10252 ;
  assign n10251 = ~n1541 & n8484 ;
  assign n10255 = n10254 ^ n10251 ;
  assign n10250 = ~n4892 & n8150 ;
  assign n10256 = n10255 ^ n10250 ;
  assign n10258 = n10257 ^ n10256 ;
  assign n10259 = n10249 & ~n10258 ;
  assign n10260 = n10259 ^ n10248 ;
  assign n10261 = n10260 ^ n9974 ;
  assign n10262 = ~n9975 & n10261 ;
  assign n10263 = n10262 ^ n9974 ;
  assign n9965 = n9834 ^ n9497 ;
  assign n10264 = n10263 ^ n9965 ;
  assign n10276 = ~n1541 & n8144 ;
  assign n10273 = n9965 ^ x8 ;
  assign n10270 = ~n4985 & n9896 ;
  assign n10271 = n10270 ^ n1670 ;
  assign n10272 = n8137 & ~n10271 ;
  assign n10274 = n10273 ^ n10272 ;
  assign n10265 = ~n1819 & n8139 ;
  assign n10275 = n10274 ^ n10265 ;
  assign n10277 = n10276 ^ n10275 ;
  assign n10278 = ~n10264 & n10277 ;
  assign n10279 = n10278 ^ n10263 ;
  assign n10280 = n10279 ^ n9958 ;
  assign n10281 = ~n9964 & ~n10280 ;
  assign n10282 = n10281 ^ n9958 ;
  assign n10283 = n10282 ^ n9948 ;
  assign n10284 = n9954 & ~n10283 ;
  assign n10285 = n10284 ^ n9948 ;
  assign n9944 = n9853 ^ n9843 ;
  assign n10286 = n10285 ^ n9944 ;
  assign n10294 = ~n1450 & n8139 ;
  assign n10290 = n9944 ^ x8 ;
  assign n10289 = ~n1345 & n8484 ;
  assign n10291 = n10290 ^ n10289 ;
  assign n10288 = ~n1751 & n8144 ;
  assign n10292 = n10291 ^ n10288 ;
  assign n10287 = n4475 & n8150 ;
  assign n10293 = n10292 ^ n10287 ;
  assign n10295 = n10294 ^ n10293 ;
  assign n10296 = n10286 & ~n10295 ;
  assign n10297 = n10296 ^ n10285 ;
  assign n9942 = n9866 ^ n9855 ;
  assign n10298 = n10297 ^ n9942 ;
  assign n10306 = ~n1450 & n8144 ;
  assign n10302 = n9942 ^ x8 ;
  assign n10301 = ~n1345 & n8139 ;
  assign n10303 = n10302 ^ n10301 ;
  assign n10300 = ~n990 & n8484 ;
  assign n10304 = n10303 ^ n10300 ;
  assign n10299 = n4307 & n8150 ;
  assign n10305 = n10304 ^ n10299 ;
  assign n10307 = n10306 ^ n10305 ;
  assign n10308 = n10298 & n10307 ;
  assign n9943 = n9942 ^ n9929 ;
  assign n10309 = n10308 ^ n9943 ;
  assign n10310 = ~n9941 & n10309 ;
  assign n10311 = n10310 ^ n9940 ;
  assign n10312 = n10311 ^ n9920 ;
  assign n10313 = n9928 & n10312 ;
  assign n10314 = n10313 ^ n9920 ;
  assign n10315 = n10314 ^ n9912 ;
  assign n10316 = n9918 & n10315 ;
  assign n10317 = n10316 ^ n9912 ;
  assign n10318 = n10317 ^ n9906 ;
  assign n10319 = n9908 & n10318 ;
  assign n10320 = n10319 ^ n10317 ;
  assign n9894 = n9889 ^ n9435 ;
  assign n10321 = n10320 ^ n9894 ;
  assign n10322 = x3 ^ x2 ;
  assign n25051 = x5 & n10322 ;
  assign n10325 = x4 & n10322 ;
  assign n10342 = n25051 ^ n10325 ;
  assign n10343 = ~n3513 & n10342 ;
  assign n10336 = n9894 ^ x5 ;
  assign n10326 = n10325 ^ x4 ;
  assign n10324 = x2 & x3 ;
  assign n10327 = n10326 ^ n10324 ;
  assign n10333 = n10327 ^ n10322 ;
  assign n10329 = x5 ^ x4 ;
  assign n10330 = x4 ^ x3 ;
  assign n10331 = ~n10322 & ~n10330 ;
  assign n10332 = ~n10329 & n10331 ;
  assign n10334 = n10333 ^ n10332 ;
  assign n10335 = ~n408 & ~n10334 ;
  assign n10337 = n10336 ^ n10335 ;
  assign n10328 = ~n3505 & n10327 ;
  assign n10338 = n10337 ^ n10328 ;
  assign n10323 = ~n368 & n10322 ;
  assign n10339 = n10338 ^ n10323 ;
  assign n10344 = n10343 ^ n10339 ;
  assign n10345 = n10321 & ~n10344 ;
  assign n10346 = n10345 ^ n10320 ;
  assign n10347 = n9893 & ~n10346 ;
  assign n10350 = ~n3505 & ~n10334 ;
  assign n10349 = ~n368 & n10327 ;
  assign n10351 = n10350 ^ n10349 ;
  assign n10352 = n10351 ^ x5 ;
  assign n10348 = n3515 & n10342 ;
  assign n10353 = n10352 ^ n10348 ;
  assign n10354 = n10347 & ~n10353 ;
  assign n10372 = ~n408 & n8139 ;
  assign n10371 = ~n3505 & n8484 ;
  assign n10373 = n10372 ^ n10371 ;
  assign n10374 = n10373 ^ x8 ;
  assign n10370 = n3840 & n8150 ;
  assign n10375 = n10374 ^ n10370 ;
  assign n10369 = ~n540 & n8144 ;
  assign n10376 = n10375 ^ n10369 ;
  assign n10368 = n8462 ^ n8178 ;
  assign n10377 = n10376 ^ n10368 ;
  assign n10365 = n8807 ^ n8805 ;
  assign n10366 = n8815 & ~n10365 ;
  assign n10367 = n10366 ^ n8807 ;
  assign n10378 = n10377 ^ n10367 ;
  assign n10379 = n10378 ^ x5 ;
  assign n10362 = ~n3509 & n10342 ;
  assign n10363 = n10362 ^ n10334 ;
  assign n10364 = ~n368 & ~n10363 ;
  assign n10380 = n10379 ^ n10364 ;
  assign n10355 = n9424 ^ n8816 ;
  assign n10356 = n8822 & ~n10355 ;
  assign n10357 = n10356 ^ n9424 ;
  assign n10381 = n10380 ^ n10357 ;
  assign n10382 = ~n10354 & ~n10381 ;
  assign n10393 = n10353 ^ n9425 ;
  assign n10394 = n10393 ^ n9892 ;
  assign n10395 = n10394 ^ n10346 ;
  assign n10385 = n9892 ^ n9425 ;
  assign n10390 = n10385 ^ n10347 ;
  assign n10386 = n10346 ^ n9892 ;
  assign n10387 = n10385 & n10386 ;
  assign n10391 = n10390 ^ n10387 ;
  assign n10392 = n10353 & n10391 ;
  assign n10396 = n10395 ^ n10392 ;
  assign n10383 = n10353 ^ n10347 ;
  assign n10384 = n10383 ^ n10354 ;
  assign n10388 = n10387 ^ n10346 ;
  assign n10389 = ~n10384 & ~n10388 ;
  assign n10397 = n10396 ^ n10389 ;
  assign n10398 = n10382 & n10397 ;
  assign n10399 = n10398 ^ n10354 ;
  assign n11755 = n10344 ^ n10320 ;
  assign n10967 = n3968 & n10342 ;
  assign n10965 = ~n698 & n10327 ;
  assign n10962 = ~n856 & ~n10334 ;
  assign n10425 = n10342 ^ n10322 ;
  assign n10961 = ~n540 & n10425 ;
  assign n10963 = n10962 ^ n10961 ;
  assign n10964 = n10963 ^ x5 ;
  assign n10966 = n10965 ^ n10964 ;
  assign n10968 = n10967 ^ n10966 ;
  assign n10420 = n10309 ^ n9940 ;
  assign n10969 = n10968 ^ n10420 ;
  assign n10426 = ~n698 & n10425 ;
  assign n10421 = n10420 ^ x5 ;
  assign n10419 = ~n3930 & n10342 ;
  assign n10422 = n10421 ^ n10419 ;
  assign n10418 = ~n1119 & ~n10334 ;
  assign n10423 = n10422 ^ n10418 ;
  assign n10417 = ~n856 & n10327 ;
  assign n10424 = n10423 ^ n10417 ;
  assign n10427 = n10426 ^ n10424 ;
  assign n10439 = ~n1119 & n10327 ;
  assign n10435 = n10307 ^ n10297 ;
  assign n10436 = n10435 ^ x5 ;
  assign n10432 = n3493 & n10329 ;
  assign n10433 = n10432 ^ n856 ;
  assign n10434 = n10322 & ~n10433 ;
  assign n10437 = n10436 ^ n10434 ;
  assign n10428 = ~n1248 & ~n10334 ;
  assign n10438 = n10437 ^ n10428 ;
  assign n10440 = n10439 ^ n10438 ;
  assign n10452 = ~n990 & ~n10334 ;
  assign n10448 = n10295 ^ n10285 ;
  assign n10449 = n10448 ^ x5 ;
  assign n10445 = n4335 & n10329 ;
  assign n10446 = n10445 ^ n1119 ;
  assign n10447 = n10322 & ~n10446 ;
  assign n10450 = n10449 ^ n10447 ;
  assign n10441 = ~n1248 & n10327 ;
  assign n10451 = n10450 ^ n10441 ;
  assign n10453 = n10452 ^ n10451 ;
  assign n10467 = ~n1345 & n10327 ;
  assign n10463 = n10279 ^ n9964 ;
  assign n10464 = n10463 ^ x5 ;
  assign n10460 = ~n3486 & n10329 ;
  assign n10461 = n10460 ^ n990 ;
  assign n10462 = n10322 & ~n10461 ;
  assign n10465 = n10464 ^ n10462 ;
  assign n10455 = ~n1450 & ~n10334 ;
  assign n10466 = n10465 ^ n10455 ;
  assign n10468 = n10467 ^ n10466 ;
  assign n10916 = ~n1450 & n10425 ;
  assign n10914 = ~n1670 & ~n10334 ;
  assign n10911 = ~n4495 & n10342 ;
  assign n10910 = ~n1751 & n10327 ;
  assign n10912 = n10911 ^ n10910 ;
  assign n10913 = n10912 ^ x5 ;
  assign n10915 = n10914 ^ n10913 ;
  assign n10917 = n10916 ^ n10915 ;
  assign n10483 = ~n1819 & ~n10334 ;
  assign n10479 = n10258 ^ n10248 ;
  assign n10480 = n10479 ^ x5 ;
  assign n10476 = ~n4492 & n10329 ;
  assign n10477 = n10476 ^ n1751 ;
  assign n10478 = n10322 & ~n10477 ;
  assign n10481 = n10480 ^ n10478 ;
  assign n10471 = ~n1670 & n10327 ;
  assign n10482 = n10481 ^ n10471 ;
  assign n10484 = n10483 ^ n10482 ;
  assign n10492 = ~n1670 & n10425 ;
  assign n10490 = ~n1541 & ~n10334 ;
  assign n10487 = n4986 & n10342 ;
  assign n10486 = ~n1819 & n10327 ;
  assign n10488 = n10487 ^ n10486 ;
  assign n10489 = n10488 ^ x5 ;
  assign n10491 = n10490 ^ n10489 ;
  assign n10493 = n10492 ^ n10491 ;
  assign n10485 = n10245 ^ n9988 ;
  assign n10494 = n10493 ^ n10485 ;
  assign n10506 = n10242 ^ n10005 ;
  assign n10503 = ~n1972 & ~n10334 ;
  assign n10502 = ~n1541 & n10327 ;
  assign n10504 = n10503 ^ n10502 ;
  assign n10495 = n1819 ^ x5 ;
  assign n10496 = n10495 ^ x4 ;
  assign n10497 = n10496 ^ n1819 ;
  assign n10498 = n4488 & n10497 ;
  assign n10499 = n10498 ^ n1819 ;
  assign n10500 = n10322 & ~n10499 ;
  assign n10501 = n10500 ^ x5 ;
  assign n10505 = n10504 ^ n10501 ;
  assign n10507 = n10506 ^ n10505 ;
  assign n10518 = n10240 ^ n10229 ;
  assign n10514 = ~n1897 & ~n10334 ;
  assign n10513 = ~n1972 & n10327 ;
  assign n10515 = n10514 ^ n10513 ;
  assign n10516 = n10515 ^ x5 ;
  assign n10510 = n4891 & ~n10329 ;
  assign n10511 = n10510 ^ n4892 ;
  assign n10512 = n10322 & ~n10511 ;
  assign n10517 = n10516 ^ n10512 ;
  assign n10519 = n10518 ^ n10517 ;
  assign n10527 = ~n1972 & n10425 ;
  assign n10525 = ~n1897 & n10327 ;
  assign n10522 = ~n5287 & n10342 ;
  assign n10521 = ~n2095 & ~n10334 ;
  assign n10523 = n10522 ^ n10521 ;
  assign n10524 = n10523 ^ x5 ;
  assign n10526 = n10525 ^ n10524 ;
  assign n10528 = n10527 ^ n10526 ;
  assign n10520 = n10226 ^ n10015 ;
  assign n10529 = n10528 ^ n10520 ;
  assign n10537 = n5824 & n10342 ;
  assign n10533 = n10224 ^ n10213 ;
  assign n10534 = n10533 ^ x5 ;
  assign n10532 = ~n2199 & ~n10334 ;
  assign n10535 = n10534 ^ n10532 ;
  assign n10531 = ~n2095 & n10327 ;
  assign n10536 = n10535 ^ n10531 ;
  assign n10538 = n10537 ^ n10536 ;
  assign n10530 = ~n1897 & n10425 ;
  assign n10539 = n10538 ^ n10530 ;
  assign n10547 = ~n2095 & n10425 ;
  assign n10545 = n5760 & n10342 ;
  assign n10542 = ~n2199 & n10327 ;
  assign n10541 = ~n2288 & ~n10334 ;
  assign n10543 = n10542 ^ n10541 ;
  assign n10544 = n10543 ^ x5 ;
  assign n10546 = n10545 ^ n10544 ;
  assign n10548 = n10547 ^ n10546 ;
  assign n10540 = n10210 ^ n10025 ;
  assign n10549 = n10548 ^ n10540 ;
  assign n10559 = ~n2288 & n10425 ;
  assign n10556 = ~n2371 & n10327 ;
  assign n10554 = ~n2467 & ~n10334 ;
  assign n10552 = n10204 ^ n10048 ;
  assign n10553 = n10552 ^ x5 ;
  assign n10555 = n10554 ^ n10553 ;
  assign n10557 = n10556 ^ n10555 ;
  assign n10551 = n6449 & n10342 ;
  assign n10558 = n10557 ^ n10551 ;
  assign n10560 = n10559 ^ n10558 ;
  assign n10570 = ~n2467 & n10425 ;
  assign n10565 = n10189 ^ n10061 ;
  assign n10566 = n10565 ^ x5 ;
  assign n10564 = ~n2552 & n10327 ;
  assign n10567 = n10566 ^ n10564 ;
  assign n10563 = ~n2589 & ~n10334 ;
  assign n10568 = n10567 ^ n10563 ;
  assign n10562 = n6008 & n10342 ;
  assign n10569 = n10568 ^ n10562 ;
  assign n10571 = n10570 ^ n10569 ;
  assign n10831 = n10183 ^ n10081 ;
  assign n10582 = ~n2712 & n10425 ;
  assign n10579 = ~n3324 & n10327 ;
  assign n10577 = ~n2748 & ~n10334 ;
  assign n10575 = n10168 ^ n10092 ;
  assign n10576 = n10575 ^ x5 ;
  assign n10578 = n10577 ^ n10576 ;
  assign n10580 = n10579 ^ n10578 ;
  assign n10574 = n6623 & n10342 ;
  assign n10581 = n10580 ^ n10574 ;
  assign n10583 = n10582 ^ n10581 ;
  assign n10595 = ~n2839 & ~n10334 ;
  assign n10591 = n10165 ^ n10105 ;
  assign n10592 = n10591 ^ x5 ;
  assign n10588 = ~n6643 & n10329 ;
  assign n10589 = n10588 ^ n3324 ;
  assign n10590 = n10322 & ~n10589 ;
  assign n10593 = n10592 ^ n10590 ;
  assign n10584 = ~n2748 & n10327 ;
  assign n10594 = n10593 ^ n10584 ;
  assign n10596 = n10595 ^ n10594 ;
  assign n10604 = ~n2839 & n10322 ;
  assign n10603 = n3439 & n10342 ;
  assign n10605 = n10604 ^ n10603 ;
  assign n10600 = ~n3248 & ~n10334 ;
  assign n10599 = ~n2935 & n10327 ;
  assign n10601 = n10600 ^ n10599 ;
  assign n10602 = n10601 ^ x5 ;
  assign n10606 = n10605 ^ n10602 ;
  assign n10598 = n10160 ^ n10148 ;
  assign n10607 = n10606 ^ n10598 ;
  assign n10617 = ~n2935 & n10425 ;
  assign n10615 = ~n3248 & n10327 ;
  assign n10612 = n6736 & n10342 ;
  assign n10611 = ~n3022 & ~n10334 ;
  assign n10613 = n10612 ^ n10611 ;
  assign n10614 = n10613 ^ x5 ;
  assign n10616 = n10615 ^ n10614 ;
  assign n10618 = n10617 ^ n10616 ;
  assign n10608 = n10145 ^ x8 ;
  assign n10609 = n10608 ^ n10122 ;
  assign n10610 = n10609 ^ n10123 ;
  assign n10619 = n10618 ^ n10610 ;
  assign n10626 = ~n3248 & n10322 ;
  assign n10625 = ~n6749 & n10342 ;
  assign n10627 = n10626 ^ n10625 ;
  assign n10622 = ~n3022 & n10327 ;
  assign n10621 = ~n3055 & ~n10334 ;
  assign n10623 = n10622 ^ n10621 ;
  assign n10624 = n10623 ^ x5 ;
  assign n10628 = n10627 ^ n10624 ;
  assign n10132 = n10131 ^ x8 ;
  assign n10620 = n10144 ^ n10132 ;
  assign n10629 = n10628 ^ n10620 ;
  assign n10656 = n6864 & n10342 ;
  assign n10653 = ~n3196 & n10327 ;
  assign n10652 = ~n3055 & n10425 ;
  assign n10654 = n10653 ^ n10652 ;
  assign n10651 = ~n3124 & ~n10334 ;
  assign n10655 = n10654 ^ n10651 ;
  assign n10657 = n10656 ^ n10655 ;
  assign n10632 = x5 & n10333 ;
  assign n10633 = ~n3124 & n10322 ;
  assign n10634 = n3429 & ~n10633 ;
  assign n10635 = n10632 & n10634 ;
  assign n10636 = n10635 ^ n10632 ;
  assign n10637 = n10636 ^ x5 ;
  assign n10646 = ~n3429 & ~n10334 ;
  assign n10645 = ~n3196 & n10322 ;
  assign n10647 = n10646 ^ n10645 ;
  assign n10642 = n3429 & n10342 ;
  assign n10643 = n10642 ^ n10327 ;
  assign n10644 = ~n3124 & n10643 ;
  assign n10648 = n10647 ^ n10644 ;
  assign n10649 = n10637 & ~n10648 ;
  assign n10658 = n10657 ^ n10649 ;
  assign n10672 = n10658 ^ x6 ;
  assign n10774 = n10672 ^ n3429 ;
  assign n10775 = n10774 ^ n10658 ;
  assign n10674 = n10658 ^ x5 ;
  assign n10776 = n10775 ^ n10674 ;
  assign n10777 = n10776 ^ x6 ;
  assign n10778 = n10777 ^ n10657 ;
  assign n10757 = n10649 ^ x6 ;
  assign n10758 = n10757 ^ n10657 ;
  assign n10678 = n10649 ^ x5 ;
  assign n10679 = n10678 ^ n3429 ;
  assign n10680 = n10679 ^ n10657 ;
  assign n10759 = n10758 ^ n10680 ;
  assign n10710 = ~n10649 & ~n10658 ;
  assign n10711 = n10710 ^ x6 ;
  assign n10712 = n10711 ^ x5 ;
  assign n10713 = n10712 ^ n10657 ;
  assign n10698 = n10674 ^ n3429 ;
  assign n10699 = n10698 ^ n10658 ;
  assign n10706 = n10699 ^ x6 ;
  assign n10714 = n10706 ^ x5 ;
  assign n10715 = n10714 ^ n10657 ;
  assign n10716 = ~n10713 & ~n10715 ;
  assign n10700 = n10699 ^ n10672 ;
  assign n10701 = n10700 ^ x5 ;
  assign n10703 = n10701 ^ n10657 ;
  assign n10677 = n10674 ^ x6 ;
  assign n10718 = n10703 ^ n10677 ;
  assign n10719 = n10701 ^ x6 ;
  assign n10720 = n10719 ^ n10703 ;
  assign n10721 = n10718 & ~n10720 ;
  assign n10722 = n10716 & n10721 ;
  assign n10723 = n10722 ^ n10710 ;
  assign n10742 = n10723 ^ n8137 ;
  assign n10688 = n3429 ^ x5 ;
  assign n10662 = n10688 ^ n10657 ;
  assign n10755 = n10742 ^ n10662 ;
  assign n10682 = n10688 ^ n10677 ;
  assign n10684 = n10682 ^ n10657 ;
  assign n10756 = n10755 ^ n10684 ;
  assign n10760 = n10759 ^ n10756 ;
  assign n10772 = n10760 ^ n10757 ;
  assign n10773 = n10772 ^ n10649 ;
  assign n10779 = n10778 ^ n10773 ;
  assign n10630 = n8136 & n10129 ;
  assign n10631 = n10630 ^ n10128 ;
  assign n10780 = n10779 ^ n10631 ;
  assign n10787 = ~n3055 & n10327 ;
  assign n10785 = n6840 & n10342 ;
  assign n10783 = ~n3196 & ~n10334 ;
  assign n10782 = n10631 ^ x5 ;
  assign n10784 = n10783 ^ n10782 ;
  assign n10786 = n10785 ^ n10784 ;
  assign n10788 = n10787 ^ n10786 ;
  assign n10781 = ~n3022 & n10425 ;
  assign n10789 = n10788 ^ n10781 ;
  assign n10790 = ~n10780 & ~n10789 ;
  assign n10791 = n10790 ^ n10779 ;
  assign n10792 = n10791 ^ n10628 ;
  assign n10793 = n10629 & ~n10792 ;
  assign n10794 = n10793 ^ n10628 ;
  assign n10795 = n10794 ^ n10618 ;
  assign n10796 = n10619 & n10795 ;
  assign n10797 = n10796 ^ n10618 ;
  assign n10798 = n10797 ^ n10606 ;
  assign n10799 = ~n10607 & n10798 ;
  assign n10800 = n10799 ^ n10606 ;
  assign n10597 = n10162 ^ n10115 ;
  assign n10801 = n10800 ^ n10597 ;
  assign n10808 = ~n2748 & n10322 ;
  assign n10806 = ~n2935 & ~n10334 ;
  assign n10804 = ~n2839 & n10327 ;
  assign n10803 = n10597 ^ x5 ;
  assign n10805 = n10804 ^ n10803 ;
  assign n10807 = n10806 ^ n10805 ;
  assign n10809 = n10808 ^ n10807 ;
  assign n10802 = n6301 & n10342 ;
  assign n10810 = n10809 ^ n10802 ;
  assign n10811 = n10801 & ~n10810 ;
  assign n10812 = n10811 ^ n10800 ;
  assign n10813 = n10812 ^ n10591 ;
  assign n10814 = n10596 & n10813 ;
  assign n10815 = n10814 ^ n10591 ;
  assign n10816 = n10815 ^ n10575 ;
  assign n10817 = n10583 & n10816 ;
  assign n10818 = n10817 ^ n10575 ;
  assign n10573 = n10181 ^ n10171 ;
  assign n10819 = n10818 ^ n10573 ;
  assign n10827 = ~n2657 & n10425 ;
  assign n10823 = n10573 ^ x5 ;
  assign n10822 = ~n3324 & ~n10334 ;
  assign n10824 = n10823 ^ n10822 ;
  assign n10821 = ~n2712 & n10327 ;
  assign n10825 = n10824 ^ n10821 ;
  assign n10820 = n6229 & n10342 ;
  assign n10826 = n10825 ^ n10820 ;
  assign n10828 = n10827 ^ n10826 ;
  assign n10829 = n10819 & ~n10828 ;
  assign n10830 = n10829 ^ n10818 ;
  assign n10832 = n10831 ^ n10830 ;
  assign n10840 = ~n2589 & n10425 ;
  assign n10836 = n10831 ^ x5 ;
  assign n10835 = ~n2712 & ~n10334 ;
  assign n10837 = n10836 ^ n10835 ;
  assign n10834 = ~n2657 & n10327 ;
  assign n10838 = n10837 ^ n10834 ;
  assign n10833 = n6079 & n10342 ;
  assign n10839 = n10838 ^ n10833 ;
  assign n10841 = n10840 ^ n10839 ;
  assign n10842 = ~n10832 & ~n10841 ;
  assign n10843 = n10842 ^ n10831 ;
  assign n10572 = n10186 ^ n10071 ;
  assign n10844 = n10843 ^ n10572 ;
  assign n10852 = ~n2552 & n10425 ;
  assign n10848 = n10572 ^ x5 ;
  assign n10847 = ~n2589 & n10327 ;
  assign n10849 = n10848 ^ n10847 ;
  assign n10846 = ~n2657 & ~n10334 ;
  assign n10850 = n10849 ^ n10846 ;
  assign n10845 = n6212 & n10342 ;
  assign n10851 = n10850 ^ n10845 ;
  assign n10853 = n10852 ^ n10851 ;
  assign n10854 = n10844 & n10853 ;
  assign n10855 = n10854 ^ n10843 ;
  assign n10856 = n10855 ^ n10565 ;
  assign n10857 = ~n10571 & n10856 ;
  assign n10858 = n10857 ^ n10565 ;
  assign n10561 = n10202 ^ n10192 ;
  assign n10859 = n10858 ^ n10561 ;
  assign n10867 = ~n2552 & ~n10334 ;
  assign n10863 = n10561 ^ x5 ;
  assign n10862 = ~n2467 & n10327 ;
  assign n10864 = n10863 ^ n10862 ;
  assign n10861 = ~n2371 & n10425 ;
  assign n10865 = n10864 ^ n10861 ;
  assign n10860 = n5696 & n10342 ;
  assign n10866 = n10865 ^ n10860 ;
  assign n10868 = n10867 ^ n10866 ;
  assign n10869 = n10859 & n10868 ;
  assign n10870 = n10869 ^ n10858 ;
  assign n10871 = n10870 ^ n10552 ;
  assign n10872 = n10560 & ~n10871 ;
  assign n10873 = n10872 ^ n10552 ;
  assign n10550 = n10207 ^ n10035 ;
  assign n10874 = n10873 ^ n10550 ;
  assign n10882 = ~n2199 & n10425 ;
  assign n10878 = n10550 ^ x5 ;
  assign n10877 = ~n2288 & n10327 ;
  assign n10879 = n10878 ^ n10877 ;
  assign n10876 = ~n2371 & ~n10334 ;
  assign n10880 = n10879 ^ n10876 ;
  assign n10875 = n5480 & n10342 ;
  assign n10881 = n10880 ^ n10875 ;
  assign n10883 = n10882 ^ n10881 ;
  assign n10884 = ~n10874 & n10883 ;
  assign n10885 = n10884 ^ n10873 ;
  assign n10886 = n10885 ^ n10540 ;
  assign n10887 = ~n10549 & n10886 ;
  assign n10888 = n10887 ^ n10548 ;
  assign n10889 = n10888 ^ n10533 ;
  assign n10890 = ~n10539 & ~n10889 ;
  assign n10891 = n10890 ^ n10533 ;
  assign n10892 = n10891 ^ n10520 ;
  assign n10893 = n10529 & n10892 ;
  assign n10894 = n10893 ^ n10528 ;
  assign n10895 = n10894 ^ n10517 ;
  assign n10896 = n10519 & ~n10895 ;
  assign n10897 = n10896 ^ n10518 ;
  assign n10898 = n10897 ^ n10505 ;
  assign n10899 = ~n10507 & ~n10898 ;
  assign n10900 = n10899 ^ n10506 ;
  assign n10901 = n10900 ^ n10493 ;
  assign n10902 = n10494 & ~n10901 ;
  assign n10903 = n10902 ^ n10493 ;
  assign n10904 = n10903 ^ n10479 ;
  assign n10905 = n10484 & n10904 ;
  assign n10906 = n10905 ^ n10479 ;
  assign n10470 = n10260 ^ n9975 ;
  assign n10909 = n10906 ^ n10470 ;
  assign n10919 = n10917 ^ n10909 ;
  assign n10918 = n10909 & ~n10917 ;
  assign n10920 = n10919 ^ n10918 ;
  assign n10907 = ~n10470 & n10906 ;
  assign n10908 = n10907 ^ n10470 ;
  assign n10921 = n10920 ^ n10908 ;
  assign n10922 = n10921 ^ n10470 ;
  assign n10469 = n10277 ^ n10263 ;
  assign n10923 = n10922 ^ n10469 ;
  assign n10932 = n10469 ^ x5 ;
  assign n10931 = ~n1450 & n10327 ;
  assign n10933 = n10932 ^ n10931 ;
  assign n10930 = ~n1751 & ~n10334 ;
  assign n10934 = n10933 ^ n10930 ;
  assign n10924 = n4475 ^ n1345 ;
  assign n10927 = ~n10329 & ~n10924 ;
  assign n10928 = n10927 ^ n4475 ;
  assign n10929 = n10322 & n10928 ;
  assign n10935 = n10934 ^ n10929 ;
  assign n10936 = ~n10923 & n10935 ;
  assign n10937 = n10936 ^ n10922 ;
  assign n10938 = n10937 ^ n10463 ;
  assign n10939 = ~n10468 & ~n10938 ;
  assign n10940 = n10939 ^ n10463 ;
  assign n10454 = n10282 ^ n9954 ;
  assign n10941 = n10940 ^ n10454 ;
  assign n10949 = ~n1248 & n10425 ;
  assign n10945 = n10454 ^ x5 ;
  assign n10944 = ~n1345 & ~n10334 ;
  assign n10946 = n10945 ^ n10944 ;
  assign n10943 = ~n990 & n10327 ;
  assign n10947 = n10946 ^ n10943 ;
  assign n10942 = n4580 & n10342 ;
  assign n10948 = n10947 ^ n10942 ;
  assign n10950 = n10949 ^ n10948 ;
  assign n10951 = n10941 & n10950 ;
  assign n10952 = n10951 ^ n10940 ;
  assign n10953 = n10952 ^ n10448 ;
  assign n10954 = n10453 & ~n10953 ;
  assign n10955 = n10954 ^ n10448 ;
  assign n10956 = n10955 ^ n10435 ;
  assign n10957 = n10440 & n10956 ;
  assign n10958 = n10957 ^ n10435 ;
  assign n10959 = n10958 ^ n10420 ;
  assign n10960 = ~n10427 & ~n10959 ;
  assign n10970 = n10969 ^ n10960 ;
  assign n10971 = n10311 ^ n9928 ;
  assign n11718 = n10971 ^ n10968 ;
  assign n11719 = n10970 & n11718 ;
  assign n11720 = n11719 ^ n10971 ;
  assign n11727 = n3812 & n10342 ;
  assign n11725 = ~n698 & ~n10334 ;
  assign n11722 = ~n540 & n10327 ;
  assign n11721 = ~n408 & n10425 ;
  assign n11723 = n11722 ^ n11721 ;
  assign n11724 = n11723 ^ x5 ;
  assign n11726 = n11725 ^ n11724 ;
  assign n11728 = n11727 ^ n11726 ;
  assign n11737 = n11720 & n11728 ;
  assign n11729 = n11728 ^ n11720 ;
  assign n11751 = n11737 ^ n11729 ;
  assign n11715 = n10317 ^ n9908 ;
  assign n11012 = x2 ^ x1 ;
  assign n11698 = ~n368 & n11012 ;
  assign n11709 = n3509 ^ x2 ;
  assign n11711 = x0 & ~n11709 ;
  assign n11712 = n11711 ^ x2 ;
  assign n11713 = n11698 & n11712 ;
  assign n11702 = ~n540 & ~n10334 ;
  assign n11701 = ~n3505 & n10425 ;
  assign n11703 = n11702 ^ n11701 ;
  assign n11704 = n11703 ^ x5 ;
  assign n11700 = n3840 & n10342 ;
  assign n11705 = n11704 ^ n11700 ;
  assign n11699 = ~n408 & n10327 ;
  assign n11706 = n11705 ^ n11699 ;
  assign n11707 = n11706 ^ x2 ;
  assign n11714 = n11713 ^ n11707 ;
  assign n11716 = n11715 ^ n11714 ;
  assign n10972 = n10971 ^ n10970 ;
  assign n10411 = x2 & ~n408 ;
  assign n10412 = n10411 ^ n3505 ;
  assign n10413 = ~x1 & ~n10412 ;
  assign n10407 = n3505 ^ x2 ;
  assign n10401 = n368 ^ x1 ;
  assign n10400 = n368 ^ x2 ;
  assign n10402 = n10401 ^ n10400 ;
  assign n10403 = n3513 & n10402 ;
  assign n10404 = n10403 ^ n10401 ;
  assign n10408 = n10407 ^ n10404 ;
  assign n10414 = n10413 ^ n10408 ;
  assign n10415 = ~x0 & n10414 ;
  assign n10416 = n10415 ^ n10404 ;
  assign n10973 = n10972 ^ n10416 ;
  assign n11632 = n10958 ^ n10427 ;
  assign n11651 = n11632 ^ n10416 ;
  assign n10990 = n10955 ^ n10440 ;
  assign n10977 = n408 ^ x1 ;
  assign n10976 = n408 ^ x2 ;
  assign n10978 = n10977 ^ n10976 ;
  assign n10979 = n3811 & n10978 ;
  assign n10980 = n10979 ^ n10977 ;
  assign n10991 = n10990 ^ n10980 ;
  assign n10985 = x2 & ~n698 ;
  assign n10986 = n10985 ^ n540 ;
  assign n10987 = ~x1 & ~n10986 ;
  assign n10981 = n540 ^ x2 ;
  assign n10982 = n10981 ^ n10980 ;
  assign n10988 = n10987 ^ n10982 ;
  assign n10989 = ~x0 & n10988 ;
  assign n10992 = n10991 ^ n10989 ;
  assign n11008 = n10952 ^ n10453 ;
  assign n10995 = n540 ^ x1 ;
  assign n10996 = n10995 ^ n10981 ;
  assign n10997 = n3955 & n10996 ;
  assign n10998 = n10997 ^ n10995 ;
  assign n11009 = n11008 ^ n10998 ;
  assign n11003 = x2 & ~n856 ;
  assign n11004 = n11003 ^ n698 ;
  assign n11005 = ~x1 & ~n11004 ;
  assign n10999 = n698 ^ x2 ;
  assign n11000 = n10999 ^ n10998 ;
  assign n11006 = n11005 ^ n11000 ;
  assign n11007 = ~x0 & n11006 ;
  assign n11010 = n11009 ^ n11007 ;
  assign n11024 = n10950 ^ n10940 ;
  assign n11013 = n3495 & n11012 ;
  assign n11014 = n11013 ^ n10999 ;
  assign n11025 = n11024 ^ n11014 ;
  assign n11016 = x2 & n1119 ;
  assign n11017 = n11016 ^ n11014 ;
  assign n11011 = n856 ^ x2 ;
  assign n11015 = n11014 ^ n11011 ;
  assign n11018 = n11017 ^ n11015 ;
  assign n11019 = n11017 ^ x1 ;
  assign n11020 = n11019 ^ n11017 ;
  assign n11021 = ~n11018 & n11020 ;
  assign n11022 = n11021 ^ n11017 ;
  assign n11023 = ~x0 & ~n11022 ;
  assign n11026 = n11025 ^ n11023 ;
  assign n11141 = ~x0 & x1 ;
  assign n11574 = n1119 ^ x2 ;
  assign n11615 = n11141 & ~n11574 ;
  assign n11138 = ~x0 & ~x1 ;
  assign n11139 = x2 & n11138 ;
  assign n11614 = n1248 & n11139 ;
  assign n11616 = n11615 ^ n11614 ;
  assign n11607 = n11011 ^ n3493 ;
  assign n11608 = n11607 ^ n11011 ;
  assign n11611 = n11012 & n11608 ;
  assign n11612 = n11611 ^ n11011 ;
  assign n11613 = x0 & ~n11612 ;
  assign n11617 = n11616 ^ n11613 ;
  assign n11622 = n11617 ^ n11024 ;
  assign n11573 = n1119 ^ x1 ;
  assign n11575 = n11574 ^ n11573 ;
  assign n11576 = ~n4335 & n11575 ;
  assign n11577 = n11576 ^ n11573 ;
  assign n11554 = n1248 ^ x2 ;
  assign n11579 = n11577 ^ n11554 ;
  assign n11580 = n11579 ^ n11577 ;
  assign n11581 = n11580 ^ n1248 ;
  assign n11582 = ~n990 & n11581 ;
  assign n11583 = n11582 ^ n1248 ;
  assign n11584 = ~x1 & ~n11583 ;
  assign n11585 = n11584 ^ n11579 ;
  assign n11586 = ~x0 & n11585 ;
  assign n11587 = n11586 ^ n11577 ;
  assign n11035 = n1345 ^ x2 ;
  assign n11545 = ~n11035 & n11141 ;
  assign n11544 = n1450 & n11139 ;
  assign n11546 = n11545 ^ n11544 ;
  assign n11541 = ~n3486 & n11012 ;
  assign n11536 = n990 ^ x2 ;
  assign n11542 = n11541 ^ n11536 ;
  assign n11543 = x0 & ~n11542 ;
  assign n11547 = n11546 ^ n11543 ;
  assign n11040 = n10900 ^ n10494 ;
  assign n11548 = n11547 ^ n11040 ;
  assign n11034 = ~n3483 & n11012 ;
  assign n11036 = n11035 ^ n11034 ;
  assign n11041 = n11040 ^ n11036 ;
  assign n11029 = n1450 ^ x2 ;
  assign n11037 = n11036 ^ n11029 ;
  assign n11031 = x2 & ~n1751 ;
  assign n11032 = n11031 ^ n1450 ;
  assign n11033 = ~x1 & ~n11032 ;
  assign n11038 = n11037 ^ n11033 ;
  assign n11039 = ~x0 & n11038 ;
  assign n11042 = n11041 ^ n11039 ;
  assign n11057 = n10897 ^ n10507 ;
  assign n11533 = n11057 ^ n11040 ;
  assign n11044 = n1450 ^ x1 ;
  assign n11045 = n11044 ^ n11029 ;
  assign n11046 = ~n4494 & n11045 ;
  assign n11047 = n11046 ^ n11044 ;
  assign n11058 = n11057 ^ n11047 ;
  assign n11052 = x2 & ~n1670 ;
  assign n11053 = n11052 ^ n1751 ;
  assign n11054 = ~x1 & ~n11053 ;
  assign n11048 = n1751 ^ x2 ;
  assign n11049 = n11048 ^ n11047 ;
  assign n11055 = n11054 ^ n11049 ;
  assign n11056 = ~x0 & n11055 ;
  assign n11059 = n11058 ^ n11056 ;
  assign n11086 = x2 & n1819 ;
  assign n11076 = ~x2 & n4492 ;
  assign n11080 = n11076 ^ n4492 ;
  assign n11081 = n11080 ^ n1751 ;
  assign n11087 = n11086 ^ n11081 ;
  assign n11088 = ~x0 & ~n11087 ;
  assign n11089 = n11088 ^ n11081 ;
  assign n11068 = n1670 ^ x2 ;
  assign n11090 = n11089 ^ n11068 ;
  assign n11077 = n11076 ^ n1751 ;
  assign n11078 = n11077 ^ n11068 ;
  assign n11079 = x0 & ~n11078 ;
  assign n11091 = n11090 ^ n11079 ;
  assign n11092 = x1 & n11091 ;
  assign n11093 = n11092 ^ n11089 ;
  assign n11530 = n11093 ^ n11057 ;
  assign n11073 = n10891 ^ n10529 ;
  assign n11067 = ~n4985 & n11012 ;
  assign n11069 = n11068 ^ n11067 ;
  assign n11074 = n11073 ^ n11069 ;
  assign n11060 = n1819 ^ x2 ;
  assign n11070 = n11069 ^ n11060 ;
  assign n11064 = x2 & ~n1541 ;
  assign n11065 = n11064 ^ n1819 ;
  assign n11066 = ~x1 & ~n11065 ;
  assign n11071 = n11070 ^ n11066 ;
  assign n11072 = ~x0 & n11071 ;
  assign n11075 = n11074 ^ n11072 ;
  assign n11111 = n10888 ^ n10539 ;
  assign n11098 = n1819 ^ x1 ;
  assign n11099 = n11098 ^ n11060 ;
  assign n11100 = ~n4488 & n11099 ;
  assign n11101 = n11100 ^ n11098 ;
  assign n11112 = n11111 ^ n11101 ;
  assign n11106 = x2 & ~n1972 ;
  assign n11107 = n11106 ^ n1541 ;
  assign n11108 = ~x1 & ~n11107 ;
  assign n11102 = n1541 ^ x2 ;
  assign n11103 = n11102 ^ n11101 ;
  assign n11109 = n11108 ^ n11103 ;
  assign n11110 = ~x0 & n11109 ;
  assign n11113 = n11112 ^ n11110 ;
  assign n11116 = n1541 ^ x1 ;
  assign n11117 = n11116 ^ n11102 ;
  assign n11118 = ~n4891 & n11117 ;
  assign n11119 = n11118 ^ n11116 ;
  assign n11114 = n10885 ^ n10549 ;
  assign n11129 = n11119 ^ n11114 ;
  assign n11124 = x2 & ~n1897 ;
  assign n11125 = n11124 ^ n1972 ;
  assign n11126 = ~x1 & ~n11125 ;
  assign n11120 = n1972 ^ x2 ;
  assign n11121 = n11120 ^ n11119 ;
  assign n11127 = n11126 ^ n11121 ;
  assign n11128 = ~x0 & n11127 ;
  assign n11130 = n11129 ^ n11128 ;
  assign n11145 = n10883 ^ n10873 ;
  assign n11142 = n1897 ^ x2 ;
  assign n11143 = n11141 & ~n11142 ;
  assign n11140 = n2095 & n11139 ;
  assign n11144 = n11143 ^ n11140 ;
  assign n11146 = n11145 ^ n11144 ;
  assign n11135 = n5286 & n11012 ;
  assign n11136 = n11135 ^ n11120 ;
  assign n11137 = x0 & ~n11136 ;
  assign n11147 = n11146 ^ n11137 ;
  assign n11157 = ~n4884 & n11012 ;
  assign n11158 = n11157 ^ n11142 ;
  assign n11148 = n10870 ^ n10560 ;
  assign n11162 = n11158 ^ n11148 ;
  assign n11152 = n2095 ^ x2 ;
  assign n11159 = n11158 ^ n11152 ;
  assign n11154 = x2 & ~n2199 ;
  assign n11155 = n11154 ^ n2095 ;
  assign n11156 = ~x1 & ~n11155 ;
  assign n11160 = n11159 ^ n11156 ;
  assign n11161 = ~x0 & n11160 ;
  assign n11163 = n11162 ^ n11161 ;
  assign n11174 = n2199 ^ x2 ;
  assign n11175 = n11141 & ~n11174 ;
  assign n11173 = n2288 & n11139 ;
  assign n11176 = n11175 ^ n11173 ;
  assign n11164 = n10868 ^ n10858 ;
  assign n11177 = n11176 ^ n11164 ;
  assign n11170 = ~n5759 & n11012 ;
  assign n11171 = n11170 ^ n11152 ;
  assign n11172 = x0 & ~n11171 ;
  assign n11178 = n11177 ^ n11172 ;
  assign n11183 = n2199 ^ x1 ;
  assign n11184 = n11183 ^ n11174 ;
  assign n11185 = n5479 & n11184 ;
  assign n11186 = n11185 ^ n11183 ;
  assign n11179 = n10855 ^ n10571 ;
  assign n11196 = n11186 ^ n11179 ;
  assign n11191 = x2 & ~n2371 ;
  assign n11192 = n11191 ^ n2288 ;
  assign n11193 = ~x1 & ~n11192 ;
  assign n11187 = n2288 ^ x2 ;
  assign n11188 = n11187 ^ n11186 ;
  assign n11194 = n11193 ^ n11188 ;
  assign n11195 = ~x0 & n11194 ;
  assign n11197 = n11196 ^ n11195 ;
  assign n11202 = n2288 ^ x1 ;
  assign n11203 = n11202 ^ n11187 ;
  assign n11204 = n5814 & n11203 ;
  assign n11205 = n11204 ^ n11202 ;
  assign n11198 = n10853 ^ n10843 ;
  assign n11215 = n11205 ^ n11198 ;
  assign n11210 = x2 & ~n2467 ;
  assign n11211 = n11210 ^ n2371 ;
  assign n11212 = ~x1 & ~n11211 ;
  assign n11206 = n2371 ^ x2 ;
  assign n11207 = n11206 ^ n11205 ;
  assign n11213 = n11212 ^ n11207 ;
  assign n11214 = ~x0 & n11213 ;
  assign n11216 = n11215 ^ n11214 ;
  assign n11245 = n10828 ^ n10818 ;
  assign n11223 = x2 & n2552 ;
  assign n11217 = n2371 ^ x1 ;
  assign n11218 = n11217 ^ n11206 ;
  assign n11219 = n5695 & n11218 ;
  assign n11220 = n11219 ^ n11217 ;
  assign n11224 = n11223 ^ n11220 ;
  assign n11221 = n2467 ^ x2 ;
  assign n11222 = n11221 ^ n11220 ;
  assign n11225 = n11224 ^ n11222 ;
  assign n11226 = n11224 ^ x1 ;
  assign n11227 = n11226 ^ n11224 ;
  assign n11228 = ~n11225 & n11227 ;
  assign n11229 = n11228 ^ n11224 ;
  assign n11230 = ~x0 & ~n11229 ;
  assign n11231 = n11230 ^ n11220 ;
  assign n11502 = n11245 ^ n11231 ;
  assign n11240 = ~n6007 & n11012 ;
  assign n11241 = n11240 ^ n11221 ;
  assign n11246 = n11245 ^ n11241 ;
  assign n11235 = n2552 ^ x2 ;
  assign n11242 = n11241 ^ n11235 ;
  assign n11237 = x2 & ~n2589 ;
  assign n11238 = n11237 ^ n2552 ;
  assign n11239 = ~x1 & ~n11238 ;
  assign n11243 = n11242 ^ n11239 ;
  assign n11244 = ~x0 & n11243 ;
  assign n11247 = n11246 ^ n11244 ;
  assign n11263 = n10815 ^ n10583 ;
  assign n11499 = n11263 ^ n11245 ;
  assign n11250 = n2552 ^ x1 ;
  assign n11251 = n11250 ^ n11235 ;
  assign n11252 = n6211 & n11251 ;
  assign n11253 = n11252 ^ n11250 ;
  assign n11264 = n11263 ^ n11253 ;
  assign n11258 = x2 & ~n2657 ;
  assign n11259 = n11258 ^ n2589 ;
  assign n11260 = ~x1 & ~n11259 ;
  assign n11254 = n2589 ^ x2 ;
  assign n11255 = n11254 ^ n11253 ;
  assign n11261 = n11260 ^ n11255 ;
  assign n11262 = ~x0 & n11261 ;
  assign n11265 = n11264 ^ n11262 ;
  assign n11270 = n2589 ^ x1 ;
  assign n11271 = n11270 ^ n11254 ;
  assign n11272 = n6078 & n11271 ;
  assign n11273 = n11272 ^ n11270 ;
  assign n11266 = n10812 ^ n10596 ;
  assign n11283 = n11273 ^ n11266 ;
  assign n11278 = x2 & ~n2712 ;
  assign n11279 = n11278 ^ n2657 ;
  assign n11280 = ~x1 & ~n11279 ;
  assign n11274 = n2657 ^ x2 ;
  assign n11275 = n11274 ^ n11273 ;
  assign n11281 = n11280 ^ n11275 ;
  assign n11282 = ~x0 & n11281 ;
  assign n11284 = n11283 ^ n11282 ;
  assign n11289 = n2657 ^ x1 ;
  assign n11290 = n11289 ^ n11274 ;
  assign n11291 = n6228 & n11290 ;
  assign n11292 = n11291 ^ n11289 ;
  assign n11285 = n10810 ^ n10800 ;
  assign n11302 = n11292 ^ n11285 ;
  assign n11297 = x2 & ~n3324 ;
  assign n11298 = n11297 ^ n2712 ;
  assign n11299 = ~x1 & ~n11298 ;
  assign n11293 = n2712 ^ x2 ;
  assign n11294 = n11293 ^ n11292 ;
  assign n11300 = n11299 ^ n11294 ;
  assign n11301 = ~x0 & n11300 ;
  assign n11303 = n11302 ^ n11301 ;
  assign n11314 = x2 & ~n2748 ;
  assign n11315 = n11314 ^ n3324 ;
  assign n11316 = ~x1 & ~n11315 ;
  assign n11310 = n3324 ^ x2 ;
  assign n11304 = n2712 ^ x1 ;
  assign n11305 = n11304 ^ n11293 ;
  assign n11306 = n6622 & n11305 ;
  assign n11307 = n11306 ^ n11304 ;
  assign n11311 = n11310 ^ n11307 ;
  assign n11317 = n11316 ^ n11311 ;
  assign n11318 = ~x0 & n11317 ;
  assign n11319 = n11318 ^ n11307 ;
  assign n11321 = n11319 ^ n10797 ;
  assign n11322 = n11321 ^ n10607 ;
  assign n11334 = x2 & ~n2839 ;
  assign n11335 = n11334 ^ n2748 ;
  assign n11336 = ~x1 & ~n11335 ;
  assign n11330 = n2748 ^ x2 ;
  assign n11323 = n3324 ^ x1 ;
  assign n11324 = n11323 ^ x2 ;
  assign n11325 = n11324 ^ n3324 ;
  assign n11326 = n6643 & n11325 ;
  assign n11327 = n11326 ^ n11323 ;
  assign n11331 = n11330 ^ n11327 ;
  assign n11337 = n11336 ^ n11331 ;
  assign n11338 = ~x0 & n11337 ;
  assign n11339 = n11338 ^ n11327 ;
  assign n11341 = n11339 ^ n10794 ;
  assign n11342 = n11341 ^ n10619 ;
  assign n11378 = n10789 ^ n10779 ;
  assign n11353 = x2 & ~n2935 ;
  assign n11354 = n11353 ^ n2839 ;
  assign n11355 = ~x1 & ~n11354 ;
  assign n11349 = n2839 ^ x2 ;
  assign n11343 = n2748 ^ x1 ;
  assign n11344 = n11343 ^ n11330 ;
  assign n11345 = ~n6301 & n11344 ;
  assign n11346 = n11345 ^ n11343 ;
  assign n11350 = n11349 ^ n11346 ;
  assign n11356 = n11355 ^ n11350 ;
  assign n11357 = ~x0 & n11356 ;
  assign n11358 = n11357 ^ n11346 ;
  assign n11484 = n11378 ^ n11358 ;
  assign n11367 = x2 & n3248 ;
  assign n11360 = x2 & ~n3439 ;
  assign n11362 = n11360 ^ n2839 ;
  assign n11368 = n11367 ^ n11362 ;
  assign n11369 = ~x0 & ~n11368 ;
  assign n11370 = n11369 ^ n11362 ;
  assign n11379 = n11378 ^ n11370 ;
  assign n11372 = n2935 ^ x2 ;
  assign n11373 = n11372 ^ n11370 ;
  assign n11361 = n11360 ^ n6695 ;
  assign n11371 = n11370 ^ n11361 ;
  assign n11374 = n11373 ^ n11371 ;
  assign n11375 = x0 & n11374 ;
  assign n11376 = n11375 ^ n11373 ;
  assign n11377 = x1 & n11376 ;
  assign n11380 = n11379 ^ n11377 ;
  assign n11456 = ~n3429 & n8137 ;
  assign n10761 = n10678 ^ n10657 ;
  assign n11457 = n11456 ^ n10761 ;
  assign n11481 = n11457 ^ n11378 ;
  assign n11436 = n3248 ^ x1 ;
  assign n11435 = n3248 ^ x2 ;
  assign n11437 = n11436 ^ n11435 ;
  assign n11438 = n6749 & n11437 ;
  assign n11439 = n11438 ^ n11436 ;
  assign n11382 = n3022 ^ x2 ;
  assign n11442 = n11439 ^ n11382 ;
  assign n11443 = n11442 ^ n11439 ;
  assign n11444 = n11443 ^ n3022 ;
  assign n11445 = ~n3055 & n11444 ;
  assign n11446 = n11445 ^ n3022 ;
  assign n11447 = ~x1 & ~n11446 ;
  assign n11448 = n11447 ^ n11442 ;
  assign n11449 = ~x0 & n11448 ;
  assign n11450 = n11449 ^ n11439 ;
  assign n11458 = n11457 ^ n11450 ;
  assign n11395 = n10324 ^ x4 ;
  assign n11396 = ~n3429 & n11395 ;
  assign n11397 = n11396 ^ n10633 ;
  assign n11451 = n11450 ^ n11397 ;
  assign n11381 = n3022 ^ x1 ;
  assign n11383 = n11382 ^ n11381 ;
  assign n11384 = n6839 & n11383 ;
  assign n11385 = n11384 ^ n11381 ;
  assign n11398 = n11397 ^ n11385 ;
  assign n11390 = x2 & ~n3196 ;
  assign n11391 = n11390 ^ n3055 ;
  assign n11392 = ~x1 & ~n11391 ;
  assign n11386 = n3055 ^ x2 ;
  assign n11387 = n11386 ^ n11385 ;
  assign n11393 = n11392 ^ n11387 ;
  assign n11394 = ~x0 & n11393 ;
  assign n11399 = n11398 ^ n11394 ;
  assign n11414 = x2 & n3124 ;
  assign n11415 = n11138 ^ n3429 ;
  assign n11404 = n3196 ^ x3 ;
  assign n11418 = n11138 & n11404 ;
  assign n11419 = n11418 ^ n3196 ;
  assign n11420 = n11415 & ~n11419 ;
  assign n11421 = n11420 ^ n3429 ;
  assign n11422 = n11414 & n11421 ;
  assign n11400 = ~x0 & n10322 ;
  assign n11401 = n11400 ^ n10322 ;
  assign n11402 = n11401 ^ x1 ;
  assign n11403 = n11402 ^ n11401 ;
  assign n11409 = n11400 & n11404 ;
  assign n11410 = n11403 & n11409 ;
  assign n11411 = n11410 ^ n11403 ;
  assign n11412 = n11411 ^ n11402 ;
  assign n11413 = ~n3429 & n11412 ;
  assign n11423 = n11422 ^ n11413 ;
  assign n11432 = n11423 ^ n11397 ;
  assign n11424 = x0 & n11423 ;
  assign n11429 = ~n6863 & n11012 ;
  assign n11430 = n11429 ^ n11386 ;
  assign n11431 = n11424 & n11430 ;
  assign n11433 = n11432 ^ n11431 ;
  assign n11434 = ~n11399 & n11433 ;
  assign n11452 = n11451 ^ n11434 ;
  assign n11453 = n11450 ^ n10648 ;
  assign n11454 = n11453 ^ n10636 ;
  assign n11455 = ~n11452 & ~n11454 ;
  assign n11459 = n11458 ^ n11455 ;
  assign n11467 = ~x1 & ~n3437 ;
  assign n11468 = n11467 ^ n2935 ;
  assign n11477 = n11468 ^ n11457 ;
  assign n11470 = n11468 ^ n3022 ;
  assign n11469 = n11468 ^ n3248 ;
  assign n11471 = n11470 ^ n11469 ;
  assign n11474 = x1 & n11471 ;
  assign n11475 = n11474 ^ n11470 ;
  assign n11476 = ~x0 & n11475 ;
  assign n11478 = n11477 ^ n11476 ;
  assign n11460 = n3437 ^ x0 ;
  assign n11461 = n11460 ^ n3437 ;
  assign n11462 = ~x1 & ~n3022 ;
  assign n11463 = n11462 ^ n3437 ;
  assign n11464 = ~n11461 & ~n11463 ;
  assign n11465 = n11464 ^ n3437 ;
  assign n11466 = ~x2 & n11465 ;
  assign n11479 = n11478 ^ n11466 ;
  assign n11480 = ~n11459 & n11479 ;
  assign n11482 = n11481 ^ n11480 ;
  assign n11483 = n11380 & ~n11482 ;
  assign n11485 = n11484 ^ n11483 ;
  assign n11486 = n11358 ^ n10629 ;
  assign n11487 = n11486 ^ n10791 ;
  assign n11488 = n11485 & n11487 ;
  assign n11359 = n11358 ^ n11339 ;
  assign n11489 = n11488 ^ n11359 ;
  assign n11490 = ~n11342 & n11489 ;
  assign n11340 = n11339 ^ n11319 ;
  assign n11491 = n11490 ^ n11340 ;
  assign n11492 = n11322 & n11491 ;
  assign n11320 = n11319 ^ n11285 ;
  assign n11493 = n11492 ^ n11320 ;
  assign n11494 = ~n11303 & ~n11493 ;
  assign n11286 = n11285 ^ n11266 ;
  assign n11495 = n11494 ^ n11286 ;
  assign n11496 = ~n11284 & n11495 ;
  assign n11267 = n11266 ^ n11263 ;
  assign n11497 = n11496 ^ n11267 ;
  assign n11498 = ~n11265 & n11497 ;
  assign n11500 = n11499 ^ n11498 ;
  assign n11501 = ~n11247 & n11500 ;
  assign n11503 = n11502 ^ n11501 ;
  assign n11504 = n11231 ^ n10841 ;
  assign n11505 = n11504 ^ n10830 ;
  assign n11506 = ~n11503 & n11505 ;
  assign n11232 = n11231 ^ n11198 ;
  assign n11507 = n11506 ^ n11232 ;
  assign n11508 = ~n11216 & ~n11507 ;
  assign n11199 = n11198 ^ n11179 ;
  assign n11509 = n11508 ^ n11199 ;
  assign n11510 = ~n11197 & n11509 ;
  assign n11180 = n11179 ^ n11164 ;
  assign n11511 = n11510 ^ n11180 ;
  assign n11512 = n11178 & n11511 ;
  assign n11165 = n11164 ^ n11148 ;
  assign n11513 = n11512 ^ n11165 ;
  assign n11514 = n11163 & ~n11513 ;
  assign n11149 = n11148 ^ n11145 ;
  assign n11515 = n11514 ^ n11149 ;
  assign n11516 = ~n11147 & n11515 ;
  assign n11517 = n11516 ^ n11145 ;
  assign n11518 = n11517 ^ n11114 ;
  assign n11519 = n11130 & n11518 ;
  assign n11115 = n11114 ^ n11111 ;
  assign n11520 = n11519 ^ n11115 ;
  assign n11521 = n11113 & n11520 ;
  assign n11522 = n11521 ^ n11111 ;
  assign n11094 = n11093 ^ n11073 ;
  assign n11095 = n11094 ^ n11093 ;
  assign n11523 = n11522 ^ n11095 ;
  assign n11524 = n11075 & n11523 ;
  assign n11525 = n11524 ^ n11094 ;
  assign n11526 = n11093 ^ n10518 ;
  assign n11527 = n11526 ^ n10517 ;
  assign n11528 = n11527 ^ n10894 ;
  assign n11529 = n11525 & ~n11528 ;
  assign n11531 = n11530 ^ n11529 ;
  assign n11532 = n11059 & n11531 ;
  assign n11534 = n11533 ^ n11532 ;
  assign n11535 = n11042 & n11534 ;
  assign n11549 = n11548 ^ n11535 ;
  assign n11550 = n11547 ^ n10903 ;
  assign n11551 = n11550 ^ n10484 ;
  assign n11552 = ~n11549 & n11551 ;
  assign n11553 = n11552 ^ n11547 ;
  assign n11555 = n1248 ^ x1 ;
  assign n11556 = n11555 ^ n11554 ;
  assign n11557 = n4333 & n11556 ;
  assign n11558 = n11557 ^ n11555 ;
  assign n11561 = n11558 ^ n11536 ;
  assign n11562 = n11561 ^ n11558 ;
  assign n11563 = n11562 ^ n990 ;
  assign n11564 = ~n1345 & n11563 ;
  assign n11565 = n11564 ^ n990 ;
  assign n11566 = ~x1 & ~n11565 ;
  assign n11567 = n11566 ^ n11561 ;
  assign n11568 = ~x0 & n11567 ;
  assign n11569 = n11568 ^ n11558 ;
  assign n11571 = n11553 & ~n11569 ;
  assign n11570 = n11569 ^ n11553 ;
  assign n11572 = n11571 ^ n11570 ;
  assign n11588 = n11587 ^ n11572 ;
  assign n11589 = n10920 & ~n10935 ;
  assign n11590 = n11589 ^ n10922 ;
  assign n11591 = n11590 ^ n11572 ;
  assign n11592 = n11591 ^ n10935 ;
  assign n11593 = n11588 & ~n11592 ;
  assign n11594 = n11593 ^ n11587 ;
  assign n11595 = n11589 ^ n11571 ;
  assign n11596 = n11587 ^ n10907 ;
  assign n11597 = n11596 ^ n10935 ;
  assign n11598 = n11587 ^ n11571 ;
  assign n11599 = n11598 ^ n10918 ;
  assign n11600 = n11598 ^ n11587 ;
  assign n11601 = n11599 & ~n11600 ;
  assign n11602 = n11597 & n11601 ;
  assign n11603 = n11602 ^ n11598 ;
  assign n11604 = ~n11595 & ~n11603 ;
  assign n11605 = n11604 ^ n11571 ;
  assign n11606 = ~n11594 & n11605 ;
  assign n11618 = n11617 ^ n11606 ;
  assign n11619 = n11606 ^ n10468 ;
  assign n11620 = n11619 ^ n10937 ;
  assign n11621 = n11618 & n11620 ;
  assign n11623 = n11622 ^ n11621 ;
  assign n11624 = ~n11026 & n11623 ;
  assign n11625 = n11624 ^ n11024 ;
  assign n11626 = n11625 ^ n11008 ;
  assign n11627 = n11010 & ~n11626 ;
  assign n11628 = n11627 ^ n11008 ;
  assign n11629 = n11628 ^ n10990 ;
  assign n11630 = ~n10992 & ~n11629 ;
  assign n11631 = n11630 ^ n10990 ;
  assign n11633 = n11632 ^ n11631 ;
  assign n11636 = n3505 ^ x1 ;
  assign n11637 = n11636 ^ n10407 ;
  assign n11638 = n3839 & n11637 ;
  assign n11639 = n11638 ^ n11636 ;
  assign n11648 = n11639 ^ n11632 ;
  assign n11640 = n11639 ^ n10976 ;
  assign n11641 = n11640 ^ n11639 ;
  assign n11642 = n11641 ^ n408 ;
  assign n11643 = ~n540 & n11642 ;
  assign n11644 = n11643 ^ n408 ;
  assign n11645 = ~x1 & ~n11644 ;
  assign n11646 = n11645 ^ n11640 ;
  assign n11647 = ~x0 & n11646 ;
  assign n11649 = n11648 ^ n11647 ;
  assign n11650 = ~n11633 & n11649 ;
  assign n11652 = n11651 ^ n11650 ;
  assign n11653 = n10973 & ~n11652 ;
  assign n11654 = n11653 ^ n10972 ;
  assign n11655 = n10314 ^ n9918 ;
  assign n11657 = x0 & x1 ;
  assign n11658 = ~n3510 & n11657 ;
  assign n11659 = n11658 ^ x2 ;
  assign n11660 = ~n368 & n11659 ;
  assign n11661 = n11660 ^ x2 ;
  assign n11662 = n3505 & n11661 ;
  assign n11663 = x0 & x2 ;
  assign n11683 = n368 & n3512 ;
  assign n11684 = n11657 & n11683 ;
  assign n11686 = x1 & x2 ;
  assign n11687 = n11684 & n11686 ;
  assign n11664 = x2 ^ x0 ;
  assign n11667 = n10400 ^ x1 ;
  assign n11665 = n11664 ^ n10400 ;
  assign n11671 = n11667 ^ n11665 ;
  assign n11675 = n11671 ^ x2 ;
  assign n11676 = n11664 & n11675 ;
  assign n11677 = n11676 ^ n11671 ;
  assign n11678 = n10400 ^ n3505 ;
  assign n11679 = n11676 ^ n11664 ;
  assign n11680 = ~n11678 & n11679 ;
  assign n11681 = n11680 ^ n10400 ;
  assign n11682 = n11677 & ~n11681 ;
  assign n11685 = n11684 ^ n11682 ;
  assign n11688 = n11687 ^ n11685 ;
  assign n11689 = n11663 & ~n11688 ;
  assign n11690 = n3510 ^ n368 ;
  assign n11691 = n11690 ^ n3510 ;
  assign n11692 = n3511 & ~n11691 ;
  assign n11693 = n11692 ^ n3510 ;
  assign n11694 = n11689 & ~n11693 ;
  assign n11695 = n11694 ^ n11688 ;
  assign n11696 = ~n11662 & ~n11695 ;
  assign n11697 = n11655 & ~n11696 ;
  assign n11717 = n11716 ^ n11697 ;
  assign n11730 = n11729 ^ n11717 ;
  assign n11731 = n11730 ^ n11717 ;
  assign n11732 = ~n11716 & ~n11720 ;
  assign n11733 = n11732 ^ n11717 ;
  assign n11734 = ~n11731 & ~n11733 ;
  assign n11735 = n11734 ^ n11717 ;
  assign n11736 = ~n11654 & ~n11735 ;
  assign n11738 = n11737 ^ n11736 ;
  assign n11739 = n11696 ^ n11655 ;
  assign n11740 = n11739 ^ n11717 ;
  assign n11741 = ~n11738 & n11740 ;
  assign n11742 = n11696 ^ n11654 ;
  assign n11747 = ~n11739 & ~n11742 ;
  assign n11748 = n11747 ^ n11655 ;
  assign n11749 = ~n11741 & ~n11748 ;
  assign n11752 = ~n11716 & n11749 ;
  assign n11753 = n11751 & n11752 ;
  assign n11750 = n11749 ^ n11741 ;
  assign n11754 = n11753 ^ n11750 ;
  assign n11756 = n11755 ^ n11754 ;
  assign n11759 = n11755 ^ n11706 ;
  assign n11757 = n11715 ^ n11706 ;
  assign n11758 = n11714 & ~n11757 ;
  assign n11760 = n11759 ^ n11758 ;
  assign n11761 = ~n11756 & n11760 ;
  assign n11762 = n11761 ^ n11755 ;
  assign n11763 = ~n10389 & ~n11762 ;
  assign n11764 = n11763 ^ n11762 ;
  assign n11765 = n11764 ^ n10381 ;
  assign n11766 = n11765 ^ n11764 ;
  assign n11769 = n11764 ^ n10392 ;
  assign n11770 = n11769 ^ n11764 ;
  assign n11771 = n11763 & ~n11770 ;
  assign n11772 = ~n11766 & n11771 ;
  assign n11773 = n11772 ^ n11766 ;
  assign n11774 = n11773 ^ n11765 ;
  assign n11775 = ~n10399 & n11774 ;
  assign n11776 = n10378 ^ n10357 ;
  assign n11777 = n10380 & n11776 ;
  assign n11778 = n11777 ^ n10378 ;
  assign n11779 = n11778 ^ n11775 ;
  assign n11780 = n8475 ^ n8465 ;
  assign n11781 = n11780 ^ n11778 ;
  assign n11782 = ~n11779 & ~n11781 ;
  assign n11783 = ~n11775 & n11782 ;
  assign n11796 = n8477 ^ n8167 ;
  assign n11808 = n11796 ^ n11782 ;
  assign n11787 = ~n408 & n8144 ;
  assign n11786 = ~n368 & n8484 ;
  assign n11788 = n11787 ^ n11786 ;
  assign n11789 = n11788 ^ x8 ;
  assign n11785 = n4398 & n8150 ;
  assign n11790 = n11789 ^ n11785 ;
  assign n11784 = ~n3505 & n8139 ;
  assign n11791 = n11790 ^ n11784 ;
  assign n11792 = n10368 ^ n10367 ;
  assign n11793 = n10377 & ~n11792 ;
  assign n11794 = n11793 ^ n10376 ;
  assign n11795 = n11791 & n11794 ;
  assign n11797 = n11796 ^ n11795 ;
  assign n11799 = n11795 ^ n11780 ;
  assign n11798 = n11795 ^ n11775 ;
  assign n11800 = n11799 ^ n11798 ;
  assign n11801 = n11799 ^ n11775 ;
  assign n11802 = n11801 ^ n11778 ;
  assign n11803 = n11802 ^ n11799 ;
  assign n11804 = n11800 & ~n11803 ;
  assign n11805 = n11804 ^ n11799 ;
  assign n11806 = n11797 & ~n11805 ;
  assign n11807 = n11806 ^ n11796 ;
  assign n11809 = n11794 ^ n11791 ;
  assign n11810 = n11809 ^ n11795 ;
  assign n11811 = ~n11807 & n11810 ;
  assign n11812 = n11808 & n11811 ;
  assign n11813 = n11812 ^ n11807 ;
  assign n11814 = n11813 ^ n11807 ;
  assign n11815 = n11783 & n11814 ;
  assign n11816 = n11815 ^ n11813 ;
  assign n11817 = n11816 ^ n8480 ;
  assign n11818 = n8481 & ~n11817 ;
  assign n11819 = n11818 ^ n8480 ;
  assign n11830 = n11829 ^ n11819 ;
  assign n11834 = n8118 ^ n8107 ;
  assign n11835 = n8115 & n11834 ;
  assign n11836 = n11835 ^ n8118 ;
  assign n11831 = n8158 ^ n8119 ;
  assign n11832 = ~n8132 & n11831 ;
  assign n11833 = n11832 ^ n8119 ;
  assign n11838 = n11836 ^ n11833 ;
  assign n11837 = n11833 & ~n11836 ;
  assign n11839 = n11838 ^ n11837 ;
  assign n11841 = n7556 ^ n7303 ;
  assign n11840 = ~n11820 & n11828 ;
  assign n11842 = n11841 ^ n11840 ;
  assign n11843 = ~n11839 & ~n11842 ;
  assign n11844 = n11830 & n11843 ;
  assign n11845 = n11841 ^ n11837 ;
  assign n11847 = n11841 ^ n11828 ;
  assign n11846 = n11841 ^ n11820 ;
  assign n11848 = n11847 ^ n11846 ;
  assign n11849 = n11841 ^ n11819 ;
  assign n11850 = n11849 ^ n11846 ;
  assign n11851 = ~n11848 & n11850 ;
  assign n11852 = n11851 ^ n11846 ;
  assign n11853 = ~n11845 & ~n11852 ;
  assign n11854 = n11853 ^ n11837 ;
  assign n11855 = ~n11844 & ~n11854 ;
  assign n11856 = n11855 ^ n7559 ;
  assign n11857 = n7560 & ~n11856 ;
  assign n11858 = n11857 ^ n7559 ;
  assign n11865 = ~n408 & ~n6547 ;
  assign n11864 = ~n3505 & ~n6529 ;
  assign n11866 = n11865 ^ n11864 ;
  assign n11861 = x13 & ~n3513 ;
  assign n11862 = n11861 ^ n368 ;
  assign n11863 = n6391 & ~n11862 ;
  assign n11867 = n11866 ^ n11863 ;
  assign n11868 = ~x14 & n11867 ;
  assign n11871 = n4398 ^ x13 ;
  assign n11872 = n11871 ^ n4398 ;
  assign n11873 = ~n3513 & n11872 ;
  assign n11874 = n11873 ^ n4398 ;
  assign n11875 = n6537 & n11874 ;
  assign n11869 = n11866 ^ x14 ;
  assign n11876 = n11875 ^ n11869 ;
  assign n11877 = ~n11868 & ~n11876 ;
  assign n11879 = n11858 & ~n11877 ;
  assign n11878 = n11877 ^ n11858 ;
  assign n11880 = n11879 ^ n11878 ;
  assign n11881 = n11879 ^ n7293 ;
  assign n11882 = n7293 ^ n7289 ;
  assign n11883 = n11882 ^ n7284 ;
  assign n11884 = n11883 ^ n7287 ;
  assign n11885 = n11884 ^ n11882 ;
  assign n11886 = n7293 ^ n7284 ;
  assign n11887 = n11886 ^ n11882 ;
  assign n11888 = n11885 & n11887 ;
  assign n11889 = n11888 ^ n11882 ;
  assign n11890 = ~n11881 & n11889 ;
  assign n11891 = n11890 ^ n11879 ;
  assign n11892 = ~n11880 & ~n11891 ;
  assign n11893 = ~n7294 & n11892 ;
  assign n11894 = n11893 ^ n11891 ;
  assign n11895 = n11894 ^ n11891 ;
  assign n11896 = n7292 & n11895 ;
  assign n11897 = n11896 ^ n11894 ;
  assign n11898 = n11897 ^ n7021 ;
  assign n11899 = n7023 & ~n11898 ;
  assign n11900 = n11899 ^ n7022 ;
  assign n11901 = n6389 ^ n6375 ;
  assign n11902 = n11901 ^ n6388 ;
  assign n11903 = n6526 ^ n6525 ;
  assign n11906 = ~n11902 & ~n11903 ;
  assign n11907 = n11906 ^ n6388 ;
  assign n11908 = n11900 & ~n11907 ;
  assign n11909 = ~n6526 & ~n11908 ;
  assign n11910 = n6389 & n11909 ;
  assign n11911 = n11900 ^ n6374 ;
  assign n11912 = n6375 & n11911 ;
  assign n11913 = n11912 ^ n6374 ;
  assign n11914 = ~n11910 & ~n11913 ;
  assign n11916 = ~n6388 & ~n11903 ;
  assign n11917 = n11914 & n11916 ;
  assign n11915 = n11914 ^ n11910 ;
  assign n11918 = n11917 ^ n11915 ;
  assign n5965 = n5964 ^ n5932 ;
  assign n5966 = ~n5937 & ~n5965 ;
  assign n5967 = n5966 ^ n5932 ;
  assign n11920 = n11918 ^ n5967 ;
  assign n11919 = n5967 & n11918 ;
  assign n11921 = n11920 ^ n11919 ;
  assign n11969 = n3840 & n5221 ;
  assign n11966 = ~n3505 & n5220 ;
  assign n11964 = ~n408 & n5426 ;
  assign n11936 = n5943 ^ n5941 ;
  assign n11937 = n5951 & n11936 ;
  assign n11938 = n11937 ^ n5943 ;
  assign n5268 = ~n4435 & n4580 ;
  assign n5266 = ~n1248 & ~n4434 ;
  assign n5263 = ~n1345 & n20603 ;
  assign n5262 = ~n990 & n4600 ;
  assign n5264 = n5263 ^ n5262 ;
  assign n5265 = n5264 ^ x26 ;
  assign n5267 = n5266 ^ n5265 ;
  assign n5269 = n5268 ^ n5267 ;
  assign n5398 = n5396 ^ n5269 ;
  assign n5407 = n5406 ^ n5398 ;
  assign n5408 = n5407 ^ n5269 ;
  assign n5409 = n5397 & ~n5408 ;
  assign n5410 = n5409 ^ n5398 ;
  assign n4904 = n4903 ^ n4856 ;
  assign n4940 = n4904 & ~n4939 ;
  assign n4862 = n4742 ^ n1879 ;
  assign n4863 = n4862 ^ n1167 ;
  assign n4859 = n1785 ^ n628 ;
  assign n4860 = n4859 ^ n903 ;
  assign n4858 = n4857 ^ n1304 ;
  assign n4861 = n4860 ^ n4858 ;
  assign n4864 = n4863 ^ n4861 ;
  assign n4865 = n4864 ^ n870 ;
  assign n4866 = n4865 ^ n538 ;
  assign n4869 = n2755 ^ n189 ;
  assign n4870 = n4869 ^ n125 ;
  assign n4868 = n2807 ^ n974 ;
  assign n4871 = n4870 ^ n4868 ;
  assign n4867 = n1404 ^ n577 ;
  assign n4872 = n4871 ^ n4867 ;
  assign n4873 = n4872 ^ n2804 ;
  assign n4874 = n4873 ^ n2997 ;
  assign n4875 = n4874 ^ n854 ;
  assign n4876 = ~n4866 & ~n4875 ;
  assign n5181 = n4940 ^ n4876 ;
  assign n5178 = ~n1751 & n3985 ;
  assign n5170 = x30 & ~n1541 ;
  assign n5156 = n5154 ^ n1541 ;
  assign n5155 = n5154 ^ n1972 ;
  assign n5157 = n5156 ^ n5155 ;
  assign n5160 = x30 & n5157 ;
  assign n5161 = n5160 ^ n5156 ;
  assign n5162 = ~n3518 & n5161 ;
  assign n5163 = n5162 ^ n5154 ;
  assign n5164 = n5163 ^ n1819 ;
  assign n5165 = n5164 ^ n5163 ;
  assign n5171 = n5170 ^ n5165 ;
  assign n5172 = ~n3518 & ~n5171 ;
  assign n5173 = n5172 ^ n5164 ;
  assign n5174 = ~x31 & n5173 ;
  assign n5175 = n5174 ^ n5163 ;
  assign n5176 = n5175 ^ x29 ;
  assign n5151 = n4494 & n5065 ;
  assign n5152 = n5151 ^ n1450 ;
  assign n5153 = n3833 & ~n5152 ;
  assign n5177 = n5176 ^ n5153 ;
  assign n5179 = n5178 ^ n5177 ;
  assign n5147 = ~n1670 & n3837 ;
  assign n5180 = n5179 ^ n5147 ;
  assign n5261 = n5181 ^ n5180 ;
  assign n11934 = n5410 ^ n5261 ;
  assign n11930 = ~n3930 & n4656 ;
  assign n11929 = ~n1119 & n4651 ;
  assign n11931 = n11930 ^ n11929 ;
  assign n11932 = n11931 ^ x23 ;
  assign n11927 = ~n698 & n4655 ;
  assign n11926 = ~n40 & ~n856 ;
  assign n11928 = n11927 ^ n11926 ;
  assign n11933 = n11932 ^ n11928 ;
  assign n11935 = n11934 ^ n11933 ;
  assign n11962 = n11938 ^ n11935 ;
  assign n11963 = n11962 ^ x20 ;
  assign n11965 = n11964 ^ n11963 ;
  assign n11967 = n11966 ^ n11965 ;
  assign n11961 = ~n540 & n13433 ;
  assign n11968 = n11967 ^ n11961 ;
  assign n11970 = n11969 ^ n11968 ;
  assign n11971 = n5963 ^ n5952 ;
  assign n11972 = ~n5960 & n11971 ;
  assign n11973 = n11972 ^ n5963 ;
  assign n11974 = n11973 ^ n11962 ;
  assign n11975 = ~n11970 & ~n11974 ;
  assign n11976 = n11975 ^ n11962 ;
  assign n11959 = n4398 & n5221 ;
  assign n11956 = ~n368 & n5220 ;
  assign n11954 = ~n408 & n13433 ;
  assign n11950 = ~n540 & n4655 ;
  assign n11947 = ~n40 & ~n698 ;
  assign n11945 = n3968 & n4656 ;
  assign n5270 = n5269 ^ n5261 ;
  assign n5411 = n5270 & ~n5410 ;
  assign n5412 = n5411 ^ n5269 ;
  assign n5259 = ~n4336 & ~n4435 ;
  assign n5256 = ~n990 & n20603 ;
  assign n5254 = ~n1248 & n4600 ;
  assign n5182 = n5181 ^ n5175 ;
  assign n5183 = n5180 & n5182 ;
  assign n5184 = n5183 ^ n5181 ;
  assign n5145 = ~n1450 & n3985 ;
  assign n5001 = ~x30 & ~n1819 ;
  assign n5002 = n5001 ^ n3465 ;
  assign n5003 = ~n3518 & n5002 ;
  assign n4988 = n4986 ^ n1541 ;
  assign n4987 = n4986 ^ n1819 ;
  assign n4989 = n4988 ^ n4987 ;
  assign n4992 = ~x30 & n4989 ;
  assign n4993 = n4992 ^ n4988 ;
  assign n4994 = ~n3518 & ~n4993 ;
  assign n4995 = n4994 ^ n4986 ;
  assign n4996 = n4995 ^ n1670 ;
  assign n5004 = n5003 ^ n4996 ;
  assign n5005 = ~x31 & ~n5004 ;
  assign n5006 = n5005 ^ n4995 ;
  assign n4957 = n1770 ^ n151 ;
  assign n4954 = n2137 ^ n1985 ;
  assign n4955 = n4954 ^ n1495 ;
  assign n4951 = n562 ^ n527 ;
  assign n4952 = n4951 ^ n240 ;
  assign n4949 = n1544 ^ n800 ;
  assign n4950 = n4949 ^ n1036 ;
  assign n4953 = n4952 ^ n4950 ;
  assign n4956 = n4955 ^ n4953 ;
  assign n4958 = n4957 ^ n4956 ;
  assign n4945 = n2510 ^ n377 ;
  assign n4946 = n4945 ^ n598 ;
  assign n4947 = n4946 ^ n4944 ;
  assign n4943 = n4942 ^ n1857 ;
  assign n4948 = n4947 ^ n4943 ;
  assign n4959 = n4958 ^ n4948 ;
  assign n4981 = n4980 ^ n4959 ;
  assign n4982 = ~n1247 & ~n4981 ;
  assign n4983 = n4982 ^ x17 ;
  assign n4877 = n4876 ^ n4856 ;
  assign n4941 = ~n4877 & n4940 ;
  assign n4984 = n4983 ^ n4941 ;
  assign n5140 = n5006 ^ n4984 ;
  assign n5141 = n5140 ^ x29 ;
  assign n5139 = ~n1345 & n4369 ;
  assign n5142 = n5141 ^ n5139 ;
  assign n5138 = ~n1751 & n3837 ;
  assign n5143 = n5142 ^ n5138 ;
  assign n5137 = n3983 & n4475 ;
  assign n5144 = n5143 ^ n5137 ;
  assign n5146 = n5145 ^ n5144 ;
  assign n5252 = n5184 ^ n5146 ;
  assign n5253 = n5252 ^ x26 ;
  assign n5255 = n5254 ^ n5253 ;
  assign n5257 = n5256 ^ n5255 ;
  assign n5251 = ~n1119 & ~n4434 ;
  assign n5258 = n5257 ^ n5251 ;
  assign n5260 = n5259 ^ n5258 ;
  assign n11943 = n5412 ^ n5260 ;
  assign n11944 = n11943 ^ x23 ;
  assign n11946 = n11945 ^ n11944 ;
  assign n11948 = n11947 ^ n11946 ;
  assign n11942 = ~n856 & n4651 ;
  assign n11949 = n11948 ^ n11942 ;
  assign n11951 = n11950 ^ n11949 ;
  assign n11939 = n11938 ^ n11933 ;
  assign n11940 = n11935 & n11939 ;
  assign n11941 = n11940 ^ n11938 ;
  assign n11952 = n11951 ^ n11941 ;
  assign n11953 = n11952 ^ x20 ;
  assign n11955 = n11954 ^ n11953 ;
  assign n11957 = n11956 ^ n11955 ;
  assign n11925 = ~n3505 & n5426 ;
  assign n11958 = n11957 ^ n11925 ;
  assign n11960 = n11959 ^ n11958 ;
  assign n11977 = n11976 ^ n11960 ;
  assign n11922 = n6382 ^ n6377 ;
  assign n11923 = n6387 & ~n11922 ;
  assign n11924 = n11923 ^ n6382 ;
  assign n11978 = n11977 ^ n11924 ;
  assign n11987 = n11973 ^ n11970 ;
  assign n11983 = ~n3509 & n6163 ;
  assign n11984 = n20437 ^ n11983 ;
  assign n11985 = ~n368 & n11984 ;
  assign n11986 = n11985 ^ x17 ;
  assign n11988 = n11987 ^ n11986 ;
  assign n11989 = n11986 ^ n11924 ;
  assign n11990 = ~n11988 & ~n11989 ;
  assign n11991 = n11990 ^ n11987 ;
  assign n11992 = n11991 ^ n11988 ;
  assign n11993 = n11992 ^ n11977 ;
  assign n11994 = ~n11978 & ~n11993 ;
  assign n11995 = n11994 ^ n11977 ;
  assign n11996 = n11921 & n11995 ;
  assign n11997 = n11977 ^ n11919 ;
  assign n11998 = n11991 ^ n11977 ;
  assign n11999 = n11997 & n11998 ;
  assign n12000 = n11999 ^ n11977 ;
  assign n12001 = ~n11996 & ~n12000 ;
  assign n5429 = n3515 & n5221 ;
  assign n5428 = ~n3505 & n13433 ;
  assign n5430 = n5429 ^ n5428 ;
  assign n5431 = n5430 ^ x20 ;
  assign n5427 = ~n368 & n5426 ;
  assign n5432 = n5431 ^ n5427 ;
  assign n12003 = n12001 ^ n5432 ;
  assign n12002 = n5432 & n12001 ;
  assign n12004 = n12003 ^ n12002 ;
  assign n5413 = n5412 ^ n5252 ;
  assign n5414 = ~n5260 & n5413 ;
  assign n5415 = n5414 ^ n5412 ;
  assign n5249 = ~n40 & ~n540 ;
  assign n5185 = n5184 ^ n5140 ;
  assign n5186 = ~n5146 & n5185 ;
  assign n5187 = n5186 ^ n5140 ;
  assign n5135 = ~n4359 & ~n4435 ;
  assign n5132 = ~n856 & ~n4434 ;
  assign n5130 = ~n1248 & n20603 ;
  assign n5019 = n4876 ^ x17 ;
  assign n5020 = n4982 ^ n4876 ;
  assign n5021 = n5019 & ~n5020 ;
  assign n5022 = n5021 ^ x17 ;
  assign n4205 = n1680 ^ n143 ;
  assign n4204 = n1418 ^ n981 ;
  assign n4206 = n4205 ^ n4204 ;
  assign n4201 = n2481 ^ n489 ;
  assign n4202 = n4201 ^ n3166 ;
  assign n4199 = n3085 ^ n507 ;
  assign n4198 = n4197 ^ n455 ;
  assign n4200 = n4199 ^ n4198 ;
  assign n4203 = n4202 ^ n4200 ;
  assign n4207 = n4206 ^ n4203 ;
  assign n4208 = n4207 ^ n2579 ;
  assign n4209 = n4208 ^ n4196 ;
  assign n3574 = n836 ^ n776 ;
  assign n4183 = n4182 ^ n3574 ;
  assign n4184 = n4183 ^ n4181 ;
  assign n4180 = n523 ^ n217 ;
  assign n4185 = n4184 ^ n4180 ;
  assign n4186 = n4185 ^ n1921 ;
  assign n4177 = n821 ^ n506 ;
  assign n4175 = n2894 ^ n417 ;
  assign n4176 = n4175 ^ n710 ;
  assign n4178 = n4177 ^ n4176 ;
  assign n4174 = n4173 ^ n3378 ;
  assign n4179 = n4178 ^ n4174 ;
  assign n4187 = n4186 ^ n4179 ;
  assign n4210 = n4209 ^ n4187 ;
  assign n4222 = n3080 ^ n575 ;
  assign n4223 = n4222 ^ n119 ;
  assign n4220 = n1997 ^ n742 ;
  assign n4219 = n2068 ^ n771 ;
  assign n4221 = n4220 ^ n4219 ;
  assign n4224 = n4223 ^ n4221 ;
  assign n4216 = n2812 ^ n192 ;
  assign n4217 = n4216 ^ n764 ;
  assign n4215 = n761 ^ n377 ;
  assign n4218 = n4217 ^ n4215 ;
  assign n4225 = n4224 ^ n4218 ;
  assign n4213 = n2849 ^ n599 ;
  assign n3631 = n2187 ^ n526 ;
  assign n4212 = n4211 ^ n3631 ;
  assign n4214 = n4213 ^ n4212 ;
  assign n4226 = n4225 ^ n4214 ;
  assign n4227 = n4226 ^ n2240 ;
  assign n4228 = ~n4210 & ~n4227 ;
  assign n5089 = n5022 ^ n4228 ;
  assign n4692 = n4690 ^ n1670 ;
  assign n4691 = n4690 ^ n1819 ;
  assign n4693 = n4692 ^ n4691 ;
  assign n4696 = x30 & n4693 ;
  assign n4697 = n4696 ^ n4692 ;
  assign n4698 = ~n3518 & ~n4697 ;
  assign n4699 = n4698 ^ n4690 ;
  assign n4700 = x31 & n4699 ;
  assign n4688 = ~n1670 & ~n3805 ;
  assign n4687 = ~n1751 & n3807 ;
  assign n4689 = n4688 ^ n4687 ;
  assign n4701 = n4700 ^ n4689 ;
  assign n5126 = n5089 ^ n4701 ;
  assign n4708 = ~n1450 & n3837 ;
  assign n4706 = ~n990 & n4369 ;
  assign n4703 = n3983 & n4307 ;
  assign n4702 = ~n1345 & n3985 ;
  assign n4704 = n4703 ^ n4702 ;
  assign n4705 = n4704 ^ x29 ;
  assign n4707 = n4706 ^ n4705 ;
  assign n4709 = n4708 ^ n4707 ;
  assign n5127 = n5126 ^ n4709 ;
  assign n5007 = n4941 ^ n4876 ;
  assign n5008 = n5007 ^ n5006 ;
  assign n5009 = n4984 & n5008 ;
  assign n5010 = n5009 ^ n5006 ;
  assign n5128 = n5127 ^ n5010 ;
  assign n5129 = n5128 ^ x26 ;
  assign n5131 = n5130 ^ n5129 ;
  assign n5133 = n5132 ^ n5131 ;
  assign n5125 = ~n1119 & n4600 ;
  assign n5134 = n5133 ^ n5125 ;
  assign n5136 = n5135 ^ n5134 ;
  assign n5245 = n5187 ^ n5136 ;
  assign n5246 = n5245 ^ x23 ;
  assign n5242 = ~n3811 & n5239 ;
  assign n5243 = n5242 ^ n408 ;
  assign n5244 = n35 & ~n5243 ;
  assign n5247 = n5246 ^ n5244 ;
  assign n5235 = ~n698 & n4651 ;
  assign n5248 = n5247 ^ n5235 ;
  assign n5250 = n5249 ^ n5248 ;
  assign n12013 = n5415 ^ n5250 ;
  assign n12010 = n11976 ^ n11952 ;
  assign n12011 = ~n11960 & ~n12010 ;
  assign n12012 = n12011 ^ n11976 ;
  assign n12014 = n12013 ^ n12012 ;
  assign n12006 = n11943 ^ n11941 ;
  assign n12007 = n11951 & n12006 ;
  assign n12008 = n12007 ^ n11943 ;
  assign n5120 = n3840 & n4656 ;
  assign n5119 = ~n540 & n4651 ;
  assign n5121 = n5120 ^ n5119 ;
  assign n5122 = n5121 ^ x23 ;
  assign n5117 = ~n40 & ~n408 ;
  assign n5116 = ~n3505 & n4655 ;
  assign n5118 = n5117 ^ n5116 ;
  assign n5123 = n5122 ^ n5118 ;
  assign n5188 = n5187 ^ n5123 ;
  assign n5189 = n5188 ^ n5128 ;
  assign n5190 = n5189 ^ n5123 ;
  assign n5191 = n5136 & n5190 ;
  assign n5192 = n5191 ^ n5188 ;
  assign n5090 = n5022 ^ n4709 ;
  assign n5087 = n5010 ^ n4701 ;
  assign n5091 = n5090 ^ n5087 ;
  assign n5092 = n5089 & ~n5091 ;
  assign n4525 = n1953 ^ n772 ;
  assign n4526 = n4525 ^ n1076 ;
  assign n4523 = n978 ^ n974 ;
  assign n4524 = n4523 ^ n1367 ;
  assign n4527 = n4526 ^ n4524 ;
  assign n4520 = n4519 ^ n485 ;
  assign n4518 = n1020 ^ n145 ;
  assign n4521 = n4520 ^ n4518 ;
  assign n4516 = n706 ^ n209 ;
  assign n4515 = n1014 ^ n764 ;
  assign n4517 = n4516 ^ n4515 ;
  assign n4522 = n4521 ^ n4517 ;
  assign n4528 = n4527 ^ n4522 ;
  assign n4511 = n1844 ^ n270 ;
  assign n4512 = n4511 ^ n603 ;
  assign n4509 = n2137 ^ n918 ;
  assign n4510 = n4509 ^ n2413 ;
  assign n4513 = n4512 ^ n4510 ;
  assign n4506 = n2783 ^ n1544 ;
  assign n4505 = n2408 ^ n793 ;
  assign n4507 = n4506 ^ n4505 ;
  assign n4508 = n4507 ^ n4504 ;
  assign n4514 = n4513 ^ n4508 ;
  assign n4529 = n4528 ^ n4514 ;
  assign n4559 = n1630 ^ n613 ;
  assign n4560 = n4559 ^ n1962 ;
  assign n4557 = n1184 ^ n800 ;
  assign n4558 = n4557 ^ n645 ;
  assign n4561 = n4560 ^ n4558 ;
  assign n4273 = n1066 ^ n395 ;
  assign n4554 = n4273 ^ n3897 ;
  assign n4555 = n4554 ^ n4098 ;
  assign n4556 = n4555 ^ n2649 ;
  assign n4562 = n4561 ^ n4556 ;
  assign n4553 = n2776 ^ n1399 ;
  assign n4563 = n4562 ^ n4553 ;
  assign n4564 = n4563 ^ n4552 ;
  assign n4565 = ~n4529 & ~n4564 ;
  assign n4673 = n4565 ^ n4228 ;
  assign n4500 = ~n1670 & n22543 ;
  assign n4499 = ~n1751 & ~n3850 ;
  assign n4501 = n4500 ^ n4499 ;
  assign n4497 = n3807 & n4494 ;
  assign n4496 = n3518 & ~n4495 ;
  assign n4498 = n4497 ^ n4496 ;
  assign n4502 = n4501 ^ n4498 ;
  assign n4686 = n4673 ^ n4502 ;
  assign n5093 = n5092 ^ n4686 ;
  assign n5011 = n5010 ^ n4709 ;
  assign n5088 = ~n5011 & ~n5087 ;
  assign n5094 = n5093 ^ n5088 ;
  assign n5085 = ~n990 & n3985 ;
  assign n5080 = ~n3930 & ~n4435 ;
  assign n5078 = ~n698 & ~n4434 ;
  assign n5075 = ~n856 & n4600 ;
  assign n5074 = ~n1119 & n20603 ;
  assign n5076 = n5075 ^ n5074 ;
  assign n5077 = n5076 ^ x26 ;
  assign n5079 = n5078 ^ n5077 ;
  assign n5081 = n5080 ^ n5079 ;
  assign n5082 = n5081 ^ x29 ;
  assign n5071 = ~n4333 & n5065 ;
  assign n5072 = n5071 ^ n1248 ;
  assign n5073 = n3833 & ~n5072 ;
  assign n5083 = n5082 ^ n5073 ;
  assign n5064 = ~n1345 & n3837 ;
  assign n5084 = n5083 ^ n5064 ;
  assign n5086 = n5085 ^ n5084 ;
  assign n5115 = n5094 ^ n5086 ;
  assign n5421 = n5192 ^ n5115 ;
  assign n5416 = n5415 ^ n5245 ;
  assign n5417 = n5250 & n5416 ;
  assign n5418 = n5417 ^ n5245 ;
  assign n5419 = n5418 ^ x20 ;
  assign n5232 = ~n3509 & n5221 ;
  assign n5233 = n13433 ^ n5232 ;
  assign n5234 = ~n368 & n5233 ;
  assign n5420 = n5419 ^ n5234 ;
  assign n12005 = n5421 ^ n5420 ;
  assign n12009 = n12008 ^ n12005 ;
  assign n12015 = n12014 ^ n12009 ;
  assign n12016 = n12015 ^ n12009 ;
  assign n12017 = n12013 ^ n12008 ;
  assign n12020 = n12016 & n12017 ;
  assign n12021 = n12020 ^ n12009 ;
  assign n12022 = ~n12004 & ~n12021 ;
  assign n12024 = n12005 ^ n12002 ;
  assign n12025 = n12024 ^ n12005 ;
  assign n12026 = ~n12008 & ~n12025 ;
  assign n12027 = n12026 ^ n12005 ;
  assign n12035 = n12025 ^ n12008 ;
  assign n12036 = n12035 ^ n12005 ;
  assign n12029 = n12013 ^ n12005 ;
  assign n12028 = n12012 ^ n12005 ;
  assign n12030 = n12029 ^ n12028 ;
  assign n12031 = n12029 ^ n12024 ;
  assign n12032 = n12031 ^ n12009 ;
  assign n12033 = n12032 ^ n12005 ;
  assign n12034 = n12030 & ~n12033 ;
  assign n12037 = n12036 ^ n12034 ;
  assign n12038 = n12027 & n12037 ;
  assign n12039 = n12038 ^ n12005 ;
  assign n12042 = ~n12022 & ~n12039 ;
  assign n5422 = n5421 ^ n5418 ;
  assign n5423 = n5420 & ~n5422 ;
  assign n5424 = n5423 ^ n5418 ;
  assign n12043 = n12042 ^ n5424 ;
  assign n5095 = n5094 ^ n5081 ;
  assign n5096 = n5086 & n5095 ;
  assign n5097 = n5096 ^ n5081 ;
  assign n5062 = n3968 & ~n4435 ;
  assign n5059 = ~n540 & ~n4434 ;
  assign n5057 = ~n856 & n20603 ;
  assign n5023 = n4701 & ~n5022 ;
  assign n5013 = ~n4709 & ~n5010 ;
  assign n5024 = ~n4228 & n5013 ;
  assign n5025 = ~n5023 & n5024 ;
  assign n5027 = n5025 ^ n5022 ;
  assign n5012 = n5011 ^ n4701 ;
  assign n5014 = n5013 ^ n5012 ;
  assign n5015 = n5014 ^ n4701 ;
  assign n5016 = n4701 ^ n4228 ;
  assign n5017 = n5016 ^ n4701 ;
  assign n5018 = ~n5015 & n5017 ;
  assign n5026 = n5025 ^ n5018 ;
  assign n5028 = n5027 ^ n5026 ;
  assign n5029 = n5025 ^ n4701 ;
  assign n5030 = n5029 ^ n5027 ;
  assign n5031 = ~n5028 & ~n5030 ;
  assign n5032 = n5031 ^ n5027 ;
  assign n5033 = n4686 & n5032 ;
  assign n5034 = n5033 ^ n5025 ;
  assign n5035 = n5022 ^ n4701 ;
  assign n5036 = n5035 ^ n5023 ;
  assign n5037 = ~n4686 & ~n5036 ;
  assign n5038 = ~n5034 & ~n5037 ;
  assign n5039 = n5010 ^ n4228 ;
  assign n5042 = ~n5011 & n5039 ;
  assign n5043 = n5042 ^ n4228 ;
  assign n5044 = n5038 & ~n5043 ;
  assign n5045 = n5044 ^ n5034 ;
  assign n4480 = ~n1450 & ~n3850 ;
  assign n4479 = ~n1751 & n22543 ;
  assign n4481 = n4480 ^ n4479 ;
  assign n4477 = ~n3483 & n3807 ;
  assign n4476 = n3518 & n4475 ;
  assign n4478 = n4477 ^ n4476 ;
  assign n4482 = n4481 ^ n4478 ;
  assign n4247 = n2843 ^ n1823 ;
  assign n4246 = n2509 ^ n510 ;
  assign n4248 = n4247 ^ n4246 ;
  assign n4244 = n1837 ^ n1630 ;
  assign n4243 = n4242 ^ n1953 ;
  assign n4245 = n4244 ^ n4243 ;
  assign n4249 = n4248 ^ n4245 ;
  assign n4239 = n1786 ^ n570 ;
  assign n4240 = n4239 ^ n476 ;
  assign n4238 = n3207 ^ n847 ;
  assign n4241 = n4240 ^ n4238 ;
  assign n4250 = n4249 ^ n4241 ;
  assign n4234 = n1135 ^ n238 ;
  assign n4236 = n4235 ^ n4234 ;
  assign n4232 = n918 ^ n243 ;
  assign n4230 = n1284 ^ n744 ;
  assign n4231 = n4230 ^ n430 ;
  assign n4233 = n4232 ^ n4231 ;
  assign n4237 = n4236 ^ n4233 ;
  assign n4251 = n4250 ^ n4237 ;
  assign n4272 = n4271 ^ n4251 ;
  assign n4296 = n4295 ^ n142 ;
  assign n4297 = n4296 ^ n603 ;
  assign n4294 = n1106 ^ n262 ;
  assign n4298 = n4297 ^ n4294 ;
  assign n4290 = n446 ^ n340 ;
  assign n4291 = n4290 ^ n710 ;
  assign n4292 = n4291 ^ n1687 ;
  assign n4288 = n969 ^ n411 ;
  assign n4289 = n4288 ^ n1236 ;
  assign n4293 = n4292 ^ n4289 ;
  assign n4299 = n4298 ^ n4293 ;
  assign n4284 = n2966 ^ n991 ;
  assign n4283 = n950 ^ n192 ;
  assign n4285 = n4284 ^ n4283 ;
  assign n4280 = n436 ^ n265 ;
  assign n4281 = n4280 ^ n1268 ;
  assign n4282 = n4281 ^ n2479 ;
  assign n4286 = n4285 ^ n4282 ;
  assign n4287 = n4286 ^ n705 ;
  assign n4300 = n4299 ^ n4287 ;
  assign n3789 = n1711 ^ n761 ;
  assign n4277 = n3789 ^ n1273 ;
  assign n4276 = n2918 ^ n318 ;
  assign n4278 = n4277 ^ n4276 ;
  assign n4274 = n4273 ^ n1065 ;
  assign n4275 = n4274 ^ n2616 ;
  assign n4279 = n4278 ^ n4275 ;
  assign n4301 = n4300 ^ n4279 ;
  assign n4302 = ~n4272 & ~n4301 ;
  assign n4474 = n4302 ^ x20 ;
  assign n4683 = n4482 ^ n4474 ;
  assign n4678 = ~n1119 & n4369 ;
  assign n4677 = ~n990 & n3837 ;
  assign n4679 = n4678 ^ n4677 ;
  assign n4680 = n4679 ^ x29 ;
  assign n4676 = n3983 & ~n4336 ;
  assign n4681 = n4680 ^ n4676 ;
  assign n4675 = ~n1248 & n3985 ;
  assign n4682 = n4681 ^ n4675 ;
  assign n4684 = n4683 ^ n4682 ;
  assign n4566 = n4565 ^ n4502 ;
  assign n4674 = n4566 & ~n4673 ;
  assign n4685 = n4684 ^ n4674 ;
  assign n5055 = n5045 ^ n4685 ;
  assign n5056 = n5055 ^ x26 ;
  assign n5058 = n5057 ^ n5056 ;
  assign n5060 = n5059 ^ n5058 ;
  assign n5054 = ~n698 & n4600 ;
  assign n5061 = n5060 ^ n5054 ;
  assign n5063 = n5062 ^ n5061 ;
  assign n5207 = n5097 ^ n5063 ;
  assign n5205 = ~n40 & ~n3505 ;
  assign n5203 = ~n408 & n4651 ;
  assign n5199 = ~n3513 & n5239 ;
  assign n5200 = n5199 ^ n368 ;
  assign n5201 = n35 & ~n5200 ;
  assign n5202 = n5201 ^ x23 ;
  assign n5204 = n5203 ^ n5202 ;
  assign n5206 = n5205 ^ n5204 ;
  assign n5208 = n5207 ^ n5206 ;
  assign n5124 = n5123 ^ n5115 ;
  assign n5193 = n5124 & ~n5192 ;
  assign n5194 = n5193 ^ n5123 ;
  assign n12225 = n5208 ^ n5194 ;
  assign n12226 = n12225 ^ n5424 ;
  assign n12227 = ~n12043 & n12226 ;
  assign n5107 = n3515 & n4656 ;
  assign n5105 = ~n3505 & n4651 ;
  assign n5103 = ~n40 & ~n368 ;
  assign n5046 = n5045 ^ n4682 ;
  assign n5047 = ~n4685 & ~n5046 ;
  assign n5048 = n5047 ^ n4682 ;
  assign n4670 = n3812 & ~n4435 ;
  assign n4668 = ~n698 & n20603 ;
  assign n4665 = ~n540 & n4600 ;
  assign n4664 = ~n408 & ~n4434 ;
  assign n4666 = n4665 ^ n4664 ;
  assign n4667 = n4666 ^ x26 ;
  assign n4669 = n4668 ^ n4667 ;
  assign n4671 = n4670 ^ n4669 ;
  assign n4483 = n4482 ^ n4228 ;
  assign n4484 = n4483 ^ n4474 ;
  assign n4569 = n4502 ^ n4482 ;
  assign n4570 = n4569 ^ n4474 ;
  assign n4571 = n4566 & n4570 ;
  assign n4572 = n4571 ^ n4474 ;
  assign n4573 = ~n4484 & n4572 ;
  assign n4574 = n4573 ^ n4482 ;
  assign n4468 = ~n1248 & n3837 ;
  assign n4467 = ~n856 & n4369 ;
  assign n4469 = n4468 ^ n4467 ;
  assign n4470 = n4469 ^ x29 ;
  assign n4466 = n3983 & ~n4359 ;
  assign n4471 = n4470 ^ n4466 ;
  assign n4465 = ~n1119 & n3985 ;
  assign n4472 = n4471 ^ n4465 ;
  assign n4319 = ~n61 & n1345 ;
  assign n4320 = n4319 ^ n990 ;
  assign n4318 = ~n61 & n990 ;
  assign n4321 = n4320 ^ n4318 ;
  assign n4322 = ~n3800 & ~n4321 ;
  assign n4309 = n4307 ^ n1345 ;
  assign n4308 = n4307 ^ n1450 ;
  assign n4310 = n4309 ^ n4308 ;
  assign n4313 = x30 & n4310 ;
  assign n4314 = n4313 ^ n4309 ;
  assign n4315 = ~n3518 & ~n4314 ;
  assign n4316 = n4315 ^ n4307 ;
  assign n4317 = x31 & n4316 ;
  assign n4323 = n4322 ^ n4317 ;
  assign n4131 = n2904 ^ n510 ;
  assign n4164 = n1630 ^ n772 ;
  assign n4165 = n4164 ^ n243 ;
  assign n4166 = n4165 ^ n589 ;
  assign n4163 = n1130 ^ n730 ;
  assign n4167 = n4166 ^ n4163 ;
  assign n4160 = n4159 ^ n845 ;
  assign n4161 = n4160 ^ n1940 ;
  assign n4156 = n831 ^ n542 ;
  assign n4157 = n4156 ^ n2500 ;
  assign n4155 = n4154 ^ n741 ;
  assign n4158 = n4157 ^ n4155 ;
  assign n4162 = n4161 ^ n4158 ;
  assign n4168 = n4167 ^ n4162 ;
  assign n4151 = n981 ^ n444 ;
  assign n4152 = n4151 ^ n1997 ;
  assign n4150 = n3038 ^ n1833 ;
  assign n4153 = n4152 ^ n4150 ;
  assign n4169 = n4168 ^ n4153 ;
  assign n4144 = n2408 ^ n199 ;
  assign n4145 = n4144 ^ n706 ;
  assign n4143 = n2519 ^ n603 ;
  assign n4146 = n4145 ^ n4143 ;
  assign n4141 = n898 ^ n578 ;
  assign n4142 = n4141 ^ n1321 ;
  assign n4147 = n4146 ^ n4142 ;
  assign n4138 = n761 ^ n137 ;
  assign n4139 = n4138 ^ n687 ;
  assign n4137 = n3713 ^ n530 ;
  assign n4140 = n4139 ^ n4137 ;
  assign n4148 = n4147 ^ n4140 ;
  assign n4133 = n2139 ^ n247 ;
  assign n4134 = n4133 ^ n414 ;
  assign n4132 = n628 ^ n494 ;
  assign n4135 = n4134 ^ n4132 ;
  assign n4136 = n4135 ^ n3364 ;
  assign n4149 = n4148 ^ n4136 ;
  assign n4170 = n4169 ^ n4149 ;
  assign n4171 = n4170 ^ n1767 ;
  assign n4172 = ~n4131 & ~n4171 ;
  assign n4461 = n4323 ^ n4172 ;
  assign n4229 = n4228 ^ x20 ;
  assign n4303 = n4302 ^ n4228 ;
  assign n4304 = n4229 & ~n4303 ;
  assign n4305 = n4304 ^ x20 ;
  assign n4464 = n4461 ^ n4305 ;
  assign n4473 = n4472 ^ n4464 ;
  assign n4663 = n4574 ^ n4473 ;
  assign n4672 = n4671 ^ n4663 ;
  assign n5053 = n5048 ^ n4672 ;
  assign n5102 = n5053 ^ x23 ;
  assign n5104 = n5103 ^ n5102 ;
  assign n5106 = n5105 ^ n5104 ;
  assign n5108 = n5107 ^ n5106 ;
  assign n5098 = n5097 ^ n5055 ;
  assign n5099 = n5063 & n5098 ;
  assign n5100 = n5099 ^ n5055 ;
  assign n12046 = n5108 ^ n5100 ;
  assign n12223 = n12046 ^ n5208 ;
  assign n12050 = n5206 ^ n5194 ;
  assign n12051 = ~n5208 & n12050 ;
  assign n12224 = n12223 ^ n12051 ;
  assign n12228 = n12227 ^ n12224 ;
  assign n12229 = n12226 ^ n12042 ;
  assign n12232 = n12017 ^ n12012 ;
  assign n12233 = ~n12003 & ~n12232 ;
  assign n12230 = n12012 ^ n12008 ;
  assign n12231 = ~n12017 & n12230 ;
  assign n12234 = n12233 ^ n12231 ;
  assign n12235 = n12234 ^ n12024 ;
  assign n12236 = n12008 ^ n5432 ;
  assign n12237 = n12236 ^ n12013 ;
  assign n12238 = n12237 ^ n12012 ;
  assign n12239 = n12238 ^ n12001 ;
  assign n12245 = n11988 & ~n11989 ;
  assign n12243 = n11988 ^ n11924 ;
  assign n12244 = ~n5967 & n12243 ;
  assign n12246 = n12245 ^ n12244 ;
  assign n12247 = n12246 ^ n11977 ;
  assign n12240 = n11988 ^ n5967 ;
  assign n12241 = n12240 ^ n11924 ;
  assign n12242 = n11918 & n12241 ;
  assign n12248 = n12247 ^ n12242 ;
  assign n12249 = n12241 ^ n11918 ;
  assign n12337 = n6526 ^ n6376 ;
  assign n12338 = n12337 ^ n6388 ;
  assign n12250 = n6525 ^ n6375 ;
  assign n12335 = n11900 ^ n6375 ;
  assign n12336 = ~n12250 & n12335 ;
  assign n12339 = n12338 ^ n12336 ;
  assign n12251 = n12250 ^ n11900 ;
  assign n12252 = n11897 ^ n7022 ;
  assign n12253 = n12252 ^ n7021 ;
  assign n12254 = n11877 ^ n7289 ;
  assign n12327 = n11878 ^ n7284 ;
  assign n12328 = n12327 ^ n7287 ;
  assign n12329 = n12254 & n12328 ;
  assign n12330 = n12329 ^ n7293 ;
  assign n12325 = n11858 ^ n7284 ;
  assign n12326 = n7288 & ~n12325 ;
  assign n12331 = n12330 ^ n12326 ;
  assign n12255 = n12254 ^ n7287 ;
  assign n12256 = n12255 ^ n7284 ;
  assign n12257 = n12256 ^ n11858 ;
  assign n12258 = n11855 ^ n7560 ;
  assign n12259 = n11833 ^ n11819 ;
  assign n12262 = n11838 & n12259 ;
  assign n12260 = n12259 ^ n11836 ;
  assign n12261 = n11829 & n12260 ;
  assign n12263 = n12262 ^ n12261 ;
  assign n12264 = n12263 ^ n11842 ;
  assign n12265 = n11833 ^ n11829 ;
  assign n12266 = n12265 ^ n11836 ;
  assign n12267 = n12266 ^ n11819 ;
  assign n12268 = n11816 ^ n8481 ;
  assign n12271 = n11794 ^ n11780 ;
  assign n12269 = n11791 ^ n11778 ;
  assign n12272 = n12269 ^ n11775 ;
  assign n12273 = n12272 ^ n11794 ;
  assign n12274 = ~n12271 & n12273 ;
  assign n12275 = n12274 ^ n11796 ;
  assign n12270 = ~n11779 & ~n12269 ;
  assign n12276 = n12275 ^ n12270 ;
  assign n12277 = n11809 ^ n11780 ;
  assign n12278 = n12277 ^ n11778 ;
  assign n12279 = n12278 ^ n11775 ;
  assign n12282 = ~n10395 & n11762 ;
  assign n12280 = n10392 ^ n10381 ;
  assign n12281 = n12280 ^ n10389 ;
  assign n12283 = n12282 ^ n12281 ;
  assign n12284 = n11762 ^ n10395 ;
  assign n12285 = n11760 ^ n11754 ;
  assign n12308 = n11728 ^ n11655 ;
  assign n12309 = n11739 ^ n11720 ;
  assign n12310 = n12309 ^ n11654 ;
  assign n12311 = ~n12308 & n12310 ;
  assign n12312 = n12311 ^ n11716 ;
  assign n12305 = n11720 ^ n11654 ;
  assign n12306 = n11720 ^ n11696 ;
  assign n12307 = n12305 & n12306 ;
  assign n12313 = n12312 ^ n12307 ;
  assign n12286 = n11728 ^ n11696 ;
  assign n12287 = n12286 ^ n11655 ;
  assign n12288 = n12287 ^ n11720 ;
  assign n12289 = n12288 ^ n11654 ;
  assign n12290 = n11652 ^ n10972 ;
  assign n12293 = n11649 ^ n11631 ;
  assign n12291 = n11625 ^ n11010 ;
  assign n12292 = n11628 ^ n10992 ;
  assign n12298 = ~n12291 & ~n12292 ;
  assign n12299 = n12298 ^ n12291 ;
  assign n12300 = n12299 ^ n12292 ;
  assign n12301 = ~n12293 & n12300 ;
  assign n12347 = ~n12290 & ~n12301 ;
  assign n12348 = ~n12289 & ~n12347 ;
  assign n12349 = n12313 & ~n12348 ;
  assign n12350 = n12285 & ~n12349 ;
  assign n12351 = ~n12284 & ~n12350 ;
  assign n12352 = n12283 & ~n12351 ;
  assign n12353 = n12279 & ~n12352 ;
  assign n12354 = n12276 & ~n12353 ;
  assign n12355 = n12268 & ~n12354 ;
  assign n12356 = n12267 & ~n12355 ;
  assign n12357 = n12264 & ~n12356 ;
  assign n12358 = n12258 & ~n12357 ;
  assign n12359 = n12257 & ~n12358 ;
  assign n12360 = ~n12331 & ~n12359 ;
  assign n12361 = n12253 & ~n12360 ;
  assign n12362 = n12251 & ~n12361 ;
  assign n12363 = n12339 & ~n12362 ;
  assign n12364 = n12249 & ~n12363 ;
  assign n12365 = n12248 & ~n12364 ;
  assign n12366 = n12239 & ~n12365 ;
  assign n12367 = n12235 & ~n12366 ;
  assign n12368 = ~n12229 & ~n12367 ;
  assign n12369 = ~n12228 & ~n12368 ;
  assign n12294 = n12293 ^ n12292 ;
  assign n12295 = n12292 & n12294 ;
  assign n12296 = ~n12291 & n12295 ;
  assign n12297 = n12296 ^ n12294 ;
  assign n12302 = n12301 ^ n12297 ;
  assign n12303 = n12290 & n12302 ;
  assign n12304 = n12289 & ~n12303 ;
  assign n12314 = ~n12304 & ~n12313 ;
  assign n12315 = ~n12285 & ~n12314 ;
  assign n12316 = n12284 & ~n12315 ;
  assign n12317 = ~n12283 & ~n12316 ;
  assign n12318 = ~n12279 & ~n12317 ;
  assign n12319 = ~n12276 & ~n12318 ;
  assign n12320 = ~n12268 & ~n12319 ;
  assign n12321 = ~n12267 & ~n12320 ;
  assign n12322 = ~n12264 & ~n12321 ;
  assign n12323 = ~n12258 & ~n12322 ;
  assign n12324 = ~n12257 & ~n12323 ;
  assign n12332 = ~n12324 & n12331 ;
  assign n12333 = ~n12253 & ~n12332 ;
  assign n12334 = ~n12251 & ~n12333 ;
  assign n12340 = ~n12334 & ~n12339 ;
  assign n12341 = ~n12249 & ~n12340 ;
  assign n12342 = ~n12248 & ~n12341 ;
  assign n12343 = ~n12239 & ~n12342 ;
  assign n12344 = ~n12235 & ~n12343 ;
  assign n12345 = n12229 & ~n12344 ;
  assign n12346 = n12228 & ~n12345 ;
  assign n12370 = n12369 ^ n12346 ;
  assign n4372 = n3812 & n3983 ;
  assign n4371 = ~n540 & n3985 ;
  assign n4373 = n4372 ^ n4371 ;
  assign n4374 = n4373 ^ x29 ;
  assign n4370 = ~n408 & n4369 ;
  assign n4375 = n4374 ^ n4370 ;
  assign n4367 = ~n698 & n3837 ;
  assign n4376 = n4375 ^ n4367 ;
  assign n4362 = ~n3492 & n3807 ;
  assign n4361 = x31 & ~n1119 ;
  assign n4363 = n4362 ^ n4361 ;
  assign n4360 = n3518 & n4359 ;
  assign n4364 = n4363 ^ n4360 ;
  assign n4356 = ~n61 & n1248 ;
  assign n4357 = n3805 & ~n4356 ;
  assign n4355 = ~n52 & n1119 ;
  assign n4358 = n4357 ^ n4355 ;
  assign n4365 = n4364 ^ n4358 ;
  assign n3687 = n1252 ^ n794 ;
  assign n3688 = n3687 ^ n3099 ;
  assign n3689 = n3688 ^ n3686 ;
  assign n3699 = n3698 ^ n3689 ;
  assign n3681 = n2576 ^ n379 ;
  assign n3680 = n3166 ^ n714 ;
  assign n3682 = n3681 ^ n3680 ;
  assign n3677 = n903 ^ n353 ;
  assign n3678 = n3677 ^ n1704 ;
  assign n3676 = n1273 ^ n862 ;
  assign n3679 = n3678 ^ n3676 ;
  assign n3683 = n3682 ^ n3679 ;
  assign n3673 = n770 ^ n452 ;
  assign n3674 = n3673 ^ n465 ;
  assign n3670 = n380 ^ n149 ;
  assign n3671 = n3670 ^ n108 ;
  assign n3672 = n3671 ^ n3407 ;
  assign n3675 = n3674 ^ n3672 ;
  assign n3684 = n3683 ^ n3675 ;
  assign n3700 = n3699 ^ n3684 ;
  assign n3728 = n3727 ^ n3700 ;
  assign n3729 = ~n2225 & ~n3728 ;
  assign n4366 = n4365 ^ n3729 ;
  assign n4609 = n4376 ^ n4366 ;
  assign n4088 = n4087 ^ n377 ;
  assign n4086 = n1360 ^ n820 ;
  assign n4089 = n4088 ^ n4086 ;
  assign n4085 = n1960 ^ n118 ;
  assign n4090 = n4089 ^ n4085 ;
  assign n4091 = n4090 ^ n1990 ;
  assign n4081 = n1330 ^ n602 ;
  assign n4082 = n4081 ^ n623 ;
  assign n4079 = n3716 ^ n1556 ;
  assign n4080 = n4079 ^ n2631 ;
  assign n4083 = n4082 ^ n4080 ;
  assign n3585 = n2187 ^ n215 ;
  assign n4077 = n3585 ^ n3048 ;
  assign n4075 = n2153 ^ n237 ;
  assign n4073 = n2988 ^ n149 ;
  assign n4074 = n4073 ^ n429 ;
  assign n4076 = n4075 ^ n4074 ;
  assign n4078 = n4077 ^ n4076 ;
  assign n4084 = n4083 ^ n4078 ;
  assign n4092 = n4091 ^ n4084 ;
  assign n4122 = n1408 ^ n706 ;
  assign n4121 = n1189 ^ n719 ;
  assign n4123 = n4122 ^ n4121 ;
  assign n4119 = n1631 ^ n546 ;
  assign n4118 = n659 ^ n596 ;
  assign n4120 = n4119 ^ n4118 ;
  assign n4124 = n4123 ^ n4120 ;
  assign n4125 = n4124 ^ n3180 ;
  assign n4114 = n4113 ^ n1314 ;
  assign n4112 = n4111 ^ n875 ;
  assign n4115 = n4114 ^ n4112 ;
  assign n4109 = n571 ^ n446 ;
  assign n4110 = n4109 ^ n766 ;
  assign n4116 = n4115 ^ n4110 ;
  assign n4117 = n4116 ^ n4108 ;
  assign n4126 = n4125 ^ n4117 ;
  assign n4127 = n4126 ^ n4102 ;
  assign n4128 = ~n4092 & ~n4127 ;
  assign n4129 = n4128 ^ x23 ;
  assign n4026 = n4025 ^ n649 ;
  assign n4027 = n4026 ^ n2949 ;
  assign n4028 = n4027 ^ n3031 ;
  assign n4022 = n2277 ^ n542 ;
  assign n4021 = n641 ^ n417 ;
  assign n4023 = n4022 ^ n4021 ;
  assign n4019 = n4018 ^ n385 ;
  assign n4017 = n900 ^ n377 ;
  assign n4020 = n4019 ^ n4017 ;
  assign n4024 = n4023 ^ n4020 ;
  assign n4029 = n4028 ^ n4024 ;
  assign n4011 = n818 ^ n706 ;
  assign n4013 = n4012 ^ n4011 ;
  assign n4010 = n484 ^ n471 ;
  assign n4014 = n4013 ^ n4010 ;
  assign n4008 = n2271 ^ n1558 ;
  assign n4007 = n1306 ^ n1277 ;
  assign n4009 = n4008 ^ n4007 ;
  assign n4015 = n4014 ^ n4009 ;
  assign n4016 = n4015 ^ n1914 ;
  assign n4030 = n4029 ^ n4016 ;
  assign n4002 = n2828 ^ n506 ;
  assign n4003 = n4002 ^ n634 ;
  assign n4001 = n3140 ^ n550 ;
  assign n4004 = n4003 ^ n4001 ;
  assign n3997 = n546 ^ n252 ;
  assign n3998 = n3997 ^ n214 ;
  assign n3999 = n3998 ^ n690 ;
  assign n3996 = n951 ^ n124 ;
  assign n4000 = n3999 ^ n3996 ;
  assign n4005 = n4004 ^ n4000 ;
  assign n4006 = n4005 ^ n2281 ;
  assign n4031 = n4030 ^ n4006 ;
  assign n4065 = n1257 ^ n877 ;
  assign n4066 = n4065 ^ n2054 ;
  assign n3664 = n3663 ^ n429 ;
  assign n3665 = n3664 ^ n842 ;
  assign n4067 = n4066 ^ n3665 ;
  assign n4063 = n1549 ^ n1160 ;
  assign n4064 = n4063 ^ n892 ;
  assign n4068 = n4067 ^ n4064 ;
  assign n4059 = n4058 ^ n2781 ;
  assign n4060 = n4059 ^ n248 ;
  assign n4056 = n1498 ^ n215 ;
  assign n4057 = n4056 ^ n272 ;
  assign n4061 = n4060 ^ n4057 ;
  assign n4053 = n1962 ^ n179 ;
  assign n4054 = n4053 ^ n956 ;
  assign n4052 = n1400 ^ n776 ;
  assign n4055 = n4054 ^ n4052 ;
  assign n4062 = n4061 ^ n4055 ;
  assign n4069 = n4068 ^ n4062 ;
  assign n4070 = n4069 ^ n4051 ;
  assign n4071 = n4070 ^ n2232 ;
  assign n4072 = ~n4031 & ~n4071 ;
  assign n4349 = n4128 ^ n4072 ;
  assign n4350 = n4129 & ~n4349 ;
  assign n4351 = n4350 ^ x23 ;
  assign n4306 = n4305 ^ n4172 ;
  assign n4324 = n4323 ^ n4128 ;
  assign n4325 = n4305 ^ n4128 ;
  assign n4326 = n4324 & ~n4325 ;
  assign n4327 = ~n4306 & n4326 ;
  assign n4328 = n4327 ^ n4128 ;
  assign n4130 = n4129 ^ n4072 ;
  assign n4329 = n4328 ^ n4130 ;
  assign n4343 = n52 ^ x31 ;
  assign n4344 = n1248 & ~n4343 ;
  assign n4340 = n4328 ^ x31 ;
  assign n4338 = n4335 ^ n1248 ;
  assign n4339 = n3807 & ~n4338 ;
  assign n4341 = n4340 ^ n4339 ;
  assign n4337 = n3518 & n4336 ;
  assign n4342 = n4341 ^ n4337 ;
  assign n4345 = n4344 ^ n4342 ;
  assign n4330 = n3805 & ~n4318 ;
  assign n4346 = n4345 ^ n4330 ;
  assign n4347 = ~n4329 & ~n4346 ;
  assign n4348 = n4347 ^ n4328 ;
  assign n4352 = n4351 ^ n4348 ;
  assign n4610 = n4609 ^ n4352 ;
  assign n4602 = ~n3505 & n20603 ;
  assign n4601 = ~n368 & n4600 ;
  assign n4603 = n4602 ^ n4601 ;
  assign n4604 = n4603 ^ x26 ;
  assign n4599 = n3515 & ~n4435 ;
  assign n4605 = n4604 ^ n4599 ;
  assign n12377 = n4610 ^ n4605 ;
  assign n4455 = ~n856 & n3837 ;
  assign n4454 = ~n540 & n4369 ;
  assign n4456 = n4455 ^ n4454 ;
  assign n4457 = n4456 ^ x29 ;
  assign n4453 = n3968 & n3983 ;
  assign n4458 = n4457 ^ n4453 ;
  assign n4452 = ~n698 & n3985 ;
  assign n4459 = n4458 ^ n4452 ;
  assign n4451 = n4346 ^ n4130 ;
  assign n4460 = n4459 ^ n4451 ;
  assign n4575 = n4574 ^ n4472 ;
  assign n4576 = ~n4473 & n4575 ;
  assign n4577 = n4576 ^ n4472 ;
  assign n4462 = ~n4306 & n4461 ;
  assign n4463 = n4462 ^ n4128 ;
  assign n4578 = n4577 ^ n4463 ;
  assign n4589 = n4318 ^ n1248 ;
  assign n4590 = n4589 ^ n4356 ;
  assign n4591 = ~n3800 & ~n4590 ;
  assign n4579 = x31 & ~n4319 ;
  assign n4588 = n4579 ^ n4463 ;
  assign n4592 = n4591 ^ n4588 ;
  assign n4581 = n4580 ^ n3518 ;
  assign n4582 = n4581 ^ n4580 ;
  assign n4583 = ~x30 & n990 ;
  assign n4584 = n4583 ^ n4580 ;
  assign n4585 = ~n4582 & ~n4584 ;
  assign n4586 = n4585 ^ n4580 ;
  assign n4587 = n4579 & ~n4586 ;
  assign n4593 = n4592 ^ n4587 ;
  assign n4594 = ~n4578 & n4593 ;
  assign n4595 = n4594 ^ n4577 ;
  assign n4596 = n4595 ^ n4459 ;
  assign n4597 = n4460 & n4596 ;
  assign n4598 = n4597 ^ n4459 ;
  assign n12378 = n12377 ^ n4598 ;
  assign n4619 = n4398 & ~n4435 ;
  assign n4616 = ~n3505 & n4600 ;
  assign n4614 = ~n408 & n20603 ;
  assign n4612 = n4595 ^ n4460 ;
  assign n4613 = n4612 ^ x26 ;
  assign n4615 = n4614 ^ n4613 ;
  assign n4617 = n4616 ^ n4615 ;
  assign n4611 = ~n368 & ~n4434 ;
  assign n4618 = n4617 ^ n4611 ;
  assign n4620 = n4619 ^ n4618 ;
  assign n4625 = ~n698 & n4369 ;
  assign n4624 = ~n1119 & n3837 ;
  assign n4626 = n4625 ^ n4624 ;
  assign n4627 = n4626 ^ x29 ;
  assign n4623 = ~n3930 & n3983 ;
  assign n4628 = n4627 ^ n4623 ;
  assign n4622 = ~n856 & n3985 ;
  assign n4629 = n4628 ^ n4622 ;
  assign n4621 = n4593 ^ n4577 ;
  assign n4630 = n4629 ^ n4621 ;
  assign n4637 = ~n540 & n20603 ;
  assign n4635 = ~n408 & n4600 ;
  assign n4633 = ~n3505 & ~n4434 ;
  assign n4632 = n4629 ^ x26 ;
  assign n4634 = n4633 ^ n4632 ;
  assign n4636 = n4635 ^ n4634 ;
  assign n4638 = n4637 ^ n4636 ;
  assign n4631 = n3840 & ~n4435 ;
  assign n4639 = n4638 ^ n4631 ;
  assign n4640 = ~n4630 & n4639 ;
  assign n4641 = n4640 ^ n4629 ;
  assign n4642 = n4641 ^ n4612 ;
  assign n4643 = n4620 & n4642 ;
  assign n4644 = n4643 ^ n4612 ;
  assign n12379 = n12378 ^ n4644 ;
  assign n4650 = n4641 ^ n4620 ;
  assign n5049 = n5048 ^ n4671 ;
  assign n5050 = ~n4672 & n5049 ;
  assign n5051 = n5050 ^ n4671 ;
  assign n4659 = ~n3509 & n4656 ;
  assign n4660 = n4659 ^ n4651 ;
  assign n4661 = ~n368 & n4660 ;
  assign n4662 = n4661 ^ x23 ;
  assign n5052 = n5051 ^ n4662 ;
  assign n5101 = n5100 ^ n5053 ;
  assign n5109 = ~n5101 & n5108 ;
  assign n5110 = n5109 ^ n5100 ;
  assign n5111 = n5110 ^ n5051 ;
  assign n5112 = ~n5052 & n5111 ;
  assign n5113 = n5112 ^ n5110 ;
  assign n5114 = ~n4650 & ~n5113 ;
  assign n12061 = n4639 ^ n4621 ;
  assign n12062 = n5113 ^ n4650 ;
  assign n12063 = n12062 ^ n5114 ;
  assign n12064 = n12061 & n12063 ;
  assign n5209 = n5207 ^ n5194 ;
  assign n5210 = ~n5208 & ~n5209 ;
  assign n5211 = ~n5194 & n5210 ;
  assign n12044 = n5424 & n12042 ;
  assign n12045 = n12044 ^ n12043 ;
  assign n12047 = n12046 ^ n5210 ;
  assign n12048 = n12046 ^ n12044 ;
  assign n12049 = n12046 ^ n5194 ;
  assign n12052 = n12051 ^ n12049 ;
  assign n12053 = ~n12048 & n12052 ;
  assign n12054 = n12053 ^ n12044 ;
  assign n12055 = ~n12047 & ~n12054 ;
  assign n12056 = n12045 & n12055 ;
  assign n12057 = n12056 ^ n12054 ;
  assign n12058 = n12057 ^ n12054 ;
  assign n12059 = n5211 & n12058 ;
  assign n12060 = n12059 ^ n12057 ;
  assign n12065 = n12064 ^ n12060 ;
  assign n12066 = ~n4662 & ~n5051 ;
  assign n12067 = ~n5110 & n12066 ;
  assign n12069 = n12067 ^ n5052 ;
  assign n12070 = n12069 ^ n5112 ;
  assign n12071 = n12070 ^ n12067 ;
  assign n12068 = n12067 ^ n12060 ;
  assign n12074 = n12068 ^ n4650 ;
  assign n12075 = n12074 ^ n12068 ;
  assign n12076 = n12071 & ~n12075 ;
  assign n12077 = n12076 ^ n12068 ;
  assign n12078 = ~n12065 & n12077 ;
  assign n12079 = n12078 ^ n12064 ;
  assign n12080 = ~n5114 & ~n12079 ;
  assign n12380 = n12379 ^ n12080 ;
  assign n12375 = n12071 ^ n4650 ;
  assign n12371 = n12061 ^ n5110 ;
  assign n12372 = n12371 ^ n5052 ;
  assign n12373 = n12061 ^ n12060 ;
  assign n12374 = ~n12372 & n12373 ;
  assign n12376 = n12375 ^ n12374 ;
  assign n12381 = n12380 ^ n12376 ;
  assign n12382 = n12372 ^ n12060 ;
  assign n12383 = n12382 ^ n12380 ;
  assign n12384 = n12381 & n12383 ;
  assign n12385 = n12370 & n12384 ;
  assign n12386 = n12384 ^ n12376 ;
  assign n12387 = n12386 ^ n12228 ;
  assign n12388 = n12385 & ~n12387 ;
  assign n12389 = n12388 ^ n12386 ;
  assign n12390 = n12389 ^ n12380 ;
  assign n13223 = n3985 & n12380 ;
  assign n13222 = n3837 & n12376 ;
  assign n13224 = n13223 ^ n13222 ;
  assign n13225 = n13224 ^ x29 ;
  assign n13226 = n13225 ^ n4368 ;
  assign n13232 = ~x28 & n13226 ;
  assign n13233 = n13232 ^ n4368 ;
  assign n13234 = n12390 & n13233 ;
  assign n13235 = n13234 ^ n4368 ;
  assign n12217 = n12080 ^ n4610 ;
  assign n12218 = n12080 ^ n4644 ;
  assign n4649 = n4605 ^ n4598 ;
  assign n12219 = n12218 ^ n4649 ;
  assign n12220 = ~n12217 & n12219 ;
  assign n4429 = ~n540 & n3837 ;
  assign n4426 = n3985 ^ x29 ;
  assign n4424 = n4368 ^ n3832 ;
  assign n4425 = n408 & n4424 ;
  assign n4427 = n4426 ^ n4425 ;
  assign n4423 = n3840 & n3983 ;
  assign n4428 = n4427 ^ n4423 ;
  assign n4430 = n4429 ^ n4428 ;
  assign n4443 = n4430 ^ x26 ;
  assign n4440 = ~n3509 & ~n4435 ;
  assign n4441 = ~n20603 ^ n4440 ;
  assign n4442 = ~n368 & ~n4441 ;
  assign n4444 = n4443 ^ n4442 ;
  assign n4417 = n4351 ^ n3729 ;
  assign n4377 = n4376 ^ n4365 ;
  assign n4418 = n4377 ^ n4351 ;
  assign n4419 = n4418 ^ n4348 ;
  assign n4420 = n4417 & n4419 ;
  assign n3929 = ~n61 & ~n856 ;
  assign n3941 = n3929 ^ n3495 ;
  assign n3932 = n3930 ^ n856 ;
  assign n3931 = n3930 ^ n1119 ;
  assign n3933 = n3932 ^ n3931 ;
  assign n3936 = x30 & n3933 ;
  assign n3937 = n3936 ^ n3932 ;
  assign n3938 = ~n3518 & n3937 ;
  assign n3939 = n3938 ^ n3930 ;
  assign n3940 = n3939 ^ n3929 ;
  assign n3942 = n3941 ^ n3940 ;
  assign n3943 = n3941 ^ n3518 ;
  assign n3944 = n3943 ^ n3941 ;
  assign n3945 = ~n3942 & ~n3944 ;
  assign n3946 = n3945 ^ n3941 ;
  assign n3947 = ~x31 & n3946 ;
  assign n3948 = n3947 ^ n3939 ;
  assign n3872 = n3185 ^ n1332 ;
  assign n3871 = n3870 ^ n3166 ;
  assign n3873 = n3872 ^ n3871 ;
  assign n3868 = n3867 ^ n385 ;
  assign n3866 = n1236 ^ n690 ;
  assign n3869 = n3868 ^ n3866 ;
  assign n3874 = n3873 ^ n3869 ;
  assign n3875 = n3874 ^ n1724 ;
  assign n3920 = n429 ^ n188 ;
  assign n3921 = n3920 ^ n746 ;
  assign n3919 = n943 ^ n362 ;
  assign n3922 = n3921 ^ n3919 ;
  assign n3916 = n513 ^ n178 ;
  assign n3917 = n3916 ^ n137 ;
  assign n3914 = n719 ^ n192 ;
  assign n3915 = n3914 ^ n272 ;
  assign n3918 = n3917 ^ n3915 ;
  assign n3923 = n3922 ^ n3918 ;
  assign n3924 = n3923 ^ n2203 ;
  assign n3910 = n3909 ^ n2898 ;
  assign n3908 = n2072 ^ n602 ;
  assign n3911 = n3910 ^ n3908 ;
  assign n3906 = n1327 ^ n346 ;
  assign n3907 = n3906 ^ n597 ;
  assign n3912 = n3911 ^ n3907 ;
  assign n3904 = n665 ^ n355 ;
  assign n3903 = n785 ^ n391 ;
  assign n3905 = n3904 ^ n3903 ;
  assign n3913 = n3912 ^ n3905 ;
  assign n3925 = n3924 ^ n3913 ;
  assign n3898 = n3897 ^ n777 ;
  assign n3895 = n1189 ^ n261 ;
  assign n3896 = n3895 ^ n3036 ;
  assign n3899 = n3898 ^ n3896 ;
  assign n3893 = n1441 ^ n1064 ;
  assign n3891 = n3890 ^ n918 ;
  assign n3892 = n3891 ^ n396 ;
  assign n3894 = n3893 ^ n3892 ;
  assign n3900 = n3899 ^ n3894 ;
  assign n3886 = n1037 ^ n211 ;
  assign n3888 = n3887 ^ n3886 ;
  assign n3884 = n1184 ^ n577 ;
  assign n3885 = n3884 ^ n2459 ;
  assign n3889 = n3888 ^ n3885 ;
  assign n3901 = n3900 ^ n3889 ;
  assign n3902 = n3901 ^ n3883 ;
  assign n3926 = n3925 ^ n3902 ;
  assign n3927 = ~n3875 & ~n3926 ;
  assign n3928 = n3927 ^ n3729 ;
  assign n4380 = n3948 ^ n3928 ;
  assign n4421 = n4420 ^ n4380 ;
  assign n4415 = n4365 ^ n4348 ;
  assign n4416 = n4377 & n4415 ;
  assign n4422 = n4421 ^ n4416 ;
  assign n4607 = n4444 ^ n4422 ;
  assign n12221 = n12220 ^ n4607 ;
  assign n12215 = n4644 ^ n4605 ;
  assign n12216 = ~n4649 & ~n12215 ;
  assign n12222 = n12221 ^ n12216 ;
  assign n13227 = ~n12222 & n13226 ;
  assign n13236 = n13235 ^ n13227 ;
  assign n13237 = n13224 ^ n3978 ;
  assign n13238 = ~n13236 & ~n13237 ;
  assign n12859 = ~n61 & n12235 ;
  assign n13186 = x31 & n12859 ;
  assign n12805 = n12368 ^ n12345 ;
  assign n12806 = x31 & ~n12805 ;
  assign n13184 = n12806 ^ n12228 ;
  assign n13185 = n3518 & ~n13184 ;
  assign n13187 = n13186 ^ n13185 ;
  assign n13183 = ~n3850 & n12229 ;
  assign n13188 = n13187 ^ n13183 ;
  assign n13181 = n3837 & ~n12382 ;
  assign n13179 = n3985 & n12376 ;
  assign n12549 = n12382 ^ n12376 ;
  assign n12552 = n12370 & n12382 ;
  assign n12553 = n12552 ^ n12346 ;
  assign n12554 = ~n12549 & ~n12553 ;
  assign n13172 = n12380 ^ x29 ;
  assign n13173 = n13172 ^ x28 ;
  assign n13174 = n13173 ^ n12380 ;
  assign n13175 = n12554 & n13174 ;
  assign n13176 = n13175 ^ n12380 ;
  assign n13177 = n3833 & n13176 ;
  assign n13178 = n13177 ^ x29 ;
  assign n13180 = n13179 ^ n13178 ;
  assign n13182 = n13181 ^ n13180 ;
  assign n13190 = n13188 ^ n13182 ;
  assign n12866 = n12367 ^ n12344 ;
  assign n12867 = n12866 ^ n12229 ;
  assign n12868 = n12867 ^ n12235 ;
  assign n12863 = n12239 ^ n12235 ;
  assign n12869 = n12868 ^ n12863 ;
  assign n12870 = n61 & n12869 ;
  assign n12871 = n12870 ^ n12863 ;
  assign n12872 = n5280 & ~n12871 ;
  assign n12873 = n12872 ^ n12235 ;
  assign n12860 = n12859 ^ n12235 ;
  assign n12800 = n3518 & n12229 ;
  assign n12861 = n12860 ^ n12800 ;
  assign n12862 = ~x31 & n12861 ;
  assign n12874 = n12873 ^ n12862 ;
  assign n12831 = n4906 ^ n3533 ;
  assign n12832 = n12831 ^ n1658 ;
  assign n12833 = n12832 ^ n3712 ;
  assign n12828 = n3008 ^ n2303 ;
  assign n12829 = n12828 ^ n2634 ;
  assign n12826 = n3621 ^ n1925 ;
  assign n12825 = n4034 ^ n396 ;
  assign n12827 = n12826 ^ n12825 ;
  assign n12830 = n12829 ^ n12827 ;
  assign n12834 = n12833 ^ n12830 ;
  assign n12822 = n2054 ^ n909 ;
  assign n12821 = n3036 ^ n1998 ;
  assign n12823 = n12822 ^ n12821 ;
  assign n12819 = n4722 ^ n1086 ;
  assign n12820 = n12819 ^ n1736 ;
  assign n12824 = n12823 ^ n12820 ;
  assign n12835 = n12834 ^ n12824 ;
  assign n12836 = n12835 ^ n3400 ;
  assign n12854 = n3061 ^ n598 ;
  assign n12848 = n469 ^ n142 ;
  assign n12849 = n12848 ^ n836 ;
  assign n12847 = n585 ^ n577 ;
  assign n12850 = n12849 ^ n12847 ;
  assign n12851 = n12850 ^ n6330 ;
  assign n12843 = n1179 ^ n910 ;
  assign n12842 = n903 ^ n252 ;
  assign n12844 = n12843 ^ n12842 ;
  assign n12840 = n476 ^ n137 ;
  assign n12841 = n12840 ^ n2187 ;
  assign n12845 = n12844 ^ n12841 ;
  assign n12837 = n567 ^ n369 ;
  assign n12838 = n12837 ^ n1384 ;
  assign n12839 = n12838 ^ n4242 ;
  assign n12846 = n12845 ^ n12839 ;
  assign n12852 = n12851 ^ n12846 ;
  assign n12853 = n12852 ^ n4720 ;
  assign n12855 = n12854 ^ n12853 ;
  assign n12856 = ~n12836 & ~n12855 ;
  assign n12875 = n12874 ^ n12856 ;
  assign n12889 = n4160 ^ n4063 ;
  assign n12886 = n236 ^ n145 ;
  assign n12887 = n12886 ^ n526 ;
  assign n12885 = n903 ^ n510 ;
  assign n12888 = n12887 ^ n12885 ;
  assign n12890 = n12889 ^ n12888 ;
  assign n12884 = n4779 ^ n1349 ;
  assign n12891 = n12890 ^ n12884 ;
  assign n12880 = n6062 ^ n178 ;
  assign n12881 = n12880 ^ n2187 ;
  assign n12879 = n1362 ^ n735 ;
  assign n12882 = n12881 ^ n12879 ;
  assign n12876 = n1544 ^ n774 ;
  assign n12877 = n12876 ^ n2035 ;
  assign n12878 = n12877 ^ n4716 ;
  assign n12883 = n12882 ^ n12878 ;
  assign n12892 = n12891 ^ n12883 ;
  assign n12893 = n12892 ^ n2490 ;
  assign n12894 = n6692 ^ n2518 ;
  assign n12895 = ~n12893 & ~n12894 ;
  assign n12896 = n12895 ^ n6546 ;
  assign n12909 = n934 ^ n592 ;
  assign n12910 = n12909 ^ n5533 ;
  assign n12902 = n585 ^ n513 ;
  assign n12903 = n12902 ^ n3270 ;
  assign n12904 = n12903 ^ n3645 ;
  assign n12900 = n1673 ^ n814 ;
  assign n12901 = n12900 ^ n1849 ;
  assign n12905 = n12904 ^ n12901 ;
  assign n12899 = n5730 ^ n519 ;
  assign n12906 = n12905 ^ n12899 ;
  assign n12907 = n12906 ^ n1965 ;
  assign n12908 = n12907 ^ n3108 ;
  assign n12911 = n12910 ^ n12908 ;
  assign n12912 = ~n1196 & ~n12911 ;
  assign n12913 = n12912 ^ n6546 ;
  assign n12914 = n12896 & n12913 ;
  assign n12897 = n12856 ^ n6546 ;
  assign n12915 = n12914 ^ n12897 ;
  assign n12916 = n12875 & ~n12915 ;
  assign n12917 = n12916 ^ n12856 ;
  assign n13240 = n13188 ^ n12917 ;
  assign n13243 = ~n13190 & ~n13240 ;
  assign n12769 = n4541 ^ n4209 ;
  assign n12782 = n1276 ^ n919 ;
  assign n12780 = n706 ^ n655 ;
  assign n12781 = n12780 ^ n435 ;
  assign n12783 = n12782 ^ n12781 ;
  assign n12778 = n751 ^ n278 ;
  assign n12777 = n4778 ^ n514 ;
  assign n12779 = n12778 ^ n12777 ;
  assign n12784 = n12783 ^ n12779 ;
  assign n12775 = n3401 ^ n982 ;
  assign n12774 = n2120 ^ n737 ;
  assign n12776 = n12775 ^ n12774 ;
  assign n12785 = n12784 ^ n12776 ;
  assign n12772 = n1084 ^ n250 ;
  assign n12771 = n3686 ^ n382 ;
  assign n12773 = n12772 ^ n12771 ;
  assign n12786 = n12785 ^ n12773 ;
  assign n12770 = n5676 ^ n1212 ;
  assign n12787 = n12786 ^ n12770 ;
  assign n12788 = n12787 ^ n2933 ;
  assign n12789 = ~n12769 & ~n12788 ;
  assign n13239 = n12856 ^ n12789 ;
  assign n13214 = n13182 ^ n12789 ;
  assign n13241 = n13240 ^ n13214 ;
  assign n13242 = n13239 & n13241 ;
  assign n13244 = n13243 ^ n13242 ;
  assign n3550 = n784 ^ n277 ;
  assign n3551 = n3550 ^ n434 ;
  assign n3552 = n3551 ^ n335 ;
  assign n3549 = n3548 ^ n3212 ;
  assign n3553 = n3552 ^ n3549 ;
  assign n3547 = n3344 ^ n1140 ;
  assign n3554 = n3553 ^ n3547 ;
  assign n3557 = n3556 ^ n3554 ;
  assign n3545 = n1008 ^ n395 ;
  assign n3546 = n3545 ^ n340 ;
  assign n3558 = n3557 ^ n3546 ;
  assign n12765 = n3558 ^ n3134 ;
  assign n12470 = n766 ^ n239 ;
  assign n12760 = n12470 ^ n1291 ;
  assign n12759 = n926 ^ n916 ;
  assign n12761 = n12760 ^ n12759 ;
  assign n12755 = n3209 ^ n493 ;
  assign n12756 = n12755 ^ n722 ;
  assign n12757 = n12756 ^ n427 ;
  assign n12758 = n12757 ^ n2352 ;
  assign n12762 = n12761 ^ n12758 ;
  assign n12753 = n6045 ^ n3227 ;
  assign n12754 = n12753 ^ n2964 ;
  assign n12763 = n12762 ^ n12754 ;
  assign n12504 = n1308 ^ n610 ;
  assign n12505 = n12504 ^ n390 ;
  assign n12506 = n12505 ^ n603 ;
  assign n12502 = n830 ^ n570 ;
  assign n12503 = n12502 ^ n675 ;
  assign n12507 = n12506 ^ n12503 ;
  assign n12500 = n4761 ^ n1330 ;
  assign n12501 = n12500 ^ n2331 ;
  assign n12508 = n12507 ^ n12501 ;
  assign n12764 = n12763 ^ n12508 ;
  assign n12766 = n12765 ^ n12764 ;
  assign n12767 = ~n5359 & ~n12766 ;
  assign n6156 = x17 & n6155 ;
  assign n6157 = ~n6153 & n6156 ;
  assign n6158 = n6157 ^ n6155 ;
  assign n12768 = n12767 ^ n6158 ;
  assign n12817 = n12789 ^ n12768 ;
  assign n12812 = n3801 ^ n52 ;
  assign n12793 = n12229 ^ n12228 ;
  assign n12809 = ~n12793 & n12806 ;
  assign n12810 = n12809 ^ n12382 ;
  assign n12811 = n3518 & n12810 ;
  assign n12813 = n12812 ^ n12811 ;
  assign n12801 = n12800 ^ n12228 ;
  assign n12802 = x31 & n12801 ;
  assign n12814 = n12813 ^ n12802 ;
  assign n12815 = n22543 ^ n12814 ;
  assign n12797 = ~n12229 & n22543 ;
  assign n12798 = n12797 ^ n12228 ;
  assign n12799 = ~n61 & ~n12798 ;
  assign n12816 = n12815 ^ n12799 ;
  assign n12818 = n12817 ^ n12816 ;
  assign n13245 = n13244 ^ n12818 ;
  assign n13246 = ~n13238 & n13245 ;
  assign n13189 = n13182 & n13188 ;
  assign n13191 = n13190 ^ n13189 ;
  assign n13170 = n12856 & ~n12917 ;
  assign n13171 = n13170 ^ n12916 ;
  assign n13192 = n13170 ^ n12789 ;
  assign n13193 = ~n13171 & ~n13192 ;
  assign n13194 = n13191 & n13193 ;
  assign n13201 = n13170 & n13189 ;
  assign n13202 = n13201 ^ n12818 ;
  assign n13203 = ~n13194 & ~n13202 ;
  assign n13206 = n12789 & n13189 ;
  assign n13207 = ~n13170 & n13206 ;
  assign n13208 = n13207 ^ n13170 ;
  assign n13197 = n13170 ^ n12818 ;
  assign n13209 = n13208 ^ n13197 ;
  assign n13210 = ~n13203 & n13209 ;
  assign n13220 = n13210 ^ n13203 ;
  assign n13211 = n13171 & n13210 ;
  assign n13217 = ~n13190 & n13214 ;
  assign n13218 = n13217 ^ n12789 ;
  assign n13219 = n13211 & n13218 ;
  assign n13221 = n13220 ^ n13219 ;
  assign n13247 = n13246 ^ n13221 ;
  assign n12857 = n12856 ^ n12816 ;
  assign n12858 = n12857 ^ n12768 ;
  assign n12918 = n12917 ^ n12816 ;
  assign n12919 = n12918 ^ n12768 ;
  assign n12920 = ~n12858 & n12919 ;
  assign n12921 = n12920 ^ n12768 ;
  assign n12922 = ~n12818 & n12921 ;
  assign n12923 = n12922 ^ n12816 ;
  assign n12790 = n12789 ^ n6158 ;
  assign n12791 = ~n12768 & n12790 ;
  assign n12792 = n12791 ^ n12789 ;
  assign n12925 = n12923 ^ n12792 ;
  assign n12474 = n5545 ^ n3203 ;
  assign n12472 = n1407 ^ n501 ;
  assign n12471 = n12470 ^ n476 ;
  assign n12473 = n12472 ^ n12471 ;
  assign n12475 = n12474 ^ n12473 ;
  assign n12467 = n2600 ^ n340 ;
  assign n12468 = n12467 ^ n243 ;
  assign n12466 = n3919 ^ n171 ;
  assign n12469 = n12468 ^ n12466 ;
  assign n12476 = n12475 ^ n12469 ;
  assign n12463 = n6669 ^ n677 ;
  assign n12462 = n4968 ^ n182 ;
  assign n12464 = n12463 ^ n12462 ;
  assign n12459 = n974 ^ n459 ;
  assign n12460 = n12459 ^ n2543 ;
  assign n12461 = n12460 ^ n2781 ;
  assign n12465 = n12464 ^ n12461 ;
  assign n12477 = n12476 ^ n12465 ;
  assign n12494 = n773 ^ n188 ;
  assign n12493 = n1107 ^ n137 ;
  assign n12495 = n12494 ^ n12493 ;
  assign n12491 = n584 ^ n114 ;
  assign n12492 = n12491 ^ n336 ;
  assign n12496 = n12495 ^ n12492 ;
  assign n12490 = n4770 ^ n910 ;
  assign n12497 = n12496 ^ n12490 ;
  assign n12486 = n867 ^ n197 ;
  assign n12487 = n12486 ^ n909 ;
  assign n12485 = n2297 ^ n1845 ;
  assign n12488 = n12487 ^ n12485 ;
  assign n12483 = n2078 ^ n628 ;
  assign n12482 = n741 ^ n145 ;
  assign n12484 = n12483 ^ n12482 ;
  assign n12489 = n12488 ^ n12484 ;
  assign n12498 = n12497 ^ n12489 ;
  assign n12479 = n4010 ^ n189 ;
  assign n12480 = n12479 ^ n2025 ;
  assign n12478 = n968 ^ n876 ;
  assign n12481 = n12480 ^ n12478 ;
  assign n12499 = n12498 ^ n12481 ;
  assign n12509 = n12508 ^ n12499 ;
  assign n12510 = ~n3159 & ~n12509 ;
  assign n12511 = ~n12477 & n12510 ;
  assign n13167 = n12925 ^ n12511 ;
  assign n12953 = n3837 & n12380 ;
  assign n12951 = n3985 & n12222 ;
  assign n12936 = ~n3849 & n12382 ;
  assign n12546 = ~n52 & n12376 ;
  assign n12939 = n3806 & ~n12546 ;
  assign n12940 = ~n12936 & n12939 ;
  assign n12928 = n12553 ^ n12376 ;
  assign n12929 = n12928 ^ n3518 ;
  assign n12930 = n12929 ^ n12928 ;
  assign n12931 = x30 & n12228 ;
  assign n12932 = n12931 ^ n12928 ;
  assign n12933 = ~n12930 & ~n12932 ;
  assign n12934 = n12933 ^ n12928 ;
  assign n12935 = x31 & ~n12934 ;
  assign n12937 = n12936 ^ n12935 ;
  assign n12941 = n12940 ^ n12937 ;
  assign n12949 = n12941 ^ x29 ;
  assign n12391 = ~n12380 & ~n12389 ;
  assign n12424 = n12222 & ~n12391 ;
  assign n12392 = n12391 ^ n12390 ;
  assign n12393 = ~n12222 & n12392 ;
  assign n12607 = n12424 ^ n12393 ;
  assign n12946 = n5065 & ~n12607 ;
  assign n4401 = n3985 ^ n408 ;
  assign n4407 = ~n3837 & ~n4401 ;
  assign n4405 = n3837 ^ n3505 ;
  assign n4406 = ~n3985 & ~n4405 ;
  assign n4408 = n4407 ^ n4406 ;
  assign n4409 = n368 & n4408 ;
  assign n4410 = n4409 ^ n4407 ;
  assign n4411 = n4410 ^ n3505 ;
  assign n4413 = n4411 ^ x29 ;
  assign n4399 = n3983 & n4398 ;
  assign n4414 = n4413 ^ n4399 ;
  assign n3967 = x31 & ~n3518 ;
  assign n3969 = n3968 ^ n698 ;
  assign n3970 = ~n3967 & ~n3969 ;
  assign n3964 = n3807 ^ n698 ;
  assign n3965 = n3964 ^ n3929 ;
  assign n3956 = n3955 ^ n3929 ;
  assign n3957 = n3956 ^ n540 ;
  assign n3958 = n3957 ^ n3956 ;
  assign n3959 = n3956 ^ n3807 ;
  assign n3960 = n3959 ^ n3956 ;
  assign n3961 = n3958 & ~n3960 ;
  assign n3962 = n3961 ^ n3956 ;
  assign n3963 = ~x31 & n3962 ;
  assign n3966 = n3965 ^ n3963 ;
  assign n3971 = n3970 ^ n3966 ;
  assign n3954 = ~n61 & ~n698 ;
  assign n3972 = n3971 ^ n3954 ;
  assign n3660 = n1092 ^ n320 ;
  assign n3659 = n1481 ^ n416 ;
  assign n3661 = n3660 ^ n3659 ;
  assign n3657 = n1176 ^ n567 ;
  assign n3656 = n3655 ^ n550 ;
  assign n3658 = n3657 ^ n3656 ;
  assign n3662 = n3661 ^ n3658 ;
  assign n3666 = n3665 ^ n3662 ;
  assign n3651 = n3226 ^ n903 ;
  assign n3650 = n2260 ^ n722 ;
  assign n3652 = n3651 ^ n3650 ;
  assign n3648 = n3647 ^ n506 ;
  assign n3649 = n3648 ^ n3646 ;
  assign n3653 = n3652 ^ n3649 ;
  assign n3641 = n1008 ^ n336 ;
  assign n3642 = n3641 ^ n1040 ;
  assign n3640 = n4722 ^ n1095 ;
  assign n3643 = n3642 ^ n3640 ;
  assign n3638 = n604 ^ n513 ;
  assign n3637 = n867 ^ n615 ;
  assign n3639 = n3638 ^ n3637 ;
  assign n3644 = n3643 ^ n3639 ;
  assign n3654 = n3653 ^ n3644 ;
  assign n3667 = n3666 ^ n3654 ;
  assign n3632 = n3631 ^ n339 ;
  assign n3630 = n836 ^ n813 ;
  assign n3633 = n3632 ^ n3630 ;
  assign n3628 = n2033 ^ n1067 ;
  assign n3627 = n3626 ^ n1321 ;
  assign n3629 = n3628 ^ n3627 ;
  assign n3634 = n3633 ^ n3629 ;
  assign n3635 = n3634 ^ n885 ;
  assign n3620 = n589 ^ n485 ;
  assign n3623 = n3622 ^ n3620 ;
  assign n3619 = n1020 ^ n908 ;
  assign n3624 = n3623 ^ n3619 ;
  assign n3625 = n3624 ^ n3618 ;
  assign n3636 = n3635 ^ n3625 ;
  assign n3668 = n3667 ^ n3636 ;
  assign n3669 = ~n3376 & ~n3668 ;
  assign n3951 = n3669 ^ x26 ;
  assign n3994 = n3972 ^ n3951 ;
  assign n3949 = n3948 ^ n3927 ;
  assign n3950 = ~n3928 & ~n3949 ;
  assign n3995 = n3994 ^ n3950 ;
  assign n12211 = n4414 ^ n3995 ;
  assign n4353 = ~n4348 & n4351 ;
  assign n4354 = n4353 ^ n4352 ;
  assign n4378 = n3949 & n4377 ;
  assign n4379 = n4366 & n4378 ;
  assign n4381 = n4380 ^ n4379 ;
  assign n4382 = ~n4354 & ~n4381 ;
  assign n4383 = n4380 ^ n4353 ;
  assign n4385 = n4380 ^ n3729 ;
  assign n4384 = n4380 ^ n4365 ;
  assign n4386 = n4385 ^ n4384 ;
  assign n4387 = n4385 ^ n4377 ;
  assign n4388 = n4387 ^ n4385 ;
  assign n4389 = ~n4386 & n4388 ;
  assign n4390 = n4389 ^ n4385 ;
  assign n4391 = ~n4383 & ~n4390 ;
  assign n4392 = n4391 ^ n4353 ;
  assign n4393 = ~n4382 & ~n4392 ;
  assign n12212 = n12211 ^ n4393 ;
  assign n4431 = n4430 ^ n4422 ;
  assign n4445 = ~n4431 & n4444 ;
  assign n4446 = n4445 ^ n4430 ;
  assign n12213 = n12212 ^ n4446 ;
  assign n4606 = ~n4598 & ~n4605 ;
  assign n4608 = n4607 ^ n4606 ;
  assign n4646 = n4644 ^ n4610 ;
  assign n4645 = ~n4610 & ~n4644 ;
  assign n4647 = n4646 ^ n4645 ;
  assign n4648 = n4608 & n4647 ;
  assign n12081 = n12080 ^ n4608 ;
  assign n12082 = n12081 ^ n4649 ;
  assign n12083 = n4648 & n12082 ;
  assign n12084 = n4645 ^ n4607 ;
  assign n12086 = n4645 ^ n4598 ;
  assign n12085 = n12080 ^ n4645 ;
  assign n12087 = n12086 ^ n12085 ;
  assign n12088 = n12086 ^ n12080 ;
  assign n12089 = n12088 ^ n4605 ;
  assign n12090 = n12089 ^ n12086 ;
  assign n12091 = n12087 & ~n12090 ;
  assign n12092 = n12091 ^ n12086 ;
  assign n12093 = n12084 & n12092 ;
  assign n12094 = n12093 ^ n4607 ;
  assign n12095 = ~n12083 & ~n12094 ;
  assign n12214 = n12213 ^ n12095 ;
  assign n12947 = n12946 ^ n12214 ;
  assign n12948 = n3833 & ~n12947 ;
  assign n12950 = n12949 ^ n12948 ;
  assign n12952 = n12951 ^ n12950 ;
  assign n12954 = n12953 ^ n12952 ;
  assign n13168 = n13167 ^ n12954 ;
  assign n13248 = n13247 ^ n13168 ;
  assign n3814 = n3812 ^ n540 ;
  assign n3813 = n3812 ^ n698 ;
  assign n3815 = n3814 ^ n3813 ;
  assign n3818 = x30 & n3815 ;
  assign n3819 = n3818 ^ n3814 ;
  assign n3820 = ~n3518 & ~n3819 ;
  assign n3821 = n3820 ^ n3812 ;
  assign n3822 = x31 & n3821 ;
  assign n3809 = ~n540 & ~n3805 ;
  assign n3808 = ~n408 & n3807 ;
  assign n3810 = n3809 ^ n3808 ;
  assign n3823 = n3822 ^ n3810 ;
  assign n3790 = n3789 ^ n230 ;
  assign n3791 = n3790 ^ n417 ;
  assign n3788 = n910 ^ n815 ;
  assign n3792 = n3791 ^ n3788 ;
  assign n3786 = n1912 ^ n563 ;
  assign n3783 = n546 ^ n94 ;
  assign n3784 = n3783 ^ n178 ;
  assign n3785 = n3784 ^ n1624 ;
  assign n3787 = n3786 ^ n3785 ;
  assign n3793 = n3792 ^ n3787 ;
  assign n3794 = n3793 ^ n973 ;
  assign n3778 = n2500 ^ n114 ;
  assign n3779 = n3778 ^ n409 ;
  assign n3776 = n1124 ^ n272 ;
  assign n3777 = n3776 ^ n523 ;
  assign n3780 = n3779 ^ n3777 ;
  assign n3781 = n3780 ^ n599 ;
  assign n3774 = n3773 ^ n571 ;
  assign n3769 = n991 ^ n737 ;
  assign n3771 = n3770 ^ n3769 ;
  assign n3768 = n3767 ^ n2865 ;
  assign n3772 = n3771 ^ n3768 ;
  assign n3775 = n3774 ^ n3772 ;
  assign n3782 = n3781 ^ n3775 ;
  assign n3795 = n3794 ^ n3782 ;
  assign n3763 = n3762 ^ n832 ;
  assign n3761 = n1190 ^ n270 ;
  assign n3764 = n3763 ^ n3761 ;
  assign n3758 = n3757 ^ n1077 ;
  assign n3759 = n3758 ^ n1052 ;
  assign n3755 = n1160 ^ n455 ;
  assign n3760 = n3759 ^ n3755 ;
  assign n3765 = n3764 ^ n3760 ;
  assign n3751 = n896 ^ n232 ;
  assign n3752 = n3751 ^ n1841 ;
  assign n3754 = n3753 ^ n3752 ;
  assign n3766 = n3765 ^ n3754 ;
  assign n3796 = n3795 ^ n3766 ;
  assign n3797 = ~n3750 & ~n3796 ;
  assign n3730 = n3729 ^ n3669 ;
  assign n3731 = n3729 ^ x26 ;
  assign n3732 = ~n3730 & n3731 ;
  assign n3733 = n3732 ^ x26 ;
  assign n3798 = n3797 ^ n3733 ;
  assign n3988 = n3823 ^ n3798 ;
  assign n3989 = n3988 ^ x29 ;
  assign n3987 = ~n3505 & n3837 ;
  assign n3990 = n3989 ^ n3987 ;
  assign n3986 = ~n368 & n3985 ;
  assign n3991 = n3990 ^ n3986 ;
  assign n3984 = n3515 & n3983 ;
  assign n3992 = n3991 ^ n3984 ;
  assign n3824 = n3823 ^ n3733 ;
  assign n3825 = ~n3798 & n3824 ;
  assign n3586 = n3585 ^ n920 ;
  assign n3582 = n2058 ^ n209 ;
  assign n3584 = n3583 ^ n3582 ;
  assign n3587 = n3586 ^ n3584 ;
  assign n3579 = n2670 ^ n339 ;
  assign n3577 = n965 ^ n318 ;
  assign n3578 = n3577 ^ n513 ;
  assign n3580 = n3579 ^ n3578 ;
  assign n3575 = n3574 ^ n3573 ;
  assign n3572 = n3571 ^ n2600 ;
  assign n3576 = n3575 ^ n3572 ;
  assign n3581 = n3580 ^ n3576 ;
  assign n3588 = n3587 ^ n3581 ;
  assign n3567 = n628 ^ n419 ;
  assign n3568 = n3567 ^ n2375 ;
  assign n3566 = n3565 ^ n331 ;
  assign n3569 = n3568 ^ n3566 ;
  assign n3564 = n3563 ^ n3562 ;
  assign n3570 = n3569 ^ n3564 ;
  assign n3589 = n3588 ^ n3570 ;
  assign n3590 = n3589 ^ n1563 ;
  assign n3591 = n3590 ^ n3558 ;
  assign n3592 = ~n1895 & ~n3591 ;
  assign n3857 = n3825 ^ n3592 ;
  assign n3852 = ~n540 & n22543 ;
  assign n3851 = ~n408 & ~n3850 ;
  assign n3853 = n3852 ^ n3851 ;
  assign n3846 = x31 & ~n3839 ;
  assign n3847 = n3846 ^ n3505 ;
  assign n3848 = n3518 & ~n3847 ;
  assign n3854 = n3853 ^ n3848 ;
  assign n3855 = n3854 ^ x29 ;
  assign n3838 = ~n368 & n3837 ;
  assign n3856 = n3855 ^ n3838 ;
  assign n12113 = n3857 ^ n3856 ;
  assign n12115 = n12113 ^ n3988 ;
  assign n3952 = n3951 ^ n3950 ;
  assign n3953 = n3950 ^ n3729 ;
  assign n3973 = n3972 ^ n3953 ;
  assign n3974 = n3952 & ~n3973 ;
  assign n3975 = n3974 ^ n3972 ;
  assign n12116 = n12115 ^ n3975 ;
  assign n12117 = n12116 ^ n12113 ;
  assign n12118 = ~n3992 & n12117 ;
  assign n12119 = n12118 ^ n12115 ;
  assign n3993 = n3992 ^ n3975 ;
  assign n4395 = n4393 ^ n3995 ;
  assign n4394 = ~n3995 & ~n4393 ;
  assign n4396 = n4395 ^ n4394 ;
  assign n4397 = ~n3993 & n4396 ;
  assign n4448 = n4414 & ~n4446 ;
  assign n4447 = n4446 ^ n4414 ;
  assign n4449 = n4448 ^ n4447 ;
  assign n4450 = n4449 ^ n3993 ;
  assign n12096 = n12095 ^ n3995 ;
  assign n12097 = n4395 & n12096 ;
  assign n12098 = n12097 ^ n3995 ;
  assign n12099 = n4450 & n12098 ;
  assign n12100 = n4394 ^ n3993 ;
  assign n12101 = n12100 ^ n4447 ;
  assign n12102 = n12101 ^ n12100 ;
  assign n12103 = ~n3993 & ~n4414 ;
  assign n12104 = n12103 ^ n12100 ;
  assign n12105 = n12102 & ~n12104 ;
  assign n12106 = n12105 ^ n12100 ;
  assign n12107 = ~n12095 & ~n12106 ;
  assign n12108 = n12107 ^ n4448 ;
  assign n12109 = ~n12099 & n12108 ;
  assign n12110 = n12109 ^ n12099 ;
  assign n12111 = n4397 & ~n12110 ;
  assign n12112 = n12111 ^ n12109 ;
  assign n12210 = n12119 ^ n12112 ;
  assign n12397 = n12095 ^ n4448 ;
  assign n12398 = ~n12213 & n12397 ;
  assign n12399 = n12398 ^ n3993 ;
  assign n12395 = n4449 ^ n4393 ;
  assign n12396 = ~n4395 & ~n12395 ;
  assign n12400 = n12399 ^ n12396 ;
  assign n12425 = n12214 & ~n12424 ;
  assign n12426 = ~n12400 & ~n12425 ;
  assign n12427 = n12210 & ~n12426 ;
  assign n12394 = ~n12214 & ~n12393 ;
  assign n12401 = ~n12394 & n12400 ;
  assign n12402 = ~n12210 & ~n12401 ;
  assign n12714 = n12427 ^ n12402 ;
  assign n12125 = n4398 ^ n408 ;
  assign n12124 = n4398 ^ n3505 ;
  assign n12126 = n12125 ^ n12124 ;
  assign n12129 = ~x30 & n12126 ;
  assign n12130 = n12129 ^ n12125 ;
  assign n12131 = ~n3518 & ~n12130 ;
  assign n12132 = n12131 ^ n4398 ;
  assign n12133 = x31 & n12132 ;
  assign n3539 = n1689 ^ n321 ;
  assign n3540 = n3539 ^ n173 ;
  assign n3594 = n3540 ^ n341 ;
  assign n310 = ~n20602 ^ n48 ;
  assign n311 = n224 & n310 ;
  assign n313 = n312 ^ n311 ;
  assign n3596 = n563 ^ n313 ;
  assign n3595 = n572 ^ n177 ;
  assign n3597 = n3596 ^ n3595 ;
  assign n3598 = n421 ^ n253 ;
  assign n3599 = n3598 ^ n2078 ;
  assign n3600 = n3599 ^ n129 ;
  assign n3601 = ~n3597 & ~n3600 ;
  assign n3602 = n3594 & n3601 ;
  assign n3605 = n3604 ^ n3603 ;
  assign n3606 = n3605 ^ n539 ;
  assign n3607 = n3602 & n3606 ;
  assign n3863 = n3607 ^ x29 ;
  assign n3864 = n3863 ^ n3592 ;
  assign n12134 = n12133 ^ n3864 ;
  assign n3826 = n3823 ^ n3592 ;
  assign n3827 = ~n3825 & n3826 ;
  assign n3828 = n3827 ^ n3823 ;
  assign n12403 = n12134 ^ n3828 ;
  assign n3858 = n3857 ^ n3854 ;
  assign n3859 = ~n3856 & ~n3858 ;
  assign n3860 = n3859 ^ n3857 ;
  assign n12404 = n12403 ^ n3860 ;
  assign n12114 = n12113 ^ n12112 ;
  assign n12120 = n12114 & n12119 ;
  assign n12121 = n12120 ^ n12113 ;
  assign n12405 = n12404 ^ n12121 ;
  assign n12715 = n12714 ^ n12405 ;
  assign n13255 = ~n4435 & n12715 ;
  assign n13253 = ~n4434 & ~n12405 ;
  assign n13250 = ~n12400 & n20603 ;
  assign n13249 = n4600 & ~n12210 ;
  assign n13251 = n13250 ^ n13249 ;
  assign n13252 = n13251 ^ x26 ;
  assign n13254 = n13253 ^ n13252 ;
  assign n13256 = n13255 ^ n13254 ;
  assign n13106 = n4600 & ~n12405 ;
  assign n13105 = ~n12210 & n20603 ;
  assign n13107 = n13106 ^ n13105 ;
  assign n13108 = n13107 ^ n97 ;
  assign n12428 = ~n12405 & ~n12427 ;
  assign n12406 = ~n12402 & n12405 ;
  assign n12650 = n12428 ^ n12406 ;
  assign n13110 = n99 ^ x25 ;
  assign n13131 = ~n12650 & ~n13110 ;
  assign n12141 = n12134 ^ n12121 ;
  assign n12407 = ~n3864 & n12133 ;
  assign n3861 = n3828 & ~n3860 ;
  assign n12413 = n12121 ^ n3861 ;
  assign n12416 = ~n12407 & n12413 ;
  assign n12142 = n3860 ^ n3828 ;
  assign n12143 = n12142 ^ n3861 ;
  assign n12408 = n12407 ^ n12143 ;
  assign n3593 = n3592 ^ x29 ;
  assign n3608 = n3607 ^ n3592 ;
  assign n3609 = n3593 & ~n3608 ;
  assign n3610 = n3609 ^ x29 ;
  assign n3524 = n1037 ^ n435 ;
  assign n3525 = n3524 ^ n195 ;
  assign n3526 = n3525 ^ n181 ;
  assign n3527 = n3526 ^ n360 ;
  assign n3537 = n3536 ^ n3527 ;
  assign n3538 = ~n1007 & n3537 ;
  assign n3542 = n282 ^ n242 ;
  assign n3541 = n3540 ^ n161 ;
  assign n3543 = n3542 ^ n3541 ;
  assign n3544 = n3538 & n3543 ;
  assign n3611 = n3610 ^ n3544 ;
  assign n3521 = n3515 & n3518 ;
  assign n3522 = n3521 ^ n368 ;
  assign n3523 = x31 & ~n3522 ;
  assign n3612 = n3611 ^ n3523 ;
  assign n12409 = n12408 ^ n3612 ;
  assign n12410 = n12409 ^ n3612 ;
  assign n12417 = n12416 ^ n12410 ;
  assign n12418 = ~n12141 & n12417 ;
  assign n12419 = n12418 ^ n12409 ;
  assign n13125 = n12419 ^ n99 ;
  assign n13111 = n13110 ^ n12419 ;
  assign n13109 = n13107 ^ x26 ;
  assign n13112 = n13111 ^ n13109 ;
  assign n13113 = n13112 ^ n99 ;
  assign n13114 = n13113 ^ n13111 ;
  assign n13119 = ~n12650 & n13110 ;
  assign n12651 = n12650 ^ n12419 ;
  assign n13120 = n13119 ^ n12651 ;
  assign n13121 = ~n13114 & n13120 ;
  assign n13126 = n13125 ^ n13121 ;
  assign n13132 = n13131 ^ n13126 ;
  assign n13133 = ~n13108 & n13132 ;
  assign n13103 = n3837 & n12222 ;
  assign n13101 = n3985 & ~n12214 ;
  assign n12961 = n12941 ^ n12511 ;
  assign n13095 = n12961 ^ n12925 ;
  assign n13096 = n12954 & n13095 ;
  assign n12592 = n2415 ^ n182 ;
  assign n12593 = n12592 ^ n999 ;
  assign n12591 = n2403 ^ n199 ;
  assign n12594 = n12593 ^ n12591 ;
  assign n12590 = n6809 ^ n2474 ;
  assign n12595 = n12594 ^ n12590 ;
  assign n12586 = n1432 ^ n510 ;
  assign n12584 = n842 ^ n592 ;
  assign n12585 = n12584 ^ n2058 ;
  assign n12587 = n12586 ^ n12585 ;
  assign n12582 = n1756 ^ n641 ;
  assign n12581 = n764 ^ n634 ;
  assign n12583 = n12582 ^ n12581 ;
  assign n12588 = n12587 ^ n12583 ;
  assign n12589 = n12588 ^ n1871 ;
  assign n12596 = n12595 ^ n12589 ;
  assign n12597 = n12596 ^ n2627 ;
  assign n12575 = n251 ^ n215 ;
  assign n12576 = n12575 ^ n1925 ;
  assign n12577 = n12576 ^ n3061 ;
  assign n12572 = n1124 ^ n145 ;
  assign n12573 = n12572 ^ n452 ;
  assign n12571 = n1643 ^ n354 ;
  assign n12574 = n12573 ^ n12571 ;
  assign n12578 = n12577 ^ n12574 ;
  assign n12568 = n2481 ^ n653 ;
  assign n12569 = n12568 ^ n2561 ;
  assign n12567 = n1140 ^ n731 ;
  assign n12570 = n12569 ^ n12567 ;
  assign n12579 = n12578 ^ n12570 ;
  assign n12580 = n12579 ^ n2613 ;
  assign n12598 = n12597 ^ n12580 ;
  assign n12599 = ~n5598 & ~n12598 ;
  assign n12734 = n12599 ^ n12511 ;
  assign n12545 = n12376 ^ n52 ;
  assign n12547 = n12546 ^ n12545 ;
  assign n12557 = n12380 ^ x31 ;
  assign n12558 = n12557 ^ n12380 ;
  assign n12559 = ~n12554 & n12558 ;
  assign n12560 = n12559 ^ n12380 ;
  assign n12561 = n3518 & n12560 ;
  assign n12562 = n12561 ^ x31 ;
  assign n12550 = n12549 & n22543 ;
  assign n12548 = ~n61 & n12376 ;
  assign n12551 = n12550 ^ n12548 ;
  assign n12563 = n12562 ^ n12551 ;
  assign n12564 = ~n12547 & n12563 ;
  assign n12927 = n12734 ^ n12564 ;
  assign n13097 = n13096 ^ n12927 ;
  assign n13092 = n12792 ^ n12511 ;
  assign n13093 = n12923 ^ n12511 ;
  assign n13094 = n13092 & ~n13093 ;
  assign n13098 = n13097 ^ n13094 ;
  assign n13099 = n13098 ^ x29 ;
  assign n12666 = n12425 ^ n12394 ;
  assign n13089 = ~n5065 & ~n12666 ;
  assign n12667 = n12666 ^ n12400 ;
  assign n13090 = n13089 ^ n12667 ;
  assign n13091 = n3833 & n13090 ;
  assign n13100 = n13099 ^ n13091 ;
  assign n13102 = n13101 ^ n13100 ;
  assign n13104 = n13103 ^ n13102 ;
  assign n13165 = n13133 ^ n13104 ;
  assign n13257 = n13256 ^ n13165 ;
  assign n13258 = n13257 ^ n13247 ;
  assign n13259 = n13258 ^ n13165 ;
  assign n13260 = n13248 & ~n13259 ;
  assign n13261 = n13260 ^ n13257 ;
  assign n315 = n314 ^ n313 ;
  assign n316 = n315 ^ n243 ;
  assign n324 = n323 ^ n316 ;
  assign n309 = ~n300 & ~n308 ;
  assign n325 = n324 ^ n309 ;
  assign n326 = n304 & n325 ;
  assign n12207 = n3544 ^ n326 ;
  assign n12152 = n3610 ^ n3523 ;
  assign n12153 = n3544 ^ n3523 ;
  assign n12205 = ~n12152 & ~n12153 ;
  assign n12206 = n12205 ^ n3610 ;
  assign n12208 = n12207 ^ n12206 ;
  assign n3862 = n3861 ^ n3612 ;
  assign n12122 = n12121 ^ n3612 ;
  assign n3865 = n3864 ^ n3612 ;
  assign n12123 = n12122 ^ n3865 ;
  assign n12137 = n12123 & n12134 ;
  assign n12138 = n12137 ^ n12122 ;
  assign n12139 = ~n3862 & ~n12138 ;
  assign n12140 = n12139 ^ n3861 ;
  assign n12144 = n12141 & ~n12143 ;
  assign n12147 = ~n3864 & ~n12121 ;
  assign n12148 = n12147 ^ n3612 ;
  assign n12149 = n12144 & ~n12148 ;
  assign n12150 = ~n12140 & ~n12149 ;
  assign n12209 = n12208 ^ n12150 ;
  assign n13161 = n4651 & ~n12209 ;
  assign n12434 = n558 & n12150 ;
  assign n12435 = n12206 & n12434 ;
  assign n13156 = n35 & ~n12435 ;
  assign n13160 = n13156 ^ x23 ;
  assign n13162 = n13161 ^ n13160 ;
  assign n244 = n243 ^ n242 ;
  assign n235 = n234 ^ n233 ;
  assign n245 = n244 ^ n235 ;
  assign n229 = n228 ^ n226 ;
  assign n246 = n245 ^ n229 ;
  assign n258 = n257 ^ n246 ;
  assign n259 = ~n222 & ~n258 ;
  assign n12151 = n12150 ^ n326 ;
  assign n12157 = n12152 & ~n12153 ;
  assign n12158 = n12157 ^ n3544 ;
  assign n12159 = n12152 ^ n326 ;
  assign n12160 = n12159 ^ n12152 ;
  assign n12161 = n12160 ^ n12151 ;
  assign n12162 = n12158 & ~n12161 ;
  assign n12163 = n12162 ^ n12152 ;
  assign n12164 = ~n12151 & n12163 ;
  assign n12165 = n12164 ^ n326 ;
  assign n12166 = ~n259 & n12165 ;
  assign n12178 = n57 & n3610 ;
  assign n12176 = ~n259 & ~n3523 ;
  assign n12177 = ~n3544 & n12176 ;
  assign n12179 = n12177 ^ n3523 ;
  assign n12180 = n12178 & ~n12179 ;
  assign n12181 = n12180 ^ n12177 ;
  assign n12182 = n12181 ^ n326 ;
  assign n12167 = n326 ^ n259 ;
  assign n12183 = n12182 ^ n12167 ;
  assign n12184 = n12207 ^ n12183 ;
  assign n12171 = n3610 ^ n326 ;
  assign n12172 = n12151 ^ n3523 ;
  assign n12173 = n12171 & ~n12172 ;
  assign n12174 = n12173 ^ n12167 ;
  assign n12175 = n12174 & n12207 ;
  assign n12185 = n12184 ^ n12175 ;
  assign n12186 = n12185 ^ n12181 ;
  assign n12197 = n12185 ^ n12184 ;
  assign n12198 = n12186 & ~n12197 ;
  assign n12199 = n326 & n12198 ;
  assign n12200 = n12199 ^ n326 ;
  assign n12192 = n12185 ^ n326 ;
  assign n12201 = n12200 ^ n12192 ;
  assign n12202 = ~n12150 & n12201 ;
  assign n12203 = n12202 ^ n12181 ;
  assign n12204 = ~n12166 & ~n12203 ;
  assign n13159 = ~n40 & ~n12204 ;
  assign n13163 = n13162 ^ n13159 ;
  assign n12429 = ~n12419 & ~n12428 ;
  assign n12430 = ~n12209 & ~n12429 ;
  assign n12431 = n12204 & ~n12430 ;
  assign n12420 = ~n12406 & n12419 ;
  assign n12421 = n12209 & ~n12420 ;
  assign n12422 = ~n12204 & n12421 ;
  assign n12423 = n12422 ^ n12204 ;
  assign n12432 = n12431 ^ n12423 ;
  assign n13157 = n5239 & n13156 ;
  assign n13158 = n12432 & n13157 ;
  assign n13164 = n13163 ^ n13158 ;
  assign n13267 = n13261 ^ n13164 ;
  assign n12736 = n12426 ^ n12401 ;
  assign n12737 = n12736 ^ n12210 ;
  assign n13277 = ~n4435 & n12737 ;
  assign n13272 = n13245 ^ n13238 ;
  assign n13273 = n13272 ^ x26 ;
  assign n13271 = n4600 & ~n12400 ;
  assign n13274 = n13273 ^ n13271 ;
  assign n13270 = ~n12214 & n20603 ;
  assign n13275 = n13274 ^ n13270 ;
  assign n13269 = ~n4434 & ~n12210 ;
  assign n13276 = n13275 ^ n13269 ;
  assign n13278 = n13277 ^ n13276 ;
  assign n13301 = n13239 ^ n13188 ;
  assign n13302 = n13301 ^ n12917 ;
  assign n13303 = n13302 ^ n13182 ;
  assign n13280 = n4600 & ~n12214 ;
  assign n13279 = n12222 & n20603 ;
  assign n13281 = n13280 ^ n13279 ;
  assign n13282 = n13281 ^ n97 ;
  assign n13283 = n13281 ^ x26 ;
  assign n13284 = n13283 ^ n99 ;
  assign n13285 = n13284 ^ x25 ;
  assign n13286 = n13285 ^ n13283 ;
  assign n13287 = n13286 ^ n12400 ;
  assign n13288 = n13287 ^ n12666 ;
  assign n13289 = n13288 ^ n13287 ;
  assign n13290 = n13283 & ~n13289 ;
  assign n13291 = n13290 ^ n13284 ;
  assign n13293 = ~n13286 & ~n13289 ;
  assign n13294 = n13293 ^ n12400 ;
  assign n13295 = ~n13284 & n13294 ;
  assign n13296 = ~n13291 & n13295 ;
  assign n13297 = n13296 ^ n13293 ;
  assign n13298 = n13297 ^ n99 ;
  assign n13299 = n13298 ^ n12400 ;
  assign n13300 = ~n13282 & ~n13299 ;
  assign n13304 = n13303 ^ n13300 ;
  assign n13317 = n12915 ^ n12874 ;
  assign n13407 = n13317 ^ n13303 ;
  assign n13315 = n3837 & ~n12228 ;
  assign n13313 = n3985 & ~n12382 ;
  assign n13306 = n12376 ^ x29 ;
  assign n13307 = n13306 ^ x28 ;
  assign n13308 = n13307 ^ n12376 ;
  assign n13309 = n12553 & n13308 ;
  assign n13310 = n13309 ^ n12376 ;
  assign n13311 = n3833 & n13310 ;
  assign n13312 = n13311 ^ x29 ;
  assign n13314 = n13313 ^ n13312 ;
  assign n13316 = n13315 ^ n13314 ;
  assign n13318 = n13317 ^ n13316 ;
  assign n13369 = n3574 ^ n1968 ;
  assign n13370 = n13369 ^ n2246 ;
  assign n13371 = n13370 ^ n1794 ;
  assign n13367 = n1499 ^ n1252 ;
  assign n13365 = n5483 ^ n464 ;
  assign n13364 = n422 ^ n369 ;
  assign n13366 = n13365 ^ n13364 ;
  assign n13368 = n13367 ^ n13366 ;
  assign n13372 = n13371 ^ n13368 ;
  assign n13361 = n1549 ^ n1146 ;
  assign n13360 = n1028 ^ n1011 ;
  assign n13362 = n13361 ^ n13360 ;
  assign n13359 = n1198 ^ n803 ;
  assign n13363 = n13362 ^ n13359 ;
  assign n13373 = n13372 ^ n13363 ;
  assign n13374 = n13373 ^ n3269 ;
  assign n13392 = n2672 ^ n1725 ;
  assign n13000 = n395 ^ n236 ;
  assign n13389 = n13000 ^ n490 ;
  assign n13390 = n13389 ^ n1994 ;
  assign n13388 = n1680 ^ n719 ;
  assign n13391 = n13390 ^ n13388 ;
  assign n13393 = n13392 ^ n13391 ;
  assign n13385 = n1036 ^ n564 ;
  assign n13386 = n13385 ^ n2879 ;
  assign n13384 = n4857 ^ n668 ;
  assign n13387 = n13386 ^ n13384 ;
  assign n13394 = n13393 ^ n13387 ;
  assign n13395 = n13394 ^ n4090 ;
  assign n13379 = n2638 ^ n215 ;
  assign n13380 = n13379 ^ n357 ;
  assign n13378 = n622 ^ n336 ;
  assign n13381 = n13380 ^ n13378 ;
  assign n13382 = n13381 ^ n4235 ;
  assign n13375 = n523 ^ n189 ;
  assign n13376 = n13375 ^ n534 ;
  assign n13377 = n13376 ^ n2543 ;
  assign n13383 = n13382 ^ n13377 ;
  assign n13396 = n13395 ^ n13383 ;
  assign n13397 = ~n13374 & ~n13396 ;
  assign n13339 = n12365 ^ n12342 ;
  assign n13320 = ~n61 & n12248 ;
  assign n13340 = n13339 ^ n13320 ;
  assign n13341 = n13340 ^ n3518 ;
  assign n13342 = n13341 ^ n13340 ;
  assign n13343 = n13339 ^ n12239 ;
  assign n13345 = n13343 ^ n12248 ;
  assign n13344 = n13343 ^ n12249 ;
  assign n13346 = n13345 ^ n13344 ;
  assign n13349 = x30 & ~n13346 ;
  assign n13350 = n13349 ^ n13345 ;
  assign n13351 = ~n3518 & n13350 ;
  assign n13352 = n13351 ^ n13343 ;
  assign n13353 = n13352 ^ n13320 ;
  assign n13354 = n13353 ^ n13340 ;
  assign n13355 = ~n13342 & ~n13354 ;
  assign n13356 = n13355 ^ n13340 ;
  assign n13357 = ~x31 & ~n13356 ;
  assign n13358 = n13357 ^ n13352 ;
  assign n13398 = n13397 ^ n13358 ;
  assign n13399 = n13358 ^ n12912 ;
  assign n13400 = n13398 & n13399 ;
  assign n13401 = n13400 ^ n12896 ;
  assign n13402 = n13400 ^ n12912 ;
  assign n13336 = ~n61 & ~n12239 ;
  assign n13332 = n12239 ^ n3807 ;
  assign n13333 = n13332 ^ n13320 ;
  assign n13319 = n12366 ^ n12343 ;
  assign n13329 = n13319 ^ n12235 ;
  assign n13330 = n13329 ^ n12239 ;
  assign n13331 = ~n3967 & n13330 ;
  assign n13334 = n13333 ^ n13331 ;
  assign n13321 = n13320 ^ n13319 ;
  assign n13322 = n13321 ^ n3807 ;
  assign n13323 = n13322 ^ n13321 ;
  assign n13324 = n13321 ^ n12235 ;
  assign n13325 = n13324 ^ n13321 ;
  assign n13326 = ~n13323 & ~n13325 ;
  assign n13327 = n13326 ^ n13321 ;
  assign n13328 = ~x31 & n13327 ;
  assign n13335 = n13334 ^ n13328 ;
  assign n13337 = n13336 ^ n13335 ;
  assign n13403 = n13402 ^ n13337 ;
  assign n13404 = n13401 & ~n13403 ;
  assign n13338 = n13337 ^ n13316 ;
  assign n13405 = n13404 ^ n13338 ;
  assign n13406 = ~n13318 & n13405 ;
  assign n13408 = n13407 ^ n13406 ;
  assign n13409 = n13304 & n13408 ;
  assign n13410 = n13409 ^ n13303 ;
  assign n13411 = n13410 ^ n13272 ;
  assign n13412 = ~n13278 & n13411 ;
  assign n13413 = n13412 ^ n13272 ;
  assign n13268 = n13256 ^ n13248 ;
  assign n13414 = n13413 ^ n13268 ;
  assign n13425 = n4651 & n12419 ;
  assign n13423 = ~n40 & ~n12209 ;
  assign n12982 = n12430 ^ n12421 ;
  assign n12983 = n12982 ^ n12204 ;
  assign n13415 = n12983 ^ n12204 ;
  assign n13416 = n12204 ^ x23 ;
  assign n13417 = n13416 ^ x22 ;
  assign n13418 = n13417 ^ n12204 ;
  assign n13419 = ~n13415 & n13418 ;
  assign n13420 = n13419 ^ n12204 ;
  assign n13421 = n35 & ~n13420 ;
  assign n13422 = n13421 ^ x23 ;
  assign n13424 = n13423 ^ n13422 ;
  assign n13426 = n13425 ^ n13424 ;
  assign n13427 = n13426 ^ n13413 ;
  assign n13428 = n13414 & ~n13427 ;
  assign n13429 = n13428 ^ n13413 ;
  assign n13430 = n13267 & n13429 ;
  assign n13051 = n12429 ^ n12420 ;
  assign n13740 = ~x22 & ~n13051 ;
  assign n13052 = n13051 ^ n12209 ;
  assign n13746 = n13740 ^ n13052 ;
  assign n13747 = n13745 & n13746 ;
  assign n13737 = ~n40 & n12419 ;
  assign n13736 = n4651 & ~n12405 ;
  assign n13738 = n13737 ^ n13736 ;
  assign n13739 = n13738 ^ x23 ;
  assign n13741 = n13740 ^ n12209 ;
  assign n13742 = n13739 & n13741 ;
  assign n13748 = n13747 ^ n13742 ;
  assign n13749 = n13743 ^ n13738 ;
  assign n13750 = ~n13748 & ~n13749 ;
  assign n13734 = n13410 ^ n13278 ;
  assign n13443 = n13408 ^ n13300 ;
  assign n13441 = ~n40 & ~n12405 ;
  assign n13439 = n4656 & ~n12651 ;
  assign n13436 = n4655 & n12419 ;
  assign n13435 = n4651 & ~n12210 ;
  assign n13437 = n13436 ^ n13435 ;
  assign n13438 = n13437 ^ x23 ;
  assign n13440 = n13439 ^ n13438 ;
  assign n13442 = n13441 ^ n13440 ;
  assign n13444 = n13443 ^ n13442 ;
  assign n13719 = n13405 ^ n13317 ;
  assign n13456 = n3837 & n12229 ;
  assign n13454 = n3985 & ~n12228 ;
  assign n13445 = n12382 ^ n12370 ;
  assign n13446 = n13445 ^ n12382 ;
  assign n13447 = n12382 ^ x29 ;
  assign n13448 = n13447 ^ x28 ;
  assign n13449 = n13448 ^ n12382 ;
  assign n13450 = ~n13446 & n13449 ;
  assign n13451 = n13450 ^ n12382 ;
  assign n13452 = n3833 & ~n13451 ;
  assign n13453 = n13452 ^ x29 ;
  assign n13455 = n13454 ^ n13453 ;
  assign n13457 = n13456 ^ n13455 ;
  assign n13458 = n13457 ^ n12896 ;
  assign n13459 = n13458 ^ n13337 ;
  assign n13460 = n13459 ^ n13400 ;
  assign n13704 = n13398 ^ n12912 ;
  assign n13542 = n3837 & ~n12239 ;
  assign n13540 = n3985 & n12235 ;
  assign n13533 = n12229 ^ x29 ;
  assign n13534 = n13533 ^ x28 ;
  assign n13535 = n13534 ^ n12229 ;
  assign n13536 = ~n12866 & n13535 ;
  assign n13537 = n13536 ^ n12229 ;
  assign n13538 = n3833 & n13537 ;
  assign n13539 = n13538 ^ x29 ;
  assign n13541 = n13540 ^ n13539 ;
  assign n13543 = n13542 ^ n13541 ;
  assign n13518 = n12364 ^ n12341 ;
  assign n13519 = n13518 ^ n12248 ;
  assign n13521 = n13519 ^ n12249 ;
  assign n13520 = n13519 ^ n12339 ;
  assign n13522 = n13521 ^ n13520 ;
  assign n13525 = x30 & ~n13522 ;
  assign n13526 = n13525 ^ n13521 ;
  assign n13527 = ~n3518 & n13526 ;
  assign n13528 = n13527 ^ n13519 ;
  assign n13529 = x31 & ~n13528 ;
  assign n13516 = n3807 & n12248 ;
  assign n13515 = ~n3805 & ~n12249 ;
  assign n13517 = n13516 ^ n13515 ;
  assign n13530 = n13529 ^ n13517 ;
  assign n13469 = n1769 ^ n237 ;
  assign n13470 = n13469 ^ n598 ;
  assign n13467 = n722 ^ n183 ;
  assign n13468 = n13467 ^ n331 ;
  assign n13471 = n13470 ^ n13468 ;
  assign n12692 = n513 ^ n251 ;
  assign n13465 = n12692 ^ n1432 ;
  assign n13464 = n1837 ^ n1038 ;
  assign n13466 = n13465 ^ n13464 ;
  assign n13472 = n13471 ^ n13466 ;
  assign n13462 = n1157 ^ n648 ;
  assign n13461 = n12490 ^ n3355 ;
  assign n13463 = n13462 ^ n13461 ;
  assign n13473 = n13472 ^ n13463 ;
  assign n13474 = n13473 ^ n854 ;
  assign n13475 = n6048 ^ n1911 ;
  assign n13476 = n13475 ^ n1320 ;
  assign n13477 = ~n13474 & ~n13476 ;
  assign n13478 = n13477 ^ n7147 ;
  assign n13484 = n805 ^ n322 ;
  assign n13485 = n13484 ^ n1442 ;
  assign n13486 = n13485 ^ n1233 ;
  assign n13481 = n664 ^ n618 ;
  assign n13482 = n13481 ^ n3295 ;
  assign n13480 = n778 ^ n250 ;
  assign n13483 = n13482 ^ n13480 ;
  assign n13487 = n13486 ^ n13483 ;
  assign n13479 = n2363 ^ n184 ;
  assign n13488 = n13487 ^ n13479 ;
  assign n13502 = n1198 ^ n957 ;
  assign n13503 = n13502 ^ n157 ;
  assign n13504 = n13503 ^ n764 ;
  assign n13501 = n800 ^ n471 ;
  assign n13505 = n13504 ^ n13501 ;
  assign n13499 = n1837 ^ n343 ;
  assign n13498 = n2677 ^ n1607 ;
  assign n13500 = n13499 ^ n13498 ;
  assign n13506 = n13505 ^ n13500 ;
  assign n13495 = n4211 ^ n2310 ;
  assign n13493 = n5543 ^ n1437 ;
  assign n13492 = n1216 ^ n435 ;
  assign n13494 = n13493 ^ n13492 ;
  assign n13496 = n13495 ^ n13494 ;
  assign n13490 = n1716 ^ n776 ;
  assign n13489 = n3604 ^ n905 ;
  assign n13491 = n13490 ^ n13489 ;
  assign n13497 = n13496 ^ n13491 ;
  assign n13507 = n13506 ^ n13497 ;
  assign n13508 = n13507 ^ n6274 ;
  assign n13509 = ~n3376 & ~n13508 ;
  assign n13510 = ~n13488 & n13509 ;
  assign n13511 = n13510 ^ n7147 ;
  assign n13512 = n13478 & n13511 ;
  assign n13513 = n13512 ^ n7147 ;
  assign n13514 = n13513 ^ n12912 ;
  assign n13531 = n13530 ^ n13514 ;
  assign n13544 = n13543 ^ n13531 ;
  assign n13567 = n13510 ^ n13478 ;
  assign n13553 = n12363 ^ n12340 ;
  assign n13554 = n13553 ^ n12249 ;
  assign n13556 = n13554 ^ n12251 ;
  assign n13555 = n13554 ^ n12339 ;
  assign n13557 = n13556 ^ n13555 ;
  assign n13560 = ~x30 & ~n13557 ;
  assign n13561 = n13560 ^ n13556 ;
  assign n13562 = ~n3518 & ~n13561 ;
  assign n13563 = n13562 ^ n13554 ;
  assign n13564 = x31 & n13563 ;
  assign n13545 = n12339 ^ n12249 ;
  assign n13550 = ~n61 & ~n13545 ;
  assign n13551 = n13550 ^ n12249 ;
  assign n13552 = ~n3800 & ~n13551 ;
  assign n13565 = n13564 ^ n13552 ;
  assign n13568 = n13567 ^ n13565 ;
  assign n13584 = n12692 ^ n2082 ;
  assign n13583 = n3714 ^ n905 ;
  assign n13585 = n13584 ^ n13583 ;
  assign n13581 = n3550 ^ n2033 ;
  assign n13582 = n13581 ^ n2153 ;
  assign n13586 = n13585 ^ n13582 ;
  assign n13578 = n1401 ^ n555 ;
  assign n13577 = n743 ^ n737 ;
  assign n13579 = n13578 ^ n13577 ;
  assign n13580 = n13579 ^ n1025 ;
  assign n13587 = n13586 ^ n13580 ;
  assign n13573 = n1864 ^ n915 ;
  assign n13574 = n13573 ^ n1106 ;
  assign n13572 = n765 ^ n269 ;
  assign n13575 = n13574 ^ n13572 ;
  assign n13570 = n1129 ^ n1095 ;
  assign n13569 = n1233 ^ n800 ;
  assign n13571 = n13570 ^ n13569 ;
  assign n13576 = n13575 ^ n13571 ;
  assign n13588 = n13587 ^ n13576 ;
  assign n13589 = n13588 ^ n2653 ;
  assign n13600 = n3362 ^ n137 ;
  assign n13598 = n2185 ^ n149 ;
  assign n13599 = n13598 ^ n314 ;
  assign n13601 = n13600 ^ n13599 ;
  assign n13602 = n13601 ^ n2995 ;
  assign n13603 = n13602 ^ n2889 ;
  assign n13595 = n13367 ^ n1361 ;
  assign n13593 = n1743 ^ n711 ;
  assign n13592 = n12584 ^ n2204 ;
  assign n13594 = n13593 ^ n13592 ;
  assign n13596 = n13595 ^ n13594 ;
  assign n13590 = n1674 ^ n1050 ;
  assign n13591 = n13590 ^ n1124 ;
  assign n13597 = n13596 ^ n13591 ;
  assign n13604 = n13603 ^ n13597 ;
  assign n13605 = n13604 ^ n4920 ;
  assign n13606 = ~n13589 & ~n13605 ;
  assign n13609 = n3636 ^ n1967 ;
  assign n13631 = n441 ^ n137 ;
  assign n13632 = n13631 ^ n677 ;
  assign n13630 = n831 ^ n436 ;
  assign n13633 = n13632 ^ n13630 ;
  assign n13627 = n805 ^ n398 ;
  assign n13628 = n13627 ^ n1254 ;
  assign n13629 = n13628 ^ n2445 ;
  assign n13634 = n13633 ^ n13629 ;
  assign n13635 = n13634 ^ n6316 ;
  assign n13624 = n2082 ^ n917 ;
  assign n13622 = n542 ^ n357 ;
  assign n13623 = n13622 ^ n1915 ;
  assign n13625 = n13624 ^ n13623 ;
  assign n13619 = n657 ^ n237 ;
  assign n13620 = n13619 ^ n1650 ;
  assign n13617 = n800 ^ n507 ;
  assign n13618 = n13617 ^ n2766 ;
  assign n13621 = n13620 ^ n13618 ;
  assign n13626 = n13625 ^ n13621 ;
  assign n13636 = n13635 ^ n13626 ;
  assign n13613 = n2363 ^ n470 ;
  assign n13614 = n13613 ^ n1384 ;
  assign n13610 = n2454 ^ n504 ;
  assign n13611 = n13610 ^ n744 ;
  assign n13612 = n13611 ^ n2320 ;
  assign n13615 = n13614 ^ n13612 ;
  assign n13616 = n13615 ^ n2698 ;
  assign n13637 = n13636 ^ n13616 ;
  assign n13638 = ~n13609 & ~n13637 ;
  assign n13607 = n19031 ^ n8143 ;
  assign n13608 = n13607 ^ n8134 ;
  assign n13639 = n13638 ^ n13608 ;
  assign n13661 = n1179 ^ n478 ;
  assign n13662 = n13661 ^ n999 ;
  assign n13663 = n13662 ^ n1987 ;
  assign n13660 = n3673 ^ n820 ;
  assign n13664 = n13663 ^ n13660 ;
  assign n13665 = n13664 ^ n4961 ;
  assign n13658 = n2807 ^ n1418 ;
  assign n13657 = n1376 ^ n1300 ;
  assign n13659 = n13658 ^ n13657 ;
  assign n13666 = n13665 ^ n13659 ;
  assign n13653 = n1252 ^ n1201 ;
  assign n13652 = n4912 ^ n857 ;
  assign n13654 = n13653 ^ n13652 ;
  assign n13655 = n13654 ^ n4218 ;
  assign n13649 = n3641 ^ n948 ;
  assign n13648 = n2631 ^ n645 ;
  assign n13650 = n13649 ^ n13648 ;
  assign n13646 = n2599 ^ n992 ;
  assign n13647 = n13646 ^ n1175 ;
  assign n13651 = n13650 ^ n13647 ;
  assign n13656 = n13655 ^ n13651 ;
  assign n13667 = n13666 ^ n13656 ;
  assign n13643 = n958 ^ n513 ;
  assign n13642 = n950 ^ n179 ;
  assign n13644 = n13643 ^ n13642 ;
  assign n13641 = n3203 ^ n1577 ;
  assign n13645 = n13644 ^ n13641 ;
  assign n13668 = n13667 ^ n13645 ;
  assign n13027 = n470 ^ n263 ;
  assign n13028 = n13027 ^ n2117 ;
  assign n13025 = n927 ^ n801 ;
  assign n13026 = n13025 ^ n357 ;
  assign n13029 = n13028 ^ n13026 ;
  assign n13023 = n4827 ^ n2297 ;
  assign n13022 = n2019 ^ n1284 ;
  assign n13024 = n13023 ^ n13022 ;
  assign n13030 = n13029 ^ n13024 ;
  assign n13640 = n13030 ^ n602 ;
  assign n13669 = n13668 ^ n13640 ;
  assign n13670 = ~n4131 & ~n13669 ;
  assign n13671 = n13670 ^ n13608 ;
  assign n13672 = n13639 & n13671 ;
  assign n13673 = n13672 ^ n13608 ;
  assign n13686 = n12253 ^ n3805 ;
  assign n13676 = n12361 ^ n12333 ;
  assign n13680 = n13676 ^ n3807 ;
  assign n13681 = n13680 ^ n13676 ;
  assign n13677 = n13676 ^ n12251 ;
  assign n13682 = n13677 ^ n13676 ;
  assign n13683 = ~n13681 & ~n13682 ;
  assign n13684 = n13683 ^ n13676 ;
  assign n13685 = ~x31 & ~n13684 ;
  assign n13687 = n13686 ^ n13685 ;
  assign n13678 = n13677 ^ n12253 ;
  assign n13679 = ~n3967 & n13678 ;
  assign n13688 = n13687 ^ n13679 ;
  assign n13675 = ~n61 & ~n12253 ;
  assign n13689 = n13688 ^ n13675 ;
  assign n13674 = ~n12331 & n22543 ;
  assign n13690 = n13689 ^ n13674 ;
  assign n13691 = ~n13673 & ~n13690 ;
  assign n13692 = ~n13510 & ~n13691 ;
  assign n13693 = ~n13606 & ~n13692 ;
  assign n13694 = n13690 ^ n13673 ;
  assign n13695 = n13694 ^ n13691 ;
  assign n13696 = n13510 & n13695 ;
  assign n13697 = n13693 & ~n13696 ;
  assign n13698 = n13697 ^ n13696 ;
  assign n13699 = n13698 ^ n13565 ;
  assign n13700 = ~n13568 & n13699 ;
  assign n13566 = n13565 ^ n13531 ;
  assign n13701 = n13700 ^ n13566 ;
  assign n13702 = ~n13544 & n13701 ;
  assign n13703 = n13702 ^ n13543 ;
  assign n13705 = n13704 ^ n13703 ;
  assign n13706 = n13703 ^ n13513 ;
  assign n13707 = n13706 ^ n13398 ;
  assign n13708 = n13530 ^ n13513 ;
  assign n13711 = ~n13707 & n13708 ;
  assign n13712 = n13711 ^ n13398 ;
  assign n13713 = ~n13705 & n13712 ;
  assign n13714 = n13713 ^ n13703 ;
  assign n13715 = n13714 ^ n13457 ;
  assign n13716 = n13460 & n13715 ;
  assign n13717 = n13716 ^ n13457 ;
  assign n13720 = n13719 ^ n13717 ;
  assign n12608 = n12607 ^ n12214 ;
  assign n13727 = ~n4435 & n12608 ;
  assign n13725 = ~n4434 & ~n12214 ;
  assign n13722 = n4600 & n12222 ;
  assign n13721 = n12380 & n20603 ;
  assign n13723 = n13722 ^ n13721 ;
  assign n13724 = n13723 ^ x26 ;
  assign n13726 = n13725 ^ n13724 ;
  assign n13728 = n13727 ^ n13726 ;
  assign n13729 = n13728 ^ n13717 ;
  assign n13730 = n13720 & n13729 ;
  assign n13718 = n13717 ^ n13443 ;
  assign n13731 = n13730 ^ n13718 ;
  assign n13732 = ~n13444 & ~n13731 ;
  assign n13733 = n13732 ^ n13443 ;
  assign n13735 = n13734 ^ n13733 ;
  assign n13762 = n13750 ^ n13735 ;
  assign n13843 = n4655 & ~n12210 ;
  assign n13842 = n4651 & ~n12214 ;
  assign n13844 = n13843 ^ n13842 ;
  assign n13845 = n13844 ^ x23 ;
  assign n13841 = n4656 & n12737 ;
  assign n13846 = n13845 ^ n13841 ;
  assign n13840 = ~n40 & ~n12400 ;
  assign n13847 = n13846 ^ n13840 ;
  assign n13791 = n3837 & n12235 ;
  assign n13789 = n3985 & n12229 ;
  assign n13783 = n12228 ^ n5065 ;
  assign n13784 = n13783 ^ n12228 ;
  assign n13785 = ~n12805 & n13784 ;
  assign n13786 = n13785 ^ n12228 ;
  assign n13787 = n3833 & ~n13786 ;
  assign n13776 = ~n13514 & n13708 ;
  assign n13775 = n13703 ^ n13398 ;
  assign n13777 = n13776 ^ n13775 ;
  assign n13778 = n13777 ^ x29 ;
  assign n13788 = n13787 ^ n13778 ;
  assign n13790 = n13789 ^ n13788 ;
  assign n13792 = n13791 ^ n13790 ;
  assign n13797 = ~x25 & n12554 ;
  assign n12555 = n12554 ^ n12380 ;
  assign n13800 = n13797 ^ n12555 ;
  assign n13801 = n99 & n13800 ;
  assign n13794 = n4600 & n12376 ;
  assign n13793 = ~n12382 & n20603 ;
  assign n13795 = n13794 ^ n13793 ;
  assign n13796 = n13795 ^ x26 ;
  assign n13798 = n13797 ^ n12380 ;
  assign n13799 = n13796 & ~n13798 ;
  assign n13802 = n13801 ^ n13799 ;
  assign n13803 = n13795 ^ n97 ;
  assign n13804 = ~n13802 & ~n13803 ;
  assign n13805 = n13804 ^ n13777 ;
  assign n13806 = n13792 & n13805 ;
  assign n13807 = n13806 ^ n13804 ;
  assign n12452 = n12389 ^ n12222 ;
  assign n13770 = n12452 ^ n12380 ;
  assign n13771 = ~n4435 & n13770 ;
  assign n13768 = ~n4434 & n12222 ;
  assign n13765 = n4600 & n12380 ;
  assign n13764 = n12376 & n20603 ;
  assign n13766 = n13765 ^ n13764 ;
  assign n13767 = n13766 ^ x26 ;
  assign n13769 = n13768 ^ n13767 ;
  assign n13772 = n13771 ^ n13769 ;
  assign n13763 = n13714 ^ n13460 ;
  assign n13773 = n13772 ^ n13763 ;
  assign n13839 = n13807 ^ n13773 ;
  assign n13848 = n13847 ^ n13839 ;
  assign n13856 = ~n40 & ~n12214 ;
  assign n13854 = n4656 & n12667 ;
  assign n13851 = n4655 & ~n12400 ;
  assign n13850 = n4651 & n12222 ;
  assign n13852 = n13851 ^ n13850 ;
  assign n13853 = n13852 ^ x23 ;
  assign n13855 = n13854 ^ n13853 ;
  assign n13857 = n13856 ^ n13855 ;
  assign n13849 = n13804 ^ n13792 ;
  assign n13858 = n13857 ^ n13849 ;
  assign n13866 = ~n4435 & n12928 ;
  assign n13864 = ~n4434 & n12376 ;
  assign n13861 = n4600 & ~n12382 ;
  assign n13860 = ~n12228 & n20603 ;
  assign n13862 = n13861 ^ n13860 ;
  assign n13863 = n13862 ^ x26 ;
  assign n13865 = n13864 ^ n13863 ;
  assign n13867 = n13866 ^ n13865 ;
  assign n13916 = n13867 ^ n13849 ;
  assign n13859 = n13701 ^ n13543 ;
  assign n13868 = n13867 ^ n13859 ;
  assign n13880 = n3837 & n12248 ;
  assign n13878 = n3985 & ~n12239 ;
  assign n13871 = n12235 ^ x29 ;
  assign n13872 = n13871 ^ x28 ;
  assign n13873 = n13872 ^ n12235 ;
  assign n13874 = ~n13319 & n13873 ;
  assign n13875 = n13874 ^ n12235 ;
  assign n13876 = n3833 & n13875 ;
  assign n13877 = n13876 ^ x29 ;
  assign n13879 = n13878 ^ n13877 ;
  assign n13881 = n13880 ^ n13879 ;
  assign n13913 = n13881 ^ n13867 ;
  assign n13869 = n13698 ^ n13568 ;
  assign n13882 = n13881 ^ n13869 ;
  assign n13893 = n13696 ^ n13692 ;
  assign n13894 = n13893 ^ n13606 ;
  assign n13884 = n12362 ^ n12334 ;
  assign n13885 = n13884 ^ n12339 ;
  assign n13889 = n5280 & ~n13885 ;
  assign n13888 = n3807 & n12339 ;
  assign n13890 = n13889 ^ n13888 ;
  assign n13886 = n13885 ^ n12253 ;
  assign n13887 = ~n13886 & n22543 ;
  assign n13891 = n13890 ^ n13887 ;
  assign n13883 = ~n3850 & ~n12251 ;
  assign n13892 = n13891 ^ n13883 ;
  assign n13895 = n13894 ^ n13892 ;
  assign n13900 = ~x28 & ~n13339 ;
  assign n13903 = n13900 ^ n13343 ;
  assign n13904 = n4368 & n13903 ;
  assign n13897 = n3985 & n12248 ;
  assign n13896 = n3837 & ~n12249 ;
  assign n13898 = n13897 ^ n13896 ;
  assign n13899 = n13898 ^ x29 ;
  assign n13901 = n13900 ^ n12239 ;
  assign n13902 = n13899 & n13901 ;
  assign n13905 = n13904 ^ n13902 ;
  assign n13906 = n13898 ^ n3978 ;
  assign n13907 = ~n13905 & ~n13906 ;
  assign n13908 = n13907 ^ n13892 ;
  assign n13909 = n13895 & n13908 ;
  assign n13910 = n13909 ^ n13894 ;
  assign n13911 = n13910 ^ n13881 ;
  assign n13912 = ~n13882 & n13911 ;
  assign n13914 = n13913 ^ n13912 ;
  assign n13915 = ~n13868 & n13914 ;
  assign n13917 = n13916 ^ n13915 ;
  assign n13918 = n13858 & ~n13917 ;
  assign n13919 = n13918 ^ n13857 ;
  assign n13920 = n13919 ^ n13847 ;
  assign n13921 = ~n13848 & n13920 ;
  assign n13922 = n13921 ^ n13847 ;
  assign n13817 = n4655 & ~n12405 ;
  assign n13816 = n4651 & ~n12400 ;
  assign n13818 = n13817 ^ n13816 ;
  assign n13819 = n13818 ^ x23 ;
  assign n13815 = n4656 & n12715 ;
  assign n13820 = n13819 ^ n13815 ;
  assign n13814 = ~n40 & ~n12210 ;
  assign n13821 = n13820 ^ n13814 ;
  assign n13774 = n13728 ^ n13720 ;
  assign n13808 = n13807 ^ n13774 ;
  assign n13809 = n13808 ^ n13772 ;
  assign n13810 = n13809 ^ n13774 ;
  assign n13811 = ~n13773 & ~n13810 ;
  assign n13812 = n13811 ^ n13808 ;
  assign n13838 = n13821 ^ n13812 ;
  assign n13923 = n13922 ^ n13838 ;
  assign n13933 = n5426 & ~n12209 ;
  assign n13931 = n12419 & n13433 ;
  assign n13924 = n12204 ^ x20 ;
  assign n13925 = n13924 ^ x19 ;
  assign n13926 = n13925 ^ n12204 ;
  assign n13927 = ~n13415 & n13926 ;
  assign n13928 = n13927 ^ n12204 ;
  assign n13929 = n5215 & ~n13928 ;
  assign n13930 = n13929 ^ x20 ;
  assign n13932 = n13931 ^ n13930 ;
  assign n13934 = n13933 ^ n13932 ;
  assign n13935 = n13934 ^ n13922 ;
  assign n13936 = ~n13923 & n13935 ;
  assign n13937 = n13936 ^ n13922 ;
  assign n13829 = n5426 & ~n12204 ;
  assign n13828 = ~n12209 & n13433 ;
  assign n13830 = n13829 ^ n13828 ;
  assign n13831 = n13830 ^ x20 ;
  assign n13827 = n5215 & ~n12435 ;
  assign n13832 = n13831 ^ n13827 ;
  assign n13833 = n13832 ^ n13831 ;
  assign n13834 = n5224 & n12432 ;
  assign n13835 = n13833 & n13834 ;
  assign n13836 = n13835 ^ n13832 ;
  assign n13813 = n13731 ^ n13442 ;
  assign n13823 = n13813 ^ n13774 ;
  assign n13822 = n13821 ^ n13813 ;
  assign n13824 = n13823 ^ n13822 ;
  assign n13825 = ~n13812 & n13824 ;
  assign n13826 = n13825 ^ n13823 ;
  assign n13837 = n13836 ^ n13826 ;
  assign n13938 = n13937 ^ n13837 ;
  assign n13939 = n13837 ^ n6158 ;
  assign n13940 = ~n13938 & n13939 ;
  assign n13941 = n13940 ^ n13937 ;
  assign n13942 = ~n13762 & ~n13941 ;
  assign n13756 = n13426 ^ n13414 ;
  assign n13751 = n13750 ^ n13733 ;
  assign n13752 = n13735 & n13751 ;
  assign n13753 = n13752 ^ n13750 ;
  assign n13754 = n13753 ^ n8619 ;
  assign n13434 = n12435 & n13433 ;
  assign n13755 = n13754 ^ n13434 ;
  assign n13761 = n13756 ^ n13755 ;
  assign n13943 = n13942 ^ n13761 ;
  assign n20458 = n13836 ^ n13813 ;
  assign n20459 = ~n13826 & ~n20458 ;
  assign n20460 = n20459 ^ n13813 ;
  assign n20461 = n20460 ^ n13761 ;
  assign n13944 = n13934 ^ n13923 ;
  assign n14145 = n6143 & ~n12435 ;
  assign n14143 = ~n12204 & n20437 ;
  assign n14140 = ~n12431 & ~n12435 ;
  assign n14141 = n6163 & ~n14140 ;
  assign n14139 = n6141 ^ x17 ;
  assign n14142 = n14141 ^ n14139 ;
  assign n14144 = n14143 ^ n14142 ;
  assign n14146 = n14145 ^ n14144 ;
  assign n14122 = n13917 ^ n13857 ;
  assign n13959 = n4655 & ~n12214 ;
  assign n13958 = n4651 & n12380 ;
  assign n13960 = n13959 ^ n13958 ;
  assign n13961 = n13960 ^ x23 ;
  assign n13957 = n4656 & n12608 ;
  assign n13962 = n13961 ^ n13957 ;
  assign n13956 = ~n40 & n12222 ;
  assign n13963 = n13962 ^ n13956 ;
  assign n13955 = n13914 ^ n13859 ;
  assign n13964 = n13963 ^ n13955 ;
  assign n13968 = n13910 ^ n13882 ;
  assign n14118 = n13968 ^ n13955 ;
  assign n13972 = n12229 & n20603 ;
  assign n13969 = n13968 ^ x26 ;
  assign n13967 = n4600 & ~n12228 ;
  assign n13970 = n13969 ^ n13967 ;
  assign n13966 = ~n4434 & ~n12382 ;
  assign n13971 = n13970 ^ n13966 ;
  assign n13973 = n13972 ^ n13971 ;
  assign n13965 = ~n4435 & n13445 ;
  assign n13974 = n13973 ^ n13965 ;
  assign n13779 = n12805 ^ n12228 ;
  assign n13982 = ~n4435 & n13779 ;
  assign n13980 = ~n4434 & ~n12228 ;
  assign n13977 = n4600 & n12229 ;
  assign n13976 = n12235 & n20603 ;
  assign n13978 = n13977 ^ n13976 ;
  assign n13979 = n13978 ^ x26 ;
  assign n13981 = n13980 ^ n13979 ;
  assign n13983 = n13982 ^ n13981 ;
  assign n13975 = n13908 ^ n13894 ;
  assign n13984 = n13983 ^ n13975 ;
  assign n13997 = n13673 ^ n13510 ;
  assign n13998 = n13997 ^ n13690 ;
  assign n14112 = n13998 ^ n13975 ;
  assign n13995 = n3837 & n12339 ;
  assign n13993 = n3985 & ~n12249 ;
  assign n13986 = n12248 ^ x29 ;
  assign n13987 = n13986 ^ x28 ;
  assign n13988 = n13987 ^ n12248 ;
  assign n13989 = ~n13518 & n13988 ;
  assign n13990 = n13989 ^ n12248 ;
  assign n13991 = n3833 & n13990 ;
  assign n13992 = n13991 ^ x29 ;
  assign n13994 = n13993 ^ n13992 ;
  assign n13996 = n13995 ^ n13994 ;
  assign n13999 = n13998 ^ n13996 ;
  assign n14010 = n4511 ^ n355 ;
  assign n14008 = n1837 ^ n1239 ;
  assign n14009 = n14008 ^ n2295 ;
  assign n14011 = n14010 ^ n14009 ;
  assign n14012 = n14011 ^ n1019 ;
  assign n14004 = n13481 ^ n195 ;
  assign n14005 = n14004 ^ n2204 ;
  assign n14002 = n12840 ^ n1968 ;
  assign n14001 = n4156 ^ n1303 ;
  assign n14003 = n14002 ^ n14001 ;
  assign n14006 = n14005 ^ n14003 ;
  assign n14007 = n14006 ^ n1101 ;
  assign n14013 = n14012 ^ n14007 ;
  assign n14014 = n14013 ^ n2498 ;
  assign n14015 = ~n2655 & ~n14014 ;
  assign n14019 = n12358 ^ n12323 ;
  assign n14020 = n14019 ^ n12257 ;
  assign n14022 = n14020 ^ n12258 ;
  assign n14021 = n14020 ^ n12264 ;
  assign n14023 = n14022 ^ n14021 ;
  assign n14026 = x30 & ~n14023 ;
  assign n14027 = n14026 ^ n14022 ;
  assign n14028 = ~n3518 & n14027 ;
  assign n14029 = n14028 ^ n14020 ;
  assign n14030 = x31 & ~n14029 ;
  assign n14017 = n3807 & n12257 ;
  assign n14016 = ~n3805 & ~n12258 ;
  assign n14018 = n14017 ^ n14016 ;
  assign n14031 = n14030 ^ n14018 ;
  assign n14033 = n10332 ^ x5 ;
  assign n14032 = ~x2 & ~n11138 ;
  assign n14034 = n14033 ^ n14032 ;
  assign n14053 = n12876 ^ n4922 ;
  assign n14054 = n14053 ^ n3918 ;
  assign n14055 = n14054 ^ n3146 ;
  assign n12528 = n277 ^ n261 ;
  assign n14049 = n12528 ^ n2185 ;
  assign n14050 = n14049 ^ n4749 ;
  assign n14051 = n14050 ^ n1059 ;
  assign n14046 = n1354 ^ n444 ;
  assign n14045 = n2383 ^ n951 ;
  assign n14047 = n14046 ^ n14045 ;
  assign n14044 = n3701 ^ n508 ;
  assign n14048 = n14047 ^ n14044 ;
  assign n14052 = n14051 ^ n14048 ;
  assign n14056 = n14055 ^ n14052 ;
  assign n14040 = n1307 ^ n1129 ;
  assign n14041 = n14040 ^ n818 ;
  assign n14042 = n14041 ^ n13574 ;
  assign n14037 = n4252 ^ n725 ;
  assign n14038 = n14037 ^ n2778 ;
  assign n14035 = n12486 ^ n1329 ;
  assign n14036 = n14035 ^ n3783 ;
  assign n14039 = n14038 ^ n14036 ;
  assign n14043 = n14042 ^ n14039 ;
  assign n14057 = n14056 ^ n14043 ;
  assign n14064 = n4256 ^ n755 ;
  assign n14065 = n14064 ^ n4098 ;
  assign n14066 = n14065 ^ n6833 ;
  assign n14067 = n14066 ^ n4024 ;
  assign n14059 = n750 ^ n468 ;
  assign n14060 = n14059 ^ n138 ;
  assign n14061 = n14060 ^ n1265 ;
  assign n14058 = n2205 ^ n543 ;
  assign n14062 = n14061 ^ n14058 ;
  assign n14063 = n14062 ^ n6285 ;
  assign n14068 = n14067 ^ n14063 ;
  assign n14069 = n14068 ^ n13488 ;
  assign n14070 = ~n14057 & ~n14069 ;
  assign n14071 = n14070 ^ n14032 ;
  assign n14072 = ~n14034 & ~n14071 ;
  assign n14073 = n14072 ^ n14033 ;
  assign n14074 = n14031 & n14073 ;
  assign n14075 = ~n13670 & ~n14074 ;
  assign n14076 = ~n14015 & ~n14075 ;
  assign n14077 = n14073 ^ n14031 ;
  assign n14078 = n14077 ^ n14074 ;
  assign n14079 = n13670 & n14078 ;
  assign n14080 = n14076 & ~n14079 ;
  assign n14081 = n14080 ^ n14079 ;
  assign n14109 = n14081 ^ n13998 ;
  assign n14000 = n13670 ^ n13639 ;
  assign n14082 = n14081 ^ n14000 ;
  assign n3803 = n3802 ^ n3800 ;
  assign n14098 = n12332 ^ n12253 ;
  assign n14101 = n52 & n14098 ;
  assign n14102 = n14101 ^ n12253 ;
  assign n14103 = n3803 & ~n14102 ;
  assign n14089 = x31 & n12257 ;
  assign n14104 = n14103 ^ n14089 ;
  assign n14086 = n12360 ^ n12324 ;
  assign n14087 = n14086 ^ n12332 ;
  assign n14088 = n14087 ^ n12324 ;
  assign n14090 = n14089 ^ n14088 ;
  assign n14095 = n52 & ~n14088 ;
  assign n14096 = n14095 ^ n3803 ;
  assign n14097 = n14090 & n14096 ;
  assign n14105 = n14104 ^ n14097 ;
  assign n14084 = n3807 & n12253 ;
  assign n14083 = ~n3805 & n12331 ;
  assign n14085 = n14084 ^ n14083 ;
  assign n14106 = n14105 ^ n14085 ;
  assign n14107 = n14106 ^ n14081 ;
  assign n14108 = ~n14082 & n14107 ;
  assign n14110 = n14109 ^ n14108 ;
  assign n14111 = n13999 & n14110 ;
  assign n14113 = n14112 ^ n14111 ;
  assign n14114 = ~n13984 & n14113 ;
  assign n14115 = n14114 ^ n13983 ;
  assign n14116 = n14115 ^ n13968 ;
  assign n14117 = ~n13974 & ~n14116 ;
  assign n14119 = n14118 ^ n14117 ;
  assign n14120 = ~n13964 & ~n14119 ;
  assign n14121 = n14120 ^ n13963 ;
  assign n14123 = n14122 ^ n14121 ;
  assign n14133 = ~n12210 & n13433 ;
  assign n14131 = n5426 & ~n12405 ;
  assign n14124 = n12651 ^ x20 ;
  assign n14125 = n14124 ^ x19 ;
  assign n14126 = n14125 ^ n12651 ;
  assign n14127 = ~n12650 & ~n14126 ;
  assign n14128 = n14127 ^ n12651 ;
  assign n14129 = n5215 & ~n14128 ;
  assign n14130 = n14129 ^ x20 ;
  assign n14132 = n14131 ^ n14130 ;
  assign n14134 = n14133 ^ n14132 ;
  assign n14135 = n14134 ^ n14121 ;
  assign n14136 = ~n14123 & n14135 ;
  assign n14137 = n14136 ^ n14134 ;
  assign n13952 = n5220 & ~n12209 ;
  assign n13948 = n13919 ^ n13848 ;
  assign n13949 = n13948 ^ x20 ;
  assign n13947 = ~n12405 & n13433 ;
  assign n13950 = n13949 ^ n13947 ;
  assign n13946 = n5221 & n13052 ;
  assign n13951 = n13950 ^ n13946 ;
  assign n13953 = n13952 ^ n13951 ;
  assign n13945 = n5426 & n12419 ;
  assign n13954 = n13953 ^ n13945 ;
  assign n14138 = n14137 ^ n13954 ;
  assign n14147 = n14146 ^ n14138 ;
  assign n14157 = n6143 & ~n12204 ;
  assign n14149 = n6141 & ~n12435 ;
  assign n14153 = n12432 & n14149 ;
  assign n14154 = x17 ^ x16 ;
  assign n14155 = n14153 & n14154 ;
  assign n14151 = ~n12209 & n20437 ;
  assign n14150 = n14149 ^ x17 ;
  assign n14152 = n14151 ^ n14150 ;
  assign n14156 = n14155 ^ n14152 ;
  assign n14158 = n14157 ^ n14156 ;
  assign n14148 = n14134 ^ n14123 ;
  assign n14159 = n14158 ^ n14148 ;
  assign n14171 = n14119 ^ n13963 ;
  assign n14394 = n14171 ^ n14148 ;
  assign n14169 = n5426 & ~n12210 ;
  assign n14167 = ~n12400 & n13433 ;
  assign n14160 = n12405 ^ x20 ;
  assign n14161 = n14160 ^ x19 ;
  assign n14162 = n14161 ^ n12405 ;
  assign n14163 = ~n12714 & n14162 ;
  assign n14164 = n14163 ^ n12405 ;
  assign n14165 = n5215 & ~n14164 ;
  assign n14166 = n14165 ^ x20 ;
  assign n14168 = n14167 ^ n14166 ;
  assign n14170 = n14169 ^ n14168 ;
  assign n14172 = n14171 ^ n14170 ;
  assign n14180 = n4651 & n12376 ;
  assign n14176 = ~n40 & n12380 ;
  assign n14175 = n4656 & n13770 ;
  assign n14177 = n14176 ^ n14175 ;
  assign n14178 = n14177 ^ x23 ;
  assign n14174 = n4655 & n12222 ;
  assign n14179 = n14178 ^ n14174 ;
  assign n14181 = n14180 ^ n14179 ;
  assign n14391 = n14181 ^ n14171 ;
  assign n14173 = n14115 ^ n13974 ;
  assign n14182 = n14181 ^ n14173 ;
  assign n14191 = n14113 ^ n13983 ;
  assign n14388 = n14191 ^ n14181 ;
  assign n14186 = n4655 & n12380 ;
  assign n14185 = n4651 & ~n12382 ;
  assign n14187 = n14186 ^ n14185 ;
  assign n14188 = n14187 ^ x23 ;
  assign n14184 = n4656 & n12555 ;
  assign n14189 = n14188 ^ n14184 ;
  assign n14183 = ~n40 & n12376 ;
  assign n14190 = n14189 ^ n14183 ;
  assign n14192 = n14191 ^ n14190 ;
  assign n14207 = n14110 ^ n13996 ;
  assign n14385 = n14207 ^ n14191 ;
  assign n14204 = n3837 & ~n12251 ;
  assign n14202 = n3985 & n12339 ;
  assign n14194 = n13554 ^ n12249 ;
  assign n14195 = n12249 ^ x29 ;
  assign n14196 = n14195 ^ x28 ;
  assign n14197 = n14196 ^ n12249 ;
  assign n14198 = ~n14194 & n14197 ;
  assign n14199 = n14198 ^ n12249 ;
  assign n14200 = n3833 & ~n14199 ;
  assign n14201 = n14200 ^ x29 ;
  assign n14203 = n14202 ^ n14201 ;
  assign n14205 = n14204 ^ n14203 ;
  assign n14193 = n14106 ^ n14082 ;
  assign n14206 = n14205 ^ n14193 ;
  assign n14219 = n12359 ^ n12324 ;
  assign n14223 = n3807 & ~n14219 ;
  assign n14220 = n14219 ^ n14089 ;
  assign n14221 = n14220 ^ n12331 ;
  assign n14222 = n3518 & ~n14221 ;
  assign n14224 = n14223 ^ n14222 ;
  assign n14225 = n14224 ^ n14089 ;
  assign n14214 = n12257 ^ n5280 ;
  assign n14215 = n14214 ^ n12257 ;
  assign n14216 = ~n12258 & n14215 ;
  assign n14217 = n14216 ^ n12257 ;
  assign n14218 = ~n61 & n14217 ;
  assign n14226 = n14225 ^ n14218 ;
  assign n14210 = n14079 ^ n14075 ;
  assign n14211 = n14210 ^ n14015 ;
  assign n14227 = n14226 ^ n14211 ;
  assign n14246 = n12264 ^ n3807 ;
  assign n14232 = ~n61 & ~n12267 ;
  assign n14247 = n14246 ^ n14232 ;
  assign n14242 = n12357 ^ n12322 ;
  assign n14243 = n14242 ^ n12258 ;
  assign n14244 = n14243 ^ n12264 ;
  assign n14245 = n14244 & n22005 ;
  assign n14248 = n14247 ^ n14245 ;
  assign n14233 = n14232 ^ n12264 ;
  assign n14234 = n14233 ^ n3807 ;
  assign n14235 = n14234 ^ n14233 ;
  assign n14236 = n14233 ^ n12258 ;
  assign n14237 = n14236 ^ n14233 ;
  assign n14238 = n14235 & n14237 ;
  assign n14239 = n14238 ^ n14233 ;
  assign n14240 = ~x31 & n14239 ;
  assign n14249 = n14248 ^ n14240 ;
  assign n14231 = ~n61 & n12264 ;
  assign n14250 = n14249 ^ n14231 ;
  assign n14230 = n14070 ^ n14034 ;
  assign n14251 = n14250 ^ n14230 ;
  assign n14260 = n4716 ^ n564 ;
  assign n14261 = n14260 ^ n3407 ;
  assign n14262 = n14261 ^ n3397 ;
  assign n14257 = n13484 ^ n2843 ;
  assign n14255 = n1299 ^ n419 ;
  assign n14256 = n14255 ^ n390 ;
  assign n14258 = n14257 ^ n14256 ;
  assign n14253 = n335 ^ n262 ;
  assign n12513 = n2566 ^ n857 ;
  assign n14252 = n12513 ^ n716 ;
  assign n14254 = n14253 ^ n14252 ;
  assign n14259 = n14258 ^ n14254 ;
  assign n14263 = n14262 ^ n14259 ;
  assign n14264 = n14263 ^ n3709 ;
  assign n14265 = n14264 ^ n652 ;
  assign n14266 = ~n4127 & ~n14265 ;
  assign n14267 = n14266 ^ n14032 ;
  assign n14280 = n1879 ^ n117 ;
  assign n14281 = n14280 ^ n6663 ;
  assign n14282 = n14281 ^ n1562 ;
  assign n14277 = n12837 ^ n928 ;
  assign n14278 = n14277 ^ n3886 ;
  assign n14279 = n14278 ^ n1421 ;
  assign n14283 = n14282 ^ n14279 ;
  assign n14273 = n4763 ^ n1020 ;
  assign n14271 = n476 ^ n114 ;
  assign n14272 = n14271 ^ n1321 ;
  assign n14274 = n14273 ^ n14272 ;
  assign n14269 = n1158 ^ n830 ;
  assign n14268 = n4857 ^ n2988 ;
  assign n14270 = n14269 ^ n14268 ;
  assign n14275 = n14274 ^ n14270 ;
  assign n12638 = n1084 ^ n149 ;
  assign n12637 = n1299 ^ n563 ;
  assign n12639 = n12638 ^ n12637 ;
  assign n14276 = n14275 ^ n12639 ;
  assign n14284 = n14283 ^ n14276 ;
  assign n14285 = ~n14057 & ~n14284 ;
  assign n14299 = n2399 ^ n741 ;
  assign n14298 = n13574 ^ n2025 ;
  assign n14300 = n14299 ^ n14298 ;
  assign n14293 = n414 ^ n211 ;
  assign n14294 = n14293 ^ n814 ;
  assign n14295 = n14294 ^ n3770 ;
  assign n14292 = n6926 ^ n2271 ;
  assign n14296 = n14295 ^ n14292 ;
  assign n14289 = n838 ^ n459 ;
  assign n14290 = n14289 ^ n2221 ;
  assign n14287 = n3297 ^ n1451 ;
  assign n14286 = n2554 ^ n1377 ;
  assign n14288 = n14287 ^ n14286 ;
  assign n14291 = n14290 ^ n14288 ;
  assign n14297 = n14296 ^ n14291 ;
  assign n14301 = n14300 ^ n14297 ;
  assign n14302 = n14301 ^ n12580 ;
  assign n14319 = n2259 ^ n627 ;
  assign n14317 = n4942 ^ n462 ;
  assign n14318 = n14317 ^ n2797 ;
  assign n14320 = n14319 ^ n14318 ;
  assign n14321 = n14320 ^ n2419 ;
  assign n14312 = n4782 ^ n562 ;
  assign n14313 = n14312 ^ n819 ;
  assign n14311 = n2267 ^ n991 ;
  assign n14314 = n14313 ^ n14311 ;
  assign n14309 = n675 ^ n348 ;
  assign n14310 = n14309 ^ n3561 ;
  assign n14315 = n14314 ^ n14310 ;
  assign n14306 = n585 ^ n377 ;
  assign n14307 = n14306 ^ n1032 ;
  assign n14308 = n14307 ^ n2139 ;
  assign n14316 = n14315 ^ n14308 ;
  assign n14322 = n14321 ^ n14316 ;
  assign n14304 = n2155 ^ n468 ;
  assign n14303 = n4973 ^ n598 ;
  assign n14305 = n14304 ^ n14303 ;
  assign n14323 = n14322 ^ n14305 ;
  assign n14324 = ~n14302 & ~n14323 ;
  assign n14336 = ~n3850 & ~n12276 ;
  assign n14335 = n3807 & n12268 ;
  assign n14337 = n14336 ^ n14335 ;
  assign n14325 = ~n61 & n12279 ;
  assign n14326 = n14325 ^ n3518 ;
  assign n14327 = n14326 ^ n14325 ;
  assign n14328 = n12354 ^ n12319 ;
  assign n14329 = n14328 ^ n12268 ;
  assign n14332 = n14327 & ~n14329 ;
  assign n14333 = n14332 ^ n14325 ;
  assign n14334 = x31 & n14333 ;
  assign n14338 = n14337 ^ n14334 ;
  assign n14339 = ~n14324 & n14338 ;
  assign n14340 = ~n14032 & ~n14339 ;
  assign n14341 = ~n14285 & ~n14340 ;
  assign n14342 = n14338 ^ n14324 ;
  assign n14343 = n14342 ^ n14339 ;
  assign n14344 = n14032 & ~n14343 ;
  assign n14345 = n14341 & ~n14344 ;
  assign n14346 = n14345 ^ n14344 ;
  assign n14347 = n14346 ^ n14266 ;
  assign n14348 = ~n14267 & n14347 ;
  assign n14349 = n14348 ^ n14032 ;
  assign n14350 = n14349 ^ n14250 ;
  assign n14351 = n14251 & n14350 ;
  assign n14352 = n14351 ^ n14250 ;
  assign n14368 = n14352 ^ n14226 ;
  assign n14228 = n14073 ^ n13670 ;
  assign n14229 = n14228 ^ n14031 ;
  assign n14353 = n14352 ^ n14229 ;
  assign n14364 = n3837 & n12331 ;
  assign n14362 = n3985 & n12253 ;
  assign n14355 = n12251 ^ x29 ;
  assign n14356 = n14355 ^ x28 ;
  assign n14357 = n14356 ^ n12251 ;
  assign n14358 = ~n13676 & n14357 ;
  assign n14359 = n14358 ^ n12251 ;
  assign n14360 = n3833 & ~n14359 ;
  assign n14361 = n14360 ^ x29 ;
  assign n14363 = n14362 ^ n14361 ;
  assign n14365 = n14364 ^ n14363 ;
  assign n14366 = n14365 ^ n14352 ;
  assign n14367 = n14353 & n14366 ;
  assign n14369 = n14368 ^ n14367 ;
  assign n14370 = n14227 & n14369 ;
  assign n14371 = n14370 ^ n14226 ;
  assign n14208 = n14207 ^ n14205 ;
  assign n14209 = n14208 ^ n14207 ;
  assign n14372 = n14371 ^ n14209 ;
  assign n14373 = ~n14206 & n14372 ;
  assign n14374 = n14373 ^ n14208 ;
  assign n14381 = ~n4435 & ~n12867 ;
  assign n14379 = ~n4434 & n12229 ;
  assign n14376 = n4600 & n12235 ;
  assign n14375 = ~n12239 & n20603 ;
  assign n14377 = n14376 ^ n14375 ;
  assign n14378 = n14377 ^ x26 ;
  assign n14380 = n14379 ^ n14378 ;
  assign n14382 = n14381 ^ n14380 ;
  assign n14383 = n14382 ^ n14207 ;
  assign n14384 = n14374 & n14383 ;
  assign n14386 = n14385 ^ n14384 ;
  assign n14387 = ~n14192 & ~n14386 ;
  assign n14389 = n14388 ^ n14387 ;
  assign n14390 = ~n14182 & ~n14389 ;
  assign n14392 = n14391 ^ n14390 ;
  assign n14393 = n14172 & n14392 ;
  assign n14395 = n14394 ^ n14393 ;
  assign n14396 = n14159 & ~n14395 ;
  assign n14397 = n14396 ^ n14158 ;
  assign n14398 = n14397 ^ n14146 ;
  assign n14399 = ~n14147 & n14398 ;
  assign n14400 = n14399 ^ n14146 ;
  assign n14401 = ~n13944 & n14400 ;
  assign n20438 = ~n12435 & n20437 ;
  assign n20439 = n20438 ^ n20433 ;
  assign n20425 = n14137 ^ n13948 ;
  assign n20426 = n13954 & ~n20425 ;
  assign n20427 = n20426 ^ n14137 ;
  assign n20399 = n14397 ^ n14147 ;
  assign n15056 = n12376 & n13433 ;
  assign n15054 = n5426 & n12380 ;
  assign n15048 = n12222 ^ n5224 ;
  assign n15049 = n15048 ^ n12222 ;
  assign n15050 = n12390 & n15049 ;
  assign n15051 = n15050 ^ n12222 ;
  assign n15052 = n5215 & n15051 ;
  assign n14968 = ~n40 & n12229 ;
  assign n14966 = n4656 & n13779 ;
  assign n14963 = n4655 & ~n12228 ;
  assign n14962 = n4651 & n12235 ;
  assign n14964 = n14963 ^ n14962 ;
  assign n14965 = n14964 ^ x23 ;
  assign n14967 = n14966 ^ n14965 ;
  assign n14969 = n14968 ^ n14967 ;
  assign n14949 = n14365 ^ n14353 ;
  assign n14425 = n3837 & n12257 ;
  assign n14423 = n3985 & n12331 ;
  assign n14416 = n12253 ^ x29 ;
  assign n14417 = n14416 ^ x28 ;
  assign n14418 = n14417 ^ n12253 ;
  assign n14419 = ~n14088 & n14418 ;
  assign n14420 = n14419 ^ n12253 ;
  assign n14421 = n3833 & n14420 ;
  assign n14422 = n14421 ^ x29 ;
  assign n14424 = n14423 ^ n14422 ;
  assign n14426 = n14425 ^ n14424 ;
  assign n14413 = n14349 ^ n14251 ;
  assign n14427 = n14426 ^ n14413 ;
  assign n14447 = n14346 ^ n14267 ;
  assign n14428 = n12356 ^ n12321 ;
  assign n14429 = n14428 ^ n12264 ;
  assign n14431 = n14429 ^ n12267 ;
  assign n14430 = n14429 ^ n12268 ;
  assign n14432 = n14431 ^ n14430 ;
  assign n14435 = x30 & ~n14432 ;
  assign n14436 = n14435 ^ n14431 ;
  assign n14437 = ~n3518 & n14436 ;
  assign n14438 = n14437 ^ n14429 ;
  assign n14448 = n14447 ^ n14438 ;
  assign n14439 = n14438 ^ n14232 ;
  assign n14442 = n14439 ^ n12264 ;
  assign n14443 = n14442 ^ n14439 ;
  assign n14444 = n3518 & n14443 ;
  assign n14445 = n14444 ^ n14439 ;
  assign n14446 = ~x31 & ~n14445 ;
  assign n14449 = n14448 ^ n14446 ;
  assign n14460 = ~n3850 & n12268 ;
  assign n14458 = ~n12276 & n22543 ;
  assign n14455 = n14344 ^ n14340 ;
  assign n14456 = n14455 ^ n14285 ;
  assign n14450 = n12355 ^ n12320 ;
  assign n14452 = n14450 ^ n12267 ;
  assign n14453 = n3518 & n14452 ;
  assign n14451 = n3807 & ~n14450 ;
  assign n14454 = n14453 ^ n14451 ;
  assign n14457 = n14456 ^ n14454 ;
  assign n14459 = n14458 ^ n14457 ;
  assign n14461 = n14460 ^ n14459 ;
  assign n14492 = n4234 ^ n413 ;
  assign n14493 = n14492 ^ n896 ;
  assign n14490 = n1424 ^ n336 ;
  assign n14491 = n14490 ^ n868 ;
  assign n14494 = n14493 ^ n14491 ;
  assign n14487 = n2894 ^ n659 ;
  assign n14488 = n14487 ^ n3377 ;
  assign n14489 = n14488 ^ n3687 ;
  assign n14495 = n14494 ^ n14489 ;
  assign n14483 = n13661 ^ n2242 ;
  assign n14482 = n3895 ^ n1565 ;
  assign n14484 = n14483 ^ n14482 ;
  assign n14485 = n14484 ^ n13491 ;
  assign n14486 = n14485 ^ n2826 ;
  assign n14496 = n14495 ^ n14486 ;
  assign n14497 = n14496 ^ n1749 ;
  assign n14498 = ~n5360 & ~n14497 ;
  assign n14465 = n12353 ^ n12318 ;
  assign n14475 = n14465 ^ n12276 ;
  assign n14478 = n14475 ^ n12279 ;
  assign n14479 = n3967 & n14478 ;
  assign n14474 = n14325 ^ n3807 ;
  assign n14476 = n14475 ^ n14474 ;
  assign n14464 = ~n61 & ~n12283 ;
  assign n14477 = n14476 ^ n14464 ;
  assign n14480 = n14479 ^ n14477 ;
  assign n14466 = n14465 ^ n14464 ;
  assign n14467 = n14466 ^ n3807 ;
  assign n14468 = n14467 ^ n14466 ;
  assign n14469 = n14466 ^ n12276 ;
  assign n14470 = n14469 ^ n14466 ;
  assign n14471 = ~n14468 & n14470 ;
  assign n14472 = n14471 ^ n14466 ;
  assign n14473 = ~x31 & n14472 ;
  assign n14481 = n14480 ^ n14473 ;
  assign n14499 = n14498 ^ n14481 ;
  assign n14514 = n12352 ^ n12317 ;
  assign n14528 = n14514 ^ n12279 ;
  assign n14529 = n14528 ^ n12283 ;
  assign n14530 = n3967 & n14529 ;
  assign n14524 = n12279 ^ n3807 ;
  assign n14525 = n14524 ^ n14464 ;
  assign n14526 = n14525 ^ n14514 ;
  assign n14515 = ~n61 & ~n12284 ;
  assign n14527 = n14526 ^ n14515 ;
  assign n14531 = n14530 ^ n14527 ;
  assign n14516 = n14515 ^ n14514 ;
  assign n14517 = n14516 ^ n3807 ;
  assign n14518 = n14517 ^ n14516 ;
  assign n14519 = n14516 ^ n12279 ;
  assign n14520 = n14519 ^ n14516 ;
  assign n14521 = ~n14518 & ~n14520 ;
  assign n14522 = n14521 ^ n14516 ;
  assign n14523 = ~x31 & n14522 ;
  assign n14532 = n14531 ^ n14523 ;
  assign n14510 = n6323 ^ n3793 ;
  assign n14505 = n2510 ^ n501 ;
  assign n14506 = n14505 ^ n1239 ;
  assign n14504 = n948 ^ n649 ;
  assign n14507 = n14506 ^ n14504 ;
  assign n14503 = n12504 ^ n2437 ;
  assign n14508 = n14507 ^ n14503 ;
  assign n14500 = n4011 ^ n3097 ;
  assign n14501 = n14500 ^ n3407 ;
  assign n14502 = n14501 ^ n2947 ;
  assign n14509 = n14508 ^ n14502 ;
  assign n14511 = n14510 ^ n14509 ;
  assign n14512 = ~n1413 & ~n14511 ;
  assign n14513 = ~n1539 & n14512 ;
  assign n14533 = n14532 ^ n14513 ;
  assign n14547 = n12351 ^ n12316 ;
  assign n14548 = n14547 ^ n12283 ;
  assign n14550 = n14548 ^ n12284 ;
  assign n14549 = n14548 ^ n12285 ;
  assign n14551 = n14550 ^ n14549 ;
  assign n14554 = x30 & n14551 ;
  assign n14555 = n14554 ^ n14550 ;
  assign n14556 = ~n3518 & ~n14555 ;
  assign n14557 = n14556 ^ n14548 ;
  assign n14558 = n14557 ^ n14515 ;
  assign n14561 = n14558 ^ n12283 ;
  assign n14562 = n14561 ^ n14558 ;
  assign n14563 = n3518 & ~n14562 ;
  assign n14564 = n14563 ^ n14558 ;
  assign n14565 = ~x31 & n14564 ;
  assign n14566 = n14565 ^ n14557 ;
  assign n14540 = n4738 ^ n420 ;
  assign n14539 = n3670 ^ n735 ;
  assign n14541 = n14540 ^ n14539 ;
  assign n14537 = n2801 ^ n2349 ;
  assign n14536 = n12584 ^ n1495 ;
  assign n14538 = n14537 ^ n14536 ;
  assign n14542 = n14541 ^ n14538 ;
  assign n14534 = n4770 ^ n2262 ;
  assign n14535 = n14534 ^ n2644 ;
  assign n14543 = n14542 ^ n14535 ;
  assign n14544 = n14543 ^ n3052 ;
  assign n14545 = n14544 ^ n2395 ;
  assign n14546 = ~n14323 & ~n14545 ;
  assign n14567 = n14566 ^ n14546 ;
  assign n14594 = ~n61 & n12313 ;
  assign n14595 = x31 & n14594 ;
  assign n14593 = ~n3850 & ~n12285 ;
  assign n14596 = n14595 ^ n14593 ;
  assign n14583 = n12350 ^ n12315 ;
  assign n14588 = n12284 ^ x31 ;
  assign n14589 = n14588 ^ n12284 ;
  assign n14590 = ~n14583 & n14589 ;
  assign n14591 = n14590 ^ n12284 ;
  assign n14592 = n3518 & ~n14591 ;
  assign n14597 = n14596 ^ n14592 ;
  assign n14576 = n5679 ^ n1077 ;
  assign n14577 = n14576 ^ n721 ;
  assign n14578 = n14577 ^ n2603 ;
  assign n14579 = n14578 ^ n4299 ;
  assign n14573 = n3774 ^ n1139 ;
  assign n14572 = n1158 ^ n935 ;
  assign n14574 = n14573 ^ n14572 ;
  assign n14569 = n1085 ^ n527 ;
  assign n14570 = n14569 ^ n1239 ;
  assign n14568 = n2262 ^ n1726 ;
  assign n14571 = n14570 ^ n14568 ;
  assign n14575 = n14574 ^ n14571 ;
  assign n14580 = n14579 ^ n14575 ;
  assign n14581 = n14580 ^ n810 ;
  assign n14582 = ~n4071 & ~n14581 ;
  assign n14598 = n14597 ^ n14582 ;
  assign n14666 = n12289 & n22543 ;
  assign n14651 = n12349 ^ n12314 ;
  assign n14652 = n14651 ^ n12285 ;
  assign n14662 = n14652 ^ n12313 ;
  assign n14663 = n3967 & n14662 ;
  assign n14653 = n14652 ^ n14651 ;
  assign n14654 = n14594 ^ n3807 ;
  assign n14655 = n14654 ^ n14652 ;
  assign n14656 = n14655 ^ n14594 ;
  assign n14657 = n14656 ^ n14651 ;
  assign n14658 = n14653 & n14657 ;
  assign n14659 = n14658 ^ n14651 ;
  assign n14660 = ~x31 & n14659 ;
  assign n14661 = n14660 ^ n14655 ;
  assign n14664 = n14663 ^ n14661 ;
  assign n14667 = n14666 ^ n14664 ;
  assign n14615 = ~n68 & n88 ;
  assign n14614 = n64 & n154 ;
  assign n14616 = n14615 ^ n14614 ;
  assign n14617 = x26 & n14616 ;
  assign n14632 = n101 ^ n86 ;
  assign n14633 = ~n68 & ~n14632 ;
  assign n14634 = ~n14617 & n14633 ;
  assign n14626 = n3773 ^ n594 ;
  assign n14627 = n14626 ^ n948 ;
  assign n14624 = n3884 ^ n1021 ;
  assign n14625 = n14624 ^ n3166 ;
  assign n14628 = n14627 ^ n14625 ;
  assign n14621 = n5581 ^ n2868 ;
  assign n14622 = n14621 ^ n3690 ;
  assign n14619 = n1009 ^ n126 ;
  assign n14618 = n1903 ^ n564 ;
  assign n14620 = n14619 ^ n14618 ;
  assign n14623 = n14622 ^ n14620 ;
  assign n14629 = n14628 ^ n14623 ;
  assign n14630 = n14629 ^ n14617 ;
  assign n14635 = n14634 ^ n14630 ;
  assign n14607 = n3677 ^ n248 ;
  assign n14608 = n14607 ^ n596 ;
  assign n14609 = n14608 ^ n2070 ;
  assign n14610 = n14609 ^ n4164 ;
  assign n14611 = n14610 ^ n3093 ;
  assign n14612 = n14611 ^ n13383 ;
  assign n14602 = n3524 ^ n213 ;
  assign n14603 = n14602 ^ n390 ;
  assign n14601 = n2415 ^ n1001 ;
  assign n14604 = n14603 ^ n14601 ;
  assign n14605 = n14604 ^ n6667 ;
  assign n14599 = n2988 ^ n178 ;
  assign n14600 = n14599 ^ n252 ;
  assign n14606 = n14605 ^ n14600 ;
  assign n14613 = n14612 ^ n14606 ;
  assign n14636 = n14635 ^ n14613 ;
  assign n14645 = n4241 ^ n1437 ;
  assign n14644 = n4182 ^ n746 ;
  assign n14646 = n14645 ^ n14644 ;
  assign n14647 = n14646 ^ n6790 ;
  assign n14640 = n4290 ^ n1277 ;
  assign n14641 = n14640 ^ n455 ;
  assign n14638 = n14306 ^ n682 ;
  assign n14639 = n14638 ^ n861 ;
  assign n14642 = n14641 ^ n14639 ;
  assign n14637 = n13384 ^ n2134 ;
  assign n14643 = n14642 ^ n14637 ;
  assign n14648 = n14647 ^ n14643 ;
  assign n14649 = n14648 ^ n1845 ;
  assign n14650 = ~n14636 & ~n14649 ;
  assign n14668 = n14667 ^ n14650 ;
  assign n14711 = n12348 ^ n12304 ;
  assign n14712 = n14711 ^ n12313 ;
  assign n14713 = x31 & n14712 ;
  assign n14710 = n12313 & ~n22005 ;
  assign n14714 = n14713 ^ n14710 ;
  assign n14707 = x31 & n12289 ;
  assign n14715 = n14714 ^ n14707 ;
  assign n14716 = n3518 & ~n14715 ;
  assign n14703 = n12290 ^ x31 ;
  assign n14702 = ~x31 & n12290 ;
  assign n14704 = n14703 ^ n14702 ;
  assign n14705 = n14704 ^ n12289 ;
  assign n14706 = ~n61 & n14705 ;
  assign n14708 = n14707 ^ n14706 ;
  assign n14709 = n14708 ^ n3807 ;
  assign n14717 = n14716 ^ n14709 ;
  assign n14681 = n13616 ^ n2063 ;
  assign n14677 = n1953 ^ n1879 ;
  assign n14676 = n3919 ^ n2965 ;
  assign n14678 = n14677 ^ n14676 ;
  assign n14673 = n1708 ^ n776 ;
  assign n14674 = n14673 ^ n876 ;
  assign n14672 = n556 ^ n526 ;
  assign n14675 = n14674 ^ n14672 ;
  assign n14679 = n14678 ^ n14675 ;
  assign n14670 = n1985 ^ n755 ;
  assign n14669 = n2519 ^ n1056 ;
  assign n14671 = n14670 ^ n14669 ;
  assign n14680 = n14679 ^ n14671 ;
  assign n14682 = n14681 ^ n14680 ;
  assign n14695 = n4946 ^ n572 ;
  assign n14696 = n14695 ^ n1060 ;
  assign n14693 = n917 ^ n94 ;
  assign n14694 = n14693 ^ n507 ;
  assign n14697 = n14696 ^ n14694 ;
  assign n14690 = n1581 ^ n241 ;
  assign n14689 = n1607 ^ n1142 ;
  assign n14691 = n14690 ^ n14689 ;
  assign n14687 = n4181 ^ n4011 ;
  assign n14688 = n14687 ^ n4046 ;
  assign n14692 = n14691 ^ n14688 ;
  assign n14698 = n14697 ^ n14692 ;
  assign n14683 = n1008 ^ n680 ;
  assign n14684 = n14683 ^ n3619 ;
  assign n14685 = n14684 ^ n13359 ;
  assign n14686 = n14685 ^ n2515 ;
  assign n14699 = n14698 ^ n14686 ;
  assign n14700 = n14699 ^ n3913 ;
  assign n14701 = ~n14682 & ~n14700 ;
  assign n14718 = n14717 ^ n14701 ;
  assign n14765 = x30 & ~n12290 ;
  assign n14748 = n12347 ^ n12303 ;
  assign n14749 = n14748 ^ n12289 ;
  assign n14751 = n14749 ^ n12290 ;
  assign n14750 = n14749 ^ n12293 ;
  assign n14752 = n14751 ^ n14750 ;
  assign n14755 = x30 & ~n14752 ;
  assign n14756 = n14755 ^ n14751 ;
  assign n14757 = ~n3518 & n14756 ;
  assign n14758 = n14757 ^ n14749 ;
  assign n14759 = n14758 ^ n12289 ;
  assign n14760 = n14759 ^ n14758 ;
  assign n14766 = n14765 ^ n14760 ;
  assign n14767 = ~n3518 & n14766 ;
  assign n14768 = n14767 ^ n14759 ;
  assign n14769 = ~x31 & ~n14768 ;
  assign n14770 = n14769 ^ n14758 ;
  assign n14731 = n3203 ^ n153 ;
  assign n14732 = n14731 ^ n991 ;
  assign n14729 = n271 ^ n211 ;
  assign n14730 = n14729 ^ n261 ;
  assign n14733 = n14732 ^ n14730 ;
  assign n14734 = n14733 ^ n13602 ;
  assign n14725 = n4242 ^ n832 ;
  assign n14724 = n13375 ^ n2444 ;
  assign n14726 = n14725 ^ n14724 ;
  assign n14722 = n12886 ^ n1719 ;
  assign n14723 = n14722 ^ n875 ;
  assign n14727 = n14726 ^ n14723 ;
  assign n14719 = n533 ^ n197 ;
  assign n14720 = n14719 ^ n750 ;
  assign n14721 = n14720 ^ n1625 ;
  assign n14728 = n14727 ^ n14721 ;
  assign n14735 = n14734 ^ n14728 ;
  assign n14740 = n3690 ^ n622 ;
  assign n14741 = n14740 ^ n386 ;
  assign n14742 = n14741 ^ n1370 ;
  assign n14739 = n5329 ^ n4868 ;
  assign n14743 = n14742 ^ n14739 ;
  assign n14736 = n2054 ^ n845 ;
  assign n14737 = n14736 ^ n1832 ;
  assign n14738 = n14737 ^ n13610 ;
  assign n14744 = n14743 ^ n14738 ;
  assign n14745 = n14744 ^ n2853 ;
  assign n14746 = ~n2225 & ~n14745 ;
  assign n14747 = ~n14735 & n14746 ;
  assign n14771 = n14770 ^ n14747 ;
  assign n12664 = n3807 ^ x31 ;
  assign n14800 = n12664 & ~n14702 ;
  assign n14796 = ~n61 & n12293 ;
  assign n14797 = n14796 ^ n12292 ;
  assign n14798 = ~n14797 & ~n22543 ;
  assign n14799 = n14798 ^ n12292 ;
  assign n14801 = n14800 ^ n14799 ;
  assign n14785 = n12297 ^ n12290 ;
  assign n14786 = n14785 ^ n3518 ;
  assign n14787 = n14786 ^ n14785 ;
  assign n14788 = ~x30 & ~n12293 ;
  assign n14789 = n14788 ^ n14785 ;
  assign n14790 = ~n14787 & n14789 ;
  assign n14791 = n14790 ^ n14785 ;
  assign n14792 = x31 & n14791 ;
  assign n14802 = n14801 ^ n14792 ;
  assign n14779 = n6718 ^ n208 ;
  assign n14780 = n14779 ^ n3184 ;
  assign n14775 = n3036 ^ n637 ;
  assign n14773 = n917 ^ n347 ;
  assign n14774 = n14773 ^ n754 ;
  assign n14776 = n14775 ^ n14774 ;
  assign n14772 = n4001 ^ n2735 ;
  assign n14777 = n14776 ^ n14772 ;
  assign n14778 = n14777 ^ n5655 ;
  assign n14781 = n14780 ^ n14778 ;
  assign n14782 = n3766 ^ n3557 ;
  assign n14783 = ~n14781 & ~n14782 ;
  assign n14784 = ~n4271 & n14783 ;
  assign n14803 = n14802 ^ n14784 ;
  assign n14821 = n3518 & n12292 ;
  assign n14820 = ~n3801 & n12291 ;
  assign n14822 = n14821 ^ n14820 ;
  assign n14833 = n14578 ^ n634 ;
  assign n14834 = n14833 ^ n1078 ;
  assign n14831 = n2163 ^ n596 ;
  assign n14832 = n14831 ^ n735 ;
  assign n14835 = n14834 ^ n14832 ;
  assign n14827 = n813 ^ n465 ;
  assign n14828 = n14827 ^ n142 ;
  assign n14829 = n14828 ^ n1332 ;
  assign n14826 = n4777 ^ n2601 ;
  assign n14830 = n14829 ^ n14826 ;
  assign n14836 = n14835 ^ n14830 ;
  assign n14824 = n13572 ^ n3639 ;
  assign n14823 = n4180 ^ n461 ;
  assign n14825 = n14824 ^ n14823 ;
  assign n14837 = n14836 ^ n14825 ;
  assign n14841 = n14309 ^ n649 ;
  assign n14840 = n355 ^ n211 ;
  assign n14842 = n14841 ^ n14840 ;
  assign n14839 = n5520 ^ n3751 ;
  assign n14843 = n14842 ^ n14839 ;
  assign n14838 = n3309 ^ n3258 ;
  assign n14844 = n14843 ^ n14838 ;
  assign n14845 = n14844 ^ n6819 ;
  assign n14846 = n14845 ^ n2961 ;
  assign n14847 = ~n14837 & ~n14846 ;
  assign n14848 = n5573 ^ n2319 ;
  assign n14849 = n14848 ^ n621 ;
  assign n14811 = n628 ^ n517 ;
  assign n14850 = n14849 ^ n14811 ;
  assign n14851 = n14847 & ~n14850 ;
  assign n14852 = n14822 & ~n14851 ;
  assign n14813 = n4763 ^ n2241 ;
  assign n14812 = n14811 ^ n874 ;
  assign n14814 = n14813 ^ n14812 ;
  assign n14809 = n805 ^ n429 ;
  assign n14807 = n3561 ^ n753 ;
  assign n14808 = n14807 ^ n609 ;
  assign n14810 = n14809 ^ n14808 ;
  assign n14815 = n14814 ^ n14810 ;
  assign n14805 = n2172 ^ n927 ;
  assign n14804 = n3908 ^ n2604 ;
  assign n14806 = n14805 ^ n14804 ;
  assign n14816 = n14815 ^ n14806 ;
  assign n14817 = n14816 ^ n14296 ;
  assign n13017 = n1689 ^ n761 ;
  assign n13018 = n13017 ^ n2493 ;
  assign n13019 = n13018 ^ n12459 ;
  assign n13020 = n13019 ^ n2294 ;
  assign n13013 = n1906 ^ n490 ;
  assign n13014 = n13013 ^ n675 ;
  assign n13012 = n1785 ^ n572 ;
  assign n13015 = n13014 ^ n13012 ;
  assign n13016 = n13015 ^ n1618 ;
  assign n13021 = n13020 ^ n13016 ;
  assign n14818 = n14817 ^ n13021 ;
  assign n14819 = ~n13589 & ~n14818 ;
  assign n14853 = n14852 ^ n14819 ;
  assign n14865 = ~n12292 & n22005 ;
  assign n14866 = n14865 ^ n5280 ;
  assign n14867 = ~n12291 & n14866 ;
  assign n14860 = n22543 ^ n12293 ;
  assign n14868 = n14867 ^ n14860 ;
  assign n14854 = n12294 ^ n12293 ;
  assign n14855 = n12293 ^ n3801 ;
  assign n14856 = n14855 ^ n12293 ;
  assign n14857 = n14854 & ~n14856 ;
  assign n14858 = n14857 ^ n12293 ;
  assign n14859 = ~n3518 & n14858 ;
  assign n14869 = n14868 ^ n14859 ;
  assign n14870 = n14869 ^ n14852 ;
  assign n14871 = ~n14853 & n14870 ;
  assign n14872 = n14871 ^ n14852 ;
  assign n14873 = n14872 ^ n14784 ;
  assign n14874 = n14803 & n14873 ;
  assign n14875 = n14874 ^ n14802 ;
  assign n14876 = n14875 ^ n14770 ;
  assign n14877 = n14771 & n14876 ;
  assign n14878 = n14877 ^ n14770 ;
  assign n14879 = n14878 ^ n14717 ;
  assign n14880 = ~n14718 & ~n14879 ;
  assign n14881 = n14880 ^ n14717 ;
  assign n14882 = n14881 ^ n14667 ;
  assign n14883 = ~n14668 & n14882 ;
  assign n14884 = n14883 ^ n14667 ;
  assign n14885 = n14884 ^ n14597 ;
  assign n14886 = ~n14598 & n14885 ;
  assign n14887 = n14886 ^ n14597 ;
  assign n14888 = n14887 ^ n14566 ;
  assign n14889 = ~n14567 & n14888 ;
  assign n14890 = n14889 ^ n14566 ;
  assign n14891 = n14890 ^ n14532 ;
  assign n14892 = n14533 & ~n14891 ;
  assign n14893 = n14892 ^ n14532 ;
  assign n14894 = n14893 ^ n14481 ;
  assign n14895 = ~n14499 & ~n14894 ;
  assign n14896 = n14895 ^ n14481 ;
  assign n14462 = n14324 ^ n14032 ;
  assign n14463 = n14462 ^ n14338 ;
  assign n14897 = n14896 ^ n14463 ;
  assign n14908 = n3837 & ~n12267 ;
  assign n14906 = n3985 & n12264 ;
  assign n14899 = n12258 ^ x29 ;
  assign n14900 = n14899 ^ x28 ;
  assign n14901 = n14900 ^ n12258 ;
  assign n14902 = ~n14242 & n14901 ;
  assign n14903 = n14902 ^ n12258 ;
  assign n14904 = n3833 & ~n14903 ;
  assign n14905 = n14904 ^ x29 ;
  assign n14907 = n14906 ^ n14905 ;
  assign n14909 = n14908 ^ n14907 ;
  assign n14910 = n14909 ^ n14896 ;
  assign n14911 = ~n14897 & n14910 ;
  assign n14912 = n14911 ^ n14896 ;
  assign n14913 = n14912 ^ n14456 ;
  assign n14914 = n14461 & n14913 ;
  assign n14915 = n14914 ^ n14456 ;
  assign n14916 = n14915 ^ n14447 ;
  assign n14917 = n14449 & ~n14916 ;
  assign n14918 = n14917 ^ n14447 ;
  assign n14919 = n14918 ^ n14426 ;
  assign n14920 = n14427 & ~n14919 ;
  assign n14921 = n14920 ^ n14426 ;
  assign n14950 = n14949 ^ n14921 ;
  assign n14957 = ~n4435 & ~n13519 ;
  assign n14955 = ~n4434 & n12248 ;
  assign n14952 = n4600 & ~n12249 ;
  assign n14951 = n12339 & n20603 ;
  assign n14953 = n14952 ^ n14951 ;
  assign n14954 = n14953 ^ x26 ;
  assign n14956 = n14955 ^ n14954 ;
  assign n14958 = n14957 ^ n14956 ;
  assign n14959 = n14958 ^ n14921 ;
  assign n14960 = n14950 & n14959 ;
  assign n14939 = ~x25 & ~n13339 ;
  assign n14942 = n14939 ^ n13343 ;
  assign n14943 = n99 & n14942 ;
  assign n14936 = n4600 & n12248 ;
  assign n14935 = ~n12249 & n20603 ;
  assign n14937 = n14936 ^ n14935 ;
  assign n14938 = n14937 ^ x26 ;
  assign n14940 = n14939 ^ n12239 ;
  assign n14941 = n14938 & n14940 ;
  assign n14944 = n14943 ^ n14941 ;
  assign n14945 = n14937 ^ n97 ;
  assign n14946 = ~n14944 & ~n14945 ;
  assign n14933 = n3837 & n12253 ;
  assign n14931 = n3985 & ~n12251 ;
  assign n14928 = n14369 ^ n14211 ;
  assign n14929 = n14928 ^ x29 ;
  assign n14922 = n13885 ^ n12339 ;
  assign n14923 = n13885 ^ n5065 ;
  assign n14924 = n14923 ^ n13885 ;
  assign n14925 = ~n14922 & ~n14924 ;
  assign n14926 = n14925 ^ n13885 ;
  assign n14927 = n3833 & ~n14926 ;
  assign n14930 = n14929 ^ n14927 ;
  assign n14932 = n14931 ^ n14930 ;
  assign n14934 = n14933 ^ n14932 ;
  assign n14947 = n14946 ^ n14934 ;
  assign n14948 = n14947 ^ n14921 ;
  assign n14961 = n14960 ^ n14948 ;
  assign n14970 = n14969 ^ n14961 ;
  assign n14411 = ~n12382 & n13433 ;
  assign n14409 = n5426 & n12376 ;
  assign n14402 = n12380 ^ x20 ;
  assign n14403 = n14402 ^ x19 ;
  assign n14404 = n14403 ^ n12380 ;
  assign n14405 = n12554 & n14404 ;
  assign n14406 = n14405 ^ n12380 ;
  assign n14407 = n5215 & n14406 ;
  assign n14408 = n14407 ^ x20 ;
  assign n14410 = n14409 ^ n14408 ;
  assign n14412 = n14411 ^ n14410 ;
  assign n14971 = n14970 ^ n14412 ;
  assign n15028 = n14958 ^ n14950 ;
  assign n15015 = ~x25 & ~n13553 ;
  assign n15018 = n15015 ^ n13554 ;
  assign n15019 = n99 & n15018 ;
  assign n15012 = n4600 & n12339 ;
  assign n15011 = ~n12251 & n20603 ;
  assign n15013 = n15012 ^ n15011 ;
  assign n15014 = n15013 ^ x26 ;
  assign n15016 = n15015 ^ n12249 ;
  assign n15017 = n15014 & n15016 ;
  assign n15020 = n15019 ^ n15017 ;
  assign n15021 = n15013 ^ n97 ;
  assign n15022 = ~n15020 & ~n15021 ;
  assign n14984 = n3837 & ~n12258 ;
  assign n14982 = n3985 & n12257 ;
  assign n14979 = n14915 ^ n14449 ;
  assign n14980 = n14979 ^ x29 ;
  assign n14972 = n14219 ^ n12331 ;
  assign n14974 = n14972 ^ n5065 ;
  assign n14975 = n14974 ^ n14972 ;
  assign n14976 = ~n14219 & ~n14975 ;
  assign n14977 = n14976 ^ n14972 ;
  assign n14978 = n3833 & ~n14977 ;
  assign n14981 = n14980 ^ n14978 ;
  assign n14983 = n14982 ^ n14981 ;
  assign n14985 = n14984 ^ n14983 ;
  assign n14987 = n4600 & ~n12251 ;
  assign n14986 = n12253 & n20603 ;
  assign n14988 = n14987 ^ n14986 ;
  assign n14989 = n14988 ^ n97 ;
  assign n14990 = n14988 ^ x26 ;
  assign n14991 = n14990 ^ n99 ;
  assign n14992 = n14991 ^ x25 ;
  assign n14993 = n14992 ^ n14990 ;
  assign n14994 = n14993 ^ n12339 ;
  assign n14995 = n14994 ^ n13884 ;
  assign n14996 = n14995 ^ n14994 ;
  assign n14997 = n14990 & ~n14996 ;
  assign n14998 = n14997 ^ n14991 ;
  assign n15000 = ~n14993 & ~n14996 ;
  assign n15001 = n15000 ^ n12339 ;
  assign n15002 = ~n14991 & ~n15001 ;
  assign n15003 = ~n14998 & n15002 ;
  assign n15004 = n15003 ^ n15000 ;
  assign n15005 = n15004 ^ n99 ;
  assign n15006 = n15005 ^ n12339 ;
  assign n15007 = ~n14989 & n15006 ;
  assign n15008 = n15007 ^ n14979 ;
  assign n15009 = ~n14985 & ~n15008 ;
  assign n15010 = n15009 ^ n15007 ;
  assign n15023 = n15022 ^ n15010 ;
  assign n15024 = n14918 ^ n14427 ;
  assign n15025 = n15024 ^ n15010 ;
  assign n15026 = ~n15023 & n15025 ;
  assign n15027 = n15026 ^ n15024 ;
  assign n15029 = n15028 ^ n15027 ;
  assign n15033 = n4655 & n12229 ;
  assign n15032 = n4651 & ~n12239 ;
  assign n15034 = n15033 ^ n15032 ;
  assign n15035 = n15034 ^ x23 ;
  assign n15031 = n4656 & ~n12867 ;
  assign n15036 = n15035 ^ n15031 ;
  assign n15030 = ~n40 & n12235 ;
  assign n15037 = n15036 ^ n15030 ;
  assign n15038 = n15037 ^ n14970 ;
  assign n15039 = n15038 ^ n14970 ;
  assign n15040 = n15039 ^ n15027 ;
  assign n15041 = n15029 & ~n15040 ;
  assign n15042 = n15041 ^ n15038 ;
  assign n15043 = ~n14971 & ~n15042 ;
  assign n15044 = n15043 ^ n14970 ;
  assign n15045 = n15044 ^ x20 ;
  assign n15053 = n15052 ^ n15045 ;
  assign n15055 = n15054 ^ n15053 ;
  assign n15057 = n15056 ^ n15055 ;
  assign n15103 = n14969 ^ n14947 ;
  assign n15104 = ~n14961 & ~n15103 ;
  assign n15105 = n15104 ^ n14947 ;
  assign n15097 = n4655 & ~n12382 ;
  assign n15096 = n4651 & n12229 ;
  assign n15098 = n15097 ^ n15096 ;
  assign n15099 = n15098 ^ x23 ;
  assign n15095 = n4656 & n13445 ;
  assign n15100 = n15099 ^ n15095 ;
  assign n15094 = ~n40 & ~n12228 ;
  assign n15101 = n15100 ^ n15094 ;
  assign n15084 = n14946 ^ n14928 ;
  assign n15085 = ~n14934 & ~n15084 ;
  assign n15086 = n15085 ^ n14946 ;
  assign n15081 = ~n4435 & ~n13329 ;
  assign n15079 = ~n4434 & n12235 ;
  assign n15076 = n4600 & ~n12239 ;
  assign n15075 = n12248 & n20603 ;
  assign n15077 = n15076 ^ n15075 ;
  assign n15078 = n15077 ^ x26 ;
  assign n15080 = n15079 ^ n15078 ;
  assign n15082 = n15081 ^ n15080 ;
  assign n15074 = n14371 ^ n14206 ;
  assign n15083 = n15082 ^ n15074 ;
  assign n15093 = n15086 ^ n15083 ;
  assign n15102 = n15101 ^ n15093 ;
  assign n15112 = n15105 ^ n15102 ;
  assign n15106 = n15105 ^ n15101 ;
  assign n15107 = n15102 & ~n15106 ;
  assign n15108 = n15107 ^ n15101 ;
  assign n15090 = n14382 ^ n14374 ;
  assign n15087 = n15086 ^ n15082 ;
  assign n15088 = ~n15083 & ~n15087 ;
  assign n15089 = n15088 ^ n15082 ;
  assign n15091 = n15090 ^ n15089 ;
  assign n15072 = ~n40 & ~n12382 ;
  assign n15070 = n4656 & n12928 ;
  assign n15067 = n4655 & n12376 ;
  assign n15066 = n4651 & ~n12228 ;
  assign n15068 = n15067 ^ n15066 ;
  assign n15069 = n15068 ^ x23 ;
  assign n15071 = n15070 ^ n15069 ;
  assign n15073 = n15072 ^ n15071 ;
  assign n15092 = n15091 ^ n15073 ;
  assign n15109 = n15108 ^ n15092 ;
  assign n15064 = n5426 & n12222 ;
  assign n15062 = n5220 & ~n12214 ;
  assign n15059 = n5221 & n12608 ;
  assign n15058 = n12380 & n13433 ;
  assign n15060 = n15059 ^ n15058 ;
  assign n15061 = n15060 ^ x20 ;
  assign n15063 = n15062 ^ n15061 ;
  assign n15065 = n15064 ^ n15063 ;
  assign n15110 = n15109 ^ n15065 ;
  assign n15113 = n15112 ^ n15110 ;
  assign n15111 = n15110 ^ n15044 ;
  assign n15114 = n15113 ^ n15111 ;
  assign n15115 = n15057 & n15114 ;
  assign n15116 = n15115 ^ n15113 ;
  assign n15144 = ~n12210 & n20437 ;
  assign n15142 = n6163 & ~n12651 ;
  assign n15139 = n6148 & n12419 ;
  assign n15138 = n6143 & ~n12405 ;
  assign n15140 = n15139 ^ n15138 ;
  assign n15141 = n15140 ^ x17 ;
  assign n15143 = n15142 ^ n15141 ;
  assign n15145 = n15144 ^ n15143 ;
  assign n15133 = n12222 & n13433 ;
  assign n15131 = n5426 & ~n12214 ;
  assign n15124 = n12667 ^ x20 ;
  assign n15125 = n15124 ^ x19 ;
  assign n15126 = n15125 ^ n12667 ;
  assign n15127 = ~n12666 & ~n15126 ;
  assign n15128 = n15127 ^ n12667 ;
  assign n15129 = n5215 & n15128 ;
  assign n15130 = n15129 ^ x20 ;
  assign n15132 = n15131 ^ n15130 ;
  assign n15134 = n15133 ^ n15132 ;
  assign n15121 = n15089 ^ n15073 ;
  assign n15122 = n15091 & n15121 ;
  assign n15119 = n14386 ^ n14190 ;
  assign n15120 = n15119 ^ n15089 ;
  assign n15123 = n15122 ^ n15120 ;
  assign n15135 = n15134 ^ n15123 ;
  assign n15136 = n15135 ^ n15108 ;
  assign n15117 = n15108 ^ n15065 ;
  assign n15118 = n15109 & n15117 ;
  assign n15137 = n15136 ^ n15118 ;
  assign n15146 = n15145 ^ n15137 ;
  assign n15156 = n15146 ^ n15110 ;
  assign n15150 = n6148 & ~n12405 ;
  assign n15149 = n6143 & ~n12210 ;
  assign n15151 = n15150 ^ n15149 ;
  assign n15152 = n15151 ^ x17 ;
  assign n15148 = n6163 & n12715 ;
  assign n15153 = n15152 ^ n15148 ;
  assign n15147 = ~n12400 & n20437 ;
  assign n15154 = n15153 ^ n15147 ;
  assign n15155 = n15154 ^ n15146 ;
  assign n15157 = n15156 ^ n15155 ;
  assign n15158 = ~n15116 & n15157 ;
  assign n15159 = n15158 ^ n15156 ;
  assign n15163 = ~n6529 & ~n12204 ;
  assign n15162 = ~n6547 & ~n12209 ;
  assign n15164 = n15163 ^ n15162 ;
  assign n15161 = n6391 & ~n12435 ;
  assign n15165 = n15164 ^ n15161 ;
  assign n15175 = n15165 ^ x14 ;
  assign n15166 = n15165 ^ n15164 ;
  assign n15160 = ~n12432 & ~n12435 ;
  assign n15167 = n15166 ^ n15160 ;
  assign n15172 = x13 & ~n15160 ;
  assign n15173 = n15172 ^ n6537 ;
  assign n15174 = n15167 & n15173 ;
  assign n15176 = n15175 ^ n15174 ;
  assign n20297 = n15176 ^ n15146 ;
  assign n20298 = ~n15159 & ~n20297 ;
  assign n20299 = n20298 ^ n15146 ;
  assign n15190 = ~n12214 & n20437 ;
  assign n15188 = n6143 & ~n12400 ;
  assign n15186 = n15112 ^ n15057 ;
  assign n15179 = n12210 ^ x17 ;
  assign n15180 = n15179 ^ x16 ;
  assign n15181 = n15180 ^ n12210 ;
  assign n15182 = ~n12736 & n15181 ;
  assign n15183 = n15182 ^ n12210 ;
  assign n15184 = n6141 & ~n15183 ;
  assign n15185 = n15184 ^ x17 ;
  assign n15187 = n15186 ^ n15185 ;
  assign n15189 = n15188 ^ n15187 ;
  assign n15191 = n15190 ^ n15189 ;
  assign n15200 = n15042 ^ n14412 ;
  assign n15198 = n12222 & n20437 ;
  assign n15196 = n6163 & n12667 ;
  assign n15193 = n6148 & ~n12400 ;
  assign n15192 = n6143 & ~n12214 ;
  assign n15194 = n15193 ^ n15192 ;
  assign n15195 = n15194 ^ x17 ;
  assign n15197 = n15196 ^ n15195 ;
  assign n15199 = n15198 ^ n15197 ;
  assign n15201 = n15200 ^ n15199 ;
  assign n15255 = n15037 ^ n15029 ;
  assign n15239 = n15024 ^ n15023 ;
  assign n15210 = n15007 ^ n14985 ;
  assign n15208 = ~n40 & n12248 ;
  assign n15206 = n4656 & n13343 ;
  assign n15203 = n4655 & ~n12239 ;
  assign n15202 = n4651 & ~n12249 ;
  assign n15204 = n15203 ^ n15202 ;
  assign n15205 = n15204 ^ x23 ;
  assign n15207 = n15206 ^ n15205 ;
  assign n15209 = n15208 ^ n15207 ;
  assign n15211 = n15210 ^ n15209 ;
  assign n15224 = n3837 & n12264 ;
  assign n15222 = n3985 & ~n12258 ;
  assign n15212 = n14912 ^ n14461 ;
  assign n15220 = n15212 ^ x29 ;
  assign n15215 = n12257 ^ n5065 ;
  assign n15216 = n15215 ^ n12257 ;
  assign n15217 = ~n14019 & n15216 ;
  assign n15218 = n15217 ^ n12257 ;
  assign n15219 = n3833 & n15218 ;
  assign n15221 = n15220 ^ n15219 ;
  assign n15223 = n15222 ^ n15221 ;
  assign n15225 = n15224 ^ n15223 ;
  assign n15232 = ~n4435 & n13677 ;
  assign n15230 = ~n4434 & ~n12251 ;
  assign n15227 = n4600 & n12253 ;
  assign n15226 = n12331 & n20603 ;
  assign n15228 = n15227 ^ n15226 ;
  assign n15229 = n15228 ^ x26 ;
  assign n15231 = n15230 ^ n15229 ;
  assign n15233 = n15232 ^ n15231 ;
  assign n15234 = n15233 ^ n15212 ;
  assign n15235 = n15225 & n15234 ;
  assign n15213 = n15212 ^ n15210 ;
  assign n15236 = n15235 ^ n15213 ;
  assign n15237 = ~n15211 & ~n15236 ;
  assign n15238 = n15237 ^ n15210 ;
  assign n15240 = n15239 ^ n15238 ;
  assign n15250 = n4651 & n12248 ;
  assign n15248 = ~n40 & ~n12239 ;
  assign n15241 = n12235 ^ x23 ;
  assign n15242 = n15241 ^ x22 ;
  assign n15243 = n15242 ^ n12235 ;
  assign n15244 = ~n13319 & n15243 ;
  assign n15245 = n15244 ^ n12235 ;
  assign n15246 = n35 & n15245 ;
  assign n15247 = n15246 ^ x23 ;
  assign n15249 = n15248 ^ n15247 ;
  assign n15251 = n15250 ^ n15249 ;
  assign n15252 = n15251 ^ n15238 ;
  assign n15253 = ~n15240 & ~n15252 ;
  assign n15254 = n15253 ^ n15251 ;
  assign n15256 = n15255 ^ n15254 ;
  assign n15266 = ~n12228 & n13433 ;
  assign n15264 = n5426 & ~n12382 ;
  assign n15257 = n12376 ^ x20 ;
  assign n15258 = n15257 ^ x19 ;
  assign n15259 = n15258 ^ n12376 ;
  assign n15260 = n12553 & n15259 ;
  assign n15261 = n15260 ^ n12376 ;
  assign n15262 = n5215 & n15261 ;
  assign n15263 = n15262 ^ x20 ;
  assign n15265 = n15264 ^ n15263 ;
  assign n15267 = n15266 ^ n15265 ;
  assign n15268 = n15267 ^ n15200 ;
  assign n15269 = n15268 ^ n15254 ;
  assign n15270 = n15269 ^ n15200 ;
  assign n15271 = n15256 & n15270 ;
  assign n15272 = n15271 ^ n15268 ;
  assign n15273 = ~n15201 & ~n15272 ;
  assign n15274 = n15273 ^ n15200 ;
  assign n15275 = n15274 ^ n15186 ;
  assign n15276 = n15191 & ~n15275 ;
  assign n15277 = n15276 ^ n15186 ;
  assign n15178 = n15154 ^ n15116 ;
  assign n15278 = n15277 ^ n15178 ;
  assign n15291 = n12209 ^ x14 ;
  assign n15280 = n12204 ^ x13 ;
  assign n15279 = n12204 ^ x14 ;
  assign n15281 = n15280 ^ n15279 ;
  assign n15282 = n12982 & n15281 ;
  assign n15283 = n15282 ^ n15280 ;
  assign n15292 = n15291 ^ n15283 ;
  assign n15284 = n12419 ^ n12209 ;
  assign n15285 = n15284 ^ n12209 ;
  assign n15286 = n12209 ^ n7310 ;
  assign n15287 = n15286 ^ n12209 ;
  assign n15288 = n15285 & n15287 ;
  assign n15289 = n15288 ^ n12209 ;
  assign n15290 = ~n6540 & ~n15289 ;
  assign n15293 = n15292 ^ n15290 ;
  assign n15294 = ~n6391 & n15293 ;
  assign n15295 = n15294 ^ n15283 ;
  assign n15296 = n15295 ^ n15277 ;
  assign n15297 = n15278 & ~n15296 ;
  assign n15298 = n15297 ^ n15295 ;
  assign n15299 = n15298 ^ n7147 ;
  assign n15177 = n15176 ^ n15159 ;
  assign n20294 = n15298 ^ n15177 ;
  assign n20295 = ~n15299 & ~n20294 ;
  assign n20296 = n20295 ^ n7147 ;
  assign n20300 = n20299 ^ n20296 ;
  assign n15573 = n6148 & ~n12214 ;
  assign n15572 = n6143 & n12222 ;
  assign n15574 = n15573 ^ n15572 ;
  assign n15575 = n15574 ^ x17 ;
  assign n15571 = n6163 & n12608 ;
  assign n15576 = n15575 ^ n15571 ;
  assign n15570 = n12380 & n20437 ;
  assign n15577 = n15576 ^ n15570 ;
  assign n15312 = n12229 & n13433 ;
  assign n15310 = n5426 & ~n12228 ;
  assign n15303 = n12382 ^ x20 ;
  assign n15304 = n15303 ^ x19 ;
  assign n15305 = n15304 ^ n12382 ;
  assign n15306 = ~n13446 & n15305 ;
  assign n15307 = n15306 ^ n12382 ;
  assign n15308 = n5215 & ~n15307 ;
  assign n15309 = n15308 ^ x20 ;
  assign n15311 = n15310 ^ n15309 ;
  assign n15313 = n15312 ^ n15311 ;
  assign n15302 = n15251 ^ n15240 ;
  assign n15314 = n15313 ^ n15302 ;
  assign n15326 = n15236 ^ n15209 ;
  assign n15324 = n12235 & n13433 ;
  assign n15322 = n5426 & n12229 ;
  assign n15315 = n12228 ^ x20 ;
  assign n15316 = n15315 ^ x19 ;
  assign n15317 = n15316 ^ n12228 ;
  assign n15318 = ~n12805 & n15317 ;
  assign n15319 = n15318 ^ n12228 ;
  assign n15320 = n5215 & ~n15319 ;
  assign n15321 = n15320 ^ x20 ;
  assign n15323 = n15322 ^ n15321 ;
  assign n15325 = n15324 ^ n15323 ;
  assign n15327 = n15326 ^ n15325 ;
  assign n15333 = n4655 & n12248 ;
  assign n15332 = n4651 & n12339 ;
  assign n15334 = n15333 ^ n15332 ;
  assign n15335 = n15334 ^ x23 ;
  assign n15331 = n4656 & ~n13519 ;
  assign n15336 = n15335 ^ n15331 ;
  assign n15330 = ~n40 & ~n12249 ;
  assign n15337 = n15336 ^ n15330 ;
  assign n15328 = n15233 ^ n15225 ;
  assign n15338 = n15337 ^ n15328 ;
  assign n15537 = n3983 & ~n14429 ;
  assign n15536 = n4369 & n12264 ;
  assign n15538 = n15537 ^ n15536 ;
  assign n15534 = n3985 & ~n12267 ;
  assign n15533 = n3837 & n12268 ;
  assign n15535 = n15534 ^ n15533 ;
  assign n15539 = n15538 ^ n15535 ;
  assign n15343 = n3983 & n14452 ;
  assign n15342 = n4369 & ~n12267 ;
  assign n15344 = n15343 ^ n15342 ;
  assign n15340 = n3837 & ~n12276 ;
  assign n15339 = n3985 & n12268 ;
  assign n15341 = n15340 ^ n15339 ;
  assign n15345 = n15344 ^ n15341 ;
  assign n15544 = n15539 ^ n15345 ;
  assign n15520 = n14893 ^ n14499 ;
  assign n15357 = n3837 & n12279 ;
  assign n15355 = n3985 & ~n12276 ;
  assign n15348 = n12268 ^ x29 ;
  assign n15349 = n15348 ^ x28 ;
  assign n15350 = n15349 ^ n12268 ;
  assign n15351 = ~n14328 & n15350 ;
  assign n15352 = n15351 ^ n12268 ;
  assign n15353 = n3833 & n15352 ;
  assign n15354 = n15353 ^ x29 ;
  assign n15356 = n15355 ^ n15354 ;
  assign n15358 = n15357 ^ n15356 ;
  assign n15346 = n14887 ^ n14567 ;
  assign n15359 = n15358 ^ n15346 ;
  assign n15371 = n3837 & ~n12283 ;
  assign n15369 = n3985 & n12279 ;
  assign n15362 = n12276 ^ x29 ;
  assign n15363 = n15362 ^ x28 ;
  assign n15364 = n15363 ^ n12276 ;
  assign n15365 = ~n14465 & n15364 ;
  assign n15366 = n15365 ^ n12276 ;
  assign n15367 = n3833 & ~n15366 ;
  assign n15368 = n15367 ^ x29 ;
  assign n15370 = n15369 ^ n15368 ;
  assign n15372 = n15371 ^ n15370 ;
  assign n15360 = n14884 ^ n14598 ;
  assign n15373 = n15372 ^ n15360 ;
  assign n15386 = n3837 & ~n12285 ;
  assign n15384 = n3985 & ~n12284 ;
  assign n15377 = n12283 ^ x29 ;
  assign n15378 = n15377 ^ x28 ;
  assign n15379 = n15378 ^ n12283 ;
  assign n15380 = ~n14547 & n15379 ;
  assign n15381 = n15380 ^ n12283 ;
  assign n15382 = n3833 & ~n15381 ;
  assign n15383 = n15382 ^ x29 ;
  assign n15385 = n15384 ^ n15383 ;
  assign n15387 = n15386 ^ n15385 ;
  assign n15375 = n14878 ^ n14718 ;
  assign n15388 = n15387 ^ n15375 ;
  assign n15399 = n3985 & ~n12285 ;
  assign n15397 = n3837 & n12313 ;
  assign n15390 = n12284 ^ x29 ;
  assign n15391 = n15390 ^ x28 ;
  assign n15392 = n15391 ^ n12284 ;
  assign n15393 = ~n14583 & n15392 ;
  assign n15394 = n15393 ^ n12284 ;
  assign n15395 = n3833 & ~n15394 ;
  assign n15396 = n15395 ^ x29 ;
  assign n15398 = n15397 ^ n15396 ;
  assign n15400 = n15399 ^ n15398 ;
  assign n15389 = n14875 ^ n14771 ;
  assign n15401 = n15400 ^ n15389 ;
  assign n15413 = n3837 & n12289 ;
  assign n15411 = n3985 & n12313 ;
  assign n15404 = n12285 ^ x29 ;
  assign n15405 = n15404 ^ x28 ;
  assign n15406 = n15405 ^ n12285 ;
  assign n15407 = ~n14651 & n15406 ;
  assign n15408 = n15407 ^ n12285 ;
  assign n15409 = n3833 & ~n15408 ;
  assign n15410 = n15409 ^ x29 ;
  assign n15412 = n15411 ^ n15410 ;
  assign n15414 = n15413 ^ n15412 ;
  assign n15402 = n14872 ^ n14803 ;
  assign n15415 = n15414 ^ n15402 ;
  assign n15418 = n3518 & n12291 ;
  assign n15423 = n12299 ^ n12293 ;
  assign n15424 = n3983 & ~n15423 ;
  assign n15422 = n3985 & n12292 ;
  assign n15425 = n15424 ^ n15422 ;
  assign n15420 = n4369 & n12293 ;
  assign n15419 = n3837 & n12291 ;
  assign n15421 = n15420 ^ n15419 ;
  assign n15426 = n15425 ^ n15421 ;
  assign n15427 = n12292 ^ n3832 ;
  assign n15428 = n3833 & ~n15427 ;
  assign n15429 = n15428 ^ n3832 ;
  assign n15430 = n12291 ^ n3833 ;
  assign n15431 = n15430 ^ x29 ;
  assign n15432 = n15429 & ~n15431 ;
  assign n15433 = n15432 ^ n3833 ;
  assign n15434 = x29 & n15433 ;
  assign n15435 = n15434 ^ x29 ;
  assign n15436 = ~n15426 & n15435 ;
  assign n15437 = ~n15418 & ~n15436 ;
  assign n15448 = n3837 & n12292 ;
  assign n15446 = n3985 & n12293 ;
  assign n15439 = n12290 ^ x29 ;
  assign n15440 = n15439 ^ x28 ;
  assign n15441 = n15440 ^ n12290 ;
  assign n15442 = n12297 & n15441 ;
  assign n15443 = n15442 ^ n12290 ;
  assign n15444 = n3833 & ~n15443 ;
  assign n15445 = n15444 ^ x29 ;
  assign n15447 = n15446 ^ n15445 ;
  assign n15449 = n15448 ^ n15447 ;
  assign n15450 = n15437 & n15449 ;
  assign n15451 = n15450 ^ n15449 ;
  assign n15417 = n14851 ^ n14822 ;
  assign n15452 = n15451 ^ n15417 ;
  assign n15463 = n3837 & n12293 ;
  assign n15461 = n3985 & ~n12290 ;
  assign n15454 = n12289 ^ x29 ;
  assign n15455 = n15454 ^ x28 ;
  assign n15456 = n15455 ^ n12289 ;
  assign n15457 = ~n14748 & n15456 ;
  assign n15458 = n15457 ^ n12289 ;
  assign n15459 = n3833 & n15458 ;
  assign n15460 = n15459 ^ x29 ;
  assign n15462 = n15461 ^ n15460 ;
  assign n15464 = n15463 ^ n15462 ;
  assign n15465 = n15464 ^ n15451 ;
  assign n15466 = ~n15452 & n15465 ;
  assign n15467 = n15466 ^ n15451 ;
  assign n15416 = n14869 ^ n14853 ;
  assign n15468 = n15467 ^ n15416 ;
  assign n15479 = n3837 & ~n12290 ;
  assign n15477 = n3985 & n12289 ;
  assign n15470 = n14712 ^ x29 ;
  assign n15471 = n15470 ^ x28 ;
  assign n15472 = n15471 ^ n14712 ;
  assign n15473 = ~n14711 & ~n15472 ;
  assign n15474 = n15473 ^ n14712 ;
  assign n15475 = n3833 & ~n15474 ;
  assign n15476 = n15475 ^ x29 ;
  assign n15478 = n15477 ^ n15476 ;
  assign n15480 = n15479 ^ n15478 ;
  assign n15481 = n15480 ^ n15416 ;
  assign n15482 = ~n15468 & n15481 ;
  assign n15483 = n15482 ^ n15467 ;
  assign n15484 = n15483 ^ n15414 ;
  assign n15485 = n15415 & n15484 ;
  assign n15486 = n15485 ^ n15414 ;
  assign n15487 = n15486 ^ n15400 ;
  assign n15488 = ~n15401 & n15487 ;
  assign n15489 = n15488 ^ n15400 ;
  assign n15490 = n15489 ^ n15387 ;
  assign n15491 = n15388 & n15490 ;
  assign n15492 = n15491 ^ n15387 ;
  assign n15374 = n14881 ^ n14668 ;
  assign n15493 = n15492 ^ n15374 ;
  assign n15504 = n3837 & ~n12284 ;
  assign n15502 = n3985 & ~n12283 ;
  assign n15500 = n15374 ^ x29 ;
  assign n15495 = n12279 ^ n5065 ;
  assign n15496 = n15495 ^ n12279 ;
  assign n15497 = ~n14514 & n15496 ;
  assign n15498 = n15497 ^ n12279 ;
  assign n15499 = n3833 & n15498 ;
  assign n15501 = n15500 ^ n15499 ;
  assign n15503 = n15502 ^ n15501 ;
  assign n15505 = n15504 ^ n15503 ;
  assign n15506 = ~n15493 & n15505 ;
  assign n15507 = n15506 ^ n15492 ;
  assign n15508 = n15507 ^ n15372 ;
  assign n15509 = ~n15373 & n15508 ;
  assign n15510 = n15509 ^ n15372 ;
  assign n15511 = n15510 ^ n15358 ;
  assign n15512 = ~n15359 & n15511 ;
  assign n15513 = n15512 ^ n15358 ;
  assign n15521 = n15520 ^ n15513 ;
  assign n15517 = n15345 ^ x29 ;
  assign n15514 = n14890 ^ n14533 ;
  assign n15518 = ~n15513 & n15514 ;
  assign n15519 = n15517 & n15518 ;
  assign n15522 = n15521 ^ n15519 ;
  assign n15545 = n15544 ^ n15522 ;
  assign n15546 = n15522 ^ n15514 ;
  assign n15547 = n15546 ^ n15522 ;
  assign n15548 = n15522 ^ n15513 ;
  assign n15549 = n15548 ^ n15522 ;
  assign n15550 = ~n15547 & n15549 ;
  assign n15551 = ~n15545 & n15550 ;
  assign n15552 = n15551 ^ n15545 ;
  assign n15553 = n15552 ^ n15544 ;
  assign n15554 = x29 & n15553 ;
  assign n15515 = n15513 & ~n15514 ;
  assign n15516 = ~n15345 & n15515 ;
  assign n15523 = n15522 ^ n15516 ;
  assign n14414 = n14088 ^ n12253 ;
  assign n15530 = ~n4435 & ~n14414 ;
  assign n15528 = ~n4434 & n12253 ;
  assign n15525 = n4600 & n12331 ;
  assign n15524 = n12257 & n20603 ;
  assign n15526 = n15525 ^ n15524 ;
  assign n15527 = n15526 ^ x26 ;
  assign n15529 = n15528 ^ n15527 ;
  assign n15531 = n15530 ^ n15529 ;
  assign n15532 = n15531 ^ n15520 ;
  assign n15540 = n15539 ^ n15532 ;
  assign n15541 = n15540 ^ n15531 ;
  assign n15542 = n15523 & n15541 ;
  assign n15543 = n15542 ^ n15532 ;
  assign n15555 = n15554 ^ n15543 ;
  assign n15558 = n14909 ^ n14897 ;
  assign n15559 = n15558 ^ n15531 ;
  assign n15560 = n15555 & ~n15559 ;
  assign n15556 = n15531 ^ n15328 ;
  assign n15561 = n15560 ^ n15556 ;
  assign n15562 = n15338 & n15561 ;
  assign n15329 = n15328 ^ n15326 ;
  assign n15563 = n15562 ^ n15329 ;
  assign n15564 = ~n15327 & ~n15563 ;
  assign n15565 = n15564 ^ n15326 ;
  assign n15566 = n15565 ^ n15313 ;
  assign n15567 = n15314 & ~n15566 ;
  assign n15568 = n15567 ^ n15313 ;
  assign n15301 = n15267 ^ n15256 ;
  assign n15569 = n15568 ^ n15301 ;
  assign n16312 = n15577 ^ n15569 ;
  assign n15943 = n15565 ^ n15314 ;
  assign n15670 = n15563 ^ n15325 ;
  assign n15665 = n6148 & n12380 ;
  assign n15664 = n6143 & n12376 ;
  assign n15666 = n15665 ^ n15664 ;
  assign n15667 = n15666 ^ x17 ;
  assign n15663 = n6163 & n12555 ;
  assign n15668 = n15667 ^ n15663 ;
  assign n15662 = ~n12382 & n20437 ;
  assign n15669 = n15668 ^ n15662 ;
  assign n15671 = n15670 ^ n15669 ;
  assign n15680 = n5426 & n12235 ;
  assign n15678 = n5220 & n12229 ;
  assign n15675 = n5221 & ~n12867 ;
  assign n15674 = ~n12239 & n13433 ;
  assign n15676 = n15675 ^ n15674 ;
  assign n15677 = n15676 ^ x20 ;
  assign n15679 = n15678 ^ n15677 ;
  assign n15681 = n15680 ^ n15679 ;
  assign n15672 = n15561 ^ n15337 ;
  assign n15682 = n15681 ^ n15672 ;
  assign n15690 = n4656 & n13554 ;
  assign n15686 = n15558 ^ n15555 ;
  assign n15687 = n15686 ^ x23 ;
  assign n15685 = n4651 & ~n12251 ;
  assign n15688 = n15687 ^ n15685 ;
  assign n15684 = n4655 & ~n12249 ;
  assign n15689 = n15688 ^ n15684 ;
  assign n15691 = n15690 ^ n15689 ;
  assign n15683 = ~n40 & n12339 ;
  assign n15692 = n15691 ^ n15683 ;
  assign n15707 = ~n4435 & ~n14972 ;
  assign n15701 = n15544 ^ n15520 ;
  assign n15698 = n15514 ^ n15513 ;
  assign n15699 = n15517 ^ n15514 ;
  assign n15700 = ~n15698 & n15699 ;
  assign n15702 = n15701 ^ n15700 ;
  assign n15703 = n15702 ^ x26 ;
  assign n15697 = n4600 & n12257 ;
  assign n15704 = n15703 ^ n15697 ;
  assign n15696 = ~n12258 & n20603 ;
  assign n15705 = n15704 ^ n15696 ;
  assign n15695 = ~n4434 & n12331 ;
  assign n15706 = n15705 ^ n15695 ;
  assign n15708 = n15707 ^ n15706 ;
  assign n15717 = ~n4435 & ~n14020 ;
  assign n15714 = n12264 & n20603 ;
  assign n15712 = n4600 & ~n12258 ;
  assign n15710 = n15698 ^ n15517 ;
  assign n15711 = n15710 ^ x26 ;
  assign n15713 = n15712 ^ n15711 ;
  assign n15715 = n15714 ^ n15713 ;
  assign n15709 = ~n4434 & n12257 ;
  assign n15716 = n15715 ^ n15709 ;
  assign n15718 = n15717 ^ n15716 ;
  assign n15727 = ~n4435 & n14243 ;
  assign n15724 = ~n12267 & n20603 ;
  assign n15722 = ~n4434 & ~n12258 ;
  assign n15720 = n15510 ^ n15359 ;
  assign n15721 = n15720 ^ x26 ;
  assign n15723 = n15722 ^ n15721 ;
  assign n15725 = n15724 ^ n15723 ;
  assign n15719 = n4600 & n12264 ;
  assign n15726 = n15725 ^ n15719 ;
  assign n15728 = n15727 ^ n15726 ;
  assign n15736 = ~n4435 & ~n14429 ;
  assign n15734 = ~n4434 & n12264 ;
  assign n15731 = n4600 & ~n12267 ;
  assign n15730 = n12268 & n20603 ;
  assign n15732 = n15731 ^ n15730 ;
  assign n15733 = n15732 ^ x26 ;
  assign n15735 = n15734 ^ n15733 ;
  assign n15737 = n15736 ^ n15735 ;
  assign n15729 = n15507 ^ n15373 ;
  assign n15738 = n15737 ^ n15729 ;
  assign n15746 = ~n4435 & n14452 ;
  assign n15744 = ~n4434 & ~n12267 ;
  assign n15741 = ~n12276 & n20603 ;
  assign n15740 = n4600 & n12268 ;
  assign n15742 = n15741 ^ n15740 ;
  assign n15743 = n15742 ^ x26 ;
  assign n15745 = n15744 ^ n15743 ;
  assign n15747 = n15746 ^ n15745 ;
  assign n15739 = n15505 ^ n15492 ;
  assign n15748 = n15747 ^ n15739 ;
  assign n15756 = ~n4435 & ~n14329 ;
  assign n15754 = n4600 & ~n12276 ;
  assign n15751 = ~n4434 & n12268 ;
  assign n15750 = n12279 & n20603 ;
  assign n15752 = n15751 ^ n15750 ;
  assign n15753 = n15752 ^ x26 ;
  assign n15755 = n15754 ^ n15753 ;
  assign n15757 = n15756 ^ n15755 ;
  assign n15749 = n15489 ^ n15388 ;
  assign n15758 = n15757 ^ n15749 ;
  assign n15765 = ~x25 & ~n14514 ;
  assign n15768 = n15765 ^ n14528 ;
  assign n15769 = n99 & ~n15768 ;
  assign n15762 = n4600 & ~n12283 ;
  assign n15761 = ~n12284 & n20603 ;
  assign n15763 = n15762 ^ n15761 ;
  assign n15764 = n15763 ^ x26 ;
  assign n15766 = n15765 ^ n12279 ;
  assign n15767 = n15764 & ~n15766 ;
  assign n15770 = n15769 ^ n15767 ;
  assign n15771 = n15763 ^ n97 ;
  assign n15772 = ~n15770 & ~n15771 ;
  assign n15760 = n15483 ^ n15415 ;
  assign n15773 = n15772 ^ n15760 ;
  assign n15781 = ~n4435 & n14548 ;
  assign n15779 = ~n4434 & ~n12283 ;
  assign n15776 = n4600 & ~n12284 ;
  assign n15775 = ~n12285 & n20603 ;
  assign n15777 = n15776 ^ n15775 ;
  assign n15778 = n15777 ^ x26 ;
  assign n15780 = n15779 ^ n15778 ;
  assign n15782 = n15781 ^ n15780 ;
  assign n15774 = n15480 ^ n15468 ;
  assign n15783 = n15782 ^ n15774 ;
  assign n15786 = n12313 & n20603 ;
  assign n15785 = n4600 & ~n12285 ;
  assign n15787 = n15786 ^ n15785 ;
  assign n15788 = n15787 ^ n97 ;
  assign n15789 = n15787 ^ x26 ;
  assign n15794 = n15789 ^ n99 ;
  assign n15790 = n13110 ^ n12284 ;
  assign n15791 = n15790 ^ n14583 ;
  assign n15792 = n15791 ^ n15790 ;
  assign n15793 = n15789 & ~n15792 ;
  assign n15795 = n15794 ^ n15793 ;
  assign n15798 = ~n13110 & ~n15792 ;
  assign n15799 = n15798 ^ n12284 ;
  assign n15800 = ~n15794 & n15799 ;
  assign n15801 = ~n15795 & n15800 ;
  assign n15802 = n15801 ^ n15798 ;
  assign n15805 = n15802 ^ n99 ;
  assign n15806 = n15805 ^ n12284 ;
  assign n15807 = ~n15788 & ~n15806 ;
  assign n15784 = n15464 ^ n15452 ;
  assign n15808 = n15807 ^ n15784 ;
  assign n15818 = n15449 ^ n15436 ;
  assign n15819 = n15818 ^ n15418 ;
  assign n15815 = ~n4435 & n14652 ;
  assign n15813 = n4600 & n12313 ;
  assign n15810 = ~n4434 & ~n12285 ;
  assign n15809 = n12289 & n20603 ;
  assign n15811 = n15810 ^ n15809 ;
  assign n15812 = n15811 ^ x26 ;
  assign n15814 = n15813 ^ n15812 ;
  assign n15816 = n15815 ^ n15814 ;
  assign n15820 = n15819 ^ n15816 ;
  assign n15829 = n15434 ^ n15426 ;
  assign n15827 = ~n4435 & ~n14712 ;
  assign n15825 = ~n4434 & n12313 ;
  assign n15822 = n4600 & n12289 ;
  assign n15821 = ~n12290 & n20603 ;
  assign n15823 = n15822 ^ n15821 ;
  assign n15824 = n15823 ^ x26 ;
  assign n15826 = n15825 ^ n15824 ;
  assign n15828 = n15827 ^ n15826 ;
  assign n15830 = n15829 ^ n15828 ;
  assign n15835 = n3833 & n12292 ;
  assign n15834 = n3832 & n12291 ;
  assign n15836 = n15835 ^ n15834 ;
  assign n15872 = n15836 ^ n15829 ;
  assign n15840 = ~n4434 & n12289 ;
  assign n15837 = n15836 ^ x26 ;
  assign n15833 = n12293 & n20603 ;
  assign n15838 = n15837 ^ n15833 ;
  assign n15832 = n4600 & ~n12290 ;
  assign n15839 = n15838 ^ n15832 ;
  assign n15841 = n15840 ^ n15839 ;
  assign n15831 = ~n4435 & ~n14749 ;
  assign n15842 = n15841 ^ n15831 ;
  assign n15843 = n3833 & n12291 ;
  assign n15844 = n96 & n12292 ;
  assign n15845 = x26 & ~n15844 ;
  assign n15846 = n12291 & n15845 ;
  assign n15847 = n7678 & n15846 ;
  assign n15848 = n15847 ^ n15845 ;
  assign n15855 = ~n4434 & n12293 ;
  assign n15853 = n4600 & n12292 ;
  assign n15852 = n12291 & n20603 ;
  assign n15854 = n15853 ^ n15852 ;
  assign n15856 = n15855 ^ n15854 ;
  assign n15851 = ~n4435 & ~n15423 ;
  assign n15857 = n15856 ^ n15851 ;
  assign n15858 = n15848 & ~n15857 ;
  assign n15859 = ~n15843 & ~n15858 ;
  assign n15866 = ~n4435 & ~n14785 ;
  assign n15864 = ~n4434 & ~n12290 ;
  assign n15861 = n4600 & n12293 ;
  assign n15860 = n12292 & n20603 ;
  assign n15862 = n15861 ^ n15860 ;
  assign n15863 = n15862 ^ x26 ;
  assign n15865 = n15864 ^ n15863 ;
  assign n15867 = n15866 ^ n15865 ;
  assign n15868 = n15859 & n15867 ;
  assign n15869 = n15868 ^ n15867 ;
  assign n15870 = n15869 ^ n15836 ;
  assign n15871 = n15842 & n15870 ;
  assign n15873 = n15872 ^ n15871 ;
  assign n15874 = n15830 & n15873 ;
  assign n15875 = n15874 ^ n15829 ;
  assign n15876 = n15875 ^ n15816 ;
  assign n15877 = n15820 & n15876 ;
  assign n15817 = n15816 ^ n15807 ;
  assign n15878 = n15877 ^ n15817 ;
  assign n15879 = n15808 & ~n15878 ;
  assign n15880 = n15879 ^ n15807 ;
  assign n15881 = n15880 ^ n15782 ;
  assign n15882 = ~n15783 & ~n15881 ;
  assign n15883 = n15882 ^ n15782 ;
  assign n15884 = n15883 ^ n15772 ;
  assign n15885 = ~n15773 & ~n15884 ;
  assign n15886 = n15885 ^ n15772 ;
  assign n15759 = n15486 ^ n15401 ;
  assign n15887 = n15886 ^ n15759 ;
  assign n15889 = n4600 & n12279 ;
  assign n15888 = ~n12283 & n20603 ;
  assign n15890 = n15889 ^ n15888 ;
  assign n15891 = n15890 ^ n97 ;
  assign n15892 = n15890 ^ x26 ;
  assign n15893 = n15892 ^ n99 ;
  assign n15894 = n13110 ^ n12276 ;
  assign n15895 = n15894 ^ n14465 ;
  assign n15896 = n15895 ^ n15894 ;
  assign n15900 = ~n13110 & ~n15896 ;
  assign n15901 = n15900 ^ n12276 ;
  assign n15902 = ~n15893 & n15901 ;
  assign n15910 = ~n15892 & n15902 ;
  assign n15903 = n15902 ^ n99 ;
  assign n15905 = n15903 ^ x25 ;
  assign n15911 = n15910 ^ n15905 ;
  assign n15912 = ~n14465 & ~n15911 ;
  assign n15904 = n15903 ^ n12276 ;
  assign n15913 = n15912 ^ n15904 ;
  assign n15914 = ~n15891 & ~n15913 ;
  assign n15915 = n15914 ^ n15886 ;
  assign n15916 = n15887 & n15915 ;
  assign n15917 = n15916 ^ n15886 ;
  assign n15918 = n15917 ^ n15757 ;
  assign n15919 = n15758 & ~n15918 ;
  assign n15920 = n15919 ^ n15757 ;
  assign n15921 = n15920 ^ n15747 ;
  assign n15922 = ~n15748 & n15921 ;
  assign n15923 = n15922 ^ n15747 ;
  assign n15924 = n15923 ^ n15737 ;
  assign n15925 = ~n15738 & n15924 ;
  assign n15926 = n15925 ^ n15737 ;
  assign n15927 = n15926 ^ n15720 ;
  assign n15928 = ~n15728 & ~n15927 ;
  assign n15929 = n15928 ^ n15720 ;
  assign n15930 = n15929 ^ n15710 ;
  assign n15931 = n15718 & ~n15930 ;
  assign n15932 = n15931 ^ n15710 ;
  assign n15933 = n15932 ^ n15702 ;
  assign n15934 = n15708 & n15933 ;
  assign n15935 = n15934 ^ n15702 ;
  assign n15693 = n15686 ^ n15672 ;
  assign n15694 = n15693 ^ n15672 ;
  assign n15936 = n15935 ^ n15694 ;
  assign n15937 = ~n15692 & ~n15936 ;
  assign n15938 = n15937 ^ n15693 ;
  assign n15939 = n15682 & ~n15938 ;
  assign n15673 = n15672 ^ n15670 ;
  assign n15940 = n15939 ^ n15673 ;
  assign n15941 = ~n15671 & ~n15940 ;
  assign n15942 = n15941 ^ n15670 ;
  assign n15944 = n15943 ^ n15942 ;
  assign n15645 = n6143 & n12380 ;
  assign n15644 = n12376 & n20437 ;
  assign n15646 = n15645 ^ n15644 ;
  assign n15647 = n15646 ^ n6145 ;
  assign n15648 = n15646 ^ x17 ;
  assign n15649 = n15648 ^ n6147 ;
  assign n15650 = ~n13770 & n15649 ;
  assign n15651 = n15650 ^ n6147 ;
  assign n15652 = n15651 ^ x16 ;
  assign n15653 = n15652 ^ n12222 ;
  assign n15654 = n15653 ^ n15651 ;
  assign n15655 = n15651 ^ n15649 ;
  assign n15656 = n15655 ^ n15651 ;
  assign n15657 = n15654 & n15656 ;
  assign n15658 = n15657 ^ n15651 ;
  assign n15659 = n12390 & n15658 ;
  assign n15660 = n15659 ^ n15651 ;
  assign n15661 = ~n15647 & ~n15660 ;
  assign n16309 = n15942 ^ n15661 ;
  assign n16310 = ~n15944 & n16309 ;
  assign n16311 = n16310 ^ n15661 ;
  assign n16313 = n16312 ^ n16311 ;
  assign n15583 = n12405 ^ x12 ;
  assign n15584 = n15583 ^ n12405 ;
  assign n15585 = ~x13 & x14 ;
  assign n15586 = ~n12210 & n15585 ;
  assign n15587 = n15586 ^ n12405 ;
  assign n15588 = ~n15584 & ~n15587 ;
  assign n15589 = n15588 ^ n12405 ;
  assign n15590 = ~n6391 & ~n15589 ;
  assign n15591 = n15590 ^ n6391 ;
  assign n15592 = ~n6534 & n15591 ;
  assign n15593 = n12405 ^ x11 ;
  assign n15594 = n15593 ^ n12405 ;
  assign n15595 = n12405 ^ n12210 ;
  assign n15596 = n15595 ^ n12405 ;
  assign n15597 = ~x14 & ~n15596 ;
  assign n15598 = n15597 ^ n12405 ;
  assign n15599 = n15594 & ~n15598 ;
  assign n15600 = n15599 ^ n12405 ;
  assign n15601 = x13 & ~n15600 ;
  assign n15602 = ~n15592 & ~n15601 ;
  assign n15603 = n15602 ^ x14 ;
  assign n15604 = n15603 ^ x13 ;
  assign n15605 = n15604 ^ n12419 ;
  assign n15606 = n15605 ^ n12650 ;
  assign n15607 = n15606 ^ n15605 ;
  assign n15608 = n15605 ^ n7310 ;
  assign n15609 = ~n12419 & ~n15608 ;
  assign n15610 = n15609 ^ n15605 ;
  assign n15611 = n15607 & ~n15610 ;
  assign n15612 = n15611 ^ n15605 ;
  assign n15613 = n6391 & ~n15612 ;
  assign n15614 = n15613 ^ n15603 ;
  assign n15581 = n15272 ^ n15199 ;
  assign n15578 = n15577 ^ n15568 ;
  assign n15579 = n15569 & n15578 ;
  assign n15580 = n15579 ^ n15577 ;
  assign n15582 = n15581 ^ n15580 ;
  assign n20212 = n15614 ^ n15582 ;
  assign n20213 = n20212 ^ n16311 ;
  assign n20214 = n20213 ^ n20212 ;
  assign n16291 = ~n6547 & ~n12400 ;
  assign n16290 = ~n6529 & ~n12210 ;
  assign n16292 = n16291 ^ n16290 ;
  assign n16293 = n16292 ^ n6537 ;
  assign n16294 = n16293 ^ x14 ;
  assign n16304 = x13 & ~n12715 ;
  assign n16303 = n8856 & ~n12405 ;
  assign n16305 = n16304 ^ n16303 ;
  assign n16306 = ~n6539 & n16305 ;
  assign n16301 = n12714 ^ n8856 ;
  assign n16295 = n16292 ^ x14 ;
  assign n16296 = n12405 ^ x13 ;
  assign n16297 = n16296 ^ n12405 ;
  assign n16298 = ~n12714 & ~n16297 ;
  assign n16299 = n16298 ^ n12405 ;
  assign n16300 = ~n16295 & n16299 ;
  assign n16302 = n16301 ^ n16300 ;
  assign n16307 = n16306 ^ n16302 ;
  assign n16308 = ~n16294 & n16307 ;
  assign n20215 = n20214 ^ n16308 ;
  assign n20216 = n16313 & n20215 ;
  assign n20217 = n20216 ^ n20213 ;
  assign n20202 = n7142 & ~n12204 ;
  assign n20201 = n7148 & ~n12209 ;
  assign n20203 = n20202 ^ n20201 ;
  assign n20200 = n7140 & ~n12435 ;
  assign n20204 = n20203 ^ n20200 ;
  assign n20205 = n20204 ^ n20203 ;
  assign n20206 = n12432 & n20205 ;
  assign n20207 = n20204 ^ x11 ;
  assign n20208 = n20207 ^ x10 ;
  assign n20209 = n20208 ^ n20204 ;
  assign n20210 = n20206 & n20209 ;
  assign n20211 = n20210 ^ n20207 ;
  assign n20218 = n20217 ^ n20211 ;
  assign n20219 = n20218 ^ n13608 ;
  assign n16314 = n16313 ^ n16308 ;
  assign n15956 = ~n6392 & n7310 ;
  assign n15957 = n12214 ^ x13 ;
  assign n15958 = n15957 ^ n12214 ;
  assign n15959 = n12400 ^ n12214 ;
  assign n15962 = ~n15958 & ~n15959 ;
  assign n15963 = n15962 ^ n12214 ;
  assign n15964 = n15956 & n15963 ;
  assign n15965 = n15964 ^ n6543 ;
  assign n15954 = ~n6541 & n6543 ;
  assign n15955 = ~n12400 & n15954 ;
  assign n15966 = n15965 ^ n15955 ;
  assign n15967 = n12214 ^ x14 ;
  assign n15968 = n15967 ^ n12214 ;
  assign n15969 = ~n12400 & n15968 ;
  assign n15970 = n15969 ^ n12214 ;
  assign n15971 = n15958 & ~n15970 ;
  assign n15972 = n15971 ^ n12214 ;
  assign n15973 = n6390 & ~n15972 ;
  assign n15974 = ~n15966 & ~n15973 ;
  assign n15947 = n12210 ^ x14 ;
  assign n15946 = n12210 ^ x13 ;
  assign n15948 = n15947 ^ n15946 ;
  assign n15949 = n15947 ^ n12736 ;
  assign n15950 = n15949 ^ n15947 ;
  assign n15951 = n15948 & ~n15950 ;
  assign n15952 = n15951 ^ n15947 ;
  assign n15953 = n6391 & n15952 ;
  assign n15975 = n15974 ^ n15953 ;
  assign n15945 = n15944 ^ n15661 ;
  assign n15976 = n15975 ^ n15945 ;
  assign n15984 = x13 ^ x11 ;
  assign n15994 = n12222 ^ n12214 ;
  assign n15995 = n15994 ^ x13 ;
  assign n15996 = ~n15984 & ~n15995 ;
  assign n15985 = n15984 ^ x14 ;
  assign n15988 = x13 & ~n12222 ;
  assign n15989 = n15988 ^ n12214 ;
  assign n15990 = n15968 & ~n15989 ;
  assign n15991 = n15990 ^ n12214 ;
  assign n15992 = n15985 & ~n15991 ;
  assign n15979 = n12400 ^ x13 ;
  assign n15980 = n15979 ^ x14 ;
  assign n15981 = n15980 ^ n12400 ;
  assign n15982 = n12666 & n15981 ;
  assign n15983 = n15982 ^ n15979 ;
  assign n15986 = n15983 ^ n12214 ;
  assign n15993 = n15992 ^ n15986 ;
  assign n15997 = n15996 ^ n15993 ;
  assign n15998 = ~n6391 & ~n15997 ;
  assign n15999 = n15998 ^ n15983 ;
  assign n16004 = ~n12214 & n15954 ;
  assign n16005 = n16004 ^ n6543 ;
  assign n16006 = ~n15999 & ~n16005 ;
  assign n15977 = n15940 ^ n15669 ;
  assign n16007 = n16006 ^ n15977 ;
  assign n16019 = n12248 & n13433 ;
  assign n16017 = n5426 & ~n12239 ;
  assign n16010 = n12235 ^ x20 ;
  assign n16011 = n16010 ^ x19 ;
  assign n16012 = n16011 ^ n12235 ;
  assign n16013 = ~n13319 & n16012 ;
  assign n16014 = n16013 ^ n12235 ;
  assign n16015 = n5215 & n16014 ;
  assign n16016 = n16015 ^ x20 ;
  assign n16018 = n16017 ^ n16016 ;
  assign n16020 = n16019 ^ n16018 ;
  assign n16009 = n15935 ^ n15692 ;
  assign n16021 = n16020 ^ n16009 ;
  assign n16029 = ~n40 & ~n12251 ;
  assign n16027 = n4656 & ~n13885 ;
  assign n16024 = n4655 & n12339 ;
  assign n16023 = n4651 & n12253 ;
  assign n16025 = n16024 ^ n16023 ;
  assign n16026 = n16025 ^ x23 ;
  assign n16028 = n16027 ^ n16026 ;
  assign n16030 = n16029 ^ n16028 ;
  assign n16022 = n15932 ^ n15708 ;
  assign n16031 = n16030 ^ n16022 ;
  assign n16036 = n4655 & ~n12251 ;
  assign n16035 = n4651 & n12331 ;
  assign n16037 = n16036 ^ n16035 ;
  assign n16038 = n16037 ^ x23 ;
  assign n16034 = n4656 & n13677 ;
  assign n16039 = n16038 ^ n16034 ;
  assign n16033 = ~n40 & n12253 ;
  assign n16040 = n16039 ^ n16033 ;
  assign n16032 = n15929 ^ n15718 ;
  assign n16041 = n16040 ^ n16032 ;
  assign n16046 = n4655 & n12253 ;
  assign n16045 = n4651 & n12257 ;
  assign n16047 = n16046 ^ n16045 ;
  assign n16048 = n16047 ^ x23 ;
  assign n16044 = n4656 & ~n14414 ;
  assign n16049 = n16048 ^ n16044 ;
  assign n16043 = ~n40 & n12331 ;
  assign n16050 = n16049 ^ n16043 ;
  assign n16042 = n15926 ^ n15728 ;
  assign n16051 = n16050 ^ n16042 ;
  assign n16059 = ~n40 & n12257 ;
  assign n16057 = n4656 & ~n14972 ;
  assign n16054 = n4655 & n12331 ;
  assign n16053 = n4651 & ~n12258 ;
  assign n16055 = n16054 ^ n16053 ;
  assign n16056 = n16055 ^ x23 ;
  assign n16058 = n16057 ^ n16056 ;
  assign n16060 = n16059 ^ n16058 ;
  assign n16052 = n15923 ^ n15738 ;
  assign n16061 = n16060 ^ n16052 ;
  assign n16069 = ~n40 & ~n12258 ;
  assign n16067 = n4656 & ~n14020 ;
  assign n16064 = n4655 & n12257 ;
  assign n16063 = n4651 & n12264 ;
  assign n16065 = n16064 ^ n16063 ;
  assign n16066 = n16065 ^ x23 ;
  assign n16068 = n16067 ^ n16066 ;
  assign n16070 = n16069 ^ n16068 ;
  assign n16062 = n15920 ^ n15748 ;
  assign n16071 = n16070 ^ n16062 ;
  assign n16079 = ~n40 & n12264 ;
  assign n16077 = n4656 & n14243 ;
  assign n16074 = n4655 & ~n12258 ;
  assign n16073 = n4651 & ~n12267 ;
  assign n16075 = n16074 ^ n16073 ;
  assign n16076 = n16075 ^ x23 ;
  assign n16078 = n16077 ^ n16076 ;
  assign n16080 = n16079 ^ n16078 ;
  assign n16072 = n15917 ^ n15758 ;
  assign n16081 = n16080 ^ n16072 ;
  assign n16089 = ~n40 & ~n12267 ;
  assign n16087 = n4656 & ~n14429 ;
  assign n16084 = n4655 & n12264 ;
  assign n16083 = n4651 & n12268 ;
  assign n16085 = n16084 ^ n16083 ;
  assign n16086 = n16085 ^ x23 ;
  assign n16088 = n16087 ^ n16086 ;
  assign n16090 = n16089 ^ n16088 ;
  assign n16082 = n15915 ^ n15759 ;
  assign n16091 = n16090 ^ n16082 ;
  assign n16096 = n4655 & ~n12267 ;
  assign n16095 = n4651 & ~n12276 ;
  assign n16097 = n16096 ^ n16095 ;
  assign n16098 = n16097 ^ x23 ;
  assign n16094 = n4656 & n14452 ;
  assign n16099 = n16098 ^ n16094 ;
  assign n16093 = ~n40 & n12268 ;
  assign n16100 = n16099 ^ n16093 ;
  assign n16092 = n15883 ^ n15773 ;
  assign n16101 = n16100 ^ n16092 ;
  assign n16112 = ~n40 & ~n12283 ;
  assign n16105 = n12279 ^ x23 ;
  assign n16106 = n16105 ^ x22 ;
  assign n16107 = n16106 ^ n12279 ;
  assign n16108 = ~n14514 & n16107 ;
  assign n16109 = n16108 ^ n12279 ;
  assign n16110 = n35 & n16109 ;
  assign n16111 = n16110 ^ x23 ;
  assign n16113 = n16112 ^ n16111 ;
  assign n16104 = n4651 & ~n12284 ;
  assign n16114 = n16113 ^ n16104 ;
  assign n16103 = n15875 ^ n15820 ;
  assign n16115 = n16114 ^ n16103 ;
  assign n16126 = n4651 & ~n12285 ;
  assign n16124 = ~n40 & ~n12284 ;
  assign n16117 = n12283 ^ x23 ;
  assign n16118 = n16117 ^ x22 ;
  assign n16119 = n16118 ^ n12283 ;
  assign n16120 = ~n14547 & n16119 ;
  assign n16121 = n16120 ^ n12283 ;
  assign n16122 = n35 & ~n16121 ;
  assign n16123 = n16122 ^ x23 ;
  assign n16125 = n16124 ^ n16123 ;
  assign n16127 = n16126 ^ n16125 ;
  assign n16116 = n15873 ^ n15828 ;
  assign n16128 = n16127 ^ n16116 ;
  assign n16138 = n15869 ^ n15842 ;
  assign n16132 = n4655 & ~n12284 ;
  assign n16131 = n4651 & n12313 ;
  assign n16133 = n16132 ^ n16131 ;
  assign n16134 = n16133 ^ x23 ;
  assign n14584 = n14583 ^ n12284 ;
  assign n16130 = n4656 & n14584 ;
  assign n16135 = n16134 ^ n16130 ;
  assign n16129 = ~n40 & ~n12285 ;
  assign n16136 = n16135 ^ n16129 ;
  assign n16139 = n16138 ^ n16136 ;
  assign n16145 = n4655 & ~n12285 ;
  assign n16144 = n4651 & n12289 ;
  assign n16146 = n16145 ^ n16144 ;
  assign n16147 = n16146 ^ x23 ;
  assign n16143 = n4656 & n14652 ;
  assign n16148 = n16147 ^ n16143 ;
  assign n16142 = ~n40 & n12313 ;
  assign n16149 = n16148 ^ n16142 ;
  assign n16140 = n15858 ^ n15843 ;
  assign n16141 = n16140 ^ n15867 ;
  assign n16150 = n16149 ^ n16141 ;
  assign n15849 = n15848 ^ x26 ;
  assign n16192 = n15857 ^ n15849 ;
  assign n16181 = n4655 & n12289 ;
  assign n16180 = n4651 & n12293 ;
  assign n16182 = n16181 ^ n16180 ;
  assign n16183 = n16182 ^ x23 ;
  assign n16179 = n4656 & ~n14749 ;
  assign n16184 = n16183 ^ n16179 ;
  assign n16178 = ~n40 & ~n12290 ;
  assign n16185 = n16184 ^ n16178 ;
  assign n16151 = n96 & n12291 ;
  assign n16152 = n35 & n12292 ;
  assign n16153 = x23 & ~n16152 ;
  assign n16154 = n12291 & n16153 ;
  assign n16155 = ~n42 & n16154 ;
  assign n16156 = n16155 ^ n16153 ;
  assign n16163 = n4656 & ~n15423 ;
  assign n16162 = n4651 & n12291 ;
  assign n16164 = n16163 ^ n16162 ;
  assign n16160 = n4655 & n12293 ;
  assign n16159 = ~n40 & n12292 ;
  assign n16161 = n16160 ^ n16159 ;
  assign n16165 = n16164 ^ n16161 ;
  assign n16166 = n16156 & ~n16165 ;
  assign n16167 = ~n16151 & ~n16166 ;
  assign n16174 = ~n40 & n12293 ;
  assign n16172 = n4656 & ~n14785 ;
  assign n16169 = n4655 & ~n12290 ;
  assign n16168 = n4651 & n12292 ;
  assign n16170 = n16169 ^ n16168 ;
  assign n16171 = n16170 ^ x23 ;
  assign n16173 = n16172 ^ n16171 ;
  assign n16175 = n16174 ^ n16173 ;
  assign n16176 = n16167 & n16175 ;
  assign n16177 = n16176 ^ n16175 ;
  assign n16186 = n16185 ^ n16177 ;
  assign n16188 = n16177 ^ n15844 ;
  assign n16187 = ~n7925 & n12291 ;
  assign n16189 = n16188 ^ n16187 ;
  assign n16190 = n16186 & ~n16189 ;
  assign n16191 = n16190 ^ n16185 ;
  assign n16193 = n16192 ^ n16191 ;
  assign n16200 = ~n40 & n12289 ;
  assign n16198 = n4656 & ~n14712 ;
  assign n16195 = n4655 & n12313 ;
  assign n16194 = n4651 & ~n12290 ;
  assign n16196 = n16195 ^ n16194 ;
  assign n16197 = n16196 ^ x23 ;
  assign n16199 = n16198 ^ n16197 ;
  assign n16201 = n16200 ^ n16199 ;
  assign n16202 = n16201 ^ n16191 ;
  assign n16203 = ~n16193 & n16202 ;
  assign n16204 = n16203 ^ n16201 ;
  assign n16205 = n16204 ^ n16141 ;
  assign n16206 = n16150 & ~n16205 ;
  assign n16207 = n16206 ^ n16149 ;
  assign n16208 = n16207 ^ n16136 ;
  assign n16209 = n16139 & n16208 ;
  assign n16137 = n16136 ^ n16127 ;
  assign n16210 = n16209 ^ n16137 ;
  assign n16211 = n16128 & n16210 ;
  assign n16212 = n16211 ^ n16127 ;
  assign n16213 = n16212 ^ n16114 ;
  assign n16214 = n16115 & n16213 ;
  assign n16215 = n16214 ^ n16114 ;
  assign n16102 = n15878 ^ n15784 ;
  assign n16217 = n16215 ^ n16102 ;
  assign n16216 = n16102 & n16215 ;
  assign n16218 = n16217 ^ n16216 ;
  assign n16223 = n4656 & n14475 ;
  assign n16222 = ~n40 & n12279 ;
  assign n16224 = n16223 ^ n16222 ;
  assign n16220 = n4655 & ~n12276 ;
  assign n16219 = n4651 & ~n12283 ;
  assign n16221 = n16220 ^ n16219 ;
  assign n16225 = n16224 ^ n16221 ;
  assign n16226 = n16225 ^ x23 ;
  assign n16234 = n15880 ^ n15783 ;
  assign n16235 = n16234 ^ n16225 ;
  assign n16231 = n4656 & ~n14329 ;
  assign n16230 = ~n40 & ~n12276 ;
  assign n16232 = n16231 ^ n16230 ;
  assign n16228 = n4655 & n12268 ;
  assign n16227 = n4651 & n12279 ;
  assign n16229 = n16228 ^ n16227 ;
  assign n16233 = n16232 ^ n16229 ;
  assign n16236 = n16235 ^ n16233 ;
  assign n16237 = n16226 & ~n16236 ;
  assign n16238 = n16218 & n16237 ;
  assign n16239 = n16234 ^ n16216 ;
  assign n16240 = n16233 ^ x23 ;
  assign n16241 = n16240 ^ n16216 ;
  assign n16242 = n16239 & n16241 ;
  assign n16243 = n16242 ^ n16216 ;
  assign n16244 = ~n16238 & ~n16243 ;
  assign n16245 = n16244 ^ n16100 ;
  assign n16246 = ~n16101 & ~n16245 ;
  assign n16247 = n16246 ^ n16100 ;
  assign n16248 = n16247 ^ n16090 ;
  assign n16249 = ~n16091 & n16248 ;
  assign n16250 = n16249 ^ n16090 ;
  assign n16251 = n16250 ^ n16080 ;
  assign n16252 = ~n16081 & n16251 ;
  assign n16253 = n16252 ^ n16080 ;
  assign n16254 = n16253 ^ n16070 ;
  assign n16255 = ~n16071 & n16254 ;
  assign n16256 = n16255 ^ n16070 ;
  assign n16257 = n16256 ^ n16060 ;
  assign n16258 = ~n16061 & n16257 ;
  assign n16259 = n16258 ^ n16060 ;
  assign n16260 = n16259 ^ n16050 ;
  assign n16261 = ~n16051 & n16260 ;
  assign n16262 = n16261 ^ n16050 ;
  assign n16263 = n16262 ^ n16040 ;
  assign n16264 = ~n16041 & n16263 ;
  assign n16265 = n16264 ^ n16040 ;
  assign n16266 = n16265 ^ n16030 ;
  assign n16267 = n16031 & n16266 ;
  assign n16268 = n16267 ^ n16030 ;
  assign n16269 = n16268 ^ n16020 ;
  assign n16270 = ~n16021 & n16269 ;
  assign n16271 = n16270 ^ n16020 ;
  assign n16008 = n15938 ^ n15681 ;
  assign n16272 = n16271 ^ n16008 ;
  assign n16280 = ~n12228 & n20437 ;
  assign n16278 = n6163 & n12928 ;
  assign n16275 = n6148 & n12376 ;
  assign n16274 = n6143 & ~n12382 ;
  assign n16276 = n16275 ^ n16274 ;
  assign n16277 = n16276 ^ x17 ;
  assign n16279 = n16278 ^ n16277 ;
  assign n16281 = n16280 ^ n16279 ;
  assign n16273 = n16271 ^ n15977 ;
  assign n16282 = n16281 ^ n16273 ;
  assign n16283 = n16282 ^ n15977 ;
  assign n16284 = ~n16272 & n16283 ;
  assign n16285 = n16284 ^ n16273 ;
  assign n16286 = ~n16007 & ~n16285 ;
  assign n15978 = n15977 ^ n15975 ;
  assign n16287 = n16286 ^ n15978 ;
  assign n16288 = ~n15976 & ~n16287 ;
  assign n16289 = n16288 ^ n15975 ;
  assign n16315 = n16314 ^ n16289 ;
  assign n15642 = n7148 & n12419 ;
  assign n15640 = n7142 & ~n12209 ;
  assign n15633 = n12204 ^ x11 ;
  assign n15634 = n15633 ^ x10 ;
  assign n15635 = n15634 ^ n12204 ;
  assign n15636 = ~n13415 & n15635 ;
  assign n15637 = n15636 ^ n12204 ;
  assign n15638 = n7140 & ~n15637 ;
  assign n15639 = n15638 ^ x11 ;
  assign n15641 = n15640 ^ n15639 ;
  assign n15643 = n15642 ^ n15641 ;
  assign n20220 = n16289 ^ n15643 ;
  assign n20221 = n16315 & n20220 ;
  assign n20222 = n20221 ^ n15643 ;
  assign n20232 = n20222 ^ n20218 ;
  assign n20233 = ~n20219 & n20232 ;
  assign n20234 = n20233 ^ n13608 ;
  assign n20223 = n20222 ^ n20219 ;
  assign n17728 = n7151 & ~n12405 ;
  assign n17727 = n7148 & ~n12400 ;
  assign n17729 = n17728 ^ n17727 ;
  assign n17730 = n17729 ^ x11 ;
  assign n17726 = n12715 & n20240 ;
  assign n17731 = n17730 ^ n17726 ;
  assign n17725 = n7142 & ~n12210 ;
  assign n17732 = n17731 ^ n17725 ;
  assign n16354 = ~n12249 & n13433 ;
  assign n16352 = n5426 & n12248 ;
  assign n16349 = n16265 ^ n16031 ;
  assign n16350 = n16349 ^ x20 ;
  assign n16344 = n12239 ^ n5224 ;
  assign n16345 = n16344 ^ n12239 ;
  assign n16346 = ~n13339 & n16345 ;
  assign n16347 = n16346 ^ n12239 ;
  assign n16348 = n5215 & ~n16347 ;
  assign n16351 = n16350 ^ n16348 ;
  assign n16353 = n16352 ^ n16351 ;
  assign n16355 = n16354 ^ n16353 ;
  assign n16363 = n5426 & ~n12249 ;
  assign n16361 = n5220 & n12248 ;
  assign n16358 = n5221 & ~n13519 ;
  assign n16357 = n12339 & n13433 ;
  assign n16359 = n16358 ^ n16357 ;
  assign n16360 = n16359 ^ x20 ;
  assign n16362 = n16361 ^ n16360 ;
  assign n16364 = n16363 ^ n16362 ;
  assign n16356 = n16262 ^ n16041 ;
  assign n16365 = n16364 ^ n16356 ;
  assign n16376 = ~n12251 & n13433 ;
  assign n16374 = n5426 & n12339 ;
  assign n16367 = n12249 ^ x20 ;
  assign n16368 = n16367 ^ x19 ;
  assign n16369 = n16368 ^ n12249 ;
  assign n16370 = ~n14194 & n16369 ;
  assign n16371 = n16370 ^ n12249 ;
  assign n16372 = n5215 & ~n16371 ;
  assign n16373 = n16372 ^ x20 ;
  assign n16375 = n16374 ^ n16373 ;
  assign n16377 = n16376 ^ n16375 ;
  assign n16366 = n16259 ^ n16051 ;
  assign n16378 = n16377 ^ n16366 ;
  assign n16651 = n16256 ^ n16061 ;
  assign n16389 = n12331 & n13433 ;
  assign n16387 = n5426 & n12253 ;
  assign n16380 = n12251 ^ x20 ;
  assign n16381 = n16380 ^ x19 ;
  assign n16382 = n16381 ^ n12251 ;
  assign n16383 = ~n13676 & n16382 ;
  assign n16384 = n16383 ^ n12251 ;
  assign n16385 = n5215 & ~n16384 ;
  assign n16386 = n16385 ^ x20 ;
  assign n16388 = n16387 ^ n16386 ;
  assign n16390 = n16389 ^ n16388 ;
  assign n16379 = n16253 ^ n16071 ;
  assign n16391 = n16390 ^ n16379 ;
  assign n16633 = n16250 ^ n16081 ;
  assign n16396 = n5215 & ~n14414 ;
  assign n16395 = n5220 & ~n14088 ;
  assign n16397 = n16396 ^ n16395 ;
  assign n16393 = n5426 & n12331 ;
  assign n16392 = n12257 & n13433 ;
  assign n16394 = n16393 ^ n16392 ;
  assign n16398 = n16397 ^ n16394 ;
  assign n16634 = n16633 ^ n16398 ;
  assign n16418 = n12264 & n13433 ;
  assign n16416 = n5426 & ~n12258 ;
  assign n16409 = n12257 ^ x20 ;
  assign n16410 = n16409 ^ x19 ;
  assign n16411 = n16410 ^ n12257 ;
  assign n16412 = ~n14019 & n16411 ;
  assign n16413 = n16412 ^ n12257 ;
  assign n16414 = n5215 & n16413 ;
  assign n16415 = n16414 ^ x20 ;
  assign n16417 = n16416 ^ n16415 ;
  assign n16419 = n16418 ^ n16417 ;
  assign n16408 = n16244 ^ n16101 ;
  assign n16420 = n16419 ^ n16408 ;
  assign n16617 = ~n12267 & n13433 ;
  assign n16615 = n5426 & n12264 ;
  assign n16608 = n12258 ^ x20 ;
  assign n16609 = n16608 ^ x19 ;
  assign n16610 = n16609 ^ n12258 ;
  assign n16611 = ~n14242 & n16610 ;
  assign n16612 = n16611 ^ n12258 ;
  assign n16613 = n5215 & ~n16612 ;
  assign n16614 = n16613 ^ x20 ;
  assign n16616 = n16615 ^ n16614 ;
  assign n16618 = n16617 ^ n16616 ;
  assign n16428 = n5426 & ~n12267 ;
  assign n16426 = n5220 & n12264 ;
  assign n16423 = n5221 & ~n14429 ;
  assign n16422 = n12268 & n13433 ;
  assign n16424 = n16423 ^ n16422 ;
  assign n16425 = n16424 ^ x20 ;
  assign n16427 = n16426 ^ n16425 ;
  assign n16429 = n16428 ^ n16427 ;
  assign n16421 = n16226 ^ n16217 ;
  assign n16430 = n16429 ^ n16421 ;
  assign n16442 = n5426 & n12268 ;
  assign n16440 = ~n12276 & n13433 ;
  assign n16433 = n12267 ^ x20 ;
  assign n16434 = n16433 ^ x19 ;
  assign n16435 = n16434 ^ n12267 ;
  assign n16436 = ~n14450 & n16435 ;
  assign n16437 = n16436 ^ n12267 ;
  assign n16438 = n5215 & ~n16437 ;
  assign n16439 = n16438 ^ x20 ;
  assign n16441 = n16440 ^ n16439 ;
  assign n16443 = n16442 ^ n16441 ;
  assign n16431 = n16212 ^ n16115 ;
  assign n16444 = n16443 ^ n16431 ;
  assign n16455 = n12279 & n13433 ;
  assign n16453 = n5426 & ~n12276 ;
  assign n16446 = n12268 ^ x20 ;
  assign n16447 = n16446 ^ x19 ;
  assign n16448 = n16447 ^ n12268 ;
  assign n16449 = ~n14328 & n16448 ;
  assign n16450 = n16449 ^ n12268 ;
  assign n16451 = n5215 & n16450 ;
  assign n16452 = n16451 ^ x20 ;
  assign n16454 = n16453 ^ n16452 ;
  assign n16456 = n16455 ^ n16454 ;
  assign n16445 = n16210 ^ n16116 ;
  assign n16457 = n16456 ^ n16445 ;
  assign n16468 = ~n12283 & n13433 ;
  assign n16466 = n5426 & n12279 ;
  assign n16459 = n12276 ^ x20 ;
  assign n16460 = n16459 ^ x19 ;
  assign n16461 = n16460 ^ n12276 ;
  assign n16462 = ~n14465 & n16461 ;
  assign n16463 = n16462 ^ n12276 ;
  assign n16464 = n5215 & ~n16463 ;
  assign n16465 = n16464 ^ x20 ;
  assign n16467 = n16466 ^ n16465 ;
  assign n16469 = n16468 ^ n16467 ;
  assign n16458 = n16207 ^ n16139 ;
  assign n16470 = n16469 ^ n16458 ;
  assign n16481 = ~n12284 & n13433 ;
  assign n16479 = n5426 & ~n12283 ;
  assign n16472 = n12279 ^ x20 ;
  assign n16473 = n16472 ^ x19 ;
  assign n16474 = n16473 ^ n12279 ;
  assign n16475 = ~n14514 & n16474 ;
  assign n16476 = n16475 ^ n12279 ;
  assign n16477 = n5215 & n16476 ;
  assign n16478 = n16477 ^ x20 ;
  assign n16480 = n16479 ^ n16478 ;
  assign n16482 = n16481 ^ n16480 ;
  assign n16471 = n16204 ^ n16150 ;
  assign n16483 = n16482 ^ n16471 ;
  assign n16494 = ~n12285 & n13433 ;
  assign n16492 = n5426 & ~n12284 ;
  assign n16485 = n12283 ^ x20 ;
  assign n16486 = n16485 ^ x19 ;
  assign n16487 = n16486 ^ n12283 ;
  assign n16488 = ~n14547 & n16487 ;
  assign n16489 = n16488 ^ n12283 ;
  assign n16490 = n5215 & ~n16489 ;
  assign n16491 = n16490 ^ x20 ;
  assign n16493 = n16492 ^ n16491 ;
  assign n16495 = n16494 ^ n16493 ;
  assign n16484 = n16201 ^ n16193 ;
  assign n16496 = n16495 ^ n16484 ;
  assign n16507 = n5426 & ~n12285 ;
  assign n16505 = n12313 & n13433 ;
  assign n16498 = n12284 ^ x20 ;
  assign n16499 = n16498 ^ x19 ;
  assign n16500 = n16499 ^ n12284 ;
  assign n16501 = ~n14583 & n16500 ;
  assign n16502 = n16501 ^ n12284 ;
  assign n16503 = n5215 & ~n16502 ;
  assign n16504 = n16503 ^ x20 ;
  assign n16506 = n16505 ^ n16504 ;
  assign n16508 = n16507 ^ n16506 ;
  assign n16497 = n16189 ^ n16185 ;
  assign n16509 = n16508 ^ n16497 ;
  assign n16521 = n12289 & n13433 ;
  assign n16519 = n5426 & n12313 ;
  assign n16512 = n12285 ^ x20 ;
  assign n16513 = n16512 ^ x19 ;
  assign n16514 = n16513 ^ n12285 ;
  assign n16515 = ~n14651 & n16514 ;
  assign n16516 = n16515 ^ n12285 ;
  assign n16517 = n5215 & ~n16516 ;
  assign n16518 = n16517 ^ x20 ;
  assign n16520 = n16519 ^ n16518 ;
  assign n16522 = n16521 ^ n16520 ;
  assign n16510 = n16166 ^ n16151 ;
  assign n16511 = n16510 ^ n16175 ;
  assign n16523 = n16522 ^ n16511 ;
  assign n16157 = n16156 ^ x23 ;
  assign n16571 = n16165 ^ n16157 ;
  assign n16563 = n12293 & n13433 ;
  assign n16561 = n5426 & ~n12290 ;
  assign n16554 = n12289 ^ x20 ;
  assign n16555 = n16554 ^ x19 ;
  assign n16556 = n16555 ^ n12289 ;
  assign n16557 = ~n14748 & n16556 ;
  assign n16558 = n16557 ^ n12289 ;
  assign n16559 = n5215 & n16558 ;
  assign n16560 = n16559 ^ x20 ;
  assign n16562 = n16561 ^ n16560 ;
  assign n16564 = n16563 ^ n16562 ;
  assign n16524 = n35 & n12291 ;
  assign n16525 = n5215 & n12292 ;
  assign n16526 = x20 & ~n16525 ;
  assign n16527 = n12291 & n16526 ;
  assign n16528 = n8316 & n16527 ;
  assign n16529 = n16528 ^ n16526 ;
  assign n16536 = n5221 & ~n15423 ;
  assign n16535 = n5426 & n12292 ;
  assign n16537 = n16536 ^ n16535 ;
  assign n16533 = n5220 & n12293 ;
  assign n16532 = n12291 & n13433 ;
  assign n16534 = n16533 ^ n16532 ;
  assign n16538 = n16537 ^ n16534 ;
  assign n16539 = n16529 & ~n16538 ;
  assign n16540 = ~n16524 & ~n16539 ;
  assign n16550 = n12292 & n13433 ;
  assign n16548 = n5426 & n12293 ;
  assign n16541 = n12290 ^ x20 ;
  assign n16542 = n16541 ^ x19 ;
  assign n16543 = n16542 ^ n12290 ;
  assign n16544 = n12297 & n16543 ;
  assign n16545 = n16544 ^ n12290 ;
  assign n16546 = n5215 & ~n16545 ;
  assign n16547 = n16546 ^ x20 ;
  assign n16549 = n16548 ^ n16547 ;
  assign n16551 = n16550 ^ n16549 ;
  assign n16552 = n16540 & n16551 ;
  assign n16553 = n16552 ^ n16551 ;
  assign n16565 = n16564 ^ n16553 ;
  assign n16567 = n16553 ^ n16152 ;
  assign n16566 = ~n8289 & n12291 ;
  assign n16568 = n16567 ^ n16566 ;
  assign n16569 = n16565 & ~n16568 ;
  assign n16570 = n16569 ^ n16564 ;
  assign n16572 = n16571 ^ n16570 ;
  assign n16577 = n5221 & ~n14712 ;
  assign n16576 = ~n12290 & n13433 ;
  assign n16578 = n16577 ^ n16576 ;
  assign n16574 = n5220 & n12313 ;
  assign n16573 = n5426 & n12289 ;
  assign n16575 = n16574 ^ n16573 ;
  assign n16579 = n16578 ^ n16575 ;
  assign n16580 = n16579 ^ x20 ;
  assign n16581 = n16580 ^ n16570 ;
  assign n16582 = n16572 & ~n16581 ;
  assign n16583 = n16582 ^ n16571 ;
  assign n16584 = n16583 ^ n16522 ;
  assign n16585 = n16523 & n16584 ;
  assign n16586 = n16585 ^ n16522 ;
  assign n16587 = n16586 ^ n16508 ;
  assign n16588 = n16509 & n16587 ;
  assign n16589 = n16588 ^ n16508 ;
  assign n16590 = n16589 ^ n16495 ;
  assign n16591 = n16496 & n16590 ;
  assign n16592 = n16591 ^ n16495 ;
  assign n16593 = n16592 ^ n16482 ;
  assign n16594 = n16483 & n16593 ;
  assign n16595 = n16594 ^ n16482 ;
  assign n16596 = n16595 ^ n16469 ;
  assign n16597 = n16470 & n16596 ;
  assign n16598 = n16597 ^ n16469 ;
  assign n16599 = n16598 ^ n16456 ;
  assign n16600 = n16457 & n16599 ;
  assign n16601 = n16600 ^ n16456 ;
  assign n16602 = n16601 ^ n16443 ;
  assign n16603 = n16444 & n16602 ;
  assign n16604 = n16603 ^ n16443 ;
  assign n16605 = n16604 ^ n16429 ;
  assign n16606 = n16430 & n16605 ;
  assign n16607 = n16606 ^ n16429 ;
  assign n16619 = n16618 ^ n16607 ;
  assign n16622 = n16618 ^ n16236 ;
  assign n16620 = n16226 ^ n16215 ;
  assign n16621 = ~n16217 & n16620 ;
  assign n16623 = n16622 ^ n16621 ;
  assign n16624 = n16619 & n16623 ;
  assign n16625 = n16624 ^ n16618 ;
  assign n16626 = n16625 ^ n16419 ;
  assign n16627 = n16420 & n16626 ;
  assign n16628 = n16627 ^ n16419 ;
  assign n16407 = n16247 ^ n16091 ;
  assign n16629 = n16628 ^ n16407 ;
  assign n16641 = n16407 ^ n16398 ;
  assign n16403 = n5215 & ~n14972 ;
  assign n16402 = n5220 & ~n14219 ;
  assign n16404 = n16403 ^ n16402 ;
  assign n16400 = n5426 & n12257 ;
  assign n16399 = ~n12258 & n13433 ;
  assign n16401 = n16400 ^ n16399 ;
  assign n16405 = n16404 ^ n16401 ;
  assign n16406 = n16405 ^ n16398 ;
  assign n16642 = n16641 ^ n16406 ;
  assign n16643 = n16629 & ~n16642 ;
  assign n16644 = n16643 ^ n16406 ;
  assign n16645 = ~n16634 & n16644 ;
  assign n16646 = n16645 ^ n16398 ;
  assign n16635 = n16634 ^ n16405 ;
  assign n16632 = n16628 ^ n16406 ;
  assign n16636 = n16635 ^ n16632 ;
  assign n16637 = n16636 ^ n16406 ;
  assign n16638 = n16629 & n16637 ;
  assign n16639 = n16638 ^ n16406 ;
  assign n16640 = x20 & ~n16639 ;
  assign n16647 = n16646 ^ n16640 ;
  assign n16648 = n16647 ^ n16390 ;
  assign n16649 = ~n16391 & n16648 ;
  assign n16650 = n16649 ^ n16390 ;
  assign n16652 = n16651 ^ n16650 ;
  assign n16662 = n12253 & n13433 ;
  assign n16660 = n5426 & ~n12251 ;
  assign n16658 = n16651 ^ x20 ;
  assign n16653 = n13885 ^ n5224 ;
  assign n16654 = n16653 ^ n13885 ;
  assign n16655 = ~n14922 & ~n16654 ;
  assign n16656 = n16655 ^ n13885 ;
  assign n16657 = n5215 & ~n16656 ;
  assign n16659 = n16658 ^ n16657 ;
  assign n16661 = n16660 ^ n16659 ;
  assign n16663 = n16662 ^ n16661 ;
  assign n16664 = ~n16652 & ~n16663 ;
  assign n16665 = n16664 ^ n16651 ;
  assign n16666 = n16665 ^ n16377 ;
  assign n16667 = ~n16378 & ~n16666 ;
  assign n16668 = n16667 ^ n16377 ;
  assign n16669 = n16668 ^ n16364 ;
  assign n16670 = ~n16365 & n16669 ;
  assign n16671 = n16670 ^ n16364 ;
  assign n16672 = n16671 ^ n16349 ;
  assign n16673 = n16355 & n16672 ;
  assign n16674 = n16673 ^ n16349 ;
  assign n16337 = n6148 & ~n12382 ;
  assign n16336 = n6143 & ~n12228 ;
  assign n16338 = n16337 ^ n16336 ;
  assign n16339 = n16338 ^ x17 ;
  assign n16335 = n6163 & n13445 ;
  assign n16340 = n16339 ^ n16335 ;
  assign n16334 = n12229 & n20437 ;
  assign n16341 = n16340 ^ n16334 ;
  assign n16333 = n16268 ^ n16021 ;
  assign n16342 = n16341 ^ n16333 ;
  assign n17057 = n16674 ^ n16342 ;
  assign n16732 = n12235 & n20437 ;
  assign n16729 = n6143 & n12229 ;
  assign n16727 = n6148 & ~n12228 ;
  assign n16725 = n16671 ^ n16355 ;
  assign n16726 = n16725 ^ x17 ;
  assign n16728 = n16727 ^ n16726 ;
  assign n16730 = n16729 ^ n16728 ;
  assign n16724 = n6163 & n13779 ;
  assign n16731 = n16730 ^ n16724 ;
  assign n16733 = n16732 ^ n16731 ;
  assign n16742 = ~n12239 & n20437 ;
  assign n16737 = n16668 ^ n16365 ;
  assign n16738 = n16737 ^ x17 ;
  assign n16736 = n6148 & n12229 ;
  assign n16739 = n16738 ^ n16736 ;
  assign n16735 = n6143 & n12235 ;
  assign n16740 = n16739 ^ n16735 ;
  assign n16734 = n6163 & ~n12867 ;
  assign n16741 = n16740 ^ n16734 ;
  assign n16743 = n16742 ^ n16741 ;
  assign n16750 = ~x16 & ~n13339 ;
  assign n16753 = n16750 ^ n13343 ;
  assign n16754 = n6147 & n16753 ;
  assign n16747 = n6143 & n12248 ;
  assign n16746 = ~n12249 & n20437 ;
  assign n16748 = n16747 ^ n16746 ;
  assign n16749 = n16748 ^ x17 ;
  assign n16751 = n16750 ^ n12239 ;
  assign n16752 = n16749 & n16751 ;
  assign n16755 = n16754 ^ n16752 ;
  assign n16756 = n16748 ^ n6145 ;
  assign n16757 = ~n16755 & ~n16756 ;
  assign n16745 = n16663 ^ n16650 ;
  assign n16758 = n16757 ^ n16745 ;
  assign n16763 = n6148 & n12248 ;
  assign n16762 = n6143 & ~n12249 ;
  assign n16764 = n16763 ^ n16762 ;
  assign n16765 = n16764 ^ x17 ;
  assign n16761 = n6163 & ~n13519 ;
  assign n16766 = n16765 ^ n16761 ;
  assign n16760 = n12339 & n20437 ;
  assign n16767 = n16766 ^ n16760 ;
  assign n16759 = n16647 ^ n16391 ;
  assign n16768 = n16767 ^ n16759 ;
  assign n16775 = n6148 & ~n12249 ;
  assign n16774 = n6143 & n12339 ;
  assign n16776 = n16775 ^ n16774 ;
  assign n16777 = n16776 ^ x17 ;
  assign n16773 = n6163 & n13554 ;
  assign n16778 = n16777 ^ n16773 ;
  assign n16772 = ~n12251 & n20437 ;
  assign n16779 = n16778 ^ n16772 ;
  assign n16780 = n16779 ^ n16635 ;
  assign n16769 = n16628 ^ x20 ;
  assign n16770 = n16769 ^ n16405 ;
  assign n16771 = n16629 & n16770 ;
  assign n16781 = n16780 ^ n16771 ;
  assign n16791 = n12253 & n20437 ;
  assign n16789 = n6163 & ~n13885 ;
  assign n16786 = n6148 & n12339 ;
  assign n16785 = n6143 & ~n12251 ;
  assign n16787 = n16786 ^ n16785 ;
  assign n16788 = n16787 ^ x17 ;
  assign n16790 = n16789 ^ n16788 ;
  assign n16792 = n16791 ^ n16790 ;
  assign n16782 = n16407 ^ x20 ;
  assign n16783 = n16782 ^ n16405 ;
  assign n16784 = n16783 ^ n16628 ;
  assign n16793 = n16792 ^ n16784 ;
  assign n16798 = n6148 & ~n12251 ;
  assign n16797 = n6143 & n12253 ;
  assign n16799 = n16798 ^ n16797 ;
  assign n16800 = n16799 ^ x17 ;
  assign n16796 = n6163 & n13677 ;
  assign n16801 = n16800 ^ n16796 ;
  assign n16795 = n12331 & n20437 ;
  assign n16802 = n16801 ^ n16795 ;
  assign n16794 = n16625 ^ n16420 ;
  assign n16803 = n16802 ^ n16794 ;
  assign n16808 = n6148 & n12253 ;
  assign n16807 = n6143 & n12331 ;
  assign n16809 = n16808 ^ n16807 ;
  assign n16810 = n16809 ^ x17 ;
  assign n16806 = n6163 & ~n14414 ;
  assign n16811 = n16810 ^ n16806 ;
  assign n16805 = n12257 & n20437 ;
  assign n16812 = n16811 ^ n16805 ;
  assign n16804 = n16623 ^ n16607 ;
  assign n16813 = n16812 ^ n16804 ;
  assign n16821 = ~n12258 & n20437 ;
  assign n16819 = n6163 & ~n14972 ;
  assign n16816 = n6148 & n12331 ;
  assign n16815 = n6143 & n12257 ;
  assign n16817 = n16816 ^ n16815 ;
  assign n16818 = n16817 ^ x17 ;
  assign n16820 = n16819 ^ n16818 ;
  assign n16822 = n16821 ^ n16820 ;
  assign n16814 = n16604 ^ n16430 ;
  assign n16823 = n16822 ^ n16814 ;
  assign n16831 = n12264 & n20437 ;
  assign n16829 = n6163 & ~n14020 ;
  assign n16826 = n6148 & n12257 ;
  assign n16825 = n6143 & ~n12258 ;
  assign n16827 = n16826 ^ n16825 ;
  assign n16828 = n16827 ^ x17 ;
  assign n16830 = n16829 ^ n16828 ;
  assign n16832 = n16831 ^ n16830 ;
  assign n16824 = n16601 ^ n16444 ;
  assign n16833 = n16832 ^ n16824 ;
  assign n16841 = ~n12267 & n20437 ;
  assign n16839 = n6163 & n14243 ;
  assign n16836 = n6148 & ~n12258 ;
  assign n16835 = n6143 & n12264 ;
  assign n16837 = n16836 ^ n16835 ;
  assign n16838 = n16837 ^ x17 ;
  assign n16840 = n16839 ^ n16838 ;
  assign n16842 = n16841 ^ n16840 ;
  assign n16834 = n16598 ^ n16457 ;
  assign n16843 = n16842 ^ n16834 ;
  assign n16852 = n6143 & ~n12267 ;
  assign n16851 = n12268 & n20437 ;
  assign n16853 = n16852 ^ n16851 ;
  assign n16854 = n16853 ^ x17 ;
  assign n16845 = ~x16 & ~n14428 ;
  assign n16848 = n16845 ^ n12264 ;
  assign n16850 = n16848 & n16849 ;
  assign n16855 = n16854 ^ n16850 ;
  assign n16846 = n16845 ^ n14429 ;
  assign n16847 = n6147 & ~n16846 ;
  assign n16856 = n16855 ^ n16847 ;
  assign n16844 = n16595 ^ n16470 ;
  assign n16857 = n16856 ^ n16844 ;
  assign n16863 = n6143 & ~n12276 ;
  assign n16862 = n6148 & n12268 ;
  assign n16864 = n16863 ^ n16862 ;
  assign n16865 = n16864 ^ x17 ;
  assign n16861 = n6163 & ~n14329 ;
  assign n16866 = n16865 ^ n16861 ;
  assign n16860 = n12279 & n20437 ;
  assign n16867 = n16866 ^ n16860 ;
  assign n16859 = n16589 ^ n16496 ;
  assign n16868 = n16867 ^ n16859 ;
  assign n16876 = ~n12283 & n20437 ;
  assign n16874 = n6163 & n14475 ;
  assign n16871 = n6148 & ~n12276 ;
  assign n16870 = n6143 & n12279 ;
  assign n16872 = n16871 ^ n16870 ;
  assign n16873 = n16872 ^ x17 ;
  assign n16875 = n16874 ^ n16873 ;
  assign n16877 = n16876 ^ n16875 ;
  assign n16869 = n16586 ^ n16509 ;
  assign n16878 = n16877 ^ n16869 ;
  assign n16883 = n6148 & n12279 ;
  assign n16882 = n6143 & ~n12283 ;
  assign n16884 = n16883 ^ n16882 ;
  assign n16885 = n16884 ^ x17 ;
  assign n16881 = n6163 & ~n14528 ;
  assign n16886 = n16885 ^ n16881 ;
  assign n16880 = ~n12284 & n20437 ;
  assign n16887 = n16886 ^ n16880 ;
  assign n16879 = n16583 ^ n16523 ;
  assign n16888 = n16887 ^ n16879 ;
  assign n16901 = ~n12285 & n20437 ;
  assign n16899 = n6143 & ~n12284 ;
  assign n16892 = n12283 ^ x17 ;
  assign n16893 = n16892 ^ x16 ;
  assign n16894 = n16893 ^ n12283 ;
  assign n16895 = ~n14547 & n16894 ;
  assign n16896 = n16895 ^ n12283 ;
  assign n16897 = n6141 & ~n16896 ;
  assign n16898 = n16897 ^ x17 ;
  assign n16900 = n16899 ^ n16898 ;
  assign n16902 = n16901 ^ n16900 ;
  assign n16889 = n16571 ^ x20 ;
  assign n16890 = n16889 ^ n16579 ;
  assign n16891 = n16890 ^ n16570 ;
  assign n16903 = n16902 ^ n16891 ;
  assign n16908 = n6148 & ~n12284 ;
  assign n16907 = n6143 & ~n12285 ;
  assign n16909 = n16908 ^ n16907 ;
  assign n16910 = n16909 ^ x17 ;
  assign n16906 = n6163 & n14584 ;
  assign n16911 = n16910 ^ n16906 ;
  assign n16905 = n12313 & n20437 ;
  assign n16912 = n16911 ^ n16905 ;
  assign n16904 = n16568 ^ n16564 ;
  assign n16913 = n16912 ^ n16904 ;
  assign n16919 = n6143 & n12313 ;
  assign n16918 = n6148 & ~n12285 ;
  assign n16920 = n16919 ^ n16918 ;
  assign n16921 = n16920 ^ x17 ;
  assign n16917 = n6163 & n14652 ;
  assign n16922 = n16921 ^ n16917 ;
  assign n16916 = n12289 & n20437 ;
  assign n16923 = n16922 ^ n16916 ;
  assign n16914 = n16539 ^ n16524 ;
  assign n16915 = n16914 ^ n16551 ;
  assign n16924 = n16923 ^ n16915 ;
  assign n16931 = n6163 & ~n14785 ;
  assign n16930 = n12292 & n20437 ;
  assign n16932 = n16931 ^ n16930 ;
  assign n16928 = n6148 & ~n12290 ;
  assign n16927 = n6143 & n12293 ;
  assign n16929 = n16928 ^ n16927 ;
  assign n16933 = n16932 ^ n16929 ;
  assign n16935 = n5215 & n12291 ;
  assign n16934 = n5212 & n12291 ;
  assign n16936 = n16935 ^ n16934 ;
  assign n16937 = n6154 & ~n12298 ;
  assign n16940 = n6163 & ~n15423 ;
  assign n16939 = n12291 & n20437 ;
  assign n16941 = n16940 ^ n16939 ;
  assign n16938 = n6148 & n12293 ;
  assign n16942 = n16941 ^ n16938 ;
  assign n16943 = x17 & ~n16942 ;
  assign n16944 = n16937 & n16943 ;
  assign n16945 = n16944 ^ n16943 ;
  assign n16948 = ~n16936 & n16945 ;
  assign n16949 = n16948 ^ n16935 ;
  assign n16950 = ~n16933 & n16949 ;
  assign n16951 = n16950 ^ n16934 ;
  assign n16952 = n16951 ^ n16525 ;
  assign n16926 = n8563 & n12291 ;
  assign n16953 = n16952 ^ n16926 ;
  assign n16957 = n6148 & n12289 ;
  assign n16956 = n6143 & ~n12290 ;
  assign n16958 = n16957 ^ n16956 ;
  assign n16959 = n16958 ^ x17 ;
  assign n16955 = n6163 & ~n14749 ;
  assign n16960 = n16959 ^ n16955 ;
  assign n16954 = n12293 & n20437 ;
  assign n16961 = n16960 ^ n16954 ;
  assign n16962 = n16961 ^ n16951 ;
  assign n16963 = n16953 & n16962 ;
  assign n16964 = n16963 ^ n16951 ;
  assign n16530 = n16529 ^ x20 ;
  assign n16925 = n16538 ^ n16530 ;
  assign n16965 = n16964 ^ n16925 ;
  assign n16972 = n6163 & ~n14712 ;
  assign n16970 = n6148 & n12313 ;
  assign n16968 = n6143 & n12289 ;
  assign n16967 = n16925 ^ x17 ;
  assign n16969 = n16968 ^ n16967 ;
  assign n16971 = n16970 ^ n16969 ;
  assign n16973 = n16972 ^ n16971 ;
  assign n16966 = ~n12290 & n20437 ;
  assign n16974 = n16973 ^ n16966 ;
  assign n16975 = n16965 & ~n16974 ;
  assign n16976 = n16975 ^ n16964 ;
  assign n16977 = n16976 ^ n16923 ;
  assign n16978 = n16924 & n16977 ;
  assign n16979 = n16978 ^ n16923 ;
  assign n16980 = n16979 ^ n16912 ;
  assign n16981 = n16913 & n16980 ;
  assign n16982 = n16981 ^ n16912 ;
  assign n16983 = n16982 ^ n16902 ;
  assign n16984 = n16903 & n16983 ;
  assign n16985 = n16984 ^ n16902 ;
  assign n16986 = n16985 ^ n16887 ;
  assign n16987 = n16888 & n16986 ;
  assign n16988 = n16987 ^ n16887 ;
  assign n16989 = n16988 ^ n16877 ;
  assign n16990 = n16878 & n16989 ;
  assign n16991 = n16990 ^ n16877 ;
  assign n16992 = n16991 ^ n16867 ;
  assign n16993 = n16868 & n16992 ;
  assign n16994 = n16993 ^ n16867 ;
  assign n16858 = n16592 ^ n16483 ;
  assign n16995 = n16994 ^ n16858 ;
  assign n17002 = ~n12276 & n20437 ;
  assign n17001 = n6143 & n12268 ;
  assign n17003 = n17002 ^ n17001 ;
  assign n17004 = n17003 ^ x17 ;
  assign n16996 = n14154 ^ n12267 ;
  assign n16997 = n16996 ^ n12267 ;
  assign n16998 = ~n14450 & n16997 ;
  assign n16999 = n16998 ^ n12267 ;
  assign n17000 = n6141 & ~n16999 ;
  assign n17005 = n17004 ^ n17000 ;
  assign n17006 = n17005 ^ n16858 ;
  assign n17007 = n16995 & ~n17006 ;
  assign n17008 = n17007 ^ n16994 ;
  assign n17009 = n17008 ^ n16844 ;
  assign n17010 = n16857 & ~n17009 ;
  assign n17011 = n17010 ^ n16856 ;
  assign n17012 = n17011 ^ n16842 ;
  assign n17013 = n16843 & n17012 ;
  assign n17014 = n17013 ^ n16842 ;
  assign n17015 = n17014 ^ n16832 ;
  assign n17016 = n16833 & n17015 ;
  assign n17017 = n17016 ^ n16832 ;
  assign n17018 = n17017 ^ n16822 ;
  assign n17019 = n16823 & n17018 ;
  assign n17020 = n17019 ^ n16822 ;
  assign n17021 = n17020 ^ n16812 ;
  assign n17022 = n16813 & n17021 ;
  assign n17023 = n17022 ^ n16812 ;
  assign n17024 = n17023 ^ n16802 ;
  assign n17025 = n16803 & n17024 ;
  assign n17026 = n17025 ^ n16802 ;
  assign n17027 = n17026 ^ n16792 ;
  assign n17028 = ~n16793 & n17027 ;
  assign n17029 = n17028 ^ n16792 ;
  assign n17030 = n17029 ^ n16779 ;
  assign n17031 = ~n16781 & n17030 ;
  assign n17032 = n17031 ^ n16779 ;
  assign n17033 = n17032 ^ n16767 ;
  assign n17034 = ~n16768 & n17033 ;
  assign n17035 = n17034 ^ n16767 ;
  assign n17036 = n17035 ^ n16757 ;
  assign n17037 = n16758 & ~n17036 ;
  assign n17038 = n17037 ^ n16757 ;
  assign n16744 = n16665 ^ n16378 ;
  assign n17039 = n17038 ^ n16744 ;
  assign n17047 = n12248 & n20437 ;
  assign n17043 = n16744 ^ x17 ;
  assign n17042 = n6148 & n12235 ;
  assign n17044 = n17043 ^ n17042 ;
  assign n17041 = n6143 & ~n12239 ;
  assign n17045 = n17044 ^ n17041 ;
  assign n17040 = n6163 & ~n13329 ;
  assign n17046 = n17045 ^ n17040 ;
  assign n17048 = n17047 ^ n17046 ;
  assign n17049 = ~n17039 & ~n17048 ;
  assign n17050 = n17049 ^ n17038 ;
  assign n17051 = n17050 ^ n16737 ;
  assign n17052 = ~n16743 & n17051 ;
  assign n17053 = n17052 ^ n16737 ;
  assign n17054 = n17053 ^ n16725 ;
  assign n17055 = n16733 & ~n17054 ;
  assign n17056 = n17055 ^ n16725 ;
  assign n17058 = n17057 ^ n17056 ;
  assign n16690 = ~n6529 & n12222 ;
  assign n16688 = ~n6547 & n12380 ;
  assign n16682 = n15967 ^ x13 ;
  assign n16683 = n16682 ^ n12214 ;
  assign n16684 = ~n12607 & n16683 ;
  assign n16685 = n16684 ^ n12214 ;
  assign n16686 = n6391 & ~n16685 ;
  assign n16687 = n16686 ^ x14 ;
  assign n16689 = n16688 ^ n16687 ;
  assign n16691 = n16690 ^ n16689 ;
  assign n16675 = n16674 ^ n16341 ;
  assign n16676 = ~n16342 & n16675 ;
  assign n16677 = n16676 ^ n16341 ;
  assign n16332 = n16281 ^ n16272 ;
  assign n16678 = n16677 ^ n16332 ;
  assign n17719 = n16691 ^ n16678 ;
  assign n16717 = ~x13 & n12390 ;
  assign n16718 = n16717 ^ n12222 ;
  assign n16721 = n16718 ^ n12390 ;
  assign n16722 = n6539 & n16721 ;
  assign n16719 = n6537 & n16718 ;
  assign n16714 = ~n6529 & n12380 ;
  assign n16713 = ~n6547 & n12376 ;
  assign n16715 = n16714 ^ n16713 ;
  assign n16716 = n16715 ^ x14 ;
  assign n16720 = n16719 ^ n16716 ;
  assign n16723 = n16722 ^ n16720 ;
  assign n17720 = n17719 ^ n16723 ;
  assign n17721 = n17720 ^ n17719 ;
  assign n17722 = n17721 ^ n17056 ;
  assign n17723 = n17058 & n17722 ;
  assign n17724 = n17723 ^ n17720 ;
  assign n17733 = n17732 ^ n17724 ;
  assign n17069 = n7148 & ~n12214 ;
  assign n17067 = n7142 & ~n12400 ;
  assign n17060 = n12210 ^ x11 ;
  assign n17061 = n17060 ^ x10 ;
  assign n17062 = n17061 ^ n12210 ;
  assign n17063 = ~n12736 & n17062 ;
  assign n17064 = n17063 ^ n12210 ;
  assign n17065 = n7140 & ~n17064 ;
  assign n17066 = n17065 ^ x11 ;
  assign n17068 = n17067 ^ n17066 ;
  assign n17070 = n17069 ^ n17068 ;
  assign n17059 = n17058 ^ n16723 ;
  assign n17071 = n17070 ^ n17059 ;
  assign n17088 = n17053 ^ n16733 ;
  assign n17073 = ~n6529 & n12376 ;
  assign n17072 = ~n6547 & ~n12382 ;
  assign n17074 = n17073 ^ n17072 ;
  assign n17075 = n17074 ^ n6537 ;
  assign n17076 = n17075 ^ x14 ;
  assign n17085 = n6539 & ~n12554 ;
  assign n17077 = n17074 ^ n6538 ;
  assign n17079 = n12555 ^ n12380 ;
  assign n17080 = n12380 ^ x13 ;
  assign n17081 = n17080 ^ n12380 ;
  assign n17082 = n17079 & ~n17081 ;
  assign n17083 = n17082 ^ n12380 ;
  assign n17084 = n17077 & ~n17083 ;
  assign n17086 = n17085 ^ n17084 ;
  assign n17087 = ~n17076 & ~n17086 ;
  assign n17089 = n17088 ^ n17087 ;
  assign n17092 = ~n6529 & ~n12382 ;
  assign n17091 = ~n6547 & ~n12228 ;
  assign n17093 = n17092 ^ n17091 ;
  assign n17094 = n17093 ^ n6537 ;
  assign n17095 = n17094 ^ x14 ;
  assign n17105 = x13 & ~n12928 ;
  assign n17104 = n8856 & n12376 ;
  assign n17106 = n17105 ^ n17104 ;
  assign n17107 = ~n6539 & n17106 ;
  assign n17102 = n12553 ^ n8856 ;
  assign n17096 = n17093 ^ x14 ;
  assign n17097 = n12376 ^ x13 ;
  assign n17098 = n17097 ^ n12376 ;
  assign n17099 = n12553 & ~n17098 ;
  assign n17100 = n17099 ^ n12376 ;
  assign n17101 = ~n17096 & ~n17100 ;
  assign n17103 = n17102 ^ n17101 ;
  assign n17108 = n17107 ^ n17103 ;
  assign n17109 = ~n17095 & ~n17108 ;
  assign n17090 = n17050 ^ n16743 ;
  assign n17110 = n17109 ^ n17090 ;
  assign n17134 = n17048 ^ n17038 ;
  assign n17112 = ~n6529 & ~n12228 ;
  assign n17111 = ~n6547 & n12229 ;
  assign n17113 = n17112 ^ n17111 ;
  assign n17114 = n17113 ^ n6537 ;
  assign n17115 = n17114 ^ x14 ;
  assign n17116 = n12382 ^ x13 ;
  assign n17117 = n17116 ^ n6539 ;
  assign n17118 = n17117 ^ n12382 ;
  assign n17119 = n12370 & ~n17118 ;
  assign n17120 = n17119 ^ n17116 ;
  assign n17121 = n17113 ^ x14 ;
  assign n17122 = n17121 ^ n12552 ;
  assign n17123 = n17122 ^ n17121 ;
  assign n17125 = n17121 ^ n17113 ;
  assign n17128 = n6391 & ~n17125 ;
  assign n17129 = ~n17123 & n17128 ;
  assign n17130 = n17129 ^ n17123 ;
  assign n17131 = n17130 ^ n17122 ;
  assign n17132 = ~n17120 & n17131 ;
  assign n17133 = ~n17115 & ~n17132 ;
  assign n17135 = n17134 ^ n17133 ;
  assign n17146 = n17035 ^ n16758 ;
  assign n17142 = ~n6529 & n12229 ;
  assign n17141 = ~n6547 & n12235 ;
  assign n17143 = n17142 ^ n17141 ;
  assign n17144 = n17143 ^ x14 ;
  assign n17136 = n12228 ^ n7310 ;
  assign n17137 = n17136 ^ n12228 ;
  assign n17138 = ~n12805 & n17137 ;
  assign n17139 = n17138 ^ n12228 ;
  assign n17140 = n6391 & ~n17139 ;
  assign n17145 = n17144 ^ n17140 ;
  assign n17147 = n17146 ^ n17145 ;
  assign n17150 = ~n6529 & n12235 ;
  assign n17149 = ~n6547 & ~n12239 ;
  assign n17151 = n17150 ^ n17149 ;
  assign n17152 = n17151 ^ n6537 ;
  assign n17153 = n17152 ^ x14 ;
  assign n17162 = n6539 & n12866 ;
  assign n17154 = n17151 ^ n6538 ;
  assign n17157 = n12229 ^ x13 ;
  assign n17158 = n17157 ^ n12229 ;
  assign n17159 = ~n12866 & ~n17158 ;
  assign n17160 = n17159 ^ n12229 ;
  assign n17161 = n17154 & ~n17160 ;
  assign n17163 = n17162 ^ n17161 ;
  assign n17164 = ~n17153 & ~n17163 ;
  assign n17148 = n17032 ^ n16768 ;
  assign n17165 = n17164 ^ n17148 ;
  assign n17168 = ~n6529 & ~n12239 ;
  assign n17167 = ~n6547 & n12248 ;
  assign n17169 = n17168 ^ n17167 ;
  assign n17170 = n17169 ^ n6537 ;
  assign n17171 = n17170 ^ x14 ;
  assign n17172 = n17169 ^ n6538 ;
  assign n17178 = ~n13319 & ~n17173 ;
  assign n17179 = n17178 ^ n12235 ;
  assign n17180 = ~n17172 & ~n17179 ;
  assign n17183 = n12235 ^ n6539 ;
  assign n17184 = n17183 ^ n17180 ;
  assign n17185 = n17184 ^ x13 ;
  assign n17186 = n17185 ^ n12235 ;
  assign n17187 = n17186 ^ x13 ;
  assign n17188 = ~n17180 & n17187 ;
  assign n17189 = n17188 ^ x13 ;
  assign n17190 = ~n13319 & ~n17189 ;
  assign n17191 = n17190 ^ n17184 ;
  assign n17192 = ~n17171 & n17191 ;
  assign n17166 = n17029 ^ n16781 ;
  assign n17193 = n17192 ^ n17166 ;
  assign n17210 = n17026 ^ n16793 ;
  assign n17195 = ~n6529 & n12248 ;
  assign n17194 = ~n6547 & ~n12249 ;
  assign n17196 = n17195 ^ n17194 ;
  assign n17197 = n17196 ^ n6537 ;
  assign n17198 = n17197 ^ x14 ;
  assign n17207 = n6539 & n13339 ;
  assign n17199 = n17196 ^ n6538 ;
  assign n17202 = n12239 ^ x13 ;
  assign n17203 = n17202 ^ n12239 ;
  assign n17204 = ~n13339 & ~n17203 ;
  assign n17205 = n17204 ^ n12239 ;
  assign n17206 = n17199 & n17205 ;
  assign n17208 = n17207 ^ n17206 ;
  assign n17209 = ~n17198 & ~n17208 ;
  assign n17211 = n17210 ^ n17209 ;
  assign n17214 = ~n6529 & ~n12249 ;
  assign n17213 = ~n6547 & n12339 ;
  assign n17215 = n17214 ^ n17213 ;
  assign n17216 = n17215 ^ n6537 ;
  assign n17217 = n17216 ^ x14 ;
  assign n17227 = x13 & n13519 ;
  assign n17226 = n8856 & n12248 ;
  assign n17228 = n17227 ^ n17226 ;
  assign n17229 = ~n6539 & n17228 ;
  assign n17224 = n13518 ^ n8856 ;
  assign n17218 = n17215 ^ x14 ;
  assign n17219 = n12248 ^ x13 ;
  assign n17220 = n17219 ^ n12248 ;
  assign n17221 = ~n13518 & ~n17220 ;
  assign n17222 = n17221 ^ n12248 ;
  assign n17223 = ~n17218 & ~n17222 ;
  assign n17225 = n17224 ^ n17223 ;
  assign n17230 = n17229 ^ n17225 ;
  assign n17231 = ~n17217 & n17230 ;
  assign n17212 = n17023 ^ n16803 ;
  assign n17232 = n17231 ^ n17212 ;
  assign n17235 = ~n6529 & n12339 ;
  assign n17234 = ~n6547 & ~n12251 ;
  assign n17236 = n17235 ^ n17234 ;
  assign n17237 = n17236 ^ n6537 ;
  assign n17238 = n17237 ^ x14 ;
  assign n17247 = n6539 & n13553 ;
  assign n17239 = n17236 ^ n6538 ;
  assign n17242 = n12249 ^ x13 ;
  assign n17243 = n17242 ^ n12249 ;
  assign n17244 = ~n14194 & ~n17243 ;
  assign n17245 = n17244 ^ n12249 ;
  assign n17246 = n17239 & n17245 ;
  assign n17248 = n17247 ^ n17246 ;
  assign n17249 = ~n17238 & ~n17248 ;
  assign n17233 = n17020 ^ n16813 ;
  assign n17250 = n17249 ^ n17233 ;
  assign n17253 = ~n6529 & ~n12251 ;
  assign n17252 = ~n6547 & n12253 ;
  assign n17254 = n17253 ^ n17252 ;
  assign n17255 = n17254 ^ n6537 ;
  assign n17256 = n17255 ^ x14 ;
  assign n17257 = n17254 ^ n6538 ;
  assign n17260 = ~n14922 & ~n17173 ;
  assign n17261 = n17260 ^ n12339 ;
  assign n17262 = ~n17257 & ~n17261 ;
  assign n17266 = n12339 ^ n6539 ;
  assign n17267 = n17266 ^ n17262 ;
  assign n17265 = n12339 ^ x13 ;
  assign n17268 = n17267 ^ n17265 ;
  assign n17269 = n17268 ^ x13 ;
  assign n17270 = ~n17262 & n17269 ;
  assign n17271 = n17270 ^ x13 ;
  assign n17272 = ~n13884 & ~n17271 ;
  assign n17273 = n17272 ^ n17267 ;
  assign n17274 = ~n17256 & n17273 ;
  assign n17251 = n17017 ^ n16823 ;
  assign n17275 = n17274 ^ n17251 ;
  assign n17278 = ~n6529 & n12253 ;
  assign n17277 = ~n6547 & n12331 ;
  assign n17279 = n17278 ^ n17277 ;
  assign n17280 = n17279 ^ n6537 ;
  assign n17281 = n17280 ^ x14 ;
  assign n17291 = x13 & ~n13677 ;
  assign n17290 = n8856 & ~n12251 ;
  assign n17292 = n17291 ^ n17290 ;
  assign n17293 = ~n6539 & n17292 ;
  assign n17288 = n13676 ^ n8856 ;
  assign n17282 = n17279 ^ x14 ;
  assign n17283 = n12251 ^ x13 ;
  assign n17284 = n17283 ^ n12251 ;
  assign n17285 = ~n13676 & ~n17284 ;
  assign n17286 = n17285 ^ n12251 ;
  assign n17287 = ~n17282 & n17286 ;
  assign n17289 = n17288 ^ n17287 ;
  assign n17294 = n17293 ^ n17289 ;
  assign n17295 = ~n17281 & n17294 ;
  assign n17276 = n17014 ^ n16833 ;
  assign n17296 = n17295 ^ n17276 ;
  assign n17299 = ~n6529 & n12331 ;
  assign n17298 = ~n6547 & n12257 ;
  assign n17300 = n17299 ^ n17298 ;
  assign n17301 = n17300 ^ n6537 ;
  assign n17302 = n17301 ^ x14 ;
  assign n17306 = n17300 ^ n6538 ;
  assign n17303 = n12253 ^ n6539 ;
  assign n17304 = n17303 ^ x13 ;
  assign n17305 = n17304 ^ n12253 ;
  assign n17307 = n17306 ^ n17305 ;
  assign n17308 = n17307 ^ n17306 ;
  assign n17310 = ~n14088 & ~n17308 ;
  assign n17311 = ~x13 & n17310 ;
  assign n17314 = n17311 ^ n17310 ;
  assign n17312 = n17311 ^ n12253 ;
  assign n17313 = n17306 & ~n17312 ;
  assign n17315 = n17314 ^ n17313 ;
  assign n17316 = n17315 ^ n6539 ;
  assign n17317 = ~n17302 & ~n17316 ;
  assign n17297 = n17011 ^ n16843 ;
  assign n17318 = n17317 ^ n17297 ;
  assign n17321 = ~n6529 & n12257 ;
  assign n17320 = ~n6547 & ~n12258 ;
  assign n17322 = n17321 ^ n17320 ;
  assign n17323 = n17322 ^ n6537 ;
  assign n17324 = n17323 ^ x14 ;
  assign n17334 = n12331 ^ n6539 ;
  assign n17325 = n17322 ^ n6538 ;
  assign n17328 = ~n14219 & ~n17173 ;
  assign n17329 = n17328 ^ n12331 ;
  assign n17330 = ~n17325 & ~n17329 ;
  assign n17335 = n17334 ^ n17330 ;
  assign n17341 = n17335 ^ n17328 ;
  assign n17342 = ~n17324 & n17341 ;
  assign n17319 = n17008 ^ n16857 ;
  assign n17343 = n17342 ^ n17319 ;
  assign n17346 = ~n6529 & ~n12258 ;
  assign n17345 = ~n6547 & n12264 ;
  assign n17347 = n17346 ^ n17345 ;
  assign n17348 = n17347 ^ n6537 ;
  assign n17349 = n17348 ^ x14 ;
  assign n17366 = n12257 ^ n6539 ;
  assign n17353 = n17347 ^ n6538 ;
  assign n17365 = ~n14019 & ~n17173 ;
  assign n17359 = n17365 ^ n12257 ;
  assign n17360 = ~n17353 & ~n17359 ;
  assign n17367 = n17366 ^ n17360 ;
  assign n17368 = n17367 ^ n17365 ;
  assign n17369 = ~n17349 & n17368 ;
  assign n17344 = n17005 ^ n16995 ;
  assign n17370 = n17369 ^ n17344 ;
  assign n17390 = n16988 ^ n16878 ;
  assign n17379 = ~n6529 & ~n12267 ;
  assign n17378 = ~n6547 & n12268 ;
  assign n17380 = n17379 ^ n17378 ;
  assign n17372 = n12264 ^ x13 ;
  assign n17373 = n17372 ^ n12264 ;
  assign n17382 = ~n14428 & ~n17373 ;
  assign n17383 = n17382 ^ n12264 ;
  assign n17384 = n6537 & ~n17383 ;
  assign n15618 = n6537 ^ x14 ;
  assign n17385 = n17384 ^ n15618 ;
  assign n17386 = n17385 ^ x14 ;
  assign n17387 = ~n17380 & ~n17386 ;
  assign n17388 = n17387 ^ x14 ;
  assign n17375 = ~n14428 & n17373 ;
  assign n17376 = n17375 ^ n12264 ;
  assign n17377 = n6539 & n17376 ;
  assign n17389 = n17388 ^ n17377 ;
  assign n17391 = n17390 ^ n17389 ;
  assign n17399 = n6391 & ~n12267 ;
  assign n17397 = n7838 & ~n14450 ;
  assign n17394 = ~n6547 & ~n12276 ;
  assign n17393 = ~n6529 & n12268 ;
  assign n17395 = n17394 ^ n17393 ;
  assign n17396 = n17395 ^ x14 ;
  assign n17398 = n17397 ^ n17396 ;
  assign n17400 = n17399 ^ n17398 ;
  assign n17392 = n16985 ^ n16888 ;
  assign n17401 = n17400 ^ n17392 ;
  assign n17404 = ~n6529 & ~n12276 ;
  assign n17403 = ~n6547 & n12279 ;
  assign n17405 = n17404 ^ n17403 ;
  assign n17406 = n17405 ^ n6537 ;
  assign n17407 = n17406 ^ x14 ;
  assign n17416 = n6539 & n14328 ;
  assign n17408 = n17405 ^ n6538 ;
  assign n17411 = n12268 ^ x13 ;
  assign n17412 = n17411 ^ n12268 ;
  assign n17413 = ~n14328 & ~n17412 ;
  assign n17414 = n17413 ^ n12268 ;
  assign n17415 = n17408 & ~n17414 ;
  assign n17417 = n17416 ^ n17415 ;
  assign n17418 = ~n17407 & ~n17417 ;
  assign n17402 = n16982 ^ n16903 ;
  assign n17419 = n17418 ^ n17402 ;
  assign n17422 = ~n6529 & n12279 ;
  assign n17421 = ~n6547 & ~n12283 ;
  assign n17423 = n17422 ^ n17421 ;
  assign n17424 = n17423 ^ n6537 ;
  assign n17425 = n17424 ^ x14 ;
  assign n17435 = x13 & ~n14475 ;
  assign n17434 = n8856 & ~n12276 ;
  assign n17436 = n17435 ^ n17434 ;
  assign n17437 = ~n6539 & n17436 ;
  assign n17432 = n14465 ^ n8856 ;
  assign n17426 = n17423 ^ x14 ;
  assign n17427 = n12276 ^ x13 ;
  assign n17428 = n17427 ^ n12276 ;
  assign n17429 = ~n14465 & ~n17428 ;
  assign n17430 = n17429 ^ n12276 ;
  assign n17431 = ~n17426 & n17430 ;
  assign n17433 = n17432 ^ n17431 ;
  assign n17438 = n17437 ^ n17433 ;
  assign n17439 = ~n17425 & n17438 ;
  assign n17420 = n16979 ^ n16913 ;
  assign n17440 = n17439 ^ n17420 ;
  assign n17458 = n16976 ^ n16924 ;
  assign n17442 = ~n6529 & ~n12283 ;
  assign n17441 = ~n6547 & ~n12284 ;
  assign n17443 = n17442 ^ n17441 ;
  assign n17444 = n17443 ^ n6537 ;
  assign n17445 = n17444 ^ x14 ;
  assign n17454 = n6539 & n14514 ;
  assign n17446 = n17443 ^ n6538 ;
  assign n17449 = n12279 ^ x13 ;
  assign n17450 = n17449 ^ n12279 ;
  assign n17451 = ~n14514 & ~n17450 ;
  assign n17452 = n17451 ^ n12279 ;
  assign n17453 = n17446 & ~n17452 ;
  assign n17455 = n17454 ^ n17453 ;
  assign n17456 = ~n17445 & ~n17455 ;
  assign n17459 = n17458 ^ n17456 ;
  assign n17462 = ~n6529 & ~n12284 ;
  assign n17461 = ~n6547 & ~n12285 ;
  assign n17463 = n17462 ^ n17461 ;
  assign n17464 = n17463 ^ n6537 ;
  assign n17465 = n17464 ^ x14 ;
  assign n17475 = x13 & ~n14548 ;
  assign n17474 = n8856 & ~n12283 ;
  assign n17476 = n17475 ^ n17474 ;
  assign n17477 = ~n6539 & n17476 ;
  assign n17472 = n14547 ^ n8856 ;
  assign n17466 = n17463 ^ x14 ;
  assign n17467 = n12283 ^ x13 ;
  assign n17468 = n17467 ^ n12283 ;
  assign n17469 = ~n14547 & ~n17468 ;
  assign n17470 = n17469 ^ n12283 ;
  assign n17471 = ~n17466 & n17470 ;
  assign n17473 = n17472 ^ n17471 ;
  assign n17478 = n17477 ^ n17473 ;
  assign n17479 = ~n17465 & n17478 ;
  assign n17460 = n16974 ^ n16964 ;
  assign n17480 = n17479 ^ n17460 ;
  assign n17483 = ~n6547 & n12313 ;
  assign n17482 = ~n6529 & ~n12285 ;
  assign n17484 = n17483 ^ n17482 ;
  assign n17485 = n17484 ^ n6537 ;
  assign n17486 = n17485 ^ x14 ;
  assign n17496 = x13 & ~n14584 ;
  assign n17495 = n8856 & ~n12284 ;
  assign n17497 = n17496 ^ n17495 ;
  assign n17498 = ~n6539 & n17497 ;
  assign n17493 = n14583 ^ n8856 ;
  assign n17487 = n17484 ^ x14 ;
  assign n17488 = n12284 ^ x13 ;
  assign n17489 = n17488 ^ n12284 ;
  assign n17490 = ~n14583 & ~n17489 ;
  assign n17491 = n17490 ^ n12284 ;
  assign n17492 = ~n17487 & n17491 ;
  assign n17494 = n17493 ^ n17492 ;
  assign n17499 = n17498 ^ n17494 ;
  assign n17500 = ~n17486 & n17499 ;
  assign n17481 = n16961 ^ n16953 ;
  assign n17501 = n17500 ^ n17481 ;
  assign n17506 = ~n6529 & n12313 ;
  assign n17505 = ~n6547 & n12289 ;
  assign n17507 = n17506 ^ n17505 ;
  assign n17508 = n17507 ^ n6537 ;
  assign n17509 = n17508 ^ x14 ;
  assign n17510 = n17507 ^ x14 ;
  assign n17511 = n17510 ^ n17507 ;
  assign n17512 = n14583 ^ n12314 ;
  assign n17513 = n6391 & n17512 ;
  assign n17514 = ~n17511 & n17513 ;
  assign n17515 = n17514 ^ n17510 ;
  assign n17517 = n12285 ^ n6539 ;
  assign n17516 = n12285 ^ x13 ;
  assign n17518 = n17517 ^ n17516 ;
  assign n17519 = n17517 ^ n14651 ;
  assign n17520 = n17519 ^ n17517 ;
  assign n17521 = ~n17518 & ~n17520 ;
  assign n17522 = n17521 ^ n17517 ;
  assign n17523 = n17515 & n17522 ;
  assign n17524 = ~n17509 & ~n17523 ;
  assign n17502 = n16935 ^ x17 ;
  assign n17503 = n17502 ^ n16945 ;
  assign n17504 = n17503 ^ n16933 ;
  assign n17525 = n17524 ^ n17504 ;
  assign n17543 = ~n6529 & n12289 ;
  assign n17542 = ~n6547 & ~n12290 ;
  assign n17544 = n17543 ^ n17542 ;
  assign n17545 = n17544 ^ n6537 ;
  assign n17546 = n17545 ^ x14 ;
  assign n17558 = x13 & n14712 ;
  assign n17557 = n8856 & n12313 ;
  assign n17559 = n17558 ^ n17557 ;
  assign n17560 = ~n6539 & n17559 ;
  assign n17555 = n14711 ^ n8856 ;
  assign n17547 = n17544 ^ x14 ;
  assign n17548 = n14712 ^ x13 ;
  assign n17549 = n17548 ^ n14712 ;
  assign n17552 = ~n14711 & n17549 ;
  assign n17553 = n17552 ^ n14712 ;
  assign n17554 = ~n17547 & n17553 ;
  assign n17556 = n17555 ^ n17554 ;
  assign n17561 = n17560 ^ n17556 ;
  assign n17562 = ~n17546 & n17561 ;
  assign n17529 = x17 & ~n12298 ;
  assign n17530 = n16942 & ~n17529 ;
  assign n17526 = n6153 ^ n6147 ;
  assign n17527 = n17526 ^ n6158 ;
  assign n17528 = n12292 & n17527 ;
  assign n17531 = n17530 ^ n17528 ;
  assign n17535 = n12292 ^ n12291 ;
  assign n17536 = n6143 & n17535 ;
  assign n17538 = n12291 & ~n16943 ;
  assign n17539 = n17536 & n17538 ;
  assign n17532 = n16942 ^ n6141 ;
  assign n17533 = n17530 ^ n17529 ;
  assign n17534 = n17532 & n17533 ;
  assign n17537 = n17536 ^ n17534 ;
  assign n17540 = n17539 ^ n17537 ;
  assign n17541 = ~n17531 & ~n17540 ;
  assign n17563 = n17562 ^ n17541 ;
  assign n17581 = n6141 & n12292 ;
  assign n17580 = n6140 & n12291 ;
  assign n17582 = n17581 ^ n17580 ;
  assign n17633 = n17582 ^ n17541 ;
  assign n17565 = ~n6529 & ~n12290 ;
  assign n17564 = ~n6547 & n12293 ;
  assign n17566 = n17565 ^ n17564 ;
  assign n17567 = n17566 ^ n6537 ;
  assign n17568 = n17567 ^ x14 ;
  assign n17577 = n6539 & n14748 ;
  assign n17569 = n17566 ^ n6538 ;
  assign n17572 = n12289 ^ x13 ;
  assign n17573 = n17572 ^ n12289 ;
  assign n17574 = ~n14748 & ~n17573 ;
  assign n17575 = n17574 ^ n12289 ;
  assign n17576 = n17569 & ~n17575 ;
  assign n17578 = n17577 ^ n17576 ;
  assign n17579 = ~n17568 & ~n17578 ;
  assign n17583 = n17582 ^ n17579 ;
  assign n17590 = ~n6529 & n12293 ;
  assign n17589 = ~n6547 & n12292 ;
  assign n17591 = n17590 ^ n17589 ;
  assign n17592 = n17591 ^ x14 ;
  assign n17584 = n12290 ^ n7310 ;
  assign n17585 = n17584 ^ n12290 ;
  assign n17586 = n12297 & n17585 ;
  assign n17587 = n17586 ^ n12290 ;
  assign n17588 = n6391 & ~n17587 ;
  assign n17593 = n17592 ^ n17588 ;
  assign n17595 = n6141 & n12291 ;
  assign n17597 = ~n6529 & n12292 ;
  assign n17596 = ~n6547 & n12291 ;
  assign n17598 = n17597 ^ n17596 ;
  assign n17599 = n17598 ^ n6537 ;
  assign n17600 = n17599 ^ x14 ;
  assign n17616 = n12293 ^ n6539 ;
  assign n17604 = n17598 ^ n6538 ;
  assign n17615 = ~n12299 & ~n17173 ;
  assign n17609 = n17615 ^ n12293 ;
  assign n17610 = ~n17604 & ~n17609 ;
  assign n17617 = n17616 ^ n17610 ;
  assign n17618 = n17617 ^ n17615 ;
  assign n17619 = ~n17600 & n17618 ;
  assign n17620 = n12292 ^ n6403 ;
  assign n17621 = ~n6391 & n17620 ;
  assign n17622 = n17621 ^ n12292 ;
  assign n17623 = n12291 ^ n6391 ;
  assign n17624 = n17623 ^ x14 ;
  assign n17625 = ~n17622 & ~n17624 ;
  assign n17626 = n17625 ^ n6391 ;
  assign n17627 = x14 & ~n17626 ;
  assign n17628 = ~n17619 & n17627 ;
  assign n17629 = ~n17595 & ~n17628 ;
  assign n17630 = n17593 & n17629 ;
  assign n17594 = n17593 ^ n17579 ;
  assign n17631 = n17630 ^ n17594 ;
  assign n17632 = ~n17583 & n17631 ;
  assign n17634 = n17633 ^ n17632 ;
  assign n17635 = n17563 & n17634 ;
  assign n17636 = n17635 ^ n17562 ;
  assign n17637 = n17636 ^ n17504 ;
  assign n17638 = ~n17525 & n17637 ;
  assign n17639 = n17638 ^ n17524 ;
  assign n17640 = n17639 ^ n17500 ;
  assign n17641 = ~n17501 & n17640 ;
  assign n17642 = n17641 ^ n17500 ;
  assign n17643 = n17642 ^ n17479 ;
  assign n17644 = ~n17480 & n17643 ;
  assign n17645 = n17644 ^ n17479 ;
  assign n17646 = n17645 ^ n17456 ;
  assign n17647 = ~n17459 & n17646 ;
  assign n17457 = n17456 ^ n17439 ;
  assign n17648 = n17647 ^ n17457 ;
  assign n17649 = ~n17440 & n17648 ;
  assign n17650 = n17649 ^ n17439 ;
  assign n17651 = n17650 ^ n17418 ;
  assign n17652 = ~n17419 & n17651 ;
  assign n17653 = n17652 ^ n17418 ;
  assign n17654 = n17653 ^ n17400 ;
  assign n17655 = n17401 & ~n17654 ;
  assign n17656 = n17655 ^ n17400 ;
  assign n17657 = n17656 ^ n17389 ;
  assign n17658 = n17391 & ~n17657 ;
  assign n17659 = n17658 ^ n17656 ;
  assign n17371 = n16991 ^ n16868 ;
  assign n17660 = n17659 ^ n17371 ;
  assign n17667 = ~n6529 & n12264 ;
  assign n17666 = ~n6547 & ~n12267 ;
  assign n17668 = n17667 ^ n17666 ;
  assign n17669 = n17668 ^ x14 ;
  assign n17661 = n12258 ^ n7310 ;
  assign n17662 = n17661 ^ n12258 ;
  assign n17663 = ~n14242 & n17662 ;
  assign n17664 = n17663 ^ n12258 ;
  assign n17665 = n6391 & ~n17664 ;
  assign n17670 = n17669 ^ n17665 ;
  assign n17671 = n17670 ^ n17371 ;
  assign n17672 = n17660 & ~n17671 ;
  assign n17673 = n17672 ^ n17659 ;
  assign n17674 = n17673 ^ n17369 ;
  assign n17675 = ~n17370 & ~n17674 ;
  assign n17676 = n17675 ^ n17369 ;
  assign n17677 = n17676 ^ n17342 ;
  assign n17678 = ~n17343 & n17677 ;
  assign n17679 = n17678 ^ n17342 ;
  assign n17680 = n17679 ^ n17317 ;
  assign n17681 = ~n17318 & n17680 ;
  assign n17682 = n17681 ^ n17317 ;
  assign n17683 = n17682 ^ n17295 ;
  assign n17684 = ~n17296 & n17683 ;
  assign n17685 = n17684 ^ n17295 ;
  assign n17686 = n17685 ^ n17274 ;
  assign n17687 = ~n17275 & n17686 ;
  assign n17688 = n17687 ^ n17274 ;
  assign n17689 = n17688 ^ n17249 ;
  assign n17690 = ~n17250 & n17689 ;
  assign n17691 = n17690 ^ n17249 ;
  assign n17692 = n17691 ^ n17231 ;
  assign n17693 = ~n17232 & n17692 ;
  assign n17694 = n17693 ^ n17231 ;
  assign n17695 = n17694 ^ n17209 ;
  assign n17696 = n17211 & n17695 ;
  assign n17697 = n17696 ^ n17209 ;
  assign n17698 = n17697 ^ n17192 ;
  assign n17699 = n17193 & n17698 ;
  assign n17700 = n17699 ^ n17192 ;
  assign n17701 = n17700 ^ n17164 ;
  assign n17702 = n17165 & n17701 ;
  assign n17703 = n17702 ^ n17164 ;
  assign n17704 = n17703 ^ n17145 ;
  assign n17705 = ~n17147 & ~n17704 ;
  assign n17706 = n17705 ^ n17703 ;
  assign n17707 = n17706 ^ n17133 ;
  assign n17708 = n17135 & n17707 ;
  assign n17709 = n17708 ^ n17133 ;
  assign n17710 = n17709 ^ n17109 ;
  assign n17711 = ~n17110 & n17710 ;
  assign n17712 = n17711 ^ n17109 ;
  assign n17713 = n17712 ^ n17087 ;
  assign n17714 = n17089 & n17713 ;
  assign n17715 = n17714 ^ n17087 ;
  assign n17716 = n17715 ^ n17070 ;
  assign n17717 = ~n17071 & ~n17716 ;
  assign n17718 = n17717 ^ n17070 ;
  assign n17734 = n17733 ^ n17718 ;
  assign n17741 = n8139 & ~n12209 ;
  assign n17739 = n8150 & n12983 ;
  assign n17736 = n8484 & ~n12204 ;
  assign n17735 = n8144 & n12419 ;
  assign n17737 = n17736 ^ n17735 ;
  assign n17738 = n17737 ^ x8 ;
  assign n17740 = n17739 ^ n17738 ;
  assign n17742 = n17741 ^ n17740 ;
  assign n17743 = n17742 ^ n17718 ;
  assign n17744 = n17734 & n17743 ;
  assign n17745 = n17744 ^ n17742 ;
  assign n17746 = n17745 ^ n14033 ;
  assign n16701 = n7142 & ~n12405 ;
  assign n16699 = ~n12651 & n20240 ;
  assign n16696 = n7151 & n12419 ;
  assign n16695 = n7148 & ~n12210 ;
  assign n16697 = n16696 ^ n16695 ;
  assign n16698 = n16697 ^ x11 ;
  assign n16700 = n16699 ^ n16698 ;
  assign n16702 = n16701 ^ n16700 ;
  assign n16679 = n16285 ^ n16006 ;
  assign n16680 = n16679 ^ n16677 ;
  assign n16681 = n16680 ^ n16679 ;
  assign n16692 = n16691 ^ n16681 ;
  assign n16693 = ~n16678 & n16692 ;
  assign n16694 = n16693 ^ n16680 ;
  assign n17759 = n16702 ^ n16694 ;
  assign n17761 = n17759 ^ n17719 ;
  assign n17760 = n17759 ^ n17732 ;
  assign n17762 = n17761 ^ n17760 ;
  assign n17763 = ~n17724 & ~n17762 ;
  assign n17764 = n17763 ^ n17761 ;
  assign n17749 = n8139 & ~n12204 ;
  assign n17748 = n8144 & ~n12209 ;
  assign n17750 = n17749 ^ n17748 ;
  assign n17747 = n8137 & ~n12435 ;
  assign n17751 = n17750 ^ n17747 ;
  assign n17752 = n17751 ^ n17750 ;
  assign n17753 = n12432 & n17752 ;
  assign n17754 = n17751 ^ x8 ;
  assign n17755 = n17754 ^ x7 ;
  assign n17756 = n17755 ^ n17751 ;
  assign n17757 = n17753 & n17756 ;
  assign n17758 = n17757 ^ n17754 ;
  assign n17765 = n17764 ^ n17758 ;
  assign n17766 = n17765 ^ n17745 ;
  assign n17767 = ~n17746 & ~n17766 ;
  assign n17768 = n17767 ^ n14033 ;
  assign n17769 = n17759 ^ n17758 ;
  assign n17770 = n17764 & ~n17769 ;
  assign n17771 = n17770 ^ n17759 ;
  assign n17773 = n17768 & n17771 ;
  assign n16325 = n7151 & ~n12209 ;
  assign n16324 = n7148 & ~n12405 ;
  assign n16326 = n16325 ^ n16324 ;
  assign n16327 = n16326 ^ x11 ;
  assign n16323 = n13052 & n20240 ;
  assign n16328 = n16327 ^ n16323 ;
  assign n16322 = n7142 & n12419 ;
  assign n16329 = n16328 ^ n16322 ;
  assign n16705 = n16679 ^ n16329 ;
  assign n16703 = n16702 ^ n16679 ;
  assign n16704 = ~n16694 & ~n16703 ;
  assign n16706 = n16705 ^ n16704 ;
  assign n16330 = n16287 ^ n15945 ;
  assign n17776 = n16706 ^ n16330 ;
  assign n17784 = n8144 & ~n12204 ;
  assign n17782 = n8484 ^ x8 ;
  assign n17779 = n8150 & ~n12431 ;
  assign n17780 = n17779 ^ n8139 ;
  assign n17781 = ~n12435 & n17780 ;
  assign n17783 = n17782 ^ n17781 ;
  assign n17785 = n17784 ^ n17783 ;
  assign n17788 = n17776 & ~n17785 ;
  assign n8140 = n8137 ^ n8134 ;
  assign n8141 = n8140 ^ n8139 ;
  assign n16709 = n8141 ^ n8135 ;
  assign n16331 = n16330 ^ n16329 ;
  assign n16707 = n16331 & n16706 ;
  assign n16708 = n16707 ^ n16330 ;
  assign n16710 = n16709 ^ n16708 ;
  assign n16317 = x7 ^ x6 ;
  assign n16318 = ~n12435 & ~n16317 ;
  assign n16319 = x8 ^ x5 ;
  assign n16320 = n9896 & n16319 ;
  assign n16321 = n16318 & n16320 ;
  assign n16711 = n16710 ^ n16321 ;
  assign n16316 = n16315 ^ n15643 ;
  assign n16712 = n16711 ^ n16316 ;
  assign n17789 = n17788 ^ n16712 ;
  assign n17790 = n17789 ^ n16712 ;
  assign n17786 = n17785 ^ n17776 ;
  assign n17772 = n17771 ^ n17768 ;
  assign n17774 = n17773 ^ n17772 ;
  assign n17775 = n17774 ^ n16712 ;
  assign n17787 = n17786 ^ n17775 ;
  assign n17791 = n17790 ^ n17787 ;
  assign n17792 = n10331 & ~n12435 ;
  assign n17793 = n10331 ^ x5 ;
  assign n17794 = n17793 ^ x4 ;
  assign n17795 = n17792 & ~n17794 ;
  assign n17796 = n17795 ^ n17793 ;
  assign n17799 = n8139 & n12419 ;
  assign n17798 = n8144 & ~n12405 ;
  assign n17800 = n17799 ^ n17798 ;
  assign n17801 = n17800 ^ n8145 ;
  assign n17802 = n17801 ^ x8 ;
  assign n17804 = ~x7 & ~n13051 ;
  assign n17807 = n17804 ^ n13052 ;
  assign n17808 = n8146 & n17807 ;
  assign n17803 = n17800 ^ x8 ;
  assign n17805 = n17804 ^ n12209 ;
  assign n17806 = n17803 & n17805 ;
  assign n17809 = n17808 ^ n17806 ;
  assign n17810 = ~n17802 & ~n17809 ;
  assign n17797 = n17715 ^ n17071 ;
  assign n17811 = n17810 ^ n17797 ;
  assign n17820 = n7142 & ~n12214 ;
  assign n17815 = n17712 ^ n17089 ;
  assign n17816 = n17815 ^ x11 ;
  assign n17814 = n7151 & ~n12400 ;
  assign n17817 = n17816 ^ n17814 ;
  assign n17813 = n7148 & n12222 ;
  assign n17818 = n17817 ^ n17813 ;
  assign n17812 = n12667 & n20240 ;
  assign n17819 = n17818 ^ n17812 ;
  assign n17821 = n17820 ^ n17819 ;
  assign n17830 = n7142 & n12222 ;
  assign n17825 = n17709 ^ n17110 ;
  assign n17826 = n17825 ^ x11 ;
  assign n17824 = n7151 & ~n12214 ;
  assign n17827 = n17826 ^ n17824 ;
  assign n17823 = n7148 & n12380 ;
  assign n17828 = n17827 ^ n17823 ;
  assign n17822 = n12608 & n20240 ;
  assign n17829 = n17828 ^ n17822 ;
  assign n17831 = n17830 ^ n17829 ;
  assign n17840 = n7148 & n12376 ;
  assign n17838 = n7151 & n12222 ;
  assign n17836 = n13770 & n20240 ;
  assign n17834 = n7142 & n12380 ;
  assign n17832 = n17706 ^ n17135 ;
  assign n17833 = n17832 ^ x11 ;
  assign n17835 = n17834 ^ n17833 ;
  assign n17837 = n17836 ^ n17835 ;
  assign n17839 = n17838 ^ n17837 ;
  assign n17841 = n17840 ^ n17839 ;
  assign n17855 = n17703 ^ n17147 ;
  assign n17843 = n7142 & n12376 ;
  assign n17842 = n7148 & ~n12382 ;
  assign n17844 = n17843 ^ n17842 ;
  assign n17845 = n17844 ^ n7149 ;
  assign n17846 = n17845 ^ x11 ;
  assign n17848 = ~x10 & n12554 ;
  assign n17851 = n17848 ^ n12555 ;
  assign n17852 = n7150 & n17851 ;
  assign n17847 = n17844 ^ x11 ;
  assign n17849 = n17848 ^ n12380 ;
  assign n17850 = n17847 & ~n17849 ;
  assign n17853 = n17852 ^ n17850 ;
  assign n17854 = ~n17846 & ~n17853 ;
  assign n17856 = n17855 ^ n17854 ;
  assign n17866 = n7142 & ~n12228 ;
  assign n17861 = n17697 ^ n17193 ;
  assign n17862 = n17861 ^ x11 ;
  assign n17860 = n7151 & ~n12382 ;
  assign n17863 = n17862 ^ n17860 ;
  assign n17859 = n7148 & n12229 ;
  assign n17864 = n17863 ^ n17859 ;
  assign n17858 = n13445 & n20240 ;
  assign n17865 = n17864 ^ n17858 ;
  assign n17867 = n17866 ^ n17865 ;
  assign n17875 = n7142 & n12229 ;
  assign n17873 = n13779 & n20240 ;
  assign n17870 = n7151 & ~n12228 ;
  assign n17869 = n7148 & n12235 ;
  assign n17871 = n17870 ^ n17869 ;
  assign n17872 = n17871 ^ x11 ;
  assign n17874 = n17873 ^ n17872 ;
  assign n17876 = n17875 ^ n17874 ;
  assign n17868 = n17694 ^ n17211 ;
  assign n17877 = n17876 ^ n17868 ;
  assign n17886 = n7142 & n12235 ;
  assign n17881 = n17691 ^ n17232 ;
  assign n17882 = n17881 ^ x11 ;
  assign n17880 = n7151 & n12229 ;
  assign n17883 = n17882 ^ n17880 ;
  assign n17879 = n7148 & ~n12239 ;
  assign n17884 = n17883 ^ n17879 ;
  assign n17878 = ~n12867 & n20240 ;
  assign n17885 = n17884 ^ n17878 ;
  assign n17887 = n17886 ^ n17885 ;
  assign n17895 = n7142 & ~n12239 ;
  assign n17893 = ~n13329 & n20240 ;
  assign n17890 = n7151 & n12235 ;
  assign n17889 = n7148 & n12248 ;
  assign n17891 = n17890 ^ n17889 ;
  assign n17892 = n17891 ^ x11 ;
  assign n17894 = n17893 ^ n17892 ;
  assign n17896 = n17895 ^ n17894 ;
  assign n17888 = n17688 ^ n17250 ;
  assign n17897 = n17896 ^ n17888 ;
  assign n17905 = n7142 & n12248 ;
  assign n17903 = n13343 & n20240 ;
  assign n17900 = n7151 & ~n12239 ;
  assign n17899 = n7148 & ~n12249 ;
  assign n17901 = n17900 ^ n17899 ;
  assign n17902 = n17901 ^ x11 ;
  assign n17904 = n17903 ^ n17902 ;
  assign n17906 = n17905 ^ n17904 ;
  assign n17898 = n17685 ^ n17275 ;
  assign n17907 = n17906 ^ n17898 ;
  assign n17912 = n7151 & n12248 ;
  assign n17911 = n7148 & n12339 ;
  assign n17913 = n17912 ^ n17911 ;
  assign n17914 = n17913 ^ x11 ;
  assign n17910 = ~n13519 & n20240 ;
  assign n17915 = n17914 ^ n17910 ;
  assign n17909 = n7142 & ~n12249 ;
  assign n17916 = n17915 ^ n17909 ;
  assign n17908 = n17682 ^ n17296 ;
  assign n17917 = n17916 ^ n17908 ;
  assign n17926 = n7142 & n12339 ;
  assign n17921 = n17679 ^ n17318 ;
  assign n17922 = n17921 ^ x11 ;
  assign n17920 = n7151 & ~n12249 ;
  assign n17923 = n17922 ^ n17920 ;
  assign n17919 = n7148 & ~n12251 ;
  assign n17924 = n17923 ^ n17919 ;
  assign n17918 = n13554 & n20240 ;
  assign n17925 = n17924 ^ n17918 ;
  assign n17927 = n17926 ^ n17925 ;
  assign n17935 = n7142 & ~n12251 ;
  assign n17933 = ~n13885 & n20240 ;
  assign n17930 = n7151 & n12339 ;
  assign n17929 = n7148 & n12253 ;
  assign n17931 = n17930 ^ n17929 ;
  assign n17932 = n17931 ^ x11 ;
  assign n17934 = n17933 ^ n17932 ;
  assign n17936 = n17935 ^ n17934 ;
  assign n17928 = n17676 ^ n17343 ;
  assign n17937 = n17936 ^ n17928 ;
  assign n17942 = n7151 & ~n12251 ;
  assign n17941 = n7148 & n12331 ;
  assign n17943 = n17942 ^ n17941 ;
  assign n17944 = n17943 ^ x11 ;
  assign n17940 = n13677 & n20240 ;
  assign n17945 = n17944 ^ n17940 ;
  assign n17939 = n7142 & n12253 ;
  assign n17946 = n17945 ^ n17939 ;
  assign n17938 = n17673 ^ n17370 ;
  assign n17947 = n17946 ^ n17938 ;
  assign n17952 = n7151 & n12253 ;
  assign n17951 = n7148 & n12257 ;
  assign n17953 = n17952 ^ n17951 ;
  assign n17954 = n17953 ^ x11 ;
  assign n17950 = ~n14414 & n20240 ;
  assign n17955 = n17954 ^ n17950 ;
  assign n17949 = n7142 & n12331 ;
  assign n17956 = n17955 ^ n17949 ;
  assign n17948 = n17671 ^ n17659 ;
  assign n17957 = n17956 ^ n17948 ;
  assign n17965 = n7142 & n12257 ;
  assign n17963 = ~n14972 & n20240 ;
  assign n17960 = n7151 & n12331 ;
  assign n17959 = n7148 & ~n12258 ;
  assign n17961 = n17960 ^ n17959 ;
  assign n17962 = n17961 ^ x11 ;
  assign n17964 = n17963 ^ n17962 ;
  assign n17966 = n17965 ^ n17964 ;
  assign n17958 = n17656 ^ n17391 ;
  assign n17967 = n17966 ^ n17958 ;
  assign n17975 = n7142 & ~n12258 ;
  assign n17973 = ~n14020 & n20240 ;
  assign n17970 = n7151 & n12257 ;
  assign n17969 = n7148 & n12264 ;
  assign n17971 = n17970 ^ n17969 ;
  assign n17972 = n17971 ^ x11 ;
  assign n17974 = n17973 ^ n17972 ;
  assign n17976 = n17975 ^ n17974 ;
  assign n17968 = n17653 ^ n17401 ;
  assign n17977 = n17976 ^ n17968 ;
  assign n17985 = n7142 & n12264 ;
  assign n17983 = n14243 & n20240 ;
  assign n17980 = n7151 & ~n12258 ;
  assign n17979 = n7148 & ~n12267 ;
  assign n17981 = n17980 ^ n17979 ;
  assign n17982 = n17981 ^ x11 ;
  assign n17984 = n17983 ^ n17982 ;
  assign n17986 = n17985 ^ n17984 ;
  assign n17978 = n17650 ^ n17419 ;
  assign n17987 = n17986 ^ n17978 ;
  assign n17993 = ~x10 & ~n14428 ;
  assign n17997 = n17993 ^ n14429 ;
  assign n17998 = n7150 & ~n17997 ;
  assign n17994 = n17993 ^ n12264 ;
  assign n17995 = n7149 & n17994 ;
  assign n17990 = n7142 & ~n12267 ;
  assign n17989 = n7148 & n12268 ;
  assign n17991 = n17990 ^ n17989 ;
  assign n17992 = n17991 ^ x11 ;
  assign n17996 = n17995 ^ n17992 ;
  assign n17999 = n17998 ^ n17996 ;
  assign n17988 = n17648 ^ n17420 ;
  assign n18000 = n17999 ^ n17988 ;
  assign n18011 = n17645 ^ n17459 ;
  assign n18007 = n7148 & ~n12276 ;
  assign n18006 = n7142 & n12268 ;
  assign n18008 = n18007 ^ n18006 ;
  assign n18009 = n18008 ^ x11 ;
  assign n18001 = n12267 ^ n9499 ;
  assign n18002 = n18001 ^ n12267 ;
  assign n18003 = ~n14450 & n18002 ;
  assign n18004 = n18003 ^ n12267 ;
  assign n18005 = n7140 & ~n18004 ;
  assign n18010 = n18009 ^ n18005 ;
  assign n18012 = n18011 ^ n18010 ;
  assign n18015 = n7142 & ~n12276 ;
  assign n18014 = n7148 & n12279 ;
  assign n18016 = n18015 ^ n18014 ;
  assign n18017 = n18016 ^ n7149 ;
  assign n18018 = n18017 ^ x11 ;
  assign n18020 = ~x10 & ~n14328 ;
  assign n18023 = n18020 ^ n14329 ;
  assign n18024 = n7150 & ~n18023 ;
  assign n18019 = n18016 ^ x11 ;
  assign n18021 = n18020 ^ n12268 ;
  assign n18022 = n18019 & ~n18021 ;
  assign n18025 = n18024 ^ n18022 ;
  assign n18026 = ~n18018 & ~n18025 ;
  assign n18013 = n17642 ^ n17480 ;
  assign n18027 = n18026 ^ n18013 ;
  assign n18039 = n17639 ^ n17501 ;
  assign n18037 = n7148 & ~n12283 ;
  assign n18035 = n7142 & n12279 ;
  assign n18028 = n12276 ^ x11 ;
  assign n18029 = n18028 ^ x10 ;
  assign n18030 = n18029 ^ n12276 ;
  assign n18031 = ~n14465 & n18030 ;
  assign n18032 = n18031 ^ n12276 ;
  assign n18033 = n7140 & ~n18032 ;
  assign n18034 = n18033 ^ x11 ;
  assign n18036 = n18035 ^ n18034 ;
  assign n18038 = n18037 ^ n18036 ;
  assign n18040 = n18039 ^ n18038 ;
  assign n18043 = n7142 & ~n12283 ;
  assign n18042 = n7148 & ~n12284 ;
  assign n18044 = n18043 ^ n18042 ;
  assign n18045 = n18044 ^ n7149 ;
  assign n18046 = n18045 ^ x11 ;
  assign n18048 = ~x10 & ~n14514 ;
  assign n18051 = n18048 ^ n14528 ;
  assign n18052 = n7150 & ~n18051 ;
  assign n18047 = n18044 ^ x11 ;
  assign n18049 = n18048 ^ n12279 ;
  assign n18050 = n18047 & ~n18049 ;
  assign n18053 = n18052 ^ n18050 ;
  assign n18054 = ~n18046 & ~n18053 ;
  assign n18164 = n18054 ^ n18039 ;
  assign n18041 = n17636 ^ n17525 ;
  assign n18055 = n18054 ^ n18041 ;
  assign n18066 = n7148 & ~n12285 ;
  assign n18064 = n7142 & ~n12284 ;
  assign n18057 = n12283 ^ x11 ;
  assign n18058 = n18057 ^ x10 ;
  assign n18059 = n18058 ^ n12283 ;
  assign n18060 = ~n14547 & n18059 ;
  assign n18061 = n18060 ^ n12283 ;
  assign n18062 = n7140 & ~n18061 ;
  assign n18063 = n18062 ^ x11 ;
  assign n18065 = n18064 ^ n18063 ;
  assign n18067 = n18066 ^ n18065 ;
  assign n18056 = n17634 ^ n17562 ;
  assign n18068 = n18067 ^ n18056 ;
  assign n18117 = n17627 ^ n17619 ;
  assign n18079 = n6391 & n12291 ;
  assign n18080 = ~n12298 & ~n20255 ;
  assign n18081 = n12301 ^ n12292 ;
  assign n18082 = ~n18081 & n20240 ;
  assign n18088 = n7151 & n12293 ;
  assign n18083 = n12293 ^ n7148 ;
  assign n18084 = n18083 ^ n7148 ;
  assign n18085 = n18084 & n20240 ;
  assign n18086 = n18085 ^ n7148 ;
  assign n18087 = n12291 & n18086 ;
  assign n18089 = n18088 ^ n18087 ;
  assign n18090 = n18082 & ~n18089 ;
  assign n18091 = n18090 ^ n18089 ;
  assign n18092 = x11 & ~n18091 ;
  assign n18093 = ~n18080 & n18092 ;
  assign n18094 = ~n18079 & ~n18093 ;
  assign n18101 = n7142 & n12293 ;
  assign n18099 = ~n14785 & n20240 ;
  assign n18096 = n7151 & ~n12290 ;
  assign n18095 = n7148 & n12292 ;
  assign n18097 = n18096 ^ n18095 ;
  assign n18098 = n18097 ^ x11 ;
  assign n18100 = n18099 ^ n18098 ;
  assign n18102 = n18101 ^ n18100 ;
  assign n18103 = n18094 & n18102 ;
  assign n18104 = n18103 ^ n18102 ;
  assign n18077 = n12291 & n15984 ;
  assign n18071 = n17535 ^ n12292 ;
  assign n18072 = n12292 ^ x12 ;
  assign n18073 = n18072 ^ n12292 ;
  assign n18074 = n18071 & ~n18073 ;
  assign n18075 = n18074 ^ n12292 ;
  assign n18076 = n6391 & n18075 ;
  assign n18078 = n18077 ^ n18076 ;
  assign n18105 = n18104 ^ n18078 ;
  assign n18113 = n7142 & ~n12290 ;
  assign n18109 = n18078 ^ x11 ;
  assign n18108 = n7151 & n12289 ;
  assign n18110 = n18109 ^ n18108 ;
  assign n18107 = n7148 & n12293 ;
  assign n18111 = n18110 ^ n18107 ;
  assign n18106 = ~n14749 & n20240 ;
  assign n18112 = n18111 ^ n18106 ;
  assign n18114 = n18113 ^ n18112 ;
  assign n18115 = n18105 & ~n18114 ;
  assign n18116 = n18115 ^ n18104 ;
  assign n18118 = n18117 ^ n18116 ;
  assign n18125 = ~n14712 & n20240 ;
  assign n18122 = n18116 ^ x11 ;
  assign n18121 = n7148 & ~n12290 ;
  assign n18123 = n18122 ^ n18121 ;
  assign n18120 = n7151 & n12313 ;
  assign n18124 = n18123 ^ n18120 ;
  assign n18126 = n18125 ^ n18124 ;
  assign n18119 = n7142 & n12289 ;
  assign n18127 = n18126 ^ n18119 ;
  assign n18128 = ~n18118 & ~n18127 ;
  assign n18129 = n18128 ^ n18117 ;
  assign n18069 = n17628 ^ n17595 ;
  assign n18070 = n18069 ^ n17593 ;
  assign n18131 = n18129 ^ n18070 ;
  assign n18130 = ~n18070 & n18129 ;
  assign n18132 = n18131 ^ n18130 ;
  assign n18137 = n14652 & n20240 ;
  assign n18136 = n7142 & n12313 ;
  assign n18138 = n18137 ^ n18136 ;
  assign n18134 = n7151 & ~n12285 ;
  assign n18133 = n7148 & n12289 ;
  assign n18135 = n18134 ^ n18133 ;
  assign n18139 = n18138 ^ n18135 ;
  assign n18140 = n18139 ^ x11 ;
  assign n18146 = n14584 & n20240 ;
  assign n18145 = n7142 & ~n12285 ;
  assign n18147 = n18146 ^ n18145 ;
  assign n18143 = n7151 & ~n12284 ;
  assign n18142 = n7148 & n12313 ;
  assign n18144 = n18143 ^ n18142 ;
  assign n18148 = n18147 ^ n18144 ;
  assign n18149 = n18148 ^ n18139 ;
  assign n18141 = n17631 ^ n17582 ;
  assign n18150 = n18149 ^ n18141 ;
  assign n18151 = ~n18140 & ~n18150 ;
  assign n18152 = ~n18132 & n18151 ;
  assign n18153 = n18141 ^ n18130 ;
  assign n18154 = n18148 ^ x11 ;
  assign n18155 = n18154 ^ n18130 ;
  assign n18156 = n18153 & ~n18155 ;
  assign n18157 = n18156 ^ n18130 ;
  assign n18158 = ~n18152 & ~n18157 ;
  assign n18159 = n18158 ^ n18067 ;
  assign n18160 = n18068 & n18159 ;
  assign n18161 = n18160 ^ n18067 ;
  assign n18162 = n18161 ^ n18041 ;
  assign n18163 = ~n18055 & ~n18162 ;
  assign n18165 = n18164 ^ n18163 ;
  assign n18166 = n18040 & ~n18165 ;
  assign n18167 = n18166 ^ n18039 ;
  assign n18168 = n18167 ^ n18013 ;
  assign n18169 = ~n18027 & ~n18168 ;
  assign n18170 = n18169 ^ n18026 ;
  assign n18171 = n18170 ^ n18010 ;
  assign n18172 = n18012 & ~n18171 ;
  assign n18173 = n18172 ^ n18010 ;
  assign n18174 = n18173 ^ n17999 ;
  assign n18175 = n18000 & n18174 ;
  assign n18176 = n18175 ^ n17999 ;
  assign n18177 = n18176 ^ n17986 ;
  assign n18178 = n17987 & n18177 ;
  assign n18179 = n18178 ^ n17986 ;
  assign n18180 = n18179 ^ n17976 ;
  assign n18181 = ~n17977 & n18180 ;
  assign n18182 = n18181 ^ n17976 ;
  assign n18183 = n18182 ^ n17966 ;
  assign n18184 = ~n17967 & n18183 ;
  assign n18185 = n18184 ^ n17966 ;
  assign n18186 = n18185 ^ n17956 ;
  assign n18187 = n17957 & n18186 ;
  assign n18188 = n18187 ^ n17956 ;
  assign n18189 = n18188 ^ n17946 ;
  assign n18190 = ~n17947 & n18189 ;
  assign n18191 = n18190 ^ n17946 ;
  assign n18192 = n18191 ^ n17936 ;
  assign n18193 = n17937 & n18192 ;
  assign n18194 = n18193 ^ n17936 ;
  assign n18195 = n18194 ^ n17921 ;
  assign n18196 = n17927 & n18195 ;
  assign n18197 = n18196 ^ n17921 ;
  assign n18198 = n18197 ^ n17916 ;
  assign n18199 = n17917 & n18198 ;
  assign n18200 = n18199 ^ n17916 ;
  assign n18201 = n18200 ^ n17906 ;
  assign n18202 = n17907 & n18201 ;
  assign n18203 = n18202 ^ n17906 ;
  assign n18204 = n18203 ^ n17896 ;
  assign n18205 = n17897 & n18204 ;
  assign n18206 = n18205 ^ n17896 ;
  assign n18207 = n18206 ^ n17881 ;
  assign n18208 = n17887 & n18207 ;
  assign n18209 = n18208 ^ n17881 ;
  assign n18210 = n18209 ^ n17876 ;
  assign n18211 = ~n17877 & n18210 ;
  assign n18212 = n18211 ^ n17876 ;
  assign n18213 = n18212 ^ n17861 ;
  assign n18214 = ~n17867 & ~n18213 ;
  assign n18215 = n18214 ^ n17861 ;
  assign n17857 = n17700 ^ n17165 ;
  assign n18216 = n18215 ^ n17857 ;
  assign n18224 = n7142 & ~n12382 ;
  assign n18220 = n17857 ^ x11 ;
  assign n18219 = n7151 & n12376 ;
  assign n18221 = n18220 ^ n18219 ;
  assign n18218 = n7148 & ~n12228 ;
  assign n18222 = n18221 ^ n18218 ;
  assign n18217 = n12928 & n20240 ;
  assign n18223 = n18222 ^ n18217 ;
  assign n18225 = n18224 ^ n18223 ;
  assign n18226 = n18216 & n18225 ;
  assign n18227 = n18226 ^ n18215 ;
  assign n18228 = n18227 ^ n17854 ;
  assign n18229 = n17856 & n18228 ;
  assign n18230 = n18229 ^ n17854 ;
  assign n18231 = n18230 ^ n17832 ;
  assign n18232 = ~n17841 & n18231 ;
  assign n18233 = n18232 ^ n17832 ;
  assign n18234 = n18233 ^ n17825 ;
  assign n18235 = n17831 & ~n18234 ;
  assign n18236 = n18235 ^ n17825 ;
  assign n18237 = n18236 ^ n17815 ;
  assign n18238 = ~n17821 & ~n18237 ;
  assign n18239 = n18238 ^ n17815 ;
  assign n18240 = n18239 ^ n17810 ;
  assign n18241 = ~n17811 & n18240 ;
  assign n18242 = n18241 ^ n17810 ;
  assign n18243 = n18242 ^ n17796 ;
  assign n18244 = n17742 ^ n17734 ;
  assign n18245 = n18244 ^ n18242 ;
  assign n18246 = ~n18243 & ~n18245 ;
  assign n18247 = ~n17796 & n18246 ;
  assign n18248 = n17765 ^ n17746 ;
  assign n20173 = n18248 ^ n18246 ;
  assign n18778 = n25051 ^ n10322 ;
  assign n18775 = ~x4 & ~n13051 ;
  assign n18779 = n18775 ^ n13052 ;
  assign n18780 = n18778 & n18779 ;
  assign n18772 = n10327 & n12419 ;
  assign n18771 = ~n10334 & ~n12405 ;
  assign n18773 = n18772 ^ n18771 ;
  assign n18774 = n18773 ^ x5 ;
  assign n18776 = n18775 ^ n12209 ;
  assign n18777 = n18774 & n18776 ;
  assign n18781 = n18780 ^ n18777 ;
  assign n10340 = x5 & ~n10322 ;
  assign n18782 = n18773 ^ n10340 ;
  assign n18783 = ~n18781 & ~n18782 ;
  assign n18289 = n8144 & n12222 ;
  assign n18287 = n8139 & ~n12214 ;
  assign n18280 = n12667 ^ x8 ;
  assign n18281 = n18280 ^ x7 ;
  assign n18282 = n18281 ^ n12667 ;
  assign n18283 = ~n12666 & ~n18282 ;
  assign n18284 = n18283 ^ n12667 ;
  assign n18285 = n8137 & n18284 ;
  assign n18286 = n18285 ^ x8 ;
  assign n18288 = n18287 ^ n18286 ;
  assign n18290 = n18289 ^ n18288 ;
  assign n18279 = n18227 ^ n17856 ;
  assign n18291 = n18290 ^ n18279 ;
  assign n18295 = n8139 & n12380 ;
  assign n18294 = n8144 & n12376 ;
  assign n18296 = n18295 ^ n18294 ;
  assign n18297 = n18296 ^ n8145 ;
  assign n18298 = n18297 ^ x8 ;
  assign n18299 = n18296 ^ x8 ;
  assign n18300 = n18299 ^ n8146 ;
  assign n18301 = ~n13770 & n18300 ;
  assign n18302 = n18301 ^ n8146 ;
  assign n18303 = n18302 ^ x7 ;
  assign n18304 = n18303 ^ n12222 ;
  assign n18305 = n18304 ^ n18302 ;
  assign n18306 = n18302 ^ n18300 ;
  assign n18307 = n18306 ^ n18302 ;
  assign n18308 = n18305 & n18307 ;
  assign n18309 = n18308 ^ n18302 ;
  assign n18310 = n12390 & n18309 ;
  assign n18311 = n18310 ^ n18302 ;
  assign n18312 = ~n18298 & ~n18311 ;
  assign n18293 = n18212 ^ n17867 ;
  assign n18313 = n18312 ^ n18293 ;
  assign n18322 = n8139 & n12376 ;
  assign n18317 = n18209 ^ n17877 ;
  assign n18318 = n18317 ^ x8 ;
  assign n18316 = n8484 & n12380 ;
  assign n18319 = n18318 ^ n18316 ;
  assign n18315 = n8144 & ~n12382 ;
  assign n18320 = n18319 ^ n18315 ;
  assign n18314 = n8150 & n12555 ;
  assign n18321 = n18320 ^ n18314 ;
  assign n18323 = n18322 ^ n18321 ;
  assign n18332 = n8139 & ~n12382 ;
  assign n18329 = n8144 & ~n12228 ;
  assign n18327 = n8484 & n12376 ;
  assign n18325 = n18206 ^ n17887 ;
  assign n18326 = n18325 ^ x8 ;
  assign n18328 = n18327 ^ n18326 ;
  assign n18330 = n18329 ^ n18328 ;
  assign n18324 = n8150 & n12928 ;
  assign n18331 = n18330 ^ n18324 ;
  assign n18333 = n18332 ^ n18331 ;
  assign n18338 = n8484 & ~n12382 ;
  assign n18337 = n8144 & n12229 ;
  assign n18339 = n18338 ^ n18337 ;
  assign n18340 = n18339 ^ x8 ;
  assign n18336 = n8150 & n13445 ;
  assign n18341 = n18340 ^ n18336 ;
  assign n18335 = n8139 & ~n12228 ;
  assign n18342 = n18341 ^ n18335 ;
  assign n18334 = n18203 ^ n17897 ;
  assign n18343 = n18342 ^ n18334 ;
  assign n18351 = n8139 & n12229 ;
  assign n18349 = n8150 & n13779 ;
  assign n18346 = n8484 & ~n12228 ;
  assign n18345 = n8144 & n12235 ;
  assign n18347 = n18346 ^ n18345 ;
  assign n18348 = n18347 ^ x8 ;
  assign n18350 = n18349 ^ n18348 ;
  assign n18352 = n18351 ^ n18350 ;
  assign n18344 = n18200 ^ n17907 ;
  assign n18353 = n18352 ^ n18344 ;
  assign n18358 = n8484 & n12229 ;
  assign n18357 = n8144 & ~n12239 ;
  assign n18359 = n18358 ^ n18357 ;
  assign n18360 = n18359 ^ x8 ;
  assign n18356 = n8150 & ~n12867 ;
  assign n18361 = n18360 ^ n18356 ;
  assign n18355 = n8139 & n12235 ;
  assign n18362 = n18361 ^ n18355 ;
  assign n18354 = n18197 ^ n17917 ;
  assign n18363 = n18362 ^ n18354 ;
  assign n18374 = n8144 & n12248 ;
  assign n18372 = n8139 & ~n12239 ;
  assign n18365 = n12235 ^ x8 ;
  assign n18366 = n18365 ^ x7 ;
  assign n18367 = n18366 ^ n12235 ;
  assign n18368 = ~n13319 & n18367 ;
  assign n18369 = n18368 ^ n12235 ;
  assign n18370 = n8137 & n18369 ;
  assign n18371 = n18370 ^ x8 ;
  assign n18373 = n18372 ^ n18371 ;
  assign n18375 = n18374 ^ n18373 ;
  assign n18364 = n18194 ^ n17927 ;
  assign n18376 = n18375 ^ n18364 ;
  assign n18390 = n18191 ^ n17937 ;
  assign n18378 = n8139 & n12248 ;
  assign n18377 = n8144 & ~n12249 ;
  assign n18379 = n18378 ^ n18377 ;
  assign n18380 = n18379 ^ n8145 ;
  assign n18381 = n18380 ^ x8 ;
  assign n18383 = ~x7 & ~n13339 ;
  assign n18386 = n18383 ^ n13343 ;
  assign n18387 = n8146 & n18386 ;
  assign n18382 = n18379 ^ x8 ;
  assign n18384 = n18383 ^ n12239 ;
  assign n18385 = n18382 & n18384 ;
  assign n18388 = n18387 ^ n18385 ;
  assign n18389 = ~n18381 & ~n18388 ;
  assign n18391 = n18390 ^ n18389 ;
  assign n18402 = n8144 & n12339 ;
  assign n18400 = n8139 & ~n12249 ;
  assign n18393 = n12248 ^ x8 ;
  assign n18394 = n18393 ^ x7 ;
  assign n18395 = n18394 ^ n12248 ;
  assign n18396 = ~n13518 & n18395 ;
  assign n18397 = n18396 ^ n12248 ;
  assign n18398 = n8137 & n18397 ;
  assign n18399 = n18398 ^ x8 ;
  assign n18401 = n18400 ^ n18399 ;
  assign n18403 = n18402 ^ n18401 ;
  assign n18392 = n18188 ^ n17947 ;
  assign n18404 = n18403 ^ n18392 ;
  assign n18407 = n8139 & n12339 ;
  assign n18406 = n8144 & ~n12251 ;
  assign n18408 = n18407 ^ n18406 ;
  assign n18409 = n18408 ^ n8145 ;
  assign n18410 = n18409 ^ x8 ;
  assign n18412 = ~x7 & ~n13553 ;
  assign n18415 = n18412 ^ n13554 ;
  assign n18416 = n8146 & n18415 ;
  assign n18411 = n18408 ^ x8 ;
  assign n18413 = n18412 ^ n12249 ;
  assign n18414 = n18411 & n18413 ;
  assign n18417 = n18416 ^ n18414 ;
  assign n18418 = ~n18410 & ~n18417 ;
  assign n18405 = n18185 ^ n17957 ;
  assign n18419 = n18418 ^ n18405 ;
  assign n18427 = n8139 & ~n12251 ;
  assign n18425 = n8150 & ~n13885 ;
  assign n18422 = n8484 & n12339 ;
  assign n18421 = n8144 & n12253 ;
  assign n18423 = n18422 ^ n18421 ;
  assign n18424 = n18423 ^ x8 ;
  assign n18426 = n18425 ^ n18424 ;
  assign n18428 = n18427 ^ n18426 ;
  assign n18420 = n18182 ^ n17967 ;
  assign n18429 = n18428 ^ n18420 ;
  assign n18440 = n8144 & n12331 ;
  assign n18438 = n8139 & n12253 ;
  assign n18431 = n12251 ^ x8 ;
  assign n18432 = n18431 ^ x7 ;
  assign n18433 = n18432 ^ n12251 ;
  assign n18434 = ~n13676 & n18433 ;
  assign n18435 = n18434 ^ n12251 ;
  assign n18436 = n8137 & ~n18435 ;
  assign n18437 = n18436 ^ x8 ;
  assign n18439 = n18438 ^ n18437 ;
  assign n18441 = n18440 ^ n18439 ;
  assign n18430 = n18179 ^ n17977 ;
  assign n18442 = n18441 ^ n18430 ;
  assign n18447 = n8484 & n12253 ;
  assign n18446 = n8144 & n12257 ;
  assign n18448 = n18447 ^ n18446 ;
  assign n18449 = n18448 ^ x8 ;
  assign n18445 = n8150 & ~n14414 ;
  assign n18450 = n18449 ^ n18445 ;
  assign n18444 = n8139 & n12331 ;
  assign n18451 = n18450 ^ n18444 ;
  assign n18443 = n18176 ^ n17987 ;
  assign n18452 = n18451 ^ n18443 ;
  assign n18455 = n8139 & n12257 ;
  assign n18454 = n8144 & ~n12258 ;
  assign n18456 = n18455 ^ n18454 ;
  assign n18457 = n18456 ^ n8145 ;
  assign n18458 = n18457 ^ x8 ;
  assign n18460 = x7 & ~n14219 ;
  assign n18463 = n18460 ^ n12331 ;
  assign n18464 = n8146 & n18463 ;
  assign n18459 = n18456 ^ x8 ;
  assign n18461 = n18460 ^ n14972 ;
  assign n18462 = n18459 & n18461 ;
  assign n18465 = n18464 ^ n18462 ;
  assign n18466 = ~n18458 & ~n18465 ;
  assign n18453 = n18173 ^ n18000 ;
  assign n18467 = n18466 ^ n18453 ;
  assign n18680 = n18170 ^ n18012 ;
  assign n18479 = n8150 & ~n14020 ;
  assign n18478 = n8139 & ~n12258 ;
  assign n18480 = n18479 ^ n18478 ;
  assign n18476 = n8484 & n12257 ;
  assign n18475 = n8144 & n12264 ;
  assign n18477 = n18476 ^ n18475 ;
  assign n18481 = n18480 ^ n18477 ;
  assign n18681 = n18680 ^ n18481 ;
  assign n18675 = n18167 ^ n18027 ;
  assign n18488 = n8484 & n12268 ;
  assign n18487 = n8144 & n12279 ;
  assign n18489 = n18488 ^ n18487 ;
  assign n18490 = n18489 ^ x8 ;
  assign n18486 = n8150 & ~n14329 ;
  assign n18491 = n18490 ^ n18486 ;
  assign n18485 = n8139 & ~n12276 ;
  assign n18492 = n18491 ^ n18485 ;
  assign n18484 = n18159 ^ n18056 ;
  assign n18493 = n18492 ^ n18484 ;
  assign n18508 = n8144 & ~n12283 ;
  assign n18506 = n8139 & n12279 ;
  assign n18499 = n12276 ^ x8 ;
  assign n18500 = n18499 ^ x7 ;
  assign n18501 = n18500 ^ n12276 ;
  assign n18502 = ~n14465 & n18501 ;
  assign n18503 = n18502 ^ n12276 ;
  assign n18504 = n8137 & ~n18503 ;
  assign n18505 = n18504 ^ x8 ;
  assign n18507 = n18506 ^ n18505 ;
  assign n18509 = n18508 ^ n18507 ;
  assign n18496 = n18148 ^ n18141 ;
  assign n18497 = n18496 ^ n18139 ;
  assign n18494 = n18140 ^ n18129 ;
  assign n18495 = n18131 & ~n18494 ;
  assign n18498 = n18497 ^ n18495 ;
  assign n18510 = n18509 ^ n18498 ;
  assign n18519 = n18140 ^ n18131 ;
  assign n18514 = n8484 & n12279 ;
  assign n18513 = n8144 & ~n12284 ;
  assign n18515 = n18514 ^ n18513 ;
  assign n18516 = n18515 ^ x8 ;
  assign n18512 = n8150 & ~n14528 ;
  assign n18517 = n18516 ^ n18512 ;
  assign n18511 = n8139 & ~n12283 ;
  assign n18518 = n18517 ^ n18511 ;
  assign n18520 = n18519 ^ n18518 ;
  assign n18529 = n8139 & ~n12284 ;
  assign n18527 = n8150 & n14548 ;
  assign n18524 = n8484 & ~n12283 ;
  assign n18523 = n8144 & ~n12285 ;
  assign n18525 = n18524 ^ n18523 ;
  assign n18526 = n18525 ^ x8 ;
  assign n18528 = n18527 ^ n18526 ;
  assign n18530 = n18529 ^ n18528 ;
  assign n18522 = n18127 ^ n18117 ;
  assign n18531 = n18530 ^ n18522 ;
  assign n18536 = n8484 & ~n12284 ;
  assign n18535 = n8144 & n12313 ;
  assign n18537 = n18536 ^ n18535 ;
  assign n18538 = n18537 ^ x8 ;
  assign n18534 = n8150 & n14584 ;
  assign n18539 = n18538 ^ n18534 ;
  assign n18533 = n8139 & ~n12285 ;
  assign n18540 = n18539 ^ n18533 ;
  assign n18532 = n18114 ^ n18104 ;
  assign n18541 = n18540 ^ n18532 ;
  assign n18547 = n8484 & ~n12285 ;
  assign n18546 = n8144 & n12289 ;
  assign n18548 = n18547 ^ n18546 ;
  assign n18549 = n18548 ^ x8 ;
  assign n18545 = n8150 & n14652 ;
  assign n18550 = n18549 ^ n18545 ;
  assign n18544 = n8139 & n12313 ;
  assign n18551 = n18550 ^ n18544 ;
  assign n18542 = n18093 ^ n18079 ;
  assign n18543 = n18542 ^ n18102 ;
  assign n18552 = n18551 ^ n18543 ;
  assign n18607 = n8144 & ~n12290 ;
  assign n18605 = n8139 & n12289 ;
  assign n18598 = n14712 ^ x8 ;
  assign n18599 = n18598 ^ x7 ;
  assign n18600 = n18599 ^ n14712 ;
  assign n18601 = ~n14711 & ~n18600 ;
  assign n18602 = n18601 ^ n14712 ;
  assign n18603 = n8137 & ~n18602 ;
  assign n18604 = n18603 ^ x8 ;
  assign n18606 = n18605 ^ n18604 ;
  assign n18608 = n18607 ^ n18606 ;
  assign n18561 = n8150 & ~n18081 ;
  assign n18567 = n8484 & n12293 ;
  assign n18564 = n8150 & n12293 ;
  assign n18565 = n18564 ^ n8144 ;
  assign n18566 = n12291 & n18565 ;
  assign n18568 = n18567 ^ n18566 ;
  assign n18569 = n18561 & ~n18568 ;
  assign n18570 = n18569 ^ n18568 ;
  assign n18571 = x8 & ~n18570 ;
  assign n18572 = ~n12298 & n19031 ;
  assign n18573 = n18571 & n18572 ;
  assign n18574 = n18573 ^ n18571 ;
  assign n18575 = n7140 & n12291 ;
  assign n18582 = n8139 & n12293 ;
  assign n18580 = n8150 & ~n14785 ;
  assign n18577 = n8484 & ~n12290 ;
  assign n18576 = n8144 & n12292 ;
  assign n18578 = n18577 ^ n18576 ;
  assign n18579 = n18578 ^ x8 ;
  assign n18581 = n18580 ^ n18579 ;
  assign n18583 = n18582 ^ n18581 ;
  assign n18584 = ~n18575 & n18583 ;
  assign n18585 = ~n18574 & n18584 ;
  assign n18586 = n18585 ^ n18583 ;
  assign n18556 = n8484 & n12289 ;
  assign n18555 = n8144 & n12293 ;
  assign n18557 = n18556 ^ n18555 ;
  assign n18558 = n18557 ^ x8 ;
  assign n18554 = n8150 & ~n14749 ;
  assign n18559 = n18558 ^ n18554 ;
  assign n18553 = n8139 & ~n12290 ;
  assign n18560 = n18559 ^ n18553 ;
  assign n18587 = n18586 ^ n18560 ;
  assign n18593 = x10 ^ x8 ;
  assign n18594 = n12291 & n18593 ;
  assign n18591 = ~x9 & n18575 ;
  assign n18589 = ~n7140 & n12292 ;
  assign n18588 = n18560 ^ n12292 ;
  assign n18590 = n18589 ^ n18588 ;
  assign n18592 = n18591 ^ n18590 ;
  assign n18595 = n18594 ^ n18592 ;
  assign n18596 = n18587 & ~n18595 ;
  assign n18597 = n18596 ^ n18586 ;
  assign n18609 = n18608 ^ n18597 ;
  assign n18610 = n18080 & n18092 ;
  assign n18615 = n18091 ^ n7142 ;
  assign n18619 = n18615 ^ n18597 ;
  assign n18616 = n18615 ^ n18091 ;
  assign n18612 = n7150 ^ n7145 ;
  assign n18613 = n12292 ^ x11 ;
  assign n18614 = n18612 & n18613 ;
  assign n18617 = n18616 ^ n18614 ;
  assign n18618 = n12299 & n18617 ;
  assign n18620 = n18619 ^ n18618 ;
  assign n18611 = n7149 & ~n12298 ;
  assign n18621 = n18620 ^ n18611 ;
  assign n18622 = n18621 ^ n18597 ;
  assign n18623 = ~n18589 & ~n18622 ;
  assign n18624 = n18610 & n18623 ;
  assign n18625 = n18624 ^ n18621 ;
  assign n18626 = n18609 & ~n18625 ;
  assign n18627 = n18626 ^ n18608 ;
  assign n18628 = n18627 ^ n18551 ;
  assign n18629 = n18552 & n18628 ;
  assign n18630 = n18629 ^ n18551 ;
  assign n18631 = n18630 ^ n18540 ;
  assign n18632 = n18541 & n18631 ;
  assign n18633 = n18632 ^ n18540 ;
  assign n18634 = n18633 ^ n18530 ;
  assign n18635 = ~n18531 & n18634 ;
  assign n18636 = n18635 ^ n18530 ;
  assign n18521 = n18518 ^ n18498 ;
  assign n18637 = n18636 ^ n18521 ;
  assign n18638 = n18637 ^ n18498 ;
  assign n18639 = ~n18520 & n18638 ;
  assign n18640 = n18639 ^ n18521 ;
  assign n18641 = ~n18510 & n18640 ;
  assign n18642 = n18641 ^ n18509 ;
  assign n18643 = n18642 ^ n18492 ;
  assign n18644 = n18493 & n18643 ;
  assign n18645 = n18644 ^ n18492 ;
  assign n18483 = n18161 ^ n18055 ;
  assign n18647 = n18645 ^ n18483 ;
  assign n18646 = ~n18483 & n18645 ;
  assign n18648 = n18647 ^ n18646 ;
  assign n18653 = n8150 & n14452 ;
  assign n18652 = n8139 & n12268 ;
  assign n18654 = n18653 ^ n18652 ;
  assign n18650 = n8484 & ~n12267 ;
  assign n18649 = n8144 & ~n12276 ;
  assign n18651 = n18650 ^ n18649 ;
  assign n18655 = n18654 ^ n18651 ;
  assign n18656 = n18655 ^ x8 ;
  assign n18664 = n18165 ^ n18038 ;
  assign n18665 = n18664 ^ n18655 ;
  assign n18661 = n8150 & ~n14429 ;
  assign n18660 = n8139 & ~n12267 ;
  assign n18662 = n18661 ^ n18660 ;
  assign n18658 = n8484 & n12264 ;
  assign n18657 = n8144 & n12268 ;
  assign n18659 = n18658 ^ n18657 ;
  assign n18663 = n18662 ^ n18659 ;
  assign n18666 = n18665 ^ n18663 ;
  assign n18667 = n18656 & n18666 ;
  assign n18668 = ~n18648 & n18667 ;
  assign n18669 = n18664 ^ n18646 ;
  assign n18670 = n18663 ^ x8 ;
  assign n18671 = n18670 ^ n18646 ;
  assign n18672 = ~n18669 & n18671 ;
  assign n18673 = n18672 ^ n18646 ;
  assign n18674 = ~n18668 & ~n18673 ;
  assign n18676 = n18675 ^ n18674 ;
  assign n18688 = n18674 ^ n18481 ;
  assign n18472 = n8150 & n14243 ;
  assign n18471 = n8139 & n12264 ;
  assign n18473 = n18472 ^ n18471 ;
  assign n18469 = n8484 & ~n12258 ;
  assign n18468 = n8144 & ~n12267 ;
  assign n18470 = n18469 ^ n18468 ;
  assign n18474 = n18473 ^ n18470 ;
  assign n18482 = n18481 ^ n18474 ;
  assign n18689 = n18688 ^ n18482 ;
  assign n18690 = ~n18676 & ~n18689 ;
  assign n18691 = n18690 ^ n18482 ;
  assign n18692 = ~n18681 & n18691 ;
  assign n18693 = n18692 ^ n18481 ;
  assign n18682 = n18681 ^ n18474 ;
  assign n18679 = n18675 ^ n18482 ;
  assign n18683 = n18682 ^ n18679 ;
  assign n18684 = n18683 ^ n18482 ;
  assign n18685 = ~n18676 & ~n18684 ;
  assign n18686 = n18685 ^ n18482 ;
  assign n18687 = x8 & ~n18686 ;
  assign n18694 = n18693 ^ n18687 ;
  assign n18695 = n18694 ^ n18466 ;
  assign n18696 = ~n18467 & ~n18695 ;
  assign n18697 = n18696 ^ n18466 ;
  assign n18698 = n18697 ^ n18451 ;
  assign n18699 = n18452 & ~n18698 ;
  assign n18700 = n18699 ^ n18451 ;
  assign n18701 = n18700 ^ n18441 ;
  assign n18702 = ~n18442 & n18701 ;
  assign n18703 = n18702 ^ n18441 ;
  assign n18704 = n18703 ^ n18428 ;
  assign n18705 = ~n18429 & n18704 ;
  assign n18706 = n18705 ^ n18428 ;
  assign n18707 = n18706 ^ n18418 ;
  assign n18708 = ~n18419 & ~n18707 ;
  assign n18709 = n18708 ^ n18418 ;
  assign n18710 = n18709 ^ n18403 ;
  assign n18711 = ~n18404 & ~n18710 ;
  assign n18712 = n18711 ^ n18403 ;
  assign n18713 = n18712 ^ n18389 ;
  assign n18714 = ~n18391 & ~n18713 ;
  assign n18715 = n18714 ^ n18389 ;
  assign n18716 = n18715 ^ n18375 ;
  assign n18717 = n18376 & ~n18716 ;
  assign n18718 = n18717 ^ n18375 ;
  assign n18719 = n18718 ^ n18362 ;
  assign n18720 = n18363 & n18719 ;
  assign n18721 = n18720 ^ n18362 ;
  assign n18722 = n18721 ^ n18352 ;
  assign n18723 = n18353 & n18722 ;
  assign n18724 = n18723 ^ n18352 ;
  assign n18725 = n18724 ^ n18342 ;
  assign n18726 = n18343 & n18725 ;
  assign n18727 = n18726 ^ n18342 ;
  assign n18728 = n18727 ^ n18325 ;
  assign n18729 = n18333 & n18728 ;
  assign n18730 = n18729 ^ n18325 ;
  assign n18731 = n18730 ^ n18317 ;
  assign n18732 = ~n18323 & ~n18731 ;
  assign n18733 = n18732 ^ n18317 ;
  assign n18734 = n18733 ^ n18312 ;
  assign n18735 = n18313 & n18734 ;
  assign n18736 = n18735 ^ n18312 ;
  assign n18292 = n18225 ^ n18215 ;
  assign n18737 = n18736 ^ n18292 ;
  assign n18745 = n8139 & n12222 ;
  assign n18741 = n18292 ^ x8 ;
  assign n18740 = n8484 & ~n12214 ;
  assign n18742 = n18741 ^ n18740 ;
  assign n18739 = n8144 & n12380 ;
  assign n18743 = n18742 ^ n18739 ;
  assign n18738 = n8150 & n12608 ;
  assign n18744 = n18743 ^ n18738 ;
  assign n18746 = n18745 ^ n18744 ;
  assign n18747 = ~n18737 & ~n18746 ;
  assign n18748 = n18747 ^ n18736 ;
  assign n18749 = n18748 ^ n18290 ;
  assign n18750 = ~n18291 & ~n18749 ;
  assign n18751 = n18750 ^ n18290 ;
  assign n18277 = n8139 & ~n12400 ;
  assign n18272 = n18230 ^ n17841 ;
  assign n18273 = n18272 ^ x8 ;
  assign n18271 = n8484 & ~n12210 ;
  assign n18274 = n18273 ^ n18271 ;
  assign n18270 = n8144 & ~n12214 ;
  assign n18275 = n18274 ^ n18270 ;
  assign n18269 = n8150 & n12737 ;
  assign n18276 = n18275 ^ n18269 ;
  assign n18278 = n18277 ^ n18276 ;
  assign n18770 = n18751 ^ n18278 ;
  assign n18784 = n18783 ^ n18770 ;
  assign n18793 = ~n10334 & ~n12210 ;
  assign n18790 = n10327 & ~n12405 ;
  assign n18788 = n10425 & n12419 ;
  assign n18786 = n18748 ^ n18291 ;
  assign n18787 = n18786 ^ x5 ;
  assign n18789 = n18788 ^ n18787 ;
  assign n18791 = n18790 ^ n18789 ;
  assign n18785 = n10342 & ~n12651 ;
  assign n18792 = n18791 ^ n18785 ;
  assign n18794 = n18793 ^ n18792 ;
  assign n18803 = n10342 & n12737 ;
  assign n18799 = n18733 ^ n18313 ;
  assign n18800 = n18799 ^ x5 ;
  assign n18798 = n10425 & ~n12210 ;
  assign n18801 = n18800 ^ n18798 ;
  assign n18797 = n10327 & ~n12400 ;
  assign n18802 = n18801 ^ n18797 ;
  assign n18804 = n18803 ^ n18802 ;
  assign n18796 = ~n10334 & ~n12214 ;
  assign n18805 = n18804 ^ n18796 ;
  assign n18813 = ~n10334 & n12222 ;
  assign n18811 = n10342 & n12667 ;
  assign n18808 = n10425 & ~n12400 ;
  assign n18807 = n10327 & ~n12214 ;
  assign n18809 = n18808 ^ n18807 ;
  assign n18810 = n18809 ^ x5 ;
  assign n18812 = n18811 ^ n18810 ;
  assign n18814 = n18813 ^ n18812 ;
  assign n18806 = n18730 ^ n18323 ;
  assign n18815 = n18814 ^ n18806 ;
  assign n18824 = ~n10334 & n12380 ;
  assign n18821 = n10327 & n12222 ;
  assign n18819 = n10425 & ~n12214 ;
  assign n18817 = n18727 ^ n18333 ;
  assign n18818 = n18817 ^ x5 ;
  assign n18820 = n18819 ^ n18818 ;
  assign n18822 = n18821 ^ n18820 ;
  assign n18816 = n10342 & n12608 ;
  assign n18823 = n18822 ^ n18816 ;
  assign n18825 = n18824 ^ n18823 ;
  assign n18830 = n10425 & n12222 ;
  assign n18829 = n10327 & n12380 ;
  assign n18831 = n18830 ^ n18829 ;
  assign n18832 = n18831 ^ x5 ;
  assign n18828 = n10342 & n13770 ;
  assign n18833 = n18832 ^ n18828 ;
  assign n18827 = ~n10334 & n12376 ;
  assign n18834 = n18833 ^ n18827 ;
  assign n18826 = n18724 ^ n18343 ;
  assign n18835 = n18834 ^ n18826 ;
  assign n19212 = n18718 ^ n18363 ;
  assign n18845 = n18715 ^ n18376 ;
  assign n18841 = n10342 & n13445 ;
  assign n18840 = ~n10334 & n12229 ;
  assign n18842 = n18841 ^ n18840 ;
  assign n18838 = n10425 & ~n12382 ;
  assign n18837 = n10327 & ~n12228 ;
  assign n18839 = n18838 ^ n18837 ;
  assign n18843 = n18842 ^ n18839 ;
  assign n18844 = n18843 ^ x5 ;
  assign n18846 = n18845 ^ n18844 ;
  assign n19196 = n18712 ^ n18391 ;
  assign n19208 = n19196 ^ n18845 ;
  assign n18851 = n10425 & n12229 ;
  assign n18850 = n10327 & n12235 ;
  assign n18852 = n18851 ^ n18850 ;
  assign n18853 = n18852 ^ x5 ;
  assign n18849 = n10342 & ~n12867 ;
  assign n18854 = n18853 ^ n18849 ;
  assign n18848 = ~n10334 & ~n12239 ;
  assign n18855 = n18854 ^ n18848 ;
  assign n18847 = n18709 ^ n18404 ;
  assign n18856 = n18855 ^ n18847 ;
  assign n18864 = ~n10334 & n12248 ;
  assign n18862 = n10342 & ~n13329 ;
  assign n18859 = n10425 & n12235 ;
  assign n18858 = n10327 & ~n12239 ;
  assign n18860 = n18859 ^ n18858 ;
  assign n18861 = n18860 ^ x5 ;
  assign n18863 = n18862 ^ n18861 ;
  assign n18865 = n18864 ^ n18863 ;
  assign n18857 = n18706 ^ n18419 ;
  assign n18866 = n18865 ^ n18857 ;
  assign n18874 = n18703 ^ n18429 ;
  assign n18875 = n18874 ^ x5 ;
  assign n18873 = ~n10334 & ~n12249 ;
  assign n18876 = n18875 ^ n18873 ;
  assign n18872 = n10327 & n12248 ;
  assign n18877 = n18876 ^ n18872 ;
  assign n18867 = n12239 ^ n10329 ;
  assign n18868 = n18867 ^ n12239 ;
  assign n18869 = ~n13339 & n18868 ;
  assign n18870 = n18869 ^ n12239 ;
  assign n18871 = n10322 & ~n18870 ;
  assign n18878 = n18877 ^ n18871 ;
  assign n18889 = ~n10334 & n12339 ;
  assign n18887 = n10327 & ~n12249 ;
  assign n18880 = n12248 ^ x5 ;
  assign n18881 = n18880 ^ x4 ;
  assign n18882 = n18881 ^ n12248 ;
  assign n18883 = ~n13518 & n18882 ;
  assign n18884 = n18883 ^ n12248 ;
  assign n18885 = n10322 & n18884 ;
  assign n18886 = n18885 ^ x5 ;
  assign n18888 = n18887 ^ n18886 ;
  assign n18890 = n18889 ^ n18888 ;
  assign n18879 = n18700 ^ n18442 ;
  assign n18891 = n18890 ^ n18879 ;
  assign n18896 = n10425 & ~n12249 ;
  assign n18895 = n10327 & n12339 ;
  assign n18897 = n18896 ^ n18895 ;
  assign n18898 = n18897 ^ x5 ;
  assign n18894 = n10342 & n13554 ;
  assign n18899 = n18898 ^ n18894 ;
  assign n18893 = ~n10334 & ~n12251 ;
  assign n18900 = n18899 ^ n18893 ;
  assign n18892 = n18697 ^ n18452 ;
  assign n18901 = n18900 ^ n18892 ;
  assign n18909 = ~n10334 & n12253 ;
  assign n18907 = n10342 & ~n13885 ;
  assign n18904 = n10425 & n12339 ;
  assign n18903 = n10327 & ~n12251 ;
  assign n18905 = n18904 ^ n18903 ;
  assign n18906 = n18905 ^ x5 ;
  assign n18908 = n18907 ^ n18906 ;
  assign n18910 = n18909 ^ n18908 ;
  assign n18902 = n18694 ^ n18467 ;
  assign n18911 = n18910 ^ n18902 ;
  assign n18926 = n10425 & n12253 ;
  assign n18925 = n10327 & n12331 ;
  assign n18927 = n18926 ^ n18925 ;
  assign n18928 = n18927 ^ x5 ;
  assign n18924 = n10342 & ~n14414 ;
  assign n18929 = n18928 ^ n18924 ;
  assign n18923 = ~n10334 & n12257 ;
  assign n18930 = n18929 ^ n18923 ;
  assign n18920 = n18675 ^ n18474 ;
  assign n18921 = n18920 ^ x8 ;
  assign n18922 = n18921 ^ n18674 ;
  assign n18931 = n18930 ^ n18922 ;
  assign n18947 = ~n10334 & n12264 ;
  assign n18945 = n10342 & ~n14020 ;
  assign n18942 = n10425 & n12257 ;
  assign n18941 = n10327 & ~n12258 ;
  assign n18943 = n18942 ^ n18941 ;
  assign n18944 = n18943 ^ x5 ;
  assign n18946 = n18945 ^ n18944 ;
  assign n18948 = n18947 ^ n18946 ;
  assign n18940 = n18656 ^ n18647 ;
  assign n18949 = n18948 ^ n18940 ;
  assign n18957 = ~n10334 & ~n12267 ;
  assign n18955 = n10342 & n14243 ;
  assign n18952 = n10425 & ~n12258 ;
  assign n18951 = n10327 & n12264 ;
  assign n18953 = n18952 ^ n18951 ;
  assign n18954 = n18953 ^ x5 ;
  assign n18956 = n18955 ^ n18954 ;
  assign n18958 = n18957 ^ n18956 ;
  assign n18950 = n18642 ^ n18493 ;
  assign n18959 = n18958 ^ n18950 ;
  assign n18967 = ~n10334 & n12268 ;
  assign n18965 = n10342 & ~n14429 ;
  assign n18962 = n10425 & n12264 ;
  assign n18961 = n10327 & ~n12267 ;
  assign n18963 = n18962 ^ n18961 ;
  assign n18964 = n18963 ^ x5 ;
  assign n18966 = n18965 ^ n18964 ;
  assign n18968 = n18967 ^ n18966 ;
  assign n18960 = n18640 ^ n18509 ;
  assign n18969 = n18968 ^ n18960 ;
  assign n18974 = n10425 & ~n12267 ;
  assign n18973 = n10327 & n12268 ;
  assign n18975 = n18974 ^ n18973 ;
  assign n18976 = n18975 ^ x5 ;
  assign n18972 = n10342 & n14452 ;
  assign n18977 = n18976 ^ n18972 ;
  assign n18971 = ~n10334 & ~n12276 ;
  assign n18978 = n18977 ^ n18971 ;
  assign n18970 = n18636 ^ n18520 ;
  assign n18979 = n18978 ^ n18970 ;
  assign n18984 = n10327 & ~n12276 ;
  assign n18983 = n10425 & n12268 ;
  assign n18985 = n18984 ^ n18983 ;
  assign n18986 = n18985 ^ x5 ;
  assign n18982 = n10342 & ~n14329 ;
  assign n18987 = n18986 ^ n18982 ;
  assign n18981 = ~n10334 & n12279 ;
  assign n18988 = n18987 ^ n18981 ;
  assign n18980 = n18633 ^ n18531 ;
  assign n18989 = n18988 ^ n18980 ;
  assign n18997 = ~n10334 & ~n12283 ;
  assign n18995 = n10342 & n14475 ;
  assign n18992 = n10425 & ~n12276 ;
  assign n18991 = n10327 & n12279 ;
  assign n18993 = n18992 ^ n18991 ;
  assign n18994 = n18993 ^ x5 ;
  assign n18996 = n18995 ^ n18994 ;
  assign n18998 = n18997 ^ n18996 ;
  assign n18990 = n18630 ^ n18541 ;
  assign n18999 = n18998 ^ n18990 ;
  assign n19127 = n10342 & ~n14528 ;
  assign n19126 = ~n10334 & ~n12284 ;
  assign n19128 = n19127 ^ n19126 ;
  assign n19124 = n10425 & n12279 ;
  assign n19123 = n10327 & ~n12283 ;
  assign n19125 = n19124 ^ n19123 ;
  assign n19129 = n19128 ^ n19125 ;
  assign n19118 = n18627 ^ n18552 ;
  assign n19137 = n19129 ^ n19118 ;
  assign n19004 = n10425 & ~n12284 ;
  assign n19003 = n10327 & ~n12285 ;
  assign n19005 = n19004 ^ n19003 ;
  assign n19006 = n19005 ^ x5 ;
  assign n19002 = n10342 & n14584 ;
  assign n19007 = n19006 ^ n19002 ;
  assign n19001 = ~n10334 & n12313 ;
  assign n19008 = n19007 ^ n19001 ;
  assign n19000 = n18595 ^ n18586 ;
  assign n19009 = n19008 ^ n19000 ;
  assign n19015 = n10327 & n12313 ;
  assign n19014 = n10425 & ~n12285 ;
  assign n19016 = n19015 ^ n19014 ;
  assign n19017 = n19016 ^ x5 ;
  assign n19013 = n10342 & n14652 ;
  assign n19018 = n19017 ^ n19013 ;
  assign n19012 = ~n10334 & n12289 ;
  assign n19019 = n19018 ^ n19012 ;
  assign n19010 = n18575 ^ n18574 ;
  assign n19011 = n19010 ^ n18583 ;
  assign n19020 = n19019 ^ n19011 ;
  assign n19037 = n13607 ^ n8146 ;
  assign n19038 = n12292 & n19037 ;
  assign n19032 = n12291 & n19031 ;
  assign n19033 = n19032 ^ n8137 ;
  assign n19034 = ~n12292 & n19033 ;
  assign n19035 = n19034 ^ n8137 ;
  assign n19036 = n18571 & n19035 ;
  assign n19039 = n19038 ^ n19036 ;
  assign n19044 = n8145 ^ n8139 ;
  assign n19045 = ~n12292 & n19044 ;
  assign n19046 = n19045 ^ n8139 ;
  assign n19047 = ~n12291 & n19046 ;
  assign n19042 = n18570 ^ n8145 ;
  assign n19048 = n19047 ^ n19042 ;
  assign n19049 = ~n19039 & ~n19048 ;
  assign n19027 = ~n10334 & ~n12290 ;
  assign n19025 = n10342 & ~n14712 ;
  assign n19022 = n10425 & n12313 ;
  assign n19021 = n10327 & n12289 ;
  assign n19023 = n19022 ^ n19021 ;
  assign n19024 = n19023 ^ x5 ;
  assign n19026 = n19025 ^ n19024 ;
  assign n19028 = n19027 ^ n19026 ;
  assign n19050 = n19049 ^ n19028 ;
  assign n19083 = n10425 & n12289 ;
  assign n19082 = n10327 & ~n12290 ;
  assign n19084 = n19083 ^ n19082 ;
  assign n19085 = n19084 ^ x5 ;
  assign n19081 = n10342 & ~n14749 ;
  assign n19086 = n19085 ^ n19081 ;
  assign n19080 = ~n10334 & n12293 ;
  assign n19087 = n19086 ^ n19080 ;
  assign n19073 = n10342 & ~n14785 ;
  assign n19072 = ~n10334 & n12292 ;
  assign n19074 = n19073 ^ n19072 ;
  assign n19070 = n10425 & ~n12290 ;
  assign n19069 = n10327 & n12293 ;
  assign n19071 = n19070 ^ n19069 ;
  assign n19075 = n19074 ^ n19071 ;
  assign n19054 = n10322 & n12292 ;
  assign n19055 = x5 & ~n19054 ;
  assign n19056 = n12291 & n19055 ;
  assign n19057 = n10333 & n19056 ;
  assign n19058 = n19057 ^ n19055 ;
  assign n19065 = n10342 & ~n12299 ;
  assign n19064 = ~n10334 & n12291 ;
  assign n19066 = n19065 ^ n19064 ;
  assign n19062 = n10322 & n12293 ;
  assign n19061 = n10327 & n12292 ;
  assign n19063 = n19062 ^ n19061 ;
  assign n19067 = n19066 ^ n19063 ;
  assign n19068 = n19058 & ~n19067 ;
  assign n19076 = n19075 ^ n19068 ;
  assign n19051 = n8137 & ~n12291 ;
  assign n19052 = n19051 ^ n8137 ;
  assign n19077 = n19068 ^ n19052 ;
  assign n19078 = n19076 & n19077 ;
  assign n19053 = x5 & n19052 ;
  assign n19079 = n19078 ^ n19053 ;
  assign n19088 = n19087 ^ n19079 ;
  assign n19093 = n8137 & n12292 ;
  assign n19090 = x7 ^ x5 ;
  assign n19091 = n12291 & n19090 ;
  assign n19089 = n19087 ^ n19053 ;
  assign n19092 = n19091 ^ n19089 ;
  assign n19094 = n19093 ^ n19092 ;
  assign n19095 = n19088 & n19094 ;
  assign n19096 = n19095 ^ n19087 ;
  assign n19097 = n19096 ^ n19028 ;
  assign n19098 = ~n19050 & ~n19097 ;
  assign n19099 = n19098 ^ n19049 ;
  assign n19100 = n19099 ^ n19011 ;
  assign n19101 = n19020 & n19100 ;
  assign n19102 = n19101 ^ n19019 ;
  assign n19103 = n19102 ^ n19008 ;
  assign n19104 = n19009 & n19103 ;
  assign n19105 = n19104 ^ n19008 ;
  assign n19119 = n19118 ^ n19105 ;
  assign n19112 = n10342 & n14548 ;
  assign n19111 = ~n10334 & ~n12285 ;
  assign n19113 = n19112 ^ n19111 ;
  assign n19109 = n10425 & ~n12283 ;
  assign n19108 = n10327 & ~n12284 ;
  assign n19110 = n19109 ^ n19108 ;
  assign n19114 = n19113 ^ n19110 ;
  assign n19115 = n19114 ^ x5 ;
  assign n19106 = n18625 ^ n18608 ;
  assign n19116 = ~n19105 & n19106 ;
  assign n19117 = n19115 & n19116 ;
  assign n19120 = n19119 ^ n19117 ;
  assign n19107 = n19105 & ~n19106 ;
  assign n19121 = n19120 ^ n19107 ;
  assign n19122 = n19121 ^ n19120 ;
  assign n19131 = n19120 ^ n19114 ;
  assign n19138 = n19131 ^ n19120 ;
  assign n19139 = n19122 & ~n19138 ;
  assign n19140 = n19139 ^ n19120 ;
  assign n19141 = n19137 & ~n19140 ;
  assign n19142 = n19141 ^ n19129 ;
  assign n19130 = n19129 ^ n19120 ;
  assign n19132 = n19131 ^ n19130 ;
  assign n19133 = n19132 ^ n19120 ;
  assign n19134 = n19122 & ~n19133 ;
  assign n19135 = n19134 ^ n19120 ;
  assign n19136 = x5 & n19135 ;
  assign n19143 = n19142 ^ n19136 ;
  assign n19144 = n19143 ^ n18990 ;
  assign n19145 = n18999 & ~n19144 ;
  assign n19146 = n19145 ^ n18998 ;
  assign n19147 = n19146 ^ n18980 ;
  assign n19148 = ~n18989 & n19147 ;
  assign n19149 = n19148 ^ n18988 ;
  assign n19150 = n19149 ^ n18978 ;
  assign n19151 = ~n18979 & n19150 ;
  assign n19152 = n19151 ^ n18978 ;
  assign n19153 = n19152 ^ n18960 ;
  assign n19154 = ~n18969 & n19153 ;
  assign n19155 = n19154 ^ n18968 ;
  assign n19156 = n19155 ^ n18950 ;
  assign n19157 = n18959 & ~n19156 ;
  assign n19158 = n19157 ^ n18958 ;
  assign n19159 = n19158 ^ n18948 ;
  assign n19160 = ~n18949 & n19159 ;
  assign n19161 = n19160 ^ n18948 ;
  assign n18938 = ~n10334 & ~n12258 ;
  assign n18936 = n10342 & ~n14972 ;
  assign n18933 = n10425 & n12331 ;
  assign n18932 = n10327 & n12257 ;
  assign n18934 = n18933 ^ n18932 ;
  assign n18935 = n18934 ^ x5 ;
  assign n18937 = n18936 ^ n18935 ;
  assign n18939 = n18938 ^ n18937 ;
  assign n19162 = n19161 ^ n18939 ;
  assign n19165 = n18939 ^ n18666 ;
  assign n19163 = n18656 ^ n18645 ;
  assign n19164 = n18647 & n19163 ;
  assign n19166 = n19165 ^ n19164 ;
  assign n19167 = n19162 & n19166 ;
  assign n19168 = n19167 ^ n19161 ;
  assign n19169 = n19168 ^ n18930 ;
  assign n19170 = n18931 & n19169 ;
  assign n19171 = n19170 ^ n18930 ;
  assign n18915 = n10425 & ~n12251 ;
  assign n18914 = n10327 & n12253 ;
  assign n18916 = n18915 ^ n18914 ;
  assign n18917 = n18916 ^ x5 ;
  assign n18913 = n10342 & n13677 ;
  assign n18918 = n18917 ^ n18913 ;
  assign n18912 = ~n10334 & n12331 ;
  assign n18919 = n18918 ^ n18912 ;
  assign n19172 = n19171 ^ n18919 ;
  assign n19174 = n18919 ^ n18682 ;
  assign n19173 = ~n18676 & ~n18921 ;
  assign n19175 = n19174 ^ n19173 ;
  assign n19176 = n19172 & n19175 ;
  assign n19177 = n19176 ^ n19171 ;
  assign n19178 = n19177 ^ n18910 ;
  assign n19179 = ~n18911 & n19178 ;
  assign n19180 = n19179 ^ n18910 ;
  assign n19181 = n19180 ^ n18900 ;
  assign n19182 = ~n18901 & n19181 ;
  assign n19183 = n19182 ^ n18900 ;
  assign n19184 = n19183 ^ n18879 ;
  assign n19185 = ~n18891 & n19184 ;
  assign n19186 = n19185 ^ n18890 ;
  assign n19187 = n19186 ^ n18874 ;
  assign n19188 = ~n18878 & ~n19187 ;
  assign n19189 = n19188 ^ n18874 ;
  assign n19190 = n19189 ^ n18865 ;
  assign n19191 = ~n18866 & ~n19190 ;
  assign n19192 = n19191 ^ n18865 ;
  assign n19193 = n19192 ^ n18855 ;
  assign n19194 = n18856 & n19193 ;
  assign n19195 = n19194 ^ n18855 ;
  assign n19197 = n19196 ^ n19195 ;
  assign n19205 = ~n10334 & n12235 ;
  assign n19201 = n19196 ^ x5 ;
  assign n19200 = n10425 & ~n12228 ;
  assign n19202 = n19201 ^ n19200 ;
  assign n19199 = n10327 & n12229 ;
  assign n19203 = n19202 ^ n19199 ;
  assign n19198 = n10342 & n13779 ;
  assign n19204 = n19203 ^ n19198 ;
  assign n19206 = n19205 ^ n19204 ;
  assign n19207 = ~n19197 & ~n19206 ;
  assign n19209 = n19208 ^ n19207 ;
  assign n19210 = ~n18846 & n19209 ;
  assign n19211 = n19210 ^ n18845 ;
  assign n19213 = n19212 ^ n19211 ;
  assign n19218 = n10342 & n12928 ;
  assign n19217 = ~n10334 & ~n12228 ;
  assign n19219 = n19218 ^ n19217 ;
  assign n19215 = n10425 & n12376 ;
  assign n19214 = n10327 & ~n12382 ;
  assign n19216 = n19215 ^ n19214 ;
  assign n19220 = n19219 ^ n19216 ;
  assign n19221 = n19220 ^ x5 ;
  assign n19222 = n19221 ^ n19211 ;
  assign n19223 = ~n19213 & n19222 ;
  assign n19224 = n19223 ^ n19212 ;
  assign n18836 = n18721 ^ n18353 ;
  assign n19225 = n19224 ^ n18836 ;
  assign n19233 = ~n10334 & ~n12382 ;
  assign n19229 = n18836 ^ x5 ;
  assign n19228 = n10425 & n12380 ;
  assign n19230 = n19229 ^ n19228 ;
  assign n19227 = n10327 & n12376 ;
  assign n19231 = n19230 ^ n19227 ;
  assign n19226 = n10342 & n12555 ;
  assign n19232 = n19231 ^ n19226 ;
  assign n19234 = n19233 ^ n19232 ;
  assign n19235 = n19225 & ~n19234 ;
  assign n19236 = n19235 ^ n19224 ;
  assign n19237 = n19236 ^ n18826 ;
  assign n19238 = n18835 & ~n19237 ;
  assign n19239 = n19238 ^ n18834 ;
  assign n19240 = n19239 ^ n18817 ;
  assign n19241 = n18825 & n19240 ;
  assign n19242 = n19241 ^ n18817 ;
  assign n19243 = n19242 ^ n18806 ;
  assign n19244 = ~n18815 & n19243 ;
  assign n19245 = n19244 ^ n18814 ;
  assign n19246 = n19245 ^ n18799 ;
  assign n19247 = ~n18805 & ~n19246 ;
  assign n19248 = n19247 ^ n18799 ;
  assign n18795 = n18746 ^ n18736 ;
  assign n19249 = n19248 ^ n18795 ;
  assign n19258 = ~n10334 & ~n12400 ;
  assign n19256 = n10327 & ~n12210 ;
  assign n19255 = n18795 ^ x5 ;
  assign n19257 = n19256 ^ n19255 ;
  assign n19259 = n19258 ^ n19257 ;
  assign n19250 = n12405 ^ n10329 ;
  assign n19251 = n19250 ^ n12405 ;
  assign n19252 = ~n12714 & n19251 ;
  assign n19253 = n19252 ^ n12405 ;
  assign n19254 = n10322 & ~n19253 ;
  assign n19260 = n19259 ^ n19254 ;
  assign n19261 = n19249 & n19260 ;
  assign n19262 = n19261 ^ n19248 ;
  assign n19263 = n19262 ^ n18786 ;
  assign n19264 = n18794 & ~n19263 ;
  assign n19265 = n19264 ^ n18786 ;
  assign n19266 = n19265 ^ n18770 ;
  assign n19267 = ~n18784 & n19266 ;
  assign n19268 = n19267 ^ n18770 ;
  assign n18768 = ~n10334 & n12419 ;
  assign n18765 = n10327 & ~n12209 ;
  assign n18763 = n10425 & ~n12204 ;
  assign n18752 = n18751 ^ n18272 ;
  assign n18753 = n18278 & n18752 ;
  assign n18754 = n18753 ^ n18272 ;
  assign n18267 = n8139 & ~n12210 ;
  assign n18262 = n18233 ^ n17831 ;
  assign n18263 = n18262 ^ x8 ;
  assign n18261 = n8484 & ~n12405 ;
  assign n18264 = n18263 ^ n18261 ;
  assign n18260 = n8144 & ~n12400 ;
  assign n18265 = n18264 ^ n18260 ;
  assign n18259 = n8150 & n12715 ;
  assign n18266 = n18265 ^ n18259 ;
  assign n18268 = n18267 ^ n18266 ;
  assign n18761 = n18754 ^ n18268 ;
  assign n18762 = n18761 ^ x5 ;
  assign n18764 = n18763 ^ n18762 ;
  assign n18766 = n18765 ^ n18764 ;
  assign n18760 = n10342 & n12983 ;
  assign n18767 = n18766 ^ n18760 ;
  assign n18769 = n18768 ^ n18767 ;
  assign n19269 = n19268 ^ n18769 ;
  assign n19270 = n19269 ^ n14032 ;
  assign n18759 = n11139 & n12435 ;
  assign n19271 = n19270 ^ n18759 ;
  assign n19284 = n19265 ^ n18784 ;
  assign n19279 = n11012 & n14140 ;
  assign n19280 = n19279 ^ x1 ;
  assign n19285 = n19284 ^ n19280 ;
  assign n19274 = n12435 ^ x2 ;
  assign n19281 = n19280 ^ n19274 ;
  assign n19272 = n12435 ^ n12204 ;
  assign n19273 = n19272 ^ n12435 ;
  assign n19275 = n19274 ^ n12435 ;
  assign n19276 = ~n19273 & n19275 ;
  assign n19277 = n19276 ^ n12435 ;
  assign n19278 = ~x1 & ~n19277 ;
  assign n19282 = n19281 ^ n19278 ;
  assign n19283 = ~x0 & n19282 ;
  assign n19286 = n19285 ^ n19283 ;
  assign n19294 = n12204 ^ x2 ;
  assign n19289 = n19274 ^ x1 ;
  assign n19290 = n12432 & n19289 ;
  assign n19291 = n19290 ^ n19274 ;
  assign n19295 = n19294 ^ n19291 ;
  assign n19296 = n19295 ^ n19291 ;
  assign n19297 = n19296 ^ n12204 ;
  assign n19298 = ~n12209 & n19297 ;
  assign n19299 = n19298 ^ n12204 ;
  assign n19300 = ~x1 & ~n19299 ;
  assign n19301 = n19300 ^ n19295 ;
  assign n19302 = ~x0 & n19301 ;
  assign n19303 = n19302 ^ n19291 ;
  assign n19287 = n19262 ^ n18794 ;
  assign n19304 = n19303 ^ n19287 ;
  assign n19324 = n12405 ^ x2 ;
  assign n19327 = n19324 ^ n12405 ;
  assign n19328 = ~n15596 & n19327 ;
  assign n19329 = n19328 ^ n12405 ;
  assign n19330 = ~x1 & ~n19329 ;
  assign n19319 = n12419 ^ x1 ;
  assign n19320 = n19319 ^ x2 ;
  assign n19321 = n19320 ^ n12419 ;
  assign n19322 = n12650 & n19321 ;
  assign n19323 = n19322 ^ n19319 ;
  assign n19325 = n19324 ^ n19323 ;
  assign n19331 = n19330 ^ n19325 ;
  assign n19332 = ~x0 & ~n19331 ;
  assign n19333 = n19332 ^ n19323 ;
  assign n19342 = n12210 ^ x2 ;
  assign n19345 = n19342 ^ n12210 ;
  assign n19346 = ~n12400 & n19345 ;
  assign n19347 = n19346 ^ n12210 ;
  assign n19348 = ~x1 & ~n19347 ;
  assign n19335 = n12405 ^ x1 ;
  assign n19336 = n19335 ^ x2 ;
  assign n19337 = n19336 ^ n12405 ;
  assign n19338 = n12714 & n19337 ;
  assign n19339 = n19338 ^ n19335 ;
  assign n19343 = n19342 ^ n19339 ;
  assign n19349 = n19348 ^ n19343 ;
  assign n19350 = ~x0 & n19349 ;
  assign n19351 = n19350 ^ n19339 ;
  assign n19334 = n19239 ^ n18825 ;
  assign n19352 = n19351 ^ n19334 ;
  assign n19368 = n19236 ^ n18835 ;
  assign n20041 = n19368 ^ n19351 ;
  assign n19357 = n15959 ^ n12400 ;
  assign n19358 = n12400 ^ x2 ;
  assign n19361 = n19358 ^ n15959 ;
  assign n19362 = ~n19357 & ~n19361 ;
  assign n19363 = n19362 ^ n15959 ;
  assign n19364 = ~x1 & n19363 ;
  assign n19353 = n12210 ^ x1 ;
  assign n19354 = n19353 ^ n19342 ;
  assign n19355 = n12736 & n19354 ;
  assign n19356 = n19355 ^ n19353 ;
  assign n19359 = n19358 ^ n19356 ;
  assign n19365 = n19364 ^ n19359 ;
  assign n19366 = ~x0 & n19365 ;
  assign n19367 = n19366 ^ n19356 ;
  assign n19369 = n19368 ^ n19367 ;
  assign n19376 = n15994 ^ n12214 ;
  assign n19377 = n12214 ^ x2 ;
  assign n19380 = n19377 ^ n12214 ;
  assign n19381 = n19376 & n19380 ;
  assign n19382 = n19381 ^ n12214 ;
  assign n19383 = ~x1 & ~n19382 ;
  assign n19371 = n12400 ^ x1 ;
  assign n19372 = n19371 ^ x2 ;
  assign n19373 = n19372 ^ n12400 ;
  assign n19374 = n12666 & n19373 ;
  assign n19375 = n19374 ^ n19371 ;
  assign n19378 = n19377 ^ n19375 ;
  assign n19384 = n19383 ^ n19378 ;
  assign n19385 = ~x0 & n19384 ;
  assign n19386 = n19385 ^ n19375 ;
  assign n19370 = n19234 ^ n19224 ;
  assign n19387 = n19386 ^ n19370 ;
  assign n19399 = n12222 ^ x2 ;
  assign n19402 = n19399 ^ n12222 ;
  assign n19403 = n12380 & n19402 ;
  assign n19404 = n19403 ^ n12222 ;
  assign n19405 = ~x1 & n19404 ;
  assign n19388 = n12214 ^ x1 ;
  assign n19389 = n19388 ^ n19377 ;
  assign n19390 = n12607 & n19389 ;
  assign n19391 = n19390 ^ n19388 ;
  assign n19400 = n19399 ^ n19391 ;
  assign n19406 = n19405 ^ n19400 ;
  assign n19407 = ~x0 & ~n19406 ;
  assign n19393 = n19211 ^ n18844 ;
  assign n19394 = n19393 ^ n18843 ;
  assign n19392 = n19220 ^ n19212 ;
  assign n19395 = n19394 ^ n19392 ;
  assign n19396 = n19395 ^ n19391 ;
  assign n19408 = n19407 ^ n19396 ;
  assign n19445 = n19192 ^ n18856 ;
  assign n19425 = n19206 ^ n19195 ;
  assign n20009 = n19445 ^ n19425 ;
  assign n19427 = n12382 ^ x2 ;
  assign n19428 = n19427 ^ n12382 ;
  assign n19429 = n12382 ^ n12228 ;
  assign n19430 = n19429 ^ n12382 ;
  assign n19431 = n19428 & ~n19430 ;
  assign n19432 = n19431 ^ n12382 ;
  assign n19433 = ~x1 & ~n19432 ;
  assign n19434 = n19433 ^ n19427 ;
  assign n19446 = n19445 ^ n19434 ;
  assign n19435 = n12376 ^ x1 ;
  assign n19436 = n19435 ^ n19434 ;
  assign n19437 = n19436 ^ x2 ;
  assign n19438 = n19437 ^ x1 ;
  assign n19439 = n19438 ^ n19436 ;
  assign n19440 = n19436 ^ n12553 ;
  assign n19441 = n19440 ^ n19436 ;
  assign n19442 = n19439 & ~n19441 ;
  assign n19443 = n19442 ^ n19436 ;
  assign n19444 = x0 & ~n19443 ;
  assign n19447 = n19446 ^ n19444 ;
  assign n19972 = n12382 ^ x1 ;
  assign n19973 = n19972 ^ x2 ;
  assign n19974 = n19973 ^ n12382 ;
  assign n19975 = n12370 & n19974 ;
  assign n19976 = n19975 ^ n19972 ;
  assign n19968 = n12228 ^ x2 ;
  assign n19977 = n19976 ^ n19968 ;
  assign n19978 = n19977 ^ n19976 ;
  assign n19979 = n19978 ^ n12228 ;
  assign n19980 = n12229 & n19979 ;
  assign n19981 = n19980 ^ n12228 ;
  assign n19982 = ~x1 & ~n19981 ;
  assign n19983 = n19982 ^ n19977 ;
  assign n19984 = ~x0 & n19983 ;
  assign n19985 = n19984 ^ n19976 ;
  assign n20006 = n19985 ^ n19445 ;
  assign n19946 = n19183 ^ n18891 ;
  assign n19947 = n19946 ^ n18878 ;
  assign n19911 = n19175 ^ n19171 ;
  assign n19898 = n12248 ^ x1 ;
  assign n19882 = n12248 ^ x2 ;
  assign n19899 = n19898 ^ n19882 ;
  assign n19900 = n13518 & n19899 ;
  assign n19901 = n19900 ^ n19898 ;
  assign n19853 = n12249 ^ x2 ;
  assign n19902 = n19901 ^ n19853 ;
  assign n19903 = n19902 ^ n19901 ;
  assign n19904 = n19903 ^ n12249 ;
  assign n19905 = n12339 & n19904 ;
  assign n19906 = n19905 ^ n12249 ;
  assign n19907 = ~x1 & ~n19906 ;
  assign n19908 = n19907 ^ n19902 ;
  assign n19909 = ~x0 & ~n19908 ;
  assign n19910 = n19909 ^ n19901 ;
  assign n19912 = n19911 ^ n19910 ;
  assign n19885 = n19882 ^ n12248 ;
  assign n19886 = ~n12249 & n19885 ;
  assign n19887 = n19886 ^ n12248 ;
  assign n19888 = ~x1 & n19887 ;
  assign n19876 = n12239 ^ x1 ;
  assign n19875 = n12239 ^ x2 ;
  assign n19877 = n19876 ^ n19875 ;
  assign n19878 = n13339 & n19877 ;
  assign n19879 = n19878 ^ n19876 ;
  assign n19883 = n19882 ^ n19879 ;
  assign n19889 = n19888 ^ n19883 ;
  assign n19890 = ~x0 & ~n19889 ;
  assign n19891 = n19890 ^ n19879 ;
  assign n19913 = n19910 ^ n19891 ;
  assign n19814 = n12251 ^ x1 ;
  assign n19813 = n12251 ^ x2 ;
  assign n19815 = n19814 ^ n19813 ;
  assign n19816 = n13676 & n19815 ;
  assign n19817 = n19816 ^ n19814 ;
  assign n19449 = n12253 ^ x2 ;
  assign n19837 = n19817 ^ n19449 ;
  assign n19838 = n19837 ^ n19817 ;
  assign n19839 = n19838 ^ n12253 ;
  assign n19840 = n12331 & n19839 ;
  assign n19841 = n19840 ^ n12253 ;
  assign n19842 = ~x1 & n19841 ;
  assign n19843 = n19842 ^ n19837 ;
  assign n19844 = ~x0 & ~n19843 ;
  assign n19823 = n12253 ^ n12251 ;
  assign n19824 = n19823 ^ n12251 ;
  assign n19818 = n12339 ^ x1 ;
  assign n19819 = n19818 ^ x2 ;
  assign n19820 = n19819 ^ n12339 ;
  assign n19821 = n13884 & n19820 ;
  assign n19822 = n19821 ^ n19818 ;
  assign n19825 = n19822 ^ n19813 ;
  assign n19826 = n19825 ^ n19822 ;
  assign n19827 = n19826 ^ n12251 ;
  assign n19828 = n19824 & n19827 ;
  assign n19829 = n19828 ^ n12251 ;
  assign n19830 = ~x1 & ~n19829 ;
  assign n19831 = n19830 ^ n19825 ;
  assign n19832 = ~x0 & ~n19831 ;
  assign n19833 = n19832 ^ n19822 ;
  assign n19834 = n19833 ^ n19817 ;
  assign n19845 = n19844 ^ n19834 ;
  assign n19846 = n19845 ^ n19833 ;
  assign n19792 = ~x2 & n14219 ;
  assign n19465 = n12257 ^ x2 ;
  assign n19795 = n19792 ^ n19465 ;
  assign n19796 = n19795 ^ n12331 ;
  assign n19797 = x0 & ~n19796 ;
  assign n19798 = n19797 ^ n19465 ;
  assign n19793 = n19792 ^ n14219 ;
  assign n19794 = n19793 ^ n12331 ;
  assign n19799 = n19798 ^ n19794 ;
  assign n19786 = n14972 ^ n12258 ;
  assign n19787 = n19786 ^ n12331 ;
  assign n19455 = n12331 ^ x2 ;
  assign n19788 = n19455 ^ n12331 ;
  assign n19789 = n19787 & n19788 ;
  assign n19790 = n19789 ^ n12331 ;
  assign n19791 = ~x0 & n19790 ;
  assign n19800 = n19799 ^ n19791 ;
  assign n19801 = ~x1 & n19800 ;
  assign n19802 = n19801 ^ n19798 ;
  assign n19490 = n12264 ^ x2 ;
  assign n19493 = n19490 ^ n12264 ;
  assign n19494 = ~n12267 & n19493 ;
  assign n19495 = n19494 ^ n12264 ;
  assign n19496 = ~x1 & n19495 ;
  assign n19482 = n12258 ^ x1 ;
  assign n19472 = n12258 ^ x2 ;
  assign n19483 = n19482 ^ n19472 ;
  assign n19484 = n14242 & n19483 ;
  assign n19485 = n19484 ^ n19482 ;
  assign n19491 = n19490 ^ n19485 ;
  assign n19497 = n19496 ^ n19491 ;
  assign n19498 = ~x0 & ~n19497 ;
  assign n19486 = n19146 ^ n18989 ;
  assign n19487 = n19486 ^ n19485 ;
  assign n19499 = n19498 ^ n19487 ;
  assign n19516 = n19143 ^ n18999 ;
  assign n19506 = n12267 ^ x2 ;
  assign n19509 = n19506 ^ n12267 ;
  assign n19510 = n12268 & n19509 ;
  assign n19511 = n19510 ^ n12267 ;
  assign n19512 = ~x1 & ~n19511 ;
  assign n19500 = n12264 ^ x1 ;
  assign n19501 = n19500 ^ n19490 ;
  assign n19502 = n14428 & n19501 ;
  assign n19503 = n19502 ^ n19500 ;
  assign n19507 = n19506 ^ n19503 ;
  assign n19513 = n19512 ^ n19507 ;
  assign n19514 = ~x0 & ~n19513 ;
  assign n19515 = n19514 ^ n19503 ;
  assign n19517 = n19516 ^ n19515 ;
  assign n19546 = n12276 ^ x2 ;
  assign n19549 = n19546 ^ n12276 ;
  assign n19550 = n12279 & n19549 ;
  assign n19551 = n19550 ^ n12276 ;
  assign n19552 = ~x1 & ~n19551 ;
  assign n19539 = n12268 ^ x1 ;
  assign n19525 = n12268 ^ x2 ;
  assign n19540 = n19539 ^ n19525 ;
  assign n19541 = n14328 & n19540 ;
  assign n19542 = n19541 ^ n19539 ;
  assign n19547 = n19546 ^ n19542 ;
  assign n19553 = n19552 ^ n19547 ;
  assign n19554 = ~x0 & ~n19553 ;
  assign n19536 = n19106 ^ n19105 ;
  assign n19537 = n19536 ^ n19115 ;
  assign n19543 = n19542 ^ n19537 ;
  assign n19555 = n19554 ^ n19543 ;
  assign n19745 = n12276 ^ x1 ;
  assign n19746 = n19745 ^ n19546 ;
  assign n19747 = n14465 & n19746 ;
  assign n19748 = n19747 ^ n19745 ;
  assign n19732 = n12279 ^ x2 ;
  assign n19751 = n19748 ^ n19732 ;
  assign n19752 = n19751 ^ n19748 ;
  assign n19753 = n19752 ^ n12279 ;
  assign n19754 = ~n12283 & n19753 ;
  assign n19755 = n19754 ^ n12279 ;
  assign n19756 = ~x1 & n19755 ;
  assign n19757 = n19756 ^ n19751 ;
  assign n19758 = ~x0 & ~n19757 ;
  assign n19759 = n19758 ^ n19748 ;
  assign n19764 = n19759 ^ n19537 ;
  assign n19721 = n19099 ^ n19020 ;
  assign n19584 = n19096 ^ n19050 ;
  assign n19722 = n19721 ^ n19584 ;
  assign n19587 = n12284 ^ x2 ;
  assign n19590 = n19587 ^ n12284 ;
  assign n19591 = ~n12285 & n19590 ;
  assign n19592 = n19591 ^ n12284 ;
  assign n19593 = ~x1 & ~n19592 ;
  assign n19557 = n14651 ^ n12313 ;
  assign n19558 = ~x2 & n19557 ;
  assign n19559 = n19558 ^ x2 ;
  assign n19560 = n19559 ^ x1 ;
  assign n19556 = ~x1 & n12285 ;
  assign n19561 = n19560 ^ n19556 ;
  assign n19562 = n12284 & n19561 ;
  assign n19563 = n19562 ^ n19559 ;
  assign n19567 = n19563 ^ n19556 ;
  assign n19564 = n19563 ^ n19558 ;
  assign n19568 = n19567 ^ n19564 ;
  assign n19569 = ~n12284 & n19568 ;
  assign n19570 = n19569 ^ n19564 ;
  assign n19571 = ~n12313 & ~n19570 ;
  assign n19572 = n19571 ^ n19563 ;
  assign n19573 = n12285 ^ n12284 ;
  assign n19575 = n12285 ^ n11012 ;
  assign n19576 = n19575 ^ n19557 ;
  assign n19577 = n19576 ^ n11012 ;
  assign n19578 = ~x1 & n19577 ;
  assign n19579 = n19578 ^ n11012 ;
  assign n19580 = n19573 & n19579 ;
  assign n19581 = n19580 ^ x2 ;
  assign n19582 = n19572 & n19581 ;
  assign n19583 = n19582 ^ n12283 ;
  assign n19588 = n19587 ^ n19583 ;
  assign n19594 = n19593 ^ n19588 ;
  assign n19595 = ~x0 & n19594 ;
  assign n19585 = n19584 ^ n19583 ;
  assign n19596 = n19595 ^ n19585 ;
  assign n19689 = n19068 ^ x6 ;
  assign n19690 = n19689 ^ n19051 ;
  assign n19691 = n19690 ^ n19075 ;
  assign n19059 = n19058 ^ x5 ;
  assign n19617 = n19067 ^ n19059 ;
  assign n19692 = n19691 ^ n19617 ;
  assign n19621 = n12289 ^ x2 ;
  assign n19624 = n19621 ^ n12289 ;
  assign n19625 = ~n12290 & n19624 ;
  assign n19626 = n19625 ^ n12289 ;
  assign n19627 = ~x1 & n19626 ;
  assign n19612 = n12313 ^ x1 ;
  assign n19613 = n19612 ^ x2 ;
  assign n19614 = n19613 ^ n12313 ;
  assign n19615 = n14711 & n19614 ;
  assign n19616 = n19615 ^ n19612 ;
  assign n19622 = n19621 ^ n19616 ;
  assign n19628 = n19627 ^ n19622 ;
  assign n19629 = ~x0 & n19628 ;
  assign n19618 = n19617 ^ n19616 ;
  assign n19630 = n19629 ^ n19618 ;
  assign n19663 = n11395 & n12291 ;
  assign n19664 = n19663 ^ n19054 ;
  assign n19636 = n12293 ^ x2 ;
  assign n19639 = n19636 ^ n12293 ;
  assign n19640 = n14854 & n19639 ;
  assign n19641 = n19640 ^ n12293 ;
  assign n19642 = ~x1 & n19641 ;
  assign n19632 = n12290 ^ x2 ;
  assign n19631 = n12290 ^ x1 ;
  assign n19633 = n19632 ^ n19631 ;
  assign n19634 = ~n12297 & n19633 ;
  assign n19635 = n19634 ^ n19631 ;
  assign n19637 = n19636 ^ n19635 ;
  assign n19643 = n19642 ^ n19637 ;
  assign n19644 = ~x0 & ~n19643 ;
  assign n19645 = n19644 ^ n19635 ;
  assign n19646 = n11663 & n12293 ;
  assign n19647 = n19646 ^ x2 ;
  assign n19648 = n19647 ^ n10322 ;
  assign n19649 = n19648 ^ n12292 ;
  assign n19650 = n19649 ^ n19648 ;
  assign n19653 = n19648 ^ n11138 ;
  assign n19654 = n19653 ^ n19648 ;
  assign n19655 = n19647 & ~n19654 ;
  assign n19656 = n19650 & n19655 ;
  assign n19657 = n19656 ^ n19650 ;
  assign n19658 = n19657 ^ n19649 ;
  assign n19659 = ~n12291 & n19658 ;
  assign n19660 = n19659 ^ n10322 ;
  assign n19661 = ~n19645 & n19660 ;
  assign n19662 = n19661 ^ n19617 ;
  assign n19665 = n19664 ^ n19662 ;
  assign n19666 = n19665 ^ n19617 ;
  assign n19671 = x2 & n12293 ;
  assign n19672 = n19671 ^ n12290 ;
  assign n19673 = ~x1 & ~n19672 ;
  assign n19674 = n19673 ^ n19632 ;
  assign n19684 = n19674 ^ n19664 ;
  assign n19667 = n12289 ^ x1 ;
  assign n19675 = n19674 ^ n19667 ;
  assign n19676 = n19675 ^ x2 ;
  assign n19677 = n19676 ^ x1 ;
  assign n19678 = n19677 ^ n19675 ;
  assign n19679 = n19675 ^ n14748 ;
  assign n19680 = n19679 ^ n19675 ;
  assign n19681 = n19678 & n19680 ;
  assign n19682 = n19681 ^ n19675 ;
  assign n19683 = x0 & ~n19682 ;
  assign n19685 = n19684 ^ n19683 ;
  assign n19686 = n19666 & n19685 ;
  assign n19687 = n19686 ^ n19662 ;
  assign n19688 = n19630 & n19687 ;
  assign n19693 = n19692 ^ n19688 ;
  assign n19699 = n12313 ^ n12289 ;
  assign n19700 = n19699 ^ n12313 ;
  assign n19701 = n12313 ^ x2 ;
  assign n19704 = n19701 ^ n12313 ;
  assign n19705 = n19700 & n19704 ;
  assign n19706 = n19705 ^ n12313 ;
  assign n19707 = ~x1 & n19706 ;
  assign n19694 = n12285 ^ x1 ;
  assign n19603 = n12285 ^ x2 ;
  assign n19695 = n19694 ^ n19603 ;
  assign n19696 = n14651 & n19695 ;
  assign n19697 = n19696 ^ n19694 ;
  assign n19702 = n19701 ^ n19697 ;
  assign n19708 = n19707 ^ n19702 ;
  assign n19709 = ~x0 & ~n19708 ;
  assign n19698 = n19697 ^ n19691 ;
  assign n19710 = n19709 ^ n19698 ;
  assign n19711 = n19693 & ~n19710 ;
  assign n19712 = n19711 ^ n19691 ;
  assign n19718 = n19712 ^ n19584 ;
  assign n19599 = n12284 ^ x1 ;
  assign n19600 = n19599 ^ n19587 ;
  assign n19601 = n14583 & n19600 ;
  assign n19602 = n19601 ^ n19599 ;
  assign n19713 = n19712 ^ n19602 ;
  assign n19597 = n12313 ^ n12285 ;
  assign n19598 = n19597 ^ n12285 ;
  assign n19606 = n19603 ^ n12285 ;
  assign n19607 = n19598 & n19606 ;
  assign n19608 = n19607 ^ n12285 ;
  assign n19609 = ~x1 & ~n19608 ;
  assign n19604 = n19603 ^ n19602 ;
  assign n19610 = n19609 ^ n19604 ;
  assign n19611 = ~x0 & n19610 ;
  assign n19714 = n19713 ^ n19611 ;
  assign n19715 = n19712 ^ n19094 ;
  assign n19716 = n19715 ^ n19079 ;
  assign n19717 = ~n19714 & n19716 ;
  assign n19719 = n19718 ^ n19717 ;
  assign n19720 = n19596 & ~n19719 ;
  assign n19723 = n19722 ^ n19720 ;
  assign n19728 = x2 & ~n12284 ;
  assign n19729 = n19728 ^ n12283 ;
  assign n19730 = ~x1 & ~n19729 ;
  assign n19726 = n12283 ^ x2 ;
  assign n19731 = n19730 ^ n19726 ;
  assign n19741 = n19731 ^ n19721 ;
  assign n19733 = n19732 ^ n19731 ;
  assign n19734 = n19733 ^ n11012 ;
  assign n19735 = n19734 ^ n19733 ;
  assign n19736 = n19733 ^ n14514 ;
  assign n19737 = n19736 ^ n19733 ;
  assign n19738 = n19735 & ~n19737 ;
  assign n19739 = n19738 ^ n19733 ;
  assign n19740 = x0 & ~n19739 ;
  assign n19742 = n19741 ^ n19740 ;
  assign n19743 = n19723 & n19742 ;
  assign n19744 = n19743 ^ n19721 ;
  assign n19760 = n19759 ^ n19744 ;
  assign n19761 = n19744 ^ n19009 ;
  assign n19762 = n19761 ^ n19102 ;
  assign n19763 = n19760 & n19762 ;
  assign n19765 = n19764 ^ n19763 ;
  assign n19766 = n19555 & ~n19765 ;
  assign n19523 = n12276 ^ n12268 ;
  assign n19524 = n19523 ^ n12268 ;
  assign n19528 = n19525 ^ n12268 ;
  assign n19529 = ~n19524 & n19528 ;
  assign n19530 = n19529 ^ n12268 ;
  assign n19531 = ~x1 & n19530 ;
  assign n19519 = n12267 ^ x1 ;
  assign n19520 = n19519 ^ n19506 ;
  assign n19521 = n14450 & n19520 ;
  assign n19522 = n19521 ^ n19519 ;
  assign n19526 = n19525 ^ n19522 ;
  assign n19532 = n19531 ^ n19526 ;
  assign n19533 = ~x0 & ~n19532 ;
  assign n19534 = n19533 ^ n19522 ;
  assign n19538 = n19537 ^ n19534 ;
  assign n19767 = n19766 ^ n19538 ;
  assign n19771 = n19115 ^ n19106 ;
  assign n19772 = ~n19536 & n19771 ;
  assign n19768 = n19118 ^ n19114 ;
  assign n19769 = n19768 ^ n19129 ;
  assign n19770 = n19769 ^ n19534 ;
  assign n19773 = n19772 ^ n19770 ;
  assign n19774 = ~n19767 & ~n19773 ;
  assign n19535 = n19534 ^ n19486 ;
  assign n19775 = n19774 ^ n19535 ;
  assign n19518 = n19515 ^ n19486 ;
  assign n19776 = n19775 ^ n19518 ;
  assign n19777 = ~n19517 & ~n19776 ;
  assign n19778 = n19777 ^ n19775 ;
  assign n19779 = n19499 & n19778 ;
  assign n19780 = n19779 ^ n19486 ;
  assign n19475 = n19472 ^ n12258 ;
  assign n19476 = n12264 & n19475 ;
  assign n19477 = n19476 ^ n12258 ;
  assign n19478 = ~x1 & ~n19477 ;
  assign n19466 = n12257 ^ x1 ;
  assign n19467 = n19466 ^ n19465 ;
  assign n19468 = n14019 & n19467 ;
  assign n19469 = n19468 ^ n19466 ;
  assign n19473 = n19472 ^ n19469 ;
  assign n19479 = n19478 ^ n19473 ;
  assign n19480 = ~x0 & ~n19479 ;
  assign n19481 = n19480 ^ n19469 ;
  assign n19781 = n19780 ^ n19481 ;
  assign n19782 = n19481 ^ n18979 ;
  assign n19783 = n19782 ^ n19149 ;
  assign n19784 = ~n19781 & n19783 ;
  assign n19785 = n19784 ^ n19780 ;
  assign n19803 = n19802 ^ n19785 ;
  assign n19804 = n19152 ^ n18969 ;
  assign n19805 = n19804 ^ n19785 ;
  assign n19806 = ~n19803 & ~n19805 ;
  assign n19807 = n19806 ^ n19802 ;
  assign n19453 = n12331 ^ n12257 ;
  assign n19454 = n19453 ^ n12331 ;
  assign n19448 = n12253 ^ x1 ;
  assign n19450 = n19449 ^ n19448 ;
  assign n19451 = n14088 & n19450 ;
  assign n19452 = n19451 ^ n19448 ;
  assign n19456 = n19455 ^ n19452 ;
  assign n19457 = n19456 ^ n19452 ;
  assign n19458 = n19457 ^ n12331 ;
  assign n19459 = n19454 & n19458 ;
  assign n19460 = n19459 ^ n12331 ;
  assign n19461 = ~x1 & n19460 ;
  assign n19462 = n19461 ^ n19456 ;
  assign n19463 = ~x0 & n19462 ;
  assign n19464 = n19463 ^ n19452 ;
  assign n19808 = n19807 ^ n19464 ;
  assign n19809 = n19464 ^ n18959 ;
  assign n19810 = n19809 ^ n19155 ;
  assign n19811 = n19808 & ~n19810 ;
  assign n19812 = n19811 ^ n19807 ;
  assign n19847 = n19846 ^ n19812 ;
  assign n19848 = n19158 ^ n18949 ;
  assign n19849 = n19848 ^ n19812 ;
  assign n19850 = ~n19847 & n19849 ;
  assign n19851 = n19850 ^ n19845 ;
  assign n19857 = n12339 ^ n12251 ;
  assign n19858 = n19857 ^ n12339 ;
  assign n19859 = n12339 ^ x2 ;
  assign n19852 = n12249 ^ x1 ;
  assign n19854 = n19853 ^ n19852 ;
  assign n19855 = n13553 & n19854 ;
  assign n19856 = n19855 ^ n19852 ;
  assign n19860 = n19859 ^ n19856 ;
  assign n19861 = n19860 ^ n19856 ;
  assign n19862 = n19861 ^ n12339 ;
  assign n19863 = ~n19858 & n19862 ;
  assign n19864 = n19863 ^ n12339 ;
  assign n19865 = ~x1 & n19864 ;
  assign n19866 = n19865 ^ n19860 ;
  assign n19867 = ~x0 & ~n19866 ;
  assign n19868 = n19867 ^ n19856 ;
  assign n19869 = n19868 ^ n19833 ;
  assign n19870 = n19869 ^ n19161 ;
  assign n19871 = n19870 ^ n19868 ;
  assign n19872 = n19871 ^ n19166 ;
  assign n19873 = ~n19851 & ~n19872 ;
  assign n19874 = n19873 ^ n19869 ;
  assign n19892 = n19891 ^ n19868 ;
  assign n19893 = n19892 ^ n19891 ;
  assign n19894 = n19893 ^ n19168 ;
  assign n19895 = n19894 ^ n18931 ;
  assign n19896 = ~n19874 & ~n19895 ;
  assign n19897 = n19896 ^ n19892 ;
  assign n19914 = n19913 ^ n19897 ;
  assign n19915 = n19912 & ~n19914 ;
  assign n19916 = n19915 ^ n19897 ;
  assign n19918 = n12235 ^ x2 ;
  assign n19917 = n12235 ^ x1 ;
  assign n19919 = n19918 ^ n19917 ;
  assign n19920 = n13319 & n19919 ;
  assign n19921 = n19920 ^ n19917 ;
  assign n19924 = n19921 ^ n19875 ;
  assign n19925 = n19924 ^ n19921 ;
  assign n19926 = n19925 ^ n12239 ;
  assign n19927 = n12248 & n19926 ;
  assign n19928 = n19927 ^ n12239 ;
  assign n19929 = ~x1 & ~n19928 ;
  assign n19930 = n19929 ^ n19924 ;
  assign n19931 = ~x0 & ~n19930 ;
  assign n19932 = n19931 ^ n19921 ;
  assign n19933 = n19932 ^ n19891 ;
  assign n19934 = n19933 ^ n18911 ;
  assign n19935 = n19934 ^ n19932 ;
  assign n19936 = n19935 ^ n19177 ;
  assign n19937 = n19916 & n19936 ;
  assign n19938 = n19937 ^ n19933 ;
  assign n19939 = n19932 ^ n18878 ;
  assign n19940 = n19939 ^ n19180 ;
  assign n19941 = n19940 ^ n18878 ;
  assign n19942 = n19941 ^ n18901 ;
  assign n19943 = ~n19938 & ~n19942 ;
  assign n19944 = n19943 ^ n19939 ;
  assign n19948 = n19947 ^ n19944 ;
  assign n19950 = n12229 ^ x1 ;
  assign n19949 = n12229 ^ x2 ;
  assign n19951 = n19950 ^ n19949 ;
  assign n19952 = n12866 & n19951 ;
  assign n19953 = n19952 ^ n19950 ;
  assign n19956 = n19953 ^ n19918 ;
  assign n19957 = n19956 ^ n19953 ;
  assign n19958 = n19957 ^ n12235 ;
  assign n19959 = ~n12239 & n19958 ;
  assign n19960 = n19959 ^ n12235 ;
  assign n19961 = ~x1 & n19960 ;
  assign n19962 = n19961 ^ n19956 ;
  assign n19963 = ~x0 & n19962 ;
  assign n19954 = n19953 ^ n19946 ;
  assign n19964 = n19963 ^ n19954 ;
  assign n19965 = ~n19948 & n19964 ;
  assign n19945 = n19944 ^ n19186 ;
  assign n19966 = n19965 ^ n19945 ;
  assign n19967 = n12228 ^ x1 ;
  assign n19969 = n19968 ^ n19967 ;
  assign n19970 = n12805 & n19969 ;
  assign n19971 = n19970 ^ n19967 ;
  assign n19989 = n19971 ^ n19949 ;
  assign n19990 = n19989 ^ n19971 ;
  assign n19991 = n19990 ^ n12229 ;
  assign n19992 = n12235 & n19991 ;
  assign n19993 = n19992 ^ n12229 ;
  assign n19994 = ~x1 & n19993 ;
  assign n19995 = n19994 ^ n19989 ;
  assign n19996 = ~x0 & ~n19995 ;
  assign n19986 = n19985 ^ n19971 ;
  assign n19997 = n19996 ^ n19986 ;
  assign n19998 = n19997 ^ n18878 ;
  assign n19999 = n19998 ^ n19186 ;
  assign n20000 = n19999 ^ n19985 ;
  assign n20001 = n19966 & n20000 ;
  assign n20002 = n20001 ^ n19997 ;
  assign n20003 = n19985 ^ n19189 ;
  assign n20004 = n20003 ^ n18866 ;
  assign n20005 = n20002 & ~n20004 ;
  assign n20007 = n20006 ^ n20005 ;
  assign n20008 = ~n19447 & ~n20007 ;
  assign n20010 = n20009 ^ n20008 ;
  assign n20016 = n12549 ^ n12376 ;
  assign n20017 = n12376 ^ x2 ;
  assign n20020 = n20017 ^ n12376 ;
  assign n20021 = ~n20016 & n20020 ;
  assign n20022 = n20021 ^ n12376 ;
  assign n20023 = ~x1 & n20022 ;
  assign n20011 = n12380 ^ x1 ;
  assign n19414 = n12380 ^ x2 ;
  assign n20012 = n20011 ^ n19414 ;
  assign n20013 = ~n12554 & n20012 ;
  assign n20014 = n20013 ^ n20011 ;
  assign n20018 = n20017 ^ n20014 ;
  assign n20024 = n20023 ^ n20018 ;
  assign n20025 = ~x0 & n20024 ;
  assign n20015 = n20014 ^ n19425 ;
  assign n20026 = n20025 ^ n20015 ;
  assign n20027 = ~n20010 & ~n20026 ;
  assign n19426 = n19425 ^ n19395 ;
  assign n20028 = n20027 ^ n19426 ;
  assign n19413 = n12381 ^ n12380 ;
  assign n19417 = n19414 ^ n12380 ;
  assign n19418 = n19413 & n19417 ;
  assign n19419 = n19418 ^ n12380 ;
  assign n19420 = ~x1 & n19419 ;
  assign n19409 = n12222 ^ x1 ;
  assign n19410 = n19409 ^ n19399 ;
  assign n19411 = ~n12390 & n19410 ;
  assign n19412 = n19411 ^ n19409 ;
  assign n19415 = n19414 ^ n19412 ;
  assign n19421 = n19420 ^ n19415 ;
  assign n19422 = ~x0 & n19421 ;
  assign n19423 = n19422 ^ n19412 ;
  assign n19424 = n19423 ^ n19395 ;
  assign n20029 = n20028 ^ n19424 ;
  assign n20030 = n19423 ^ n18844 ;
  assign n20031 = n20030 ^ n19209 ;
  assign n20032 = ~n20029 & ~n20031 ;
  assign n20033 = n20032 ^ n20028 ;
  assign n20034 = n19408 & n20033 ;
  assign n20035 = n20034 ^ n19395 ;
  assign n20036 = n20035 ^ n19386 ;
  assign n20037 = ~n19387 & n20036 ;
  assign n20038 = n20037 ^ n19386 ;
  assign n20039 = n20038 ^ n19367 ;
  assign n20040 = ~n19369 & ~n20039 ;
  assign n20042 = n20041 ^ n20040 ;
  assign n20043 = ~n19352 & ~n20042 ;
  assign n20044 = n20043 ^ n19351 ;
  assign n20045 = n19333 & ~n20044 ;
  assign n20058 = ~n18814 & ~n19242 ;
  assign n20060 = n20058 ^ n18805 ;
  assign n20073 = ~n20045 & ~n20060 ;
  assign n20046 = n20044 ^ n19333 ;
  assign n20047 = n20046 ^ n20045 ;
  assign n20065 = n19242 ^ n18814 ;
  assign n20066 = n20065 ^ n20058 ;
  assign n20067 = n20066 ^ n19245 ;
  assign n20068 = n20066 ^ n18805 ;
  assign n20069 = n20068 ^ n20066 ;
  assign n20070 = n20067 & n20069 ;
  assign n20071 = n20070 ^ n20066 ;
  assign n20072 = n20047 & ~n20071 ;
  assign n20074 = n19243 ^ n18814 ;
  assign n20075 = ~n20072 & n20074 ;
  assign n20076 = n20073 & n20075 ;
  assign n20077 = n20076 ^ n20072 ;
  assign n20094 = n20077 ^ x2 ;
  assign n20048 = n19242 ^ n18815 ;
  assign n20049 = ~n20047 & ~n20048 ;
  assign n20054 = ~n18806 & n19242 ;
  assign n20055 = n20054 ^ n18805 ;
  assign n20056 = n20049 & ~n20055 ;
  assign n20078 = n20077 ^ n20056 ;
  assign n20057 = n20045 & ~n20056 ;
  assign n20059 = n20058 ^ n19245 ;
  assign n20061 = n20060 ^ n20058 ;
  assign n20062 = n20059 & n20061 ;
  assign n20063 = n20062 ^ n20058 ;
  assign n20064 = n20057 & n20063 ;
  assign n20079 = n20078 ^ n20064 ;
  assign n20081 = n11012 & ~n13051 ;
  assign n20082 = n20081 ^ n12209 ;
  assign n20090 = n20082 ^ x2 ;
  assign n20083 = n20082 ^ n12419 ;
  assign n20084 = n20083 ^ n20082 ;
  assign n20087 = x1 & n20084 ;
  assign n20088 = n20087 ^ n20082 ;
  assign n20089 = ~x0 & ~n20088 ;
  assign n20091 = n20090 ^ n20089 ;
  assign n20080 = n11139 & ~n12405 ;
  assign n20092 = n20091 ^ n20080 ;
  assign n20093 = ~n20079 & n20092 ;
  assign n20095 = n20094 ^ n20093 ;
  assign n19311 = n12209 ^ x2 ;
  assign n19312 = n19311 ^ n12209 ;
  assign n19313 = n15285 & n19312 ;
  assign n19314 = n19313 ^ n12209 ;
  assign n19315 = ~x1 & ~n19314 ;
  assign n19305 = n11012 & ~n12982 ;
  assign n19306 = n19305 ^ n12204 ;
  assign n19307 = n19306 ^ n12209 ;
  assign n19316 = n19315 ^ n19307 ;
  assign n19317 = ~x0 & n19316 ;
  assign n19318 = n19317 ^ n19306 ;
  assign n20096 = n20095 ^ n19318 ;
  assign n20098 = n19260 ^ n19248 ;
  assign n20099 = n20098 ^ n19318 ;
  assign n20100 = n20099 ^ n20095 ;
  assign n20097 = n19318 ^ x2 ;
  assign n20101 = n20100 ^ n20097 ;
  assign n20102 = ~n20096 & n20101 ;
  assign n20103 = n20102 ^ n20100 ;
  assign n20104 = n20103 ^ n19303 ;
  assign n20105 = n19304 & n20104 ;
  assign n20106 = n20105 ^ n19303 ;
  assign n20107 = n20106 ^ n19284 ;
  assign n20108 = n19286 & n20107 ;
  assign n20109 = n20108 ^ n19284 ;
  assign n20110 = n20109 ^ n19269 ;
  assign n20111 = ~n19271 & n20110 ;
  assign n20112 = n20111 ^ n19269 ;
  assign n18755 = n18754 ^ n18262 ;
  assign n18756 = ~n18268 & ~n18755 ;
  assign n18757 = n18756 ^ n18262 ;
  assign n18257 = n8139 & ~n12405 ;
  assign n18254 = n8144 & ~n12210 ;
  assign n18252 = n8484 & n12419 ;
  assign n18250 = n18236 ^ n17821 ;
  assign n18251 = n18250 ^ x8 ;
  assign n18253 = n18252 ^ n18251 ;
  assign n18255 = n18254 ^ n18253 ;
  assign n18249 = n8150 & ~n12651 ;
  assign n18256 = n18255 ^ n18249 ;
  assign n18258 = n18257 ^ n18256 ;
  assign n18758 = n18757 ^ n18258 ;
  assign n20114 = n20112 ^ n18758 ;
  assign n20113 = n18758 & ~n20112 ;
  assign n20115 = n20114 ^ n20113 ;
  assign n20125 = n10327 & ~n12435 ;
  assign n20122 = ~n10334 & ~n12204 ;
  assign n20121 = n10322 ^ x5 ;
  assign n20123 = n20122 ^ n20121 ;
  assign n20120 = n10342 & ~n14140 ;
  assign n20124 = n20123 ^ n20120 ;
  assign n20126 = n20125 ^ n20124 ;
  assign n20119 = n18239 ^ n17811 ;
  assign n20127 = n20126 ^ n20119 ;
  assign n20116 = n18757 ^ n18250 ;
  assign n20117 = n18258 & n20116 ;
  assign n20118 = n20117 ^ n18757 ;
  assign n20128 = n20127 ^ n20118 ;
  assign n20129 = n20128 ^ n14032 ;
  assign n20132 = n10327 & ~n12204 ;
  assign n20131 = ~n10334 & ~n12209 ;
  assign n20133 = n20132 ^ n20131 ;
  assign n20134 = n20133 ^ x5 ;
  assign n20130 = n10322 & ~n12435 ;
  assign n20135 = n20134 ^ n20130 ;
  assign n20136 = n20135 ^ n20134 ;
  assign n20137 = n10329 & n12432 ;
  assign n20138 = n20136 & n20137 ;
  assign n20139 = n20138 ^ n20135 ;
  assign n20140 = n20139 ^ n20128 ;
  assign n20141 = ~n20129 & ~n20140 ;
  assign n20142 = n19268 ^ n18761 ;
  assign n20143 = n18769 & ~n20142 ;
  assign n20144 = n20143 ^ n19268 ;
  assign n20145 = n20144 ^ n20139 ;
  assign n20146 = n20141 & ~n20145 ;
  assign n20147 = n20146 ^ n20128 ;
  assign n20148 = ~n20115 & ~n20147 ;
  assign n20149 = n20128 ^ n20113 ;
  assign n20152 = n20140 ^ n20129 ;
  assign n20153 = ~n20145 & n20152 ;
  assign n20154 = n20153 ^ n20129 ;
  assign n20155 = ~n20149 & n20154 ;
  assign n20156 = n20155 ^ n20113 ;
  assign n20157 = ~n20148 & ~n20156 ;
  assign n20158 = n20126 ^ n20118 ;
  assign n20159 = n20127 & ~n20158 ;
  assign n20160 = n20159 ^ n20126 ;
  assign n20161 = n20157 & ~n20160 ;
  assign n20162 = n20161 ^ n18248 ;
  assign n20164 = n18248 ^ n18242 ;
  assign n20163 = n18248 ^ n17796 ;
  assign n20165 = n20164 ^ n20163 ;
  assign n20166 = n18244 ^ n17796 ;
  assign n20169 = n20165 & ~n20166 ;
  assign n20170 = n20169 ^ n20164 ;
  assign n20171 = n20162 & ~n20170 ;
  assign n20172 = n20171 ^ n20161 ;
  assign n20174 = n20160 ^ n20157 ;
  assign n20175 = n20174 ^ n20161 ;
  assign n20176 = ~n20172 & ~n20175 ;
  assign n20177 = n20173 & n20176 ;
  assign n20178 = n20177 ^ n20172 ;
  assign n20179 = n20178 ^ n20172 ;
  assign n20180 = n18247 & n20179 ;
  assign n20181 = n20180 ^ n20178 ;
  assign n20184 = ~n17775 & n17789 ;
  assign n20185 = n20184 ^ n17790 ;
  assign n20186 = n20181 & ~n20185 ;
  assign n20187 = n17791 & n20186 ;
  assign n20188 = n20187 ^ n20184 ;
  assign n20189 = n20188 ^ n17788 ;
  assign n20190 = ~n17773 & n20189 ;
  assign n20191 = n20181 ^ n17789 ;
  assign n20192 = n20190 & n20191 ;
  assign n20195 = n17788 ^ n17786 ;
  assign n20196 = n20181 ^ n17788 ;
  assign n20197 = ~n20195 & ~n20196 ;
  assign n20198 = n20192 & n20197 ;
  assign n20193 = n20192 ^ n20189 ;
  assign n20199 = n20198 ^ n20193 ;
  assign n20224 = n20223 ^ n20199 ;
  assign n20225 = n20223 ^ n16316 ;
  assign n20226 = n20225 ^ n20223 ;
  assign n20227 = n20226 ^ n16708 ;
  assign n20228 = ~n16711 & ~n20227 ;
  assign n20229 = n20228 ^ n20225 ;
  assign n20230 = n20224 & n20229 ;
  assign n20231 = n20230 ^ n20223 ;
  assign n20235 = n20234 ^ n20231 ;
  assign n15631 = n15274 ^ n15191 ;
  assign n15624 = ~x13 & ~n13051 ;
  assign n15628 = n15624 ^ n13052 ;
  assign n15629 = n6539 & n15628 ;
  assign n15625 = n15624 ^ n12209 ;
  assign n15626 = n6537 & n15625 ;
  assign n15622 = ~n6529 & n12419 ;
  assign n15620 = ~n6547 & ~n12405 ;
  assign n15615 = n15614 ^ n15580 ;
  assign n15616 = n15582 & ~n15615 ;
  assign n15617 = n15616 ^ n15614 ;
  assign n15619 = n15618 ^ n15617 ;
  assign n15621 = n15620 ^ n15619 ;
  assign n15623 = n15622 ^ n15621 ;
  assign n15627 = n15626 ^ n15623 ;
  assign n15630 = n15629 ^ n15627 ;
  assign n15632 = n15631 ^ n15630 ;
  assign n20236 = n20235 ^ n15632 ;
  assign n20248 = n20212 ^ n20211 ;
  assign n20249 = ~n20217 & n20248 ;
  assign n20250 = n20249 ^ n20212 ;
  assign n20246 = n7148 & ~n12204 ;
  assign n20244 = n7151 ^ x11 ;
  assign n20241 = ~n12431 & n20240 ;
  assign n20242 = n20241 ^ n7142 ;
  assign n20243 = ~n12435 & n20242 ;
  assign n20245 = n20244 ^ n20243 ;
  assign n20247 = n20246 ^ n20245 ;
  assign n20252 = n20250 ^ n20247 ;
  assign n20251 = n20247 & n20250 ;
  assign n20253 = n20252 ^ n20251 ;
  assign n20264 = n15631 ^ n15617 ;
  assign n20265 = n15630 & n20264 ;
  assign n20266 = n20265 ^ n15631 ;
  assign n20256 = ~n12435 & n20255 ;
  assign n20258 = n15295 ^ n15278 ;
  assign n20259 = n20258 ^ n20257 ;
  assign n20260 = n20259 ^ x10 ;
  assign n20261 = n20260 ^ n20258 ;
  assign n20262 = n20256 & ~n20261 ;
  assign n20263 = n20262 ^ n20259 ;
  assign n20267 = n20266 ^ n20263 ;
  assign n20268 = n20267 ^ n15632 ;
  assign n20269 = n20268 ^ n20267 ;
  assign n20270 = n20267 ^ n20234 ;
  assign n20271 = n20270 ^ n20267 ;
  assign n20272 = n20269 & n20271 ;
  assign n20273 = n20272 ^ n20267 ;
  assign n20274 = n20253 & n20273 ;
  assign n20275 = ~n20236 & n20274 ;
  assign n20276 = n20267 ^ n20251 ;
  assign n20277 = n20267 ^ n20231 ;
  assign n20278 = n20277 ^ n20268 ;
  assign n20279 = n20268 ^ n20235 ;
  assign n20280 = n20279 ^ n20268 ;
  assign n20281 = ~n20278 & n20280 ;
  assign n20282 = n20281 ^ n20268 ;
  assign n20283 = n20276 & ~n20282 ;
  assign n20284 = n20283 ^ n20251 ;
  assign n20285 = ~n20275 & ~n20284 ;
  assign n15300 = n15299 ^ n15177 ;
  assign n20286 = n20285 ^ n15300 ;
  assign n20288 = n20258 ^ n15300 ;
  assign n20287 = n20266 ^ n15300 ;
  assign n20289 = n20288 ^ n20287 ;
  assign n20290 = ~n20263 & ~n20289 ;
  assign n20291 = n20290 ^ n20288 ;
  assign n20292 = ~n20286 & ~n20291 ;
  assign n20293 = n20292 ^ n20285 ;
  assign n20301 = n20300 ^ n20293 ;
  assign n20330 = ~n12214 & n13433 ;
  assign n20328 = n5426 & ~n12400 ;
  assign n20321 = n12210 ^ x20 ;
  assign n20322 = n20321 ^ x19 ;
  assign n20323 = n20322 ^ n12210 ;
  assign n20324 = ~n12736 & n20323 ;
  assign n20325 = n20324 ^ n12210 ;
  assign n20326 = n5215 & ~n20325 ;
  assign n20327 = n20326 ^ x20 ;
  assign n20329 = n20328 ^ n20327 ;
  assign n20331 = n20330 ^ n20329 ;
  assign n20320 = n14389 ^ n14173 ;
  assign n20332 = n20331 ^ n20320 ;
  assign n20317 = n15134 ^ n15119 ;
  assign n20318 = ~n15123 & ~n20317 ;
  assign n20319 = n20318 ^ n15119 ;
  assign n20333 = n20332 ^ n20319 ;
  assign n20314 = n15145 ^ n15135 ;
  assign n20315 = ~n15137 & ~n20314 ;
  assign n20316 = n20315 ^ n15135 ;
  assign n20334 = n20333 ^ n20316 ;
  assign n20306 = ~x16 & ~n13051 ;
  assign n20309 = n20306 ^ n13052 ;
  assign n20310 = n6147 & n20309 ;
  assign n20303 = n6143 & n12419 ;
  assign n20302 = ~n12405 & n20437 ;
  assign n20304 = n20303 ^ n20302 ;
  assign n20305 = n20304 ^ x17 ;
  assign n20307 = n20306 ^ n12209 ;
  assign n20308 = n20305 & n20307 ;
  assign n20311 = n20310 ^ n20308 ;
  assign n20312 = n20304 ^ n6145 ;
  assign n20313 = ~n20311 & ~n20312 ;
  assign n20335 = n20334 ^ n20313 ;
  assign n20338 = ~n6547 & ~n12204 ;
  assign n20337 = ~n6529 & ~n12435 ;
  assign n20339 = n20338 ^ n20337 ;
  assign n20340 = n20339 ^ n6536 ;
  assign n20336 = n7838 & ~n14140 ;
  assign n20341 = n20340 ^ n20336 ;
  assign n20343 = n20335 & ~n20341 ;
  assign n20342 = n20341 ^ n20335 ;
  assign n20344 = n20343 ^ n20342 ;
  assign n20368 = n20331 ^ n20319 ;
  assign n20369 = n20332 & ~n20368 ;
  assign n20370 = n20369 ^ n20331 ;
  assign n20367 = n14392 ^ n14170 ;
  assign n20371 = n20370 ^ n20367 ;
  assign n20365 = n12419 & n20437 ;
  assign n20363 = n6143 & ~n12209 ;
  assign n20356 = n12204 ^ x17 ;
  assign n20357 = n20356 ^ x16 ;
  assign n20358 = n20357 ^ n12204 ;
  assign n20359 = ~n13415 & n20358 ;
  assign n20360 = n20359 ^ n12204 ;
  assign n20361 = n6141 & ~n20360 ;
  assign n20362 = n20361 ^ x17 ;
  assign n20364 = n20363 ^ n20362 ;
  assign n20366 = n20365 ^ n20364 ;
  assign n20372 = n20371 ^ n20366 ;
  assign n20346 = n6532 & ~n12435 ;
  assign n20348 = n20316 ^ n20313 ;
  assign n20349 = ~n20334 & n20348 ;
  assign n20350 = n20349 ^ n20313 ;
  assign n20351 = n20350 ^ n20347 ;
  assign n20352 = n20351 ^ x13 ;
  assign n20353 = n20352 ^ n20350 ;
  assign n20354 = n20346 & ~n20353 ;
  assign n20355 = n20354 ^ n20351 ;
  assign n20373 = n20372 ^ n20355 ;
  assign n20374 = n20373 ^ n20296 ;
  assign n20375 = n20374 ^ n20373 ;
  assign n20376 = n20373 ^ n20299 ;
  assign n20377 = n20376 ^ n20373 ;
  assign n20378 = ~n20375 & n20377 ;
  assign n20379 = n20378 ^ n20373 ;
  assign n20380 = ~n20344 & ~n20379 ;
  assign n20381 = ~n20301 & n20380 ;
  assign n20382 = n20373 ^ n20343 ;
  assign n20383 = n20376 ^ n20296 ;
  assign n20384 = n20383 ^ n20293 ;
  assign n20385 = n20384 ^ n20376 ;
  assign n20386 = n20343 ^ n20296 ;
  assign n20387 = n20386 ^ n20376 ;
  assign n20388 = n20385 & ~n20387 ;
  assign n20389 = n20388 ^ n20376 ;
  assign n20390 = ~n20382 & ~n20389 ;
  assign n20391 = n20390 ^ n20373 ;
  assign n20392 = ~n20381 & n20391 ;
  assign n20393 = n20370 ^ n20366 ;
  assign n20394 = n20371 & n20393 ;
  assign n20395 = n20394 ^ n20370 ;
  assign n20397 = ~n20392 & ~n20395 ;
  assign n20396 = n20395 ^ n20392 ;
  assign n20398 = n20397 ^ n20396 ;
  assign n20400 = n20399 ^ n20398 ;
  assign n20405 = n14395 ^ n14158 ;
  assign n20401 = n20372 ^ n20350 ;
  assign n20402 = n20355 & ~n20401 ;
  assign n20403 = n20402 ^ n20350 ;
  assign n20406 = n20405 ^ n20403 ;
  assign n20409 = n20405 ^ n6546 ;
  assign n20404 = n20403 ^ n20398 ;
  assign n20410 = n20409 ^ n20404 ;
  assign n20411 = n20410 ^ n20404 ;
  assign n20412 = ~n20406 & ~n20411 ;
  assign n20413 = n20412 ^ n20404 ;
  assign n20414 = n20400 & ~n20413 ;
  assign n20415 = n20414 ^ n20399 ;
  assign n20416 = n20399 ^ n6546 ;
  assign n20417 = n20403 ^ n20399 ;
  assign n20418 = n20405 ^ n20399 ;
  assign n20419 = n20417 & ~n20418 ;
  assign n20420 = ~n20416 & n20419 ;
  assign n20421 = n20420 ^ n20416 ;
  assign n20422 = n20421 ^ n6546 ;
  assign n20423 = ~n20397 & ~n20422 ;
  assign n20424 = n20415 & ~n20423 ;
  assign n20429 = n20427 ^ n20424 ;
  assign n20428 = n20424 & ~n20427 ;
  assign n20430 = n20429 ^ n20428 ;
  assign n20444 = n13937 ^ n6158 ;
  assign n20445 = n20444 ^ n13837 ;
  assign n20440 = n20439 ^ n13944 ;
  assign n20441 = n14400 ^ n13944 ;
  assign n20442 = n20440 & ~n20441 ;
  assign n20443 = n20442 ^ n20440 ;
  assign n20446 = n20445 ^ n20443 ;
  assign n20447 = ~n20430 & n20446 ;
  assign n20448 = n20439 & n20447 ;
  assign n20449 = n14401 & n20448 ;
  assign n20450 = n20449 ^ n20447 ;
  assign n20451 = n20445 ^ n20428 ;
  assign n20452 = n20442 ^ n14400 ;
  assign n20453 = n20452 ^ n20428 ;
  assign n20454 = n20451 & ~n20453 ;
  assign n20455 = n20454 ^ n20428 ;
  assign n20456 = ~n20450 & ~n20455 ;
  assign n20457 = n20456 ^ n13761 ;
  assign n20462 = n20461 ^ n20457 ;
  assign n20468 = n5426 & ~n12435 ;
  assign n20466 = n5221 & ~n14140 ;
  assign n20464 = ~n12204 & n13433 ;
  assign n20463 = n5215 ^ x20 ;
  assign n20465 = n20464 ^ n20463 ;
  assign n20467 = n20466 ^ n20465 ;
  assign n20469 = n20468 ^ n20467 ;
  assign n20470 = n20469 ^ n13761 ;
  assign n20471 = n20470 ^ n20461 ;
  assign n20472 = ~n20462 & ~n20471 ;
  assign n20473 = n20472 ^ n20461 ;
  assign n20474 = n13943 & ~n20473 ;
  assign n20475 = n20474 ^ n13942 ;
  assign n20476 = n13941 ^ n13762 ;
  assign n20477 = n20476 ^ n13942 ;
  assign n20478 = ~n20457 & n20461 ;
  assign n20479 = ~n20470 & n20478 ;
  assign n20480 = n20479 ^ n20470 ;
  assign n20481 = n20480 ^ n20469 ;
  assign n20482 = n20477 & n20481 ;
  assign n20483 = ~n20475 & ~n20482 ;
  assign n13757 = n13756 ^ n13753 ;
  assign n13758 = n13755 & ~n13757 ;
  assign n13759 = n13758 ^ n13756 ;
  assign n13760 = n13759 ^ n8619 ;
  assign n20484 = n20483 ^ n13760 ;
  assign n20485 = ~n13430 & n20484 ;
  assign n20488 = ~n8619 & ~n13759 ;
  assign n13166 = n13165 ^ n13164 ;
  assign n13262 = ~n13166 & ~n13261 ;
  assign n13263 = n13262 ^ n13165 ;
  assign n13152 = n4655 ^ x23 ;
  assign n13142 = ~x25 & ~n13051 ;
  assign n13145 = n13142 ^ n13052 ;
  assign n13146 = n99 & n13145 ;
  assign n13139 = n4600 & n12419 ;
  assign n13138 = ~n12405 & n20603 ;
  assign n13140 = n13139 ^ n13138 ;
  assign n13141 = n13140 ^ x26 ;
  assign n13143 = n13142 ^ n12209 ;
  assign n13144 = n13141 & n13143 ;
  assign n13147 = n13146 ^ n13144 ;
  assign n13148 = n13140 ^ n97 ;
  assign n13149 = ~n13147 & ~n13148 ;
  assign n12924 = ~n12792 & n12923 ;
  assign n12926 = n12925 ^ n12924 ;
  assign n12942 = n12941 ^ n12927 ;
  assign n12600 = n12599 ^ n12564 ;
  assign n12955 = ~n12600 & n12954 ;
  assign n12956 = n12942 & n12955 ;
  assign n12957 = n12956 ^ n12927 ;
  assign n12958 = ~n12926 & ~n12957 ;
  assign n12959 = n12927 ^ n12924 ;
  assign n12960 = n12941 ^ n12924 ;
  assign n12964 = n12960 ^ n12954 ;
  assign n12965 = n12964 ^ n12960 ;
  assign n12966 = ~n12961 & ~n12965 ;
  assign n12967 = n12966 ^ n12960 ;
  assign n12968 = ~n12959 & n12967 ;
  assign n12969 = n12968 ^ n12927 ;
  assign n12970 = ~n12958 & n12969 ;
  assign n12539 = n3425 ^ n1458 ;
  assign n12534 = n1298 ^ n791 ;
  assign n12535 = n12534 ^ n462 ;
  assign n12536 = n12535 ^ n1615 ;
  assign n12532 = n4256 ^ n453 ;
  assign n12533 = n12532 ^ n722 ;
  assign n12537 = n12536 ^ n12533 ;
  assign n12530 = n1711 ^ n1303 ;
  assign n12529 = n12528 ^ n1376 ;
  assign n12531 = n12530 ^ n12529 ;
  assign n12538 = n12537 ^ n12531 ;
  assign n12540 = n12539 ^ n12538 ;
  assign n12522 = n1307 ^ n687 ;
  assign n12523 = n12522 ^ n903 ;
  assign n12521 = n803 ^ n735 ;
  assign n12524 = n12523 ^ n12521 ;
  assign n12520 = n1314 ^ n751 ;
  assign n12525 = n12524 ^ n12520 ;
  assign n12526 = n12525 ^ n2047 ;
  assign n12517 = n5496 ^ n1329 ;
  assign n12515 = n2689 ^ n2058 ;
  assign n12516 = n12515 ^ n1283 ;
  assign n12518 = n12517 ^ n12516 ;
  assign n12514 = n12513 ^ n3129 ;
  assign n12519 = n12518 ^ n12514 ;
  assign n12527 = n12526 ^ n12519 ;
  assign n12541 = n12540 ^ n12527 ;
  assign n12542 = ~n2465 & ~n12541 ;
  assign n12543 = n12542 ^ n8619 ;
  assign n12455 = n5280 & n12376 ;
  assign n12453 = n12452 ^ n12376 ;
  assign n12454 = n12453 & n22005 ;
  assign n12456 = n12455 ^ n12454 ;
  assign n12451 = n3807 & n12222 ;
  assign n12457 = n12456 ^ n12451 ;
  assign n12450 = ~n3801 & n12380 ;
  assign n12458 = n12457 ^ n12450 ;
  assign n12750 = n12543 ^ n12458 ;
  assign n12748 = n3837 & ~n12214 ;
  assign n12746 = n3985 & ~n12400 ;
  assign n12739 = n12210 ^ x29 ;
  assign n12740 = n12739 ^ x28 ;
  assign n12741 = n12740 ^ n12210 ;
  assign n12742 = ~n12736 & n12741 ;
  assign n12743 = n12742 ^ n12210 ;
  assign n12744 = n3833 & ~n12743 ;
  assign n12745 = n12744 ^ x29 ;
  assign n12747 = n12746 ^ n12745 ;
  assign n12749 = n12748 ^ n12747 ;
  assign n12751 = n12750 ^ n12749 ;
  assign n12735 = n12600 & ~n12734 ;
  assign n12752 = n12751 ^ n12735 ;
  assign n13137 = n12970 ^ n12752 ;
  assign n13150 = n13149 ^ n13137 ;
  assign n13134 = n13133 ^ n13098 ;
  assign n13135 = ~n13104 & ~n13134 ;
  assign n13136 = n13135 ^ n13133 ;
  assign n13151 = n13150 ^ n13136 ;
  assign n13153 = n13152 ^ n13151 ;
  assign n13084 = n4656 & ~n12431 ;
  assign n13085 = n13084 ^ n40 ;
  assign n13086 = ~n12435 & ~n13085 ;
  assign n13154 = n13153 ^ n13086 ;
  assign n13081 = n4651 & ~n12204 ;
  assign n13155 = n13154 ^ n13081 ;
  assign n20486 = n13263 ^ n13155 ;
  assign n20487 = n20486 ^ n13760 ;
  assign n20489 = n20488 ^ n20487 ;
  assign n20490 = n20485 & n20489 ;
  assign n20491 = n13429 ^ n13267 ;
  assign n20492 = n20491 ^ n13430 ;
  assign n20493 = n20492 ^ n20486 ;
  assign n20496 = n20488 ^ n13760 ;
  assign n20497 = ~n20483 & n20496 ;
  assign n20498 = n20497 ^ n20493 ;
  assign n20499 = ~n20488 & n20498 ;
  assign n20500 = n20499 ^ n20486 ;
  assign n20501 = n20493 & ~n20500 ;
  assign n20502 = n20501 ^ n20486 ;
  assign n20503 = ~n20490 & ~n20502 ;
  assign n20504 = n20503 ^ n20490 ;
  assign n13264 = n13263 ^ n13151 ;
  assign n13265 = ~n13155 & ~n13264 ;
  assign n13266 = n13265 ^ n13263 ;
  assign n20505 = n20504 ^ n13266 ;
  assign n20510 = n13137 ^ n13136 ;
  assign n20511 = ~n13150 & ~n20510 ;
  assign n20512 = n20511 ^ n13137 ;
  assign n20518 = n20512 ^ n13266 ;
  assign n20531 = n20505 & n20518 ;
  assign n12984 = ~n4435 & n12983 ;
  assign n12980 = ~n4434 & ~n12204 ;
  assign n12977 = n12419 & n20603 ;
  assign n12976 = n4600 & ~n12209 ;
  assign n12978 = n12977 ^ n12976 ;
  assign n12979 = n12978 ^ x26 ;
  assign n12981 = n12980 ^ n12979 ;
  assign n12985 = n12984 ^ n12981 ;
  assign n12726 = n3985 & ~n12210 ;
  assign n12724 = n3837 & ~n12400 ;
  assign n12717 = n12405 ^ x29 ;
  assign n12718 = n12717 ^ x28 ;
  assign n12719 = n12718 ^ n12405 ;
  assign n12720 = ~n12714 & n12719 ;
  assign n12721 = n12720 ^ n12405 ;
  assign n12722 = n3833 & ~n12721 ;
  assign n12723 = n12722 ^ x29 ;
  assign n12725 = n12724 ^ n12723 ;
  assign n12727 = n12726 ^ n12725 ;
  assign n12644 = n12511 ^ n8619 ;
  assign n12645 = n12543 & n12644 ;
  assign n12646 = n12645 ^ n8619 ;
  assign n12634 = n906 ^ n819 ;
  assign n12635 = n12634 ^ n2454 ;
  assign n12636 = n12635 ^ n3391 ;
  assign n12640 = n12639 ^ n12636 ;
  assign n12631 = n3013 ^ n108 ;
  assign n12630 = n5333 ^ n517 ;
  assign n12632 = n12631 ^ n12630 ;
  assign n12626 = n772 ^ n398 ;
  assign n12627 = n12626 ^ n215 ;
  assign n12628 = n12627 ^ n240 ;
  assign n12629 = n12628 ^ n12568 ;
  assign n12633 = n12632 ^ n12629 ;
  assign n12641 = n12640 ^ n12633 ;
  assign n12642 = n12641 ^ n3875 ;
  assign n12643 = ~n2257 & ~n12642 ;
  assign n12647 = n12646 ^ n12643 ;
  assign n12620 = ~n61 & n12222 ;
  assign n12618 = n12214 ^ n3518 ;
  assign n12617 = ~n3518 & n12214 ;
  assign n12619 = n12618 ^ n12617 ;
  assign n12621 = n12620 ^ n12619 ;
  assign n12622 = n12621 ^ n12608 ;
  assign n12610 = n12608 ^ n12222 ;
  assign n12609 = n12608 ^ n12380 ;
  assign n12611 = n12610 ^ n12609 ;
  assign n12614 = x30 & n12611 ;
  assign n12615 = n12614 ^ n12610 ;
  assign n12616 = ~n3518 & n12615 ;
  assign n12623 = n12622 ^ n12616 ;
  assign n12624 = x31 & n12623 ;
  assign n12625 = n12624 ^ n12621 ;
  assign n12648 = n12647 ^ n12625 ;
  assign n12512 = n12511 ^ n12458 ;
  assign n12544 = n12543 ^ n12512 ;
  assign n12565 = n12564 ^ n12458 ;
  assign n12566 = n12565 ^ n12543 ;
  assign n12601 = n12600 ^ n12543 ;
  assign n12602 = n12601 ^ n12543 ;
  assign n12603 = n12566 & n12602 ;
  assign n12604 = n12603 ^ n12543 ;
  assign n12605 = ~n12544 & n12604 ;
  assign n12606 = n12605 ^ n12458 ;
  assign n12649 = n12648 ^ n12606 ;
  assign n12974 = n12727 ^ n12649 ;
  assign n12971 = n12970 ^ n12749 ;
  assign n12972 = ~n12752 & ~n12971 ;
  assign n12973 = n12972 ^ n12749 ;
  assign n12975 = n12974 ^ n12973 ;
  assign n20506 = n12985 ^ n12975 ;
  assign n20514 = n20506 ^ n44 ;
  assign n20513 = n4651 & ~n12435 ;
  assign n20515 = n20514 ^ n20513 ;
  assign n20528 = n20506 ^ n20505 ;
  assign n20529 = n20528 ^ n20512 ;
  assign n20530 = ~n20515 & n20529 ;
  assign n20532 = n20531 ^ n20530 ;
  assign n12988 = n12985 ^ n12973 ;
  assign n12989 = n12975 & n12988 ;
  assign n12710 = x31 & n12620 ;
  assign n12706 = ~n61 & ~n12214 ;
  assign n12696 = n1067 ^ n209 ;
  assign n12697 = n12696 ^ n900 ;
  assign n12695 = n2484 ^ n575 ;
  assign n12698 = n12697 ^ n12695 ;
  assign n12693 = n12692 ^ n3877 ;
  assign n12694 = n12693 ^ n4763 ;
  assign n12699 = n12698 ^ n12694 ;
  assign n12690 = n1459 ^ n568 ;
  assign n12691 = n12690 ^ n1322 ;
  assign n12700 = n12699 ^ n12691 ;
  assign n12686 = n3783 ^ n1811 ;
  assign n12687 = n12686 ^ n886 ;
  assign n12684 = n6682 ^ n1048 ;
  assign n12683 = n1143 ^ n1014 ;
  assign n12685 = n12684 ^ n12683 ;
  assign n12688 = n12687 ^ n12685 ;
  assign n12689 = n12688 ^ n6036 ;
  assign n12701 = n12700 ^ n12689 ;
  assign n12702 = n12701 ^ n12477 ;
  assign n12681 = n952 ^ n529 ;
  assign n12682 = n12681 ^ n837 ;
  assign n12703 = n12702 ^ n12682 ;
  assign n12704 = ~n4748 & ~n12703 ;
  assign n12676 = n12643 & n12646 ;
  assign n12679 = ~n12625 & n12676 ;
  assign n12677 = n12676 ^ n12647 ;
  assign n12678 = n12625 & ~n12677 ;
  assign n12680 = n12679 ^ n12678 ;
  assign n12705 = n12704 ^ n12680 ;
  assign n12707 = n12706 ^ n12705 ;
  assign n12671 = n12667 ^ x31 ;
  assign n12672 = n12671 ^ n12667 ;
  assign n12673 = ~n12666 & ~n12672 ;
  assign n12674 = n12673 ^ n12667 ;
  assign n12675 = n3518 & ~n12674 ;
  assign n12708 = n12707 ^ n12675 ;
  assign n12665 = ~n12617 & n12664 ;
  assign n12709 = n12708 ^ n12665 ;
  assign n12711 = n12710 ^ n12709 ;
  assign n12662 = n3837 & ~n12210 ;
  assign n12660 = n3985 & ~n12405 ;
  assign n12653 = n12651 ^ x29 ;
  assign n12654 = n12653 ^ x28 ;
  assign n12655 = n12654 ^ n12651 ;
  assign n12656 = ~n12650 & ~n12655 ;
  assign n12657 = n12656 ^ n12651 ;
  assign n12658 = n3833 & ~n12657 ;
  assign n12659 = n12658 ^ x29 ;
  assign n12661 = n12660 ^ n12659 ;
  assign n12663 = n12662 ^ n12661 ;
  assign n12712 = n12711 ^ n12663 ;
  assign n12713 = n12712 ^ n12606 ;
  assign n12728 = n12727 ^ n12713 ;
  assign n12729 = n12728 ^ n12712 ;
  assign n12730 = ~n12649 & n12729 ;
  assign n12731 = n12730 ^ n12713 ;
  assign n12440 = n4600 & ~n12204 ;
  assign n12439 = ~n12209 & n20603 ;
  assign n12441 = n12440 ^ n12439 ;
  assign n12438 = n96 & ~n12435 ;
  assign n12442 = n12441 ^ n12438 ;
  assign n12443 = n12442 ^ n12441 ;
  assign n12444 = n12432 & n12443 ;
  assign n12448 = n285 & n12444 ;
  assign n12445 = n12442 ^ x26 ;
  assign n12449 = n12448 ^ n12445 ;
  assign n12732 = n12731 ^ n12449 ;
  assign n12986 = n12985 ^ n12732 ;
  assign n12990 = n12989 ^ n12986 ;
  assign n46 = n45 ^ x23 ;
  assign n47 = n46 ^ n41 ;
  assign n20533 = n12990 ^ n47 ;
  assign n20534 = ~n20532 & ~n20533 ;
  assign n20507 = n20506 ^ n20504 ;
  assign n20508 = ~n20505 & ~n20507 ;
  assign n20509 = n20508 ^ n20504 ;
  assign n20522 = n20507 ^ n20505 ;
  assign n20523 = n20522 ^ n20504 ;
  assign n20516 = n20515 ^ n20506 ;
  assign n20517 = n20516 ^ n20512 ;
  assign n20519 = n20518 ^ n20506 ;
  assign n20520 = n20519 ^ n20504 ;
  assign n20521 = n20517 & n20520 ;
  assign n20524 = n20523 ^ n20521 ;
  assign n20525 = ~n20509 & ~n20524 ;
  assign n20535 = n20534 ^ n20525 ;
  assign n13076 = ~n12204 & n20603 ;
  assign n13074 = n4434 ^ x26 ;
  assign n13071 = ~n4435 & ~n12431 ;
  assign n13072 = n13071 ^ n4600 ;
  assign n13073 = ~n12435 & n13072 ;
  assign n13075 = n13074 ^ n13073 ;
  assign n13077 = n13076 ^ n13075 ;
  assign n13063 = n3837 & ~n12405 ;
  assign n13061 = n3985 & n12419 ;
  assign n13054 = n12209 ^ x29 ;
  assign n13055 = n13054 ^ x28 ;
  assign n13056 = n13055 ^ n12209 ;
  assign n13057 = ~n13051 & n13056 ;
  assign n13058 = n13057 ^ n12209 ;
  assign n13059 = n3833 & ~n13058 ;
  assign n13060 = n13059 ^ x29 ;
  assign n13062 = n13061 ^ n13060 ;
  assign n13064 = n13063 ^ n13062 ;
  assign n13065 = n13064 ^ n12678 ;
  assign n13045 = ~n12736 & n22005 ;
  assign n13046 = n13045 ^ n12210 ;
  assign n13043 = ~n3518 & n12210 ;
  assign n13044 = n13043 ^ n3518 ;
  assign n13047 = n13046 ^ n13044 ;
  assign n13042 = ~n61 & ~n12400 ;
  assign n13048 = n13047 ^ n13042 ;
  assign n13035 = n12706 ^ n12400 ;
  assign n13036 = n13035 ^ n12706 ;
  assign n13037 = n12706 ^ n3518 ;
  assign n13038 = n13037 ^ n12706 ;
  assign n13039 = ~n13036 & ~n13038 ;
  assign n13040 = n13039 ^ n12706 ;
  assign n13041 = x31 & n13040 ;
  assign n13049 = n13048 ^ n13041 ;
  assign n13008 = n4512 ^ n662 ;
  assign n13005 = n4011 ^ n478 ;
  assign n13006 = n13005 ^ n1549 ;
  assign n13003 = n1233 ^ n784 ;
  assign n13004 = n13003 ^ n915 ;
  assign n13007 = n13006 ^ n13004 ;
  assign n13009 = n13008 ^ n13007 ;
  assign n13001 = n13000 ^ n3565 ;
  assign n13002 = n13001 ^ n2884 ;
  assign n13010 = n13009 ^ n13002 ;
  assign n13011 = n13010 ^ n12853 ;
  assign n13031 = n13030 ^ n13021 ;
  assign n13032 = n13031 ^ n5332 ;
  assign n13033 = ~n13011 & ~n13032 ;
  assign n13034 = n13033 ^ n47 ;
  assign n13050 = n13049 ^ n13034 ;
  assign n13066 = n13065 ^ n13050 ;
  assign n12999 = n12680 & n12704 ;
  assign n13067 = n13066 ^ n12999 ;
  assign n12996 = n12705 ^ n12663 ;
  assign n12997 = ~n12711 & ~n12996 ;
  assign n12998 = n12997 ^ n12705 ;
  assign n13068 = n13067 ^ n12998 ;
  assign n13078 = n13077 ^ n13068 ;
  assign n12993 = n12712 ^ n12449 ;
  assign n12994 = ~n12731 & ~n12993 ;
  assign n12995 = n12994 ^ n12712 ;
  assign n13079 = n13078 ^ n12995 ;
  assign n12733 = n12732 ^ n47 ;
  assign n12991 = n12733 & ~n12990 ;
  assign n12992 = n12991 ^ n12732 ;
  assign n13080 = n13079 ^ n12992 ;
  assign n20613 = n20535 ^ n13080 ;
  assign n20606 = n13064 ^ n12998 ;
  assign n20607 = n13067 & ~n20606 ;
  assign n20608 = n20607 ^ n13064 ;
  assign n20604 = ~n12435 & n20603 ;
  assign n20598 = n107 ^ n86 ;
  assign n20599 = n20598 ^ n135 ;
  assign n20605 = n20604 ^ n20599 ;
  assign n20609 = n20608 ^ n20605 ;
  assign n20584 = n4843 ^ n528 ;
  assign n20582 = n999 ^ n514 ;
  assign n20581 = n429 ^ n251 ;
  assign n20583 = n20582 ^ n20581 ;
  assign n20585 = n20584 ^ n20583 ;
  assign n20586 = n20585 ^ n6901 ;
  assign n20589 = n2829 ^ n1167 ;
  assign n20587 = n2053 ^ n343 ;
  assign n20588 = n20587 ^ n1188 ;
  assign n20590 = n20589 ^ n20588 ;
  assign n20591 = n20590 ^ n553 ;
  assign n20592 = n3540 & ~n20591 ;
  assign n20593 = ~n20586 & n20592 ;
  assign n20594 = ~n855 & n20593 ;
  assign n20568 = n13049 ^ n12704 ;
  assign n20569 = n20568 ^ n13034 ;
  assign n20570 = n13049 ^ n12679 ;
  assign n20571 = n20570 ^ n13049 ;
  assign n20572 = n20570 ^ n12678 ;
  assign n20573 = n20572 ^ n20570 ;
  assign n20574 = n20570 ^ n13034 ;
  assign n20575 = ~n20573 & n20574 ;
  assign n20576 = ~n20571 & n20575 ;
  assign n20577 = n20576 ^ n20571 ;
  assign n20578 = n20577 ^ n13049 ;
  assign n20579 = n20569 & ~n20578 ;
  assign n20580 = n20579 ^ n13049 ;
  assign n20595 = n20594 ^ n20580 ;
  assign n20564 = n12704 ^ n47 ;
  assign n20565 = n13034 & ~n20564 ;
  assign n20566 = n20565 ^ n12704 ;
  assign n20562 = x31 & n13042 ;
  assign n20560 = n12664 & ~n13043 ;
  assign n20558 = ~n61 & ~n12210 ;
  assign n20555 = x31 & ~n12714 ;
  assign n20556 = n20555 ^ n12405 ;
  assign n20557 = n3518 & n20556 ;
  assign n20559 = n20558 ^ n20557 ;
  assign n20561 = n20560 ^ n20559 ;
  assign n20563 = n20562 ^ n20561 ;
  assign n20567 = n20566 ^ n20563 ;
  assign n20596 = n20595 ^ n20567 ;
  assign n20551 = n3985 & ~n12209 ;
  assign n20549 = n3837 & n12419 ;
  assign n20542 = n12204 ^ x29 ;
  assign n20543 = n20542 ^ x28 ;
  assign n20544 = n20543 ^ n12204 ;
  assign n20545 = ~n13415 & n20544 ;
  assign n20546 = n20545 ^ n12204 ;
  assign n20547 = n3833 & ~n20546 ;
  assign n20548 = n20547 ^ x29 ;
  assign n20550 = n20549 ^ n20548 ;
  assign n20552 = n20551 ^ n20550 ;
  assign n20597 = n20596 ^ n20552 ;
  assign n20610 = n20609 ^ n20597 ;
  assign n20539 = n13077 ^ n12995 ;
  assign n20540 = n13078 & n20539 ;
  assign n20541 = n20540 ^ n13077 ;
  assign n20611 = n20610 ^ n20541 ;
  assign n20536 = n20535 ^ n12992 ;
  assign n20537 = ~n13080 & n20536 ;
  assign n20538 = n20537 ^ n20535 ;
  assign n20612 = n20611 ^ n20538 ;
  assign n24104 = n20612 ^ x2 ;
  assign n24107 = n24104 ^ n20612 ;
  assign n24108 = ~n20613 & n24107 ;
  assign n24109 = n24108 ^ n20612 ;
  assign n24110 = ~x1 & ~n24109 ;
  assign n20614 = n20533 ^ n20532 ;
  assign n20615 = n20515 ^ n20512 ;
  assign n20616 = n20615 ^ n13266 ;
  assign n20617 = n20616 ^ n20504 ;
  assign n20618 = n20491 ^ n20488 ;
  assign n20619 = n20484 & n20618 ;
  assign n20620 = n20619 ^ n20498 ;
  assign n20621 = n13267 ^ n8619 ;
  assign n20622 = n20621 ^ n13429 ;
  assign n20623 = n20622 ^ n13759 ;
  assign n20624 = n20623 ^ n20483 ;
  assign n20625 = n20469 ^ n13762 ;
  assign n20823 = n20460 ^ n13941 ;
  assign n20825 = n20823 ^ n20469 ;
  assign n20826 = n20825 ^ n20456 ;
  assign n20827 = ~n20625 & ~n20826 ;
  assign n20828 = n20827 ^ n13761 ;
  assign n20822 = n20456 ^ n13941 ;
  assign n20824 = ~n20822 & n20823 ;
  assign n20829 = n20828 ^ n20824 ;
  assign n20626 = n20625 ^ n20460 ;
  assign n20627 = n20626 ^ n13941 ;
  assign n20628 = n20627 ^ n20456 ;
  assign n20816 = n20440 ^ n14400 ;
  assign n20817 = n20816 ^ n20427 ;
  assign n20818 = n20429 & ~n20817 ;
  assign n20819 = n20818 ^ n20446 ;
  assign n20629 = n20440 ^ n20427 ;
  assign n20630 = n20629 ^ n14400 ;
  assign n20631 = n20630 ^ n20424 ;
  assign n20656 = n20403 ^ n6546 ;
  assign n20655 = n20395 ^ n6546 ;
  assign n20657 = n20656 ^ n20655 ;
  assign n20658 = n20655 ^ n20392 ;
  assign n20659 = n20658 ^ n20656 ;
  assign n20662 = ~n20657 & n20659 ;
  assign n20663 = n20662 ^ n20656 ;
  assign n20673 = n20659 ^ n20657 ;
  assign n20674 = n20673 ^ n20656 ;
  assign n20667 = n20658 ^ n20395 ;
  assign n20664 = n20656 ^ n20405 ;
  assign n20665 = n20664 ^ n20658 ;
  assign n20668 = n20667 ^ n20665 ;
  assign n20670 = n20655 ^ n20395 ;
  assign n20671 = n20670 ^ n20656 ;
  assign n20672 = ~n20668 & n20671 ;
  assign n20675 = n20674 ^ n20672 ;
  assign n20676 = n20663 & ~n20675 ;
  assign n20632 = n20405 ^ n20395 ;
  assign n20633 = n20632 ^ n20406 ;
  assign n20634 = n20632 ^ n20392 ;
  assign n20635 = n20634 ^ n6546 ;
  assign n20636 = n20635 ^ n20406 ;
  assign n20639 = n20636 ^ n20632 ;
  assign n20640 = ~n20633 & n20639 ;
  assign n20641 = n20640 ^ n20632 ;
  assign n20652 = n20635 ^ n20632 ;
  assign n20644 = n20406 ^ n20405 ;
  assign n20645 = n20644 ^ n20636 ;
  assign n20642 = n20406 ^ n6546 ;
  assign n20643 = n20642 ^ n20636 ;
  assign n20646 = n20645 ^ n20643 ;
  assign n20649 = n20632 ^ n20405 ;
  assign n20650 = ~n20646 & ~n20649 ;
  assign n20653 = n20652 ^ n20650 ;
  assign n20654 = ~n20641 & n20653 ;
  assign n20679 = n20676 ^ n20654 ;
  assign n20680 = n20679 ^ n20399 ;
  assign n20681 = n20409 ^ n20395 ;
  assign n20682 = n20681 ^ n20403 ;
  assign n20683 = n20682 ^ n20392 ;
  assign n20684 = n20342 ^ n20296 ;
  assign n20687 = n20342 ^ n20293 ;
  assign n20688 = ~n20684 & n20687 ;
  assign n20685 = n20684 ^ n20293 ;
  assign n20686 = ~n20299 & n20685 ;
  assign n20689 = n20688 ^ n20686 ;
  assign n20690 = n20689 ^ n20382 ;
  assign n20691 = n20342 ^ n20299 ;
  assign n20692 = n20691 ^ n20296 ;
  assign n20693 = n20692 ^ n20293 ;
  assign n20694 = n20291 ^ n20285 ;
  assign n20697 = n20250 ^ n20234 ;
  assign n20701 = n20235 & ~n20697 ;
  assign n20695 = n20247 ^ n15632 ;
  assign n20696 = n20247 ^ n20231 ;
  assign n20698 = n20697 ^ n20696 ;
  assign n20699 = ~n20695 & ~n20698 ;
  assign n20700 = n20699 ^ n20267 ;
  assign n20702 = n20701 ^ n20700 ;
  assign n20703 = n20695 ^ n20250 ;
  assign n20704 = n20703 ^ n20234 ;
  assign n20705 = n20704 ^ n20231 ;
  assign n20706 = n20229 ^ n20199 ;
  assign n20711 = n20181 ^ n17768 ;
  assign n20712 = ~n17772 & ~n20711 ;
  assign n20707 = n17776 ^ n17772 ;
  assign n20708 = n20707 ^ n20181 ;
  assign n20709 = n17786 & n20708 ;
  assign n20710 = n20709 ^ n16712 ;
  assign n20713 = n20712 ^ n20710 ;
  assign n20714 = n17786 ^ n17771 ;
  assign n20715 = n20714 ^ n17768 ;
  assign n20716 = n20715 ^ n20181 ;
  assign n20720 = n20157 ^ n18244 ;
  assign n20721 = n20157 ^ n18243 ;
  assign n20722 = n20721 ^ n20160 ;
  assign n20723 = ~n20720 & ~n20722 ;
  assign n20724 = n20723 ^ n18248 ;
  assign n20717 = n20160 ^ n17796 ;
  assign n20718 = n20160 ^ n18242 ;
  assign n20719 = n20717 & n20718 ;
  assign n20725 = n20724 ^ n20719 ;
  assign n20726 = n20725 ^ n20716 ;
  assign n20727 = n20166 ^ n18242 ;
  assign n20728 = n20727 ^ n20160 ;
  assign n20729 = n20728 ^ n20157 ;
  assign n20730 = n20729 ^ n20725 ;
  assign n20738 = n20103 ^ n19304 ;
  assign n20733 = n18758 ^ n14032 ;
  assign n20734 = n20145 ^ n20114 ;
  assign n20735 = ~n20733 & ~n20734 ;
  assign n20736 = n20735 ^ n20128 ;
  assign n20731 = n20139 ^ n20112 ;
  assign n20732 = ~n20145 & n20731 ;
  assign n20737 = n20736 ^ n20732 ;
  assign n20745 = n20109 ^ n19271 ;
  assign n20746 = n20092 ^ n20079 ;
  assign n20747 = n20042 ^ n19334 ;
  assign n20749 = n20074 ^ n19333 ;
  assign n20750 = n20749 ^ n20044 ;
  assign n20748 = n20038 ^ n19369 ;
  assign n20757 = n20035 ^ n19387 ;
  assign n20763 = n19351 ^ n18825 ;
  assign n20758 = n19367 ^ n18834 ;
  assign n20761 = n20758 ^ n19236 ;
  assign n20762 = ~n18826 & ~n20761 ;
  assign n20764 = n20763 ^ n20762 ;
  assign n20759 = n19367 ^ n19236 ;
  assign n20760 = n20758 & n20759 ;
  assign n20765 = n20764 ^ n20760 ;
  assign n20766 = ~n20757 & ~n20765 ;
  assign n20767 = n20748 & ~n20766 ;
  assign n20768 = n20750 & ~n20767 ;
  assign n20769 = n20747 & n20768 ;
  assign n20770 = n20769 ^ n20750 ;
  assign n20771 = ~n20746 & ~n20770 ;
  assign n20772 = n20100 & ~n20771 ;
  assign n20773 = n20738 & ~n20772 ;
  assign n20751 = n20748 & ~n20750 ;
  assign n20752 = ~n20747 & n20751 ;
  assign n20753 = n20752 ^ n20750 ;
  assign n20754 = n20746 & n20753 ;
  assign n20755 = ~n20100 & ~n20754 ;
  assign n20756 = ~n20738 & ~n20755 ;
  assign n20774 = n20773 ^ n20756 ;
  assign n20775 = n20774 ^ n20738 ;
  assign n20776 = n20745 & n20775 ;
  assign n20777 = n20737 & n20776 ;
  assign n20739 = n20106 ^ n19286 ;
  assign n20740 = n20139 ^ n18758 ;
  assign n20741 = n20740 ^ n14032 ;
  assign n20742 = n20741 ^ n20144 ;
  assign n20743 = n20742 ^ n20112 ;
  assign n20744 = ~n20739 & ~n20743 ;
  assign n20778 = n20777 ^ n20744 ;
  assign n20779 = ~n20738 & n20778 ;
  assign n20780 = n20743 ^ n20737 ;
  assign n20781 = n20745 ^ n20743 ;
  assign n20782 = n20743 ^ n20739 ;
  assign n20783 = ~n20781 & ~n20782 ;
  assign n20784 = n20783 ^ n20745 ;
  assign n20785 = n20784 ^ n20737 ;
  assign n20786 = n20785 ^ n20775 ;
  assign n20788 = n20785 ^ n20784 ;
  assign n20791 = n20783 & ~n20788 ;
  assign n20792 = n20786 & n20791 ;
  assign n20793 = n20792 ^ n20786 ;
  assign n20794 = n20793 ^ n20775 ;
  assign n20795 = ~n20780 & ~n20794 ;
  assign n20796 = n20795 ^ n20743 ;
  assign n20797 = ~n20779 & n20796 ;
  assign n20798 = n20797 ^ n20737 ;
  assign n20799 = n20797 ^ n20729 ;
  assign n20800 = n20798 & ~n20799 ;
  assign n20801 = n20730 & ~n20800 ;
  assign n20802 = n20726 & ~n20801 ;
  assign n20803 = n20802 ^ n20716 ;
  assign n20804 = ~n20716 & ~n20803 ;
  assign n21149 = n20713 & ~n20804 ;
  assign n21150 = n20706 & ~n21149 ;
  assign n21151 = ~n20705 & ~n21150 ;
  assign n21152 = n20702 & ~n21151 ;
  assign n21153 = ~n20694 & ~n21152 ;
  assign n21154 = n20693 & ~n21153 ;
  assign n21155 = ~n20690 & ~n21154 ;
  assign n21156 = n20683 & ~n21155 ;
  assign n21157 = n20680 & ~n21156 ;
  assign n21158 = ~n20631 & ~n21157 ;
  assign n21159 = n20819 & ~n21158 ;
  assign n21160 = n20628 & ~n21159 ;
  assign n21161 = n20829 & ~n21160 ;
  assign n21162 = ~n20624 & ~n21161 ;
  assign n21163 = ~n20620 & ~n21162 ;
  assign n21164 = n20617 & ~n21163 ;
  assign n21165 = ~n20614 & ~n21164 ;
  assign n21166 = n20613 & ~n21165 ;
  assign n21167 = ~n20612 & ~n21166 ;
  assign n20805 = n20804 ^ n20802 ;
  assign n20806 = ~n20713 & n20805 ;
  assign n20807 = ~n20706 & ~n20806 ;
  assign n20808 = n20705 & ~n20807 ;
  assign n20809 = ~n20702 & ~n20808 ;
  assign n20810 = n20694 & ~n20809 ;
  assign n20811 = ~n20693 & ~n20810 ;
  assign n20812 = n20690 & ~n20811 ;
  assign n20813 = ~n20683 & ~n20812 ;
  assign n20814 = ~n20680 & ~n20813 ;
  assign n20815 = n20631 & ~n20814 ;
  assign n20820 = ~n20815 & ~n20819 ;
  assign n20821 = ~n20628 & ~n20820 ;
  assign n20830 = ~n20821 & ~n20829 ;
  assign n20831 = n20624 & ~n20830 ;
  assign n20832 = n20620 & ~n20831 ;
  assign n20833 = ~n20617 & ~n20832 ;
  assign n20834 = n20614 & ~n20833 ;
  assign n20835 = ~n20613 & ~n20834 ;
  assign n20836 = n20612 & ~n20835 ;
  assign n24096 = n21167 ^ n20836 ;
  assign n20899 = ~n20541 & ~n20597 ;
  assign n20888 = n20597 ^ n20541 ;
  assign n20900 = n20899 ^ n20888 ;
  assign n20901 = ~n20538 & n20900 ;
  assign n20902 = n20899 ^ n20605 ;
  assign n20903 = n20609 & ~n20902 ;
  assign n20904 = n20903 ^ n20608 ;
  assign n20905 = n20901 & n20904 ;
  assign n20837 = n20605 ^ n20597 ;
  assign n20838 = n20837 ^ n20608 ;
  assign n20839 = n20838 ^ n20541 ;
  assign n20881 = n20563 ^ n20552 ;
  assign n20884 = n20567 & n20881 ;
  assign n20880 = n20580 ^ n20566 ;
  assign n20882 = n20881 ^ n20880 ;
  assign n20883 = n20595 & n20882 ;
  assign n20885 = n20884 ^ n20883 ;
  assign n20873 = n12405 ^ n3807 ;
  assign n20874 = n20873 ^ n20558 ;
  assign n20872 = ~n61 & ~n12405 ;
  assign n20875 = n20874 ^ n20872 ;
  assign n20870 = n12651 ^ n12405 ;
  assign n20871 = n20870 & n22005 ;
  assign n20876 = n20875 ^ n20871 ;
  assign n20862 = n20558 ^ n12405 ;
  assign n20863 = n20862 ^ n12419 ;
  assign n20864 = n20863 ^ n20862 ;
  assign n20865 = n20862 ^ n3807 ;
  assign n20866 = n20865 ^ n20862 ;
  assign n20867 = ~n20864 & n20866 ;
  assign n20868 = n20867 ^ n20862 ;
  assign n20869 = ~x31 & ~n20868 ;
  assign n20877 = n20876 ^ n20869 ;
  assign n20855 = n14293 ^ n327 ;
  assign n20854 = n533 ^ n355 ;
  assign n20856 = n20855 ^ n20854 ;
  assign n20852 = n2780 ^ n362 ;
  assign n20853 = n20852 ^ n975 ;
  assign n20857 = n20856 ^ n20853 ;
  assign n20858 = n20857 ^ n499 ;
  assign n20859 = n20858 ^ n376 ;
  assign n20860 = n3594 & ~n20859 ;
  assign n20861 = ~n697 & n20860 ;
  assign n20878 = n20877 ^ n20861 ;
  assign n20879 = n20878 ^ n20552 ;
  assign n20886 = n20885 ^ n20879 ;
  assign n20849 = n3837 & ~n12209 ;
  assign n20847 = n3985 & ~n12204 ;
  assign n20841 = n3833 & ~n12435 ;
  assign n20842 = n12432 & n20841 ;
  assign n20843 = n20841 ^ x29 ;
  assign n20844 = n20843 ^ x28 ;
  assign n20845 = n20842 & ~n20844 ;
  assign n20846 = n20845 ^ n20843 ;
  assign n20848 = n20847 ^ n20846 ;
  assign n20850 = n20849 ^ n20848 ;
  assign n20851 = n20850 ^ n20600 ;
  assign n20887 = n20886 ^ n20851 ;
  assign n20889 = n20888 ^ n20887 ;
  assign n20840 = ~n20609 & ~n20837 ;
  assign n20890 = n20889 ^ n20840 ;
  assign n20891 = n20890 ^ n20887 ;
  assign n20892 = n20891 ^ n20838 ;
  assign n20893 = n20838 ^ n20538 ;
  assign n20894 = n20893 ^ n20838 ;
  assign n20895 = ~n20892 & ~n20894 ;
  assign n20896 = n20895 ^ n20838 ;
  assign n20897 = n20839 & n20896 ;
  assign n20898 = n20897 ^ n20890 ;
  assign n20906 = n20898 ^ n20887 ;
  assign n20907 = n20905 & n20906 ;
  assign n20908 = n20907 ^ n20898 ;
  assign n24097 = n20908 ^ x1 ;
  assign n24098 = n24097 ^ x2 ;
  assign n24099 = n24098 ^ n20908 ;
  assign n24100 = n24096 & n24099 ;
  assign n24101 = n24100 ^ n24097 ;
  assign n24105 = n24104 ^ n24101 ;
  assign n24111 = n24110 ^ n24105 ;
  assign n24112 = ~x0 & ~n24111 ;
  assign n24113 = n24112 ^ n24101 ;
  assign n21226 = n21165 ^ n20834 ;
  assign n24728 = n20613 ^ x1 ;
  assign n24114 = n20613 ^ x2 ;
  assign n24729 = n24728 ^ n24114 ;
  assign n24730 = n21226 & n24729 ;
  assign n24731 = n24730 ^ n24728 ;
  assign n24135 = n20614 ^ x2 ;
  assign n24734 = n24731 ^ n24135 ;
  assign n24735 = n24734 ^ n24731 ;
  assign n24736 = n24735 ^ n20614 ;
  assign n24737 = ~n20617 & n24736 ;
  assign n24738 = n24737 ^ n20614 ;
  assign n24739 = ~x1 & ~n24738 ;
  assign n24740 = n24739 ^ n24734 ;
  assign n24741 = ~x0 & n24740 ;
  assign n24742 = n24741 ^ n24731 ;
  assign n23016 = n8139 & ~n20693 ;
  assign n22734 = n7151 & ~n20705 ;
  assign n22733 = n7148 & n20713 ;
  assign n22735 = n22734 ^ n22733 ;
  assign n22736 = n22735 ^ x11 ;
  assign n21769 = n21150 ^ n20807 ;
  assign n21770 = n21769 ^ n20705 ;
  assign n22732 = n20240 & n21770 ;
  assign n22737 = n22736 ^ n22732 ;
  assign n22731 = n7142 & ~n20706 ;
  assign n22738 = n22737 ^ n22731 ;
  assign n22233 = ~x13 & n20800 ;
  assign n22234 = n22233 ^ n20725 ;
  assign n22241 = n6537 & n22234 ;
  assign n22238 = ~n6529 & n20729 ;
  assign n22237 = ~n6547 & n20737 ;
  assign n22239 = n22238 ^ n22237 ;
  assign n22240 = n22239 ^ x14 ;
  assign n22242 = n22241 ^ n22240 ;
  assign n22235 = n22234 ^ n20800 ;
  assign n22236 = n6539 & n22235 ;
  assign n22243 = n22242 ^ n22236 ;
  assign n21834 = n20437 & ~n20738 ;
  assign n21427 = ~n20739 & ~n20773 ;
  assign n21426 = n20739 & ~n20756 ;
  assign n21428 = n21427 ^ n21426 ;
  assign n21429 = n21428 ^ n20745 ;
  assign n21832 = n6163 & ~n21429 ;
  assign n21829 = n6148 & n20745 ;
  assign n21828 = n6143 & ~n20739 ;
  assign n21830 = n21829 ^ n21828 ;
  assign n21831 = n21830 ^ x17 ;
  assign n21833 = n21832 ^ n21831 ;
  assign n21835 = n21834 ^ n21833 ;
  assign n21284 = ~n20748 & ~n20757 ;
  assign n21521 = n8316 & ~n21284 ;
  assign n21285 = n21284 ^ n20757 ;
  assign n21522 = n21285 ^ n20748 ;
  assign n21523 = n20747 & n21522 ;
  assign n21524 = n21523 ^ n20748 ;
  assign n21525 = n5221 & ~n21524 ;
  assign n21531 = n5220 & ~n20747 ;
  assign n21528 = n5221 & ~n20747 ;
  assign n21529 = n21528 ^ n13433 ;
  assign n21530 = n20757 & n21529 ;
  assign n21532 = n21531 ^ n21530 ;
  assign n21533 = n21525 & ~n21532 ;
  assign n21534 = n21533 ^ n21532 ;
  assign n21535 = n21521 & ~n21534 ;
  assign n21536 = n21535 ^ n21534 ;
  assign n21275 = n20767 ^ n20747 ;
  assign n21541 = n5220 & ~n21275 ;
  assign n21276 = n21275 ^ n20750 ;
  assign n21540 = n5215 & ~n21276 ;
  assign n21542 = n21541 ^ n21540 ;
  assign n21538 = n5426 & ~n20747 ;
  assign n21537 = n13433 & n20748 ;
  assign n21539 = n21538 ^ n21537 ;
  assign n21543 = n21542 ^ n21539 ;
  assign n21544 = n35 & n20757 ;
  assign n21545 = n21543 ^ x20 ;
  assign n21546 = ~n21544 & n21545 ;
  assign n21547 = ~n21543 & n21546 ;
  assign n21548 = ~n21536 & n21547 ;
  assign n21549 = n21548 ^ n21546 ;
  assign n21550 = n21549 ^ n21545 ;
  assign n21518 = n13433 & ~n20747 ;
  assign n21516 = n5426 & n20750 ;
  assign n21307 = n20770 ^ n20753 ;
  assign n21509 = n20746 ^ x20 ;
  assign n21510 = n21509 ^ x19 ;
  assign n21511 = n21510 ^ n20746 ;
  assign n21512 = n21307 & n21511 ;
  assign n21513 = n21512 ^ n20746 ;
  assign n21514 = n5215 & n21513 ;
  assign n21515 = n21514 ^ x20 ;
  assign n21517 = n21516 ^ n21515 ;
  assign n21519 = n21518 ^ n21517 ;
  assign n21551 = n21550 ^ n21519 ;
  assign n21346 = n35 & n20748 ;
  assign n21553 = n21550 ^ n21346 ;
  assign n21552 = ~n8289 & n20757 ;
  assign n21554 = n21553 ^ n21552 ;
  assign n21555 = n21551 & ~n21554 ;
  assign n21347 = x23 & ~n21346 ;
  assign n21348 = ~n42 & n20757 ;
  assign n21349 = n21347 & n21348 ;
  assign n21350 = n21349 ^ n21347 ;
  assign n21493 = n21350 ^ x23 ;
  assign n21286 = n21285 ^ n20747 ;
  assign n21355 = n4656 & n21286 ;
  assign n21354 = n4651 & n20757 ;
  assign n21356 = n21355 ^ n21354 ;
  assign n21352 = n4655 & ~n20747 ;
  assign n21351 = ~n40 & n20748 ;
  assign n21353 = n21352 ^ n21351 ;
  assign n21357 = n21356 ^ n21353 ;
  assign n21494 = n21493 ^ n21357 ;
  assign n21520 = n21519 ^ n21494 ;
  assign n21556 = n21555 ^ n21520 ;
  assign n21505 = n13433 & n20750 ;
  assign n21503 = n5426 & n20746 ;
  assign n21380 = n20771 ^ n20754 ;
  assign n21496 = n20100 ^ x20 ;
  assign n21497 = n21496 ^ x19 ;
  assign n21498 = n21497 ^ n20100 ;
  assign n21499 = ~n21380 & n21498 ;
  assign n21500 = n21499 ^ n20100 ;
  assign n21501 = n5215 & n21500 ;
  assign n21502 = n21501 ^ x20 ;
  assign n21504 = n21503 ^ n21502 ;
  assign n21506 = n21505 ^ n21504 ;
  assign n21827 = n21556 ^ n21506 ;
  assign n21836 = n21835 ^ n21827 ;
  assign n21844 = n20100 & n20437 ;
  assign n21316 = n20774 ^ n20739 ;
  assign n21842 = n6163 & n21316 ;
  assign n21839 = n6148 & ~n20739 ;
  assign n21838 = n6143 & ~n20738 ;
  assign n21840 = n21839 ^ n21838 ;
  assign n21841 = n21840 ^ x17 ;
  assign n21843 = n21842 ^ n21841 ;
  assign n21845 = n21844 ^ n21843 ;
  assign n21837 = n21554 ^ n21519 ;
  assign n21846 = n21845 ^ n21837 ;
  assign n21917 = n20437 & n20746 ;
  assign n21328 = n20772 ^ n20755 ;
  assign n21329 = n21328 ^ n20738 ;
  assign n21915 = n6163 & n21329 ;
  assign n21912 = n6148 & ~n20738 ;
  assign n21911 = n6143 & n20100 ;
  assign n21913 = n21912 ^ n21911 ;
  assign n21914 = n21913 ^ x17 ;
  assign n21916 = n21915 ^ n21914 ;
  assign n21918 = n21917 ^ n21916 ;
  assign n21858 = n5215 & n20757 ;
  assign n21859 = n6141 & n20748 ;
  assign n21860 = x17 & ~n21859 ;
  assign n21861 = n20757 & n21860 ;
  assign n21862 = n6154 & n21861 ;
  assign n21863 = n21862 ^ n21860 ;
  assign n21870 = n6163 & n21286 ;
  assign n21869 = n20437 & n20757 ;
  assign n21871 = n21870 ^ n21869 ;
  assign n21867 = n6148 & ~n20747 ;
  assign n21866 = n6143 & n20748 ;
  assign n21868 = n21867 ^ n21866 ;
  assign n21872 = n21871 ^ n21868 ;
  assign n21873 = n21863 & ~n21872 ;
  assign n21874 = ~n21858 & ~n21873 ;
  assign n21881 = n20437 & n20748 ;
  assign n21879 = n6163 & ~n21276 ;
  assign n21876 = n6148 & n20750 ;
  assign n21875 = n6143 & ~n20747 ;
  assign n21877 = n21876 ^ n21875 ;
  assign n21878 = n21877 ^ x17 ;
  assign n21880 = n21879 ^ n21878 ;
  assign n21882 = n21881 ^ n21880 ;
  assign n21883 = n21874 & n21882 ;
  assign n21884 = n21883 ^ n21882 ;
  assign n21856 = n5215 & n20748 ;
  assign n21855 = n8563 & n20757 ;
  assign n21857 = n21856 ^ n21855 ;
  assign n21885 = n21884 ^ n21857 ;
  assign n21892 = n20437 & ~n20747 ;
  assign n21308 = n21307 ^ n20746 ;
  assign n21890 = n6163 & n21308 ;
  assign n21887 = n6148 & n20746 ;
  assign n21886 = n6143 & n20750 ;
  assign n21888 = n21887 ^ n21886 ;
  assign n21889 = n21888 ^ x17 ;
  assign n21891 = n21890 ^ n21889 ;
  assign n21893 = n21892 ^ n21891 ;
  assign n21894 = n21893 ^ n21884 ;
  assign n21895 = n21885 & n21894 ;
  assign n21896 = n21895 ^ n21884 ;
  assign n21853 = n20437 & n20750 ;
  assign n21381 = n21380 ^ n20100 ;
  assign n21851 = n6163 & ~n21381 ;
  assign n21848 = n6148 & n20100 ;
  assign n21847 = n6143 & n20746 ;
  assign n21849 = n21848 ^ n21847 ;
  assign n21850 = n21849 ^ x17 ;
  assign n21852 = n21851 ^ n21850 ;
  assign n21854 = n21853 ^ n21852 ;
  assign n21897 = n21896 ^ n21854 ;
  assign n21901 = n20757 ^ n20748 ;
  assign n21898 = n8620 ^ n5426 ;
  assign n21899 = n20748 & ~n21898 ;
  assign n21902 = n21899 ^ n8620 ;
  assign n21903 = n21901 & ~n21902 ;
  assign n21900 = n21899 ^ n21534 ;
  assign n21904 = n21903 ^ n21900 ;
  assign n21907 = n21904 ^ n21854 ;
  assign n21905 = n20748 & n21903 ;
  assign n21906 = ~n21904 & n21905 ;
  assign n21908 = n21907 ^ n21906 ;
  assign n21909 = n21897 & ~n21908 ;
  assign n21910 = n21909 ^ n21896 ;
  assign n21919 = n21918 ^ n21910 ;
  assign n21921 = n21544 ^ n21543 ;
  assign n21922 = n21921 ^ n21918 ;
  assign n21920 = x20 & n21536 ;
  assign n21923 = n21922 ^ n21920 ;
  assign n21924 = n21919 & n21923 ;
  assign n21925 = n21924 ^ n21918 ;
  assign n21926 = n21925 ^ n21845 ;
  assign n21927 = n21846 & n21926 ;
  assign n21928 = n21927 ^ n21845 ;
  assign n21929 = n21928 ^ n21835 ;
  assign n21930 = n21836 & n21929 ;
  assign n21931 = n21930 ^ n21835 ;
  assign n21824 = n20437 & ~n20739 ;
  assign n21438 = ~n20745 & ~n21427 ;
  assign n21437 = n20745 & ~n21426 ;
  assign n21439 = n21438 ^ n21437 ;
  assign n21440 = n21439 ^ n20743 ;
  assign n21822 = n6163 & n21440 ;
  assign n21819 = n6148 & ~n20743 ;
  assign n21818 = n6143 & n20745 ;
  assign n21820 = n21819 ^ n21818 ;
  assign n21821 = n21820 ^ x17 ;
  assign n21823 = n21822 ^ n21821 ;
  assign n21825 = n21824 ^ n21823 ;
  assign n21507 = n21506 ^ n21494 ;
  assign n21557 = n21507 & ~n21556 ;
  assign n21558 = n21557 ^ n21506 ;
  assign n21490 = n13433 & n20746 ;
  assign n21488 = n5426 & n20100 ;
  assign n21481 = n20738 ^ x20 ;
  assign n21482 = n21481 ^ x19 ;
  assign n21483 = n21482 ^ n20738 ;
  assign n21484 = ~n21328 & n21483 ;
  assign n21485 = n21484 ^ n20738 ;
  assign n21486 = n5215 & ~n21485 ;
  assign n21487 = n21486 ^ x20 ;
  assign n21489 = n21488 ^ n21487 ;
  assign n21491 = n21490 ^ n21489 ;
  assign n21358 = n21350 & ~n21357 ;
  assign n21345 = n96 & n20757 ;
  assign n21478 = n21358 ^ n21345 ;
  assign n21343 = ~n40 & ~n20747 ;
  assign n21341 = n4656 & ~n21276 ;
  assign n21338 = n4655 & n20750 ;
  assign n21337 = n4651 & n20748 ;
  assign n21339 = n21338 ^ n21337 ;
  assign n21340 = n21339 ^ x23 ;
  assign n21342 = n21341 ^ n21340 ;
  assign n21344 = n21343 ^ n21342 ;
  assign n21479 = n21478 ^ n21344 ;
  assign n21492 = n21491 ^ n21479 ;
  assign n21817 = n21558 ^ n21492 ;
  assign n21826 = n21825 ^ n21817 ;
  assign n22232 = n21931 ^ n21826 ;
  assign n22244 = n22243 ^ n22232 ;
  assign n22447 = n21928 ^ n21836 ;
  assign n22248 = ~n6529 & n20745 ;
  assign n22247 = ~n6547 & ~n20739 ;
  assign n22249 = n22248 ^ n22247 ;
  assign n22250 = n22249 ^ n6537 ;
  assign n22251 = n22250 ^ x14 ;
  assign n22261 = x13 & ~n21440 ;
  assign n22260 = n8856 & ~n20743 ;
  assign n22262 = n22261 ^ n22260 ;
  assign n22263 = ~n6539 & n22262 ;
  assign n22258 = n21439 ^ n8856 ;
  assign n22252 = n22249 ^ x14 ;
  assign n22253 = n20743 ^ x13 ;
  assign n22254 = n22253 ^ n20743 ;
  assign n22255 = ~n21439 & ~n22254 ;
  assign n22256 = n22255 ^ n20743 ;
  assign n22257 = ~n22252 & n22256 ;
  assign n22259 = n22258 ^ n22257 ;
  assign n22264 = n22263 ^ n22259 ;
  assign n22265 = ~n22251 & n22264 ;
  assign n22246 = n21923 ^ n21910 ;
  assign n22266 = n22265 ^ n22246 ;
  assign n22269 = ~n6529 & ~n20739 ;
  assign n22268 = ~n6547 & ~n20738 ;
  assign n22270 = n22269 ^ n22268 ;
  assign n22271 = n22270 ^ n6537 ;
  assign n22272 = n22271 ^ x14 ;
  assign n22281 = n6539 & n21428 ;
  assign n22273 = n22270 ^ n6538 ;
  assign n22276 = n20745 ^ x13 ;
  assign n22277 = n22276 ^ n20745 ;
  assign n22278 = ~n21428 & ~n22277 ;
  assign n22279 = n22278 ^ n20745 ;
  assign n22280 = n22273 & ~n22279 ;
  assign n22282 = n22281 ^ n22280 ;
  assign n22283 = ~n22272 & ~n22282 ;
  assign n22267 = n21908 ^ n21896 ;
  assign n22284 = n22283 ^ n22267 ;
  assign n22287 = ~n6529 & ~n20738 ;
  assign n22286 = ~n6547 & n20100 ;
  assign n22288 = n22287 ^ n22286 ;
  assign n22289 = n22288 ^ n6537 ;
  assign n22290 = n22289 ^ x14 ;
  assign n22291 = n22288 ^ x14 ;
  assign n22292 = n22291 ^ n6539 ;
  assign n22294 = n20739 ^ x13 ;
  assign n22295 = n22294 ^ n22291 ;
  assign n22296 = n22295 ^ n20739 ;
  assign n22297 = ~n20774 & n22296 ;
  assign n22298 = n22297 ^ n20739 ;
  assign n22299 = n22292 & n22298 ;
  assign n22300 = n22299 ^ n6539 ;
  assign n22301 = ~n22290 & ~n22300 ;
  assign n22285 = n21893 ^ n21885 ;
  assign n22302 = n22301 ^ n22285 ;
  assign n22399 = n21873 ^ n21858 ;
  assign n22400 = n22399 ^ n21882 ;
  assign n22376 = ~n6529 & n20746 ;
  assign n22375 = ~n6547 & n20750 ;
  assign n22377 = n22376 ^ n22375 ;
  assign n22378 = n22377 ^ n6537 ;
  assign n22379 = n22378 ^ x14 ;
  assign n22389 = x13 & n21381 ;
  assign n22388 = n8856 & n20100 ;
  assign n22390 = n22389 ^ n22388 ;
  assign n22391 = ~n6539 & n22390 ;
  assign n22386 = n21380 ^ n8856 ;
  assign n22380 = n22377 ^ x14 ;
  assign n22381 = n20100 ^ x13 ;
  assign n22382 = n22381 ^ n20100 ;
  assign n22383 = ~n21380 & ~n22382 ;
  assign n22384 = n22383 ^ n20100 ;
  assign n22385 = ~n22380 & ~n22384 ;
  assign n22387 = n22386 ^ n22385 ;
  assign n22392 = n22391 ^ n22387 ;
  assign n22393 = ~n22379 & n22392 ;
  assign n22305 = ~n6529 & ~n20747 ;
  assign n22304 = ~n6547 & n20748 ;
  assign n22306 = n22305 ^ n22304 ;
  assign n22307 = n22306 ^ n6537 ;
  assign n22308 = n22307 ^ x14 ;
  assign n22317 = n6539 & n21275 ;
  assign n22309 = n22306 ^ n6538 ;
  assign n22312 = n20750 ^ x13 ;
  assign n22313 = n22312 ^ n20750 ;
  assign n22314 = ~n21275 & ~n22313 ;
  assign n22315 = n22314 ^ n20750 ;
  assign n22316 = n22309 & ~n22315 ;
  assign n22318 = n22317 ^ n22316 ;
  assign n22319 = ~n22308 & ~n22318 ;
  assign n22321 = ~n6529 & n20748 ;
  assign n22320 = ~n6547 & n20757 ;
  assign n22322 = n22321 ^ n22320 ;
  assign n22323 = n22322 ^ n6537 ;
  assign n22324 = n22323 ^ x14 ;
  assign n22325 = n22322 ^ x14 ;
  assign n22330 = n22325 ^ n6539 ;
  assign n22326 = n20747 ^ n17173 ;
  assign n22327 = n22326 ^ n21285 ;
  assign n22328 = n22327 ^ n22326 ;
  assign n22329 = n22325 & ~n22328 ;
  assign n22331 = n22330 ^ n22329 ;
  assign n22332 = n22326 ^ n20747 ;
  assign n22333 = ~n22328 & ~n22332 ;
  assign n22334 = n22333 ^ n20747 ;
  assign n22335 = ~n22330 & n22334 ;
  assign n22336 = ~n22331 & n22335 ;
  assign n22337 = n22336 ^ n22333 ;
  assign n22338 = n22337 ^ n6539 ;
  assign n22339 = n22338 ^ n20747 ;
  assign n22340 = ~n22324 & ~n22339 ;
  assign n22341 = n6391 & n20748 ;
  assign n22342 = x14 & ~n22341 ;
  assign n22343 = ~n6532 & n20757 ;
  assign n22344 = n22342 & n22343 ;
  assign n22345 = n22344 ^ n22342 ;
  assign n22346 = ~n22340 & n22345 ;
  assign n22347 = n6141 & n20757 ;
  assign n22348 = ~n22346 & ~n22347 ;
  assign n22349 = ~n22319 & n22348 ;
  assign n22350 = n22349 ^ n22319 ;
  assign n22351 = n22350 ^ n21859 ;
  assign n22303 = n6140 & n20757 ;
  assign n22352 = n22351 ^ n22303 ;
  assign n22354 = ~n6529 & n20750 ;
  assign n22353 = ~n6547 & ~n20747 ;
  assign n22355 = n22354 ^ n22353 ;
  assign n22356 = n22355 ^ n6537 ;
  assign n22357 = n22356 ^ x14 ;
  assign n22367 = x13 & ~n21308 ;
  assign n22366 = n8856 & n20746 ;
  assign n22368 = n22367 ^ n22366 ;
  assign n22369 = ~n6539 & n22368 ;
  assign n22364 = n21307 ^ n8856 ;
  assign n22358 = n22355 ^ x14 ;
  assign n22359 = n20746 ^ x13 ;
  assign n22360 = n22359 ^ n20746 ;
  assign n22361 = n21307 & ~n22360 ;
  assign n22362 = n22361 ^ n20746 ;
  assign n22363 = ~n22358 & ~n22362 ;
  assign n22365 = n22364 ^ n22363 ;
  assign n22370 = n22369 ^ n22365 ;
  assign n22371 = ~n22357 & ~n22370 ;
  assign n22372 = n22371 ^ n22350 ;
  assign n22373 = ~n22352 & n22372 ;
  assign n22374 = n22373 ^ n22350 ;
  assign n22394 = n22393 ^ n22374 ;
  assign n21864 = n21863 ^ x17 ;
  assign n22395 = n21872 ^ n21864 ;
  assign n22396 = n22395 ^ n22393 ;
  assign n22397 = n22394 & ~n22396 ;
  assign n22398 = n22397 ^ n22393 ;
  assign n22401 = n22400 ^ n22398 ;
  assign n22410 = n22400 ^ x14 ;
  assign n22409 = n6537 & ~n21328 ;
  assign n22411 = n22410 ^ n22409 ;
  assign n22408 = ~n6529 & n20100 ;
  assign n22412 = n22411 ^ n22408 ;
  assign n22407 = ~n6547 & n20746 ;
  assign n22413 = n22412 ^ n22407 ;
  assign n22402 = n20738 ^ x13 ;
  assign n22403 = n22402 ^ n20738 ;
  assign n22404 = ~n21328 & n22403 ;
  assign n22405 = n22404 ^ n20738 ;
  assign n22406 = n6391 & ~n22405 ;
  assign n22414 = n22413 ^ n22406 ;
  assign n22415 = ~n22401 & n22414 ;
  assign n22416 = n22415 ^ n22400 ;
  assign n22417 = n22416 ^ n22301 ;
  assign n22418 = ~n22302 & ~n22417 ;
  assign n22419 = n22418 ^ n22301 ;
  assign n22420 = n22419 ^ n22283 ;
  assign n22421 = ~n22284 & n22420 ;
  assign n22422 = n22421 ^ n22283 ;
  assign n22423 = n22422 ^ n22265 ;
  assign n22424 = ~n22266 & n22423 ;
  assign n22425 = n22424 ^ n22265 ;
  assign n22245 = n21925 ^ n21846 ;
  assign n22426 = n22425 ^ n22245 ;
  assign n22433 = ~n6529 & ~n20743 ;
  assign n22432 = ~n6547 & n20745 ;
  assign n22434 = n22433 ^ n22432 ;
  assign n22435 = n22434 ^ x14 ;
  assign n22436 = n22434 ^ n15618 ;
  assign n22437 = x14 & ~n22436 ;
  assign n21573 = n20743 & n21439 ;
  assign n21574 = n21573 ^ n21438 ;
  assign n21575 = n21574 ^ n20737 ;
  assign n22427 = n21575 ^ x13 ;
  assign n22428 = n22427 ^ n21575 ;
  assign n22438 = n21574 & n22428 ;
  assign n22439 = n22438 ^ n21575 ;
  assign n22440 = n22437 & ~n22439 ;
  assign n22441 = n22440 ^ n22436 ;
  assign n22442 = n22435 & n22441 ;
  assign n22429 = n21574 & ~n22428 ;
  assign n22430 = n22429 ^ n21575 ;
  assign n22431 = n6539 & n22430 ;
  assign n22443 = n22442 ^ n22431 ;
  assign n22444 = n22443 ^ n22425 ;
  assign n22445 = ~n22426 & ~n22444 ;
  assign n22446 = n22445 ^ n22425 ;
  assign n22448 = n22447 ^ n22446 ;
  assign n22457 = ~n6529 & n20737 ;
  assign n22456 = ~n6547 & ~n20743 ;
  assign n22458 = n22457 ^ n22456 ;
  assign n22459 = n22458 ^ x14 ;
  assign n22460 = n22459 ^ n6391 ;
  assign n21592 = n20737 ^ n20729 ;
  assign n21593 = n21592 ^ n20797 ;
  assign n21594 = n21593 ^ n20729 ;
  assign n22449 = n20729 ^ x13 ;
  assign n22450 = n22449 ^ n20729 ;
  assign n22461 = ~n21594 & ~n22450 ;
  assign n22462 = n22461 ^ n20729 ;
  assign n22463 = x14 & ~n22462 ;
  assign n22464 = n22463 ^ n22459 ;
  assign n22465 = ~n22460 & n22464 ;
  assign n22466 = ~n22458 & ~n22465 ;
  assign n22467 = n22466 ^ x14 ;
  assign n22453 = ~n20798 & n22450 ;
  assign n22454 = n22453 ^ n20729 ;
  assign n22455 = n6539 & n22454 ;
  assign n22468 = n22467 ^ n22455 ;
  assign n22469 = n22468 ^ n22446 ;
  assign n22470 = ~n22448 & n22469 ;
  assign n22471 = n22470 ^ n22446 ;
  assign n22472 = n22471 ^ n22232 ;
  assign n22473 = n22244 & n22472 ;
  assign n22474 = n22473 ^ n22243 ;
  assign n22213 = ~n6529 & n20725 ;
  assign n22212 = ~n6547 & n20729 ;
  assign n22214 = n22213 ^ n22212 ;
  assign n22215 = n22214 ^ n6537 ;
  assign n22216 = n22215 ^ x14 ;
  assign n22226 = n8856 & n20716 ;
  assign n21754 = n20801 ^ n20716 ;
  assign n22225 = x13 & ~n21754 ;
  assign n22227 = n22226 ^ n22225 ;
  assign n22228 = ~n6539 & n22227 ;
  assign n22223 = n20801 ^ n8856 ;
  assign n22217 = n22214 ^ x14 ;
  assign n22218 = n20716 ^ x13 ;
  assign n22219 = n22218 ^ n20716 ;
  assign n22220 = n20801 & ~n22219 ;
  assign n22221 = n22220 ^ n20716 ;
  assign n22222 = ~n22217 & ~n22221 ;
  assign n22224 = n22223 ^ n22222 ;
  assign n22229 = n22228 ^ n22224 ;
  assign n22230 = ~n22216 & ~n22229 ;
  assign n21559 = n21558 ^ n21491 ;
  assign n21560 = n21492 & n21559 ;
  assign n21561 = n21560 ^ n21491 ;
  assign n21475 = n5426 & ~n20738 ;
  assign n21473 = n5220 & ~n20739 ;
  assign n21470 = n5221 & n21316 ;
  assign n21469 = n13433 & n20100 ;
  assign n21471 = n21470 ^ n21469 ;
  assign n21472 = n21471 ^ x20 ;
  assign n21474 = n21473 ^ n21472 ;
  assign n21476 = n21475 ^ n21474 ;
  assign n21370 = ~n40 & n20750 ;
  assign n21368 = n4656 & n21308 ;
  assign n21365 = n4655 & n20746 ;
  assign n21364 = n4651 & ~n20747 ;
  assign n21366 = n21365 ^ n21364 ;
  assign n21367 = n21366 ^ x23 ;
  assign n21369 = n21368 ^ n21367 ;
  assign n21371 = n21370 ^ n21369 ;
  assign n21359 = ~n21345 & ~n21358 ;
  assign n21360 = n21344 & n21359 ;
  assign n21361 = n21360 ^ n21344 ;
  assign n21279 = n96 & n20748 ;
  assign n21362 = n21361 ^ n21279 ;
  assign n21336 = ~n7925 & n20757 ;
  assign n21363 = n21362 ^ n21336 ;
  assign n21468 = n21371 ^ n21363 ;
  assign n21477 = n21476 ^ n21468 ;
  assign n21943 = n21561 ^ n21477 ;
  assign n21940 = n6163 & n21575 ;
  assign n21938 = n6148 & n20737 ;
  assign n21936 = n6143 & ~n20743 ;
  assign n21932 = n21931 ^ n21825 ;
  assign n21933 = n21826 & n21932 ;
  assign n21934 = n21933 ^ n21825 ;
  assign n21935 = n21934 ^ x17 ;
  assign n21937 = n21936 ^ n21935 ;
  assign n21939 = n21938 ^ n21937 ;
  assign n21941 = n21940 ^ n21939 ;
  assign n21816 = n20437 & n20745 ;
  assign n21942 = n21941 ^ n21816 ;
  assign n22211 = n21943 ^ n21942 ;
  assign n22231 = n22230 ^ n22211 ;
  assign n22730 = n22474 ^ n22231 ;
  assign n22739 = n22738 ^ n22730 ;
  assign n22744 = n7151 & ~n20706 ;
  assign n22743 = n7148 & n20716 ;
  assign n22745 = n22744 ^ n22743 ;
  assign n22746 = n22745 ^ x11 ;
  assign n21781 = n21149 ^ n20806 ;
  assign n21782 = n21781 ^ n20706 ;
  assign n22742 = n20240 & n21782 ;
  assign n22747 = n22746 ^ n22742 ;
  assign n22741 = n7142 & n20713 ;
  assign n22748 = n22747 ^ n22741 ;
  assign n22740 = n22471 ^ n22244 ;
  assign n22749 = n22748 ^ n22740 ;
  assign n22754 = n7151 & n20713 ;
  assign n22753 = n7148 & n20725 ;
  assign n22755 = n22754 ^ n22753 ;
  assign n22756 = n22755 ^ x11 ;
  assign n21793 = n20802 ^ n20713 ;
  assign n22752 = n20240 & n21793 ;
  assign n22757 = n22756 ^ n22752 ;
  assign n22751 = n7142 & n20716 ;
  assign n22758 = n22757 ^ n22751 ;
  assign n22750 = n22468 ^ n22448 ;
  assign n22759 = n22758 ^ n22750 ;
  assign n22764 = n7151 & n20716 ;
  assign n22763 = n7148 & n20729 ;
  assign n22765 = n22764 ^ n22763 ;
  assign n22766 = n22765 ^ x11 ;
  assign n22762 = n20240 & n21754 ;
  assign n22767 = n22766 ^ n22762 ;
  assign n22761 = n7142 & n20725 ;
  assign n22768 = n22767 ^ n22761 ;
  assign n22760 = n22443 ^ n22426 ;
  assign n22769 = n22768 ^ n22760 ;
  assign n22899 = n7142 & n20737 ;
  assign n22897 = n20240 & ~n21593 ;
  assign n22895 = n7151 & n20729 ;
  assign n22893 = n7148 & ~n20743 ;
  assign n22879 = n22416 ^ n22302 ;
  assign n22778 = n7142 & n20745 ;
  assign n22776 = n20240 & n21440 ;
  assign n22773 = n7151 & ~n20743 ;
  assign n22772 = n7148 & ~n20739 ;
  assign n22774 = n22773 ^ n22772 ;
  assign n22775 = n22774 ^ x11 ;
  assign n22777 = n22776 ^ n22775 ;
  assign n22779 = n22778 ^ n22777 ;
  assign n22771 = n22414 ^ n22398 ;
  assign n22780 = n22779 ^ n22771 ;
  assign n22788 = n7142 & ~n20739 ;
  assign n22786 = n20240 & ~n21429 ;
  assign n22783 = n7151 & n20745 ;
  assign n22782 = n7148 & ~n20738 ;
  assign n22784 = n22783 ^ n22782 ;
  assign n22785 = n22784 ^ x11 ;
  assign n22787 = n22786 ^ n22785 ;
  assign n22789 = n22788 ^ n22787 ;
  assign n22781 = n22396 ^ n22374 ;
  assign n22790 = n22789 ^ n22781 ;
  assign n22798 = n7142 & ~n20738 ;
  assign n22796 = n20240 & n21316 ;
  assign n22793 = n7151 & ~n20739 ;
  assign n22792 = n7148 & n20100 ;
  assign n22794 = n22793 ^ n22792 ;
  assign n22795 = n22794 ^ x11 ;
  assign n22797 = n22796 ^ n22795 ;
  assign n22799 = n22798 ^ n22797 ;
  assign n22791 = n22371 ^ n22352 ;
  assign n22800 = n22799 ^ n22791 ;
  assign n22809 = n7142 & n20100 ;
  assign n22807 = n20240 & n21329 ;
  assign n22804 = n7151 & ~n20738 ;
  assign n22803 = n7148 & n20746 ;
  assign n22805 = n22804 ^ n22803 ;
  assign n22806 = n22805 ^ x11 ;
  assign n22808 = n22807 ^ n22806 ;
  assign n22810 = n22809 ^ n22808 ;
  assign n22801 = n22347 ^ n22346 ;
  assign n22802 = n22801 ^ n22319 ;
  assign n22811 = n22810 ^ n22802 ;
  assign n22854 = n22345 ^ n22340 ;
  assign n22846 = n7142 & n20750 ;
  assign n22844 = n20240 & n21308 ;
  assign n22841 = n7151 & n20746 ;
  assign n22840 = n7148 & ~n20747 ;
  assign n22842 = n22841 ^ n22840 ;
  assign n22843 = n22842 ^ x11 ;
  assign n22845 = n22844 ^ n22843 ;
  assign n22847 = n22846 ^ n22845 ;
  assign n22812 = n6391 & n20757 ;
  assign n22813 = ~n20255 & ~n21284 ;
  assign n22816 = n20240 & ~n20747 ;
  assign n22817 = n22816 ^ n7148 ;
  assign n22818 = n20757 & n22817 ;
  assign n22819 = n7140 & ~n22818 ;
  assign n22820 = n21524 ^ n20747 ;
  assign n22821 = n20747 ^ n9499 ;
  assign n22822 = n22821 ^ n20747 ;
  assign n22823 = n22820 & n22822 ;
  assign n22824 = n22823 ^ n20747 ;
  assign n22825 = n22819 & ~n22824 ;
  assign n22826 = n22825 ^ n22818 ;
  assign n22827 = x11 & ~n22826 ;
  assign n22828 = ~n22813 & n22827 ;
  assign n22829 = ~n22812 & ~n22828 ;
  assign n22836 = n7142 & ~n20747 ;
  assign n22834 = n20240 & ~n21276 ;
  assign n22831 = n7151 & n20750 ;
  assign n22830 = n7148 & n20748 ;
  assign n22832 = n22831 ^ n22830 ;
  assign n22833 = n22832 ^ x11 ;
  assign n22835 = n22834 ^ n22833 ;
  assign n22837 = n22836 ^ n22835 ;
  assign n22838 = n22829 & n22837 ;
  assign n22839 = n22838 ^ n22837 ;
  assign n22848 = n22847 ^ n22839 ;
  assign n22850 = n22839 ^ n22341 ;
  assign n22849 = ~n6531 & n20757 ;
  assign n22851 = n22850 ^ n22849 ;
  assign n22852 = n22848 & ~n22851 ;
  assign n22853 = n22852 ^ n22847 ;
  assign n22855 = n22854 ^ n22853 ;
  assign n22862 = n7142 & n20746 ;
  assign n22860 = n20240 & ~n21381 ;
  assign n22857 = n7151 & n20100 ;
  assign n22856 = n7148 & n20750 ;
  assign n22858 = n22857 ^ n22856 ;
  assign n22859 = n22858 ^ x11 ;
  assign n22861 = n22860 ^ n22859 ;
  assign n22863 = n22862 ^ n22861 ;
  assign n22864 = n22863 ^ n22853 ;
  assign n22865 = n22855 & n22864 ;
  assign n22866 = n22865 ^ n22863 ;
  assign n22867 = n22866 ^ n22810 ;
  assign n22868 = ~n22811 & n22867 ;
  assign n22869 = n22868 ^ n22810 ;
  assign n22870 = n22869 ^ n22799 ;
  assign n22871 = n22800 & n22870 ;
  assign n22872 = n22871 ^ n22799 ;
  assign n22873 = n22872 ^ n22789 ;
  assign n22874 = n22790 & n22873 ;
  assign n22875 = n22874 ^ n22789 ;
  assign n22876 = n22875 ^ n22779 ;
  assign n22877 = ~n22780 & n22876 ;
  assign n22878 = n22877 ^ n22779 ;
  assign n22880 = n22879 ^ n22878 ;
  assign n22887 = n20240 & n21575 ;
  assign n22885 = n7151 & n20737 ;
  assign n22883 = n7148 & n20745 ;
  assign n22882 = n22878 ^ x11 ;
  assign n22884 = n22883 ^ n22882 ;
  assign n22886 = n22885 ^ n22884 ;
  assign n22888 = n22887 ^ n22886 ;
  assign n22881 = n7142 & ~n20743 ;
  assign n22889 = n22888 ^ n22881 ;
  assign n22890 = ~n22880 & ~n22889 ;
  assign n22891 = n22890 ^ n22879 ;
  assign n22892 = n22891 ^ x11 ;
  assign n22894 = n22893 ^ n22892 ;
  assign n22896 = n22895 ^ n22894 ;
  assign n22898 = n22897 ^ n22896 ;
  assign n22900 = n22899 ^ n22898 ;
  assign n22901 = n22419 ^ n22284 ;
  assign n22902 = n22901 ^ n22891 ;
  assign n22903 = n22900 & ~n22902 ;
  assign n22904 = n22903 ^ n22901 ;
  assign n22770 = n22422 ^ n22266 ;
  assign n22905 = n22904 ^ n22770 ;
  assign n22915 = n7148 & n20737 ;
  assign n22913 = n7142 & n20729 ;
  assign n21736 = n20800 ^ n20725 ;
  assign n22906 = n21736 ^ x11 ;
  assign n22907 = n22906 ^ x10 ;
  assign n22908 = n22907 ^ n21736 ;
  assign n22909 = n20800 & ~n22908 ;
  assign n22910 = n22909 ^ n21736 ;
  assign n22911 = n7140 & n22910 ;
  assign n22912 = n22911 ^ x11 ;
  assign n22914 = n22913 ^ n22912 ;
  assign n22916 = n22915 ^ n22914 ;
  assign n22917 = n22916 ^ n22904 ;
  assign n22918 = n22905 & n22917 ;
  assign n22919 = n22918 ^ n22904 ;
  assign n22920 = n22919 ^ n22768 ;
  assign n22921 = ~n22769 & n22920 ;
  assign n22922 = n22921 ^ n22768 ;
  assign n22923 = n22922 ^ n22758 ;
  assign n22924 = n22759 & n22923 ;
  assign n22925 = n22924 ^ n22758 ;
  assign n22926 = n22925 ^ n22748 ;
  assign n22927 = ~n22749 & n22926 ;
  assign n22928 = n22927 ^ n22748 ;
  assign n22929 = n22928 ^ n22738 ;
  assign n22930 = ~n22739 & n22929 ;
  assign n22931 = n22930 ^ n22738 ;
  assign n22728 = n7142 & ~n20705 ;
  assign n22475 = n22474 ^ n22230 ;
  assign n22476 = ~n22231 & ~n22475 ;
  assign n22477 = n22476 ^ n22230 ;
  assign n21951 = n6148 & n20729 ;
  assign n21950 = n6143 & n20737 ;
  assign n21952 = n21951 ^ n21950 ;
  assign n21953 = n21952 ^ x17 ;
  assign n21949 = n6163 & ~n21593 ;
  assign n21954 = n21953 ^ n21949 ;
  assign n21948 = n20437 & ~n20743 ;
  assign n21955 = n21954 ^ n21948 ;
  assign n21944 = n21943 ^ n21934 ;
  assign n21945 = n21942 & n21944 ;
  assign n21946 = n21945 ^ n21934 ;
  assign n21562 = n21561 ^ n21476 ;
  assign n21563 = ~n21477 & n21562 ;
  assign n21564 = n21563 ^ n21561 ;
  assign n21465 = n13433 & ~n20738 ;
  assign n21463 = n5426 & ~n20739 ;
  assign n21456 = n20745 ^ x20 ;
  assign n21457 = n21456 ^ x19 ;
  assign n21458 = n21457 ^ n20745 ;
  assign n21459 = ~n21428 & n21458 ;
  assign n21460 = n21459 ^ n20745 ;
  assign n21461 = n5215 & n21460 ;
  assign n21462 = n21461 ^ x20 ;
  assign n21464 = n21463 ^ n21462 ;
  assign n21466 = n21465 ^ n21464 ;
  assign n21280 = x26 & ~n21279 ;
  assign n21281 = n7678 & n20757 ;
  assign n21282 = n21280 & n21281 ;
  assign n21283 = n21282 ^ n21280 ;
  assign n21385 = n21283 ^ x26 ;
  assign n21291 = ~n4434 & ~n20747 ;
  assign n21289 = n4600 & n20748 ;
  assign n21288 = n20603 & n20757 ;
  assign n21290 = n21289 ^ n21288 ;
  assign n21292 = n21291 ^ n21290 ;
  assign n21287 = ~n4435 & n21286 ;
  assign n21293 = n21292 ^ n21287 ;
  assign n21386 = n21385 ^ n21293 ;
  assign n21382 = n4656 & ~n21381 ;
  assign n21378 = n4655 & n20100 ;
  assign n21376 = n4651 & n20750 ;
  assign n21372 = n21371 ^ n21361 ;
  assign n21373 = ~n21363 & n21372 ;
  assign n21374 = n21373 ^ n21371 ;
  assign n21375 = n21374 ^ x23 ;
  assign n21377 = n21376 ^ n21375 ;
  assign n21379 = n21378 ^ n21377 ;
  assign n21383 = n21382 ^ n21379 ;
  assign n21335 = ~n40 & n20746 ;
  assign n21384 = n21383 ^ n21335 ;
  assign n21454 = n21386 ^ n21384 ;
  assign n21467 = n21466 ^ n21454 ;
  assign n21815 = n21564 ^ n21467 ;
  assign n21947 = n21946 ^ n21815 ;
  assign n22209 = n21955 ^ n21947 ;
  assign n22206 = n21793 ^ x13 ;
  assign n22195 = n20802 ^ n7310 ;
  assign n22196 = n22195 ^ n20802 ;
  assign n22199 = n22195 ^ n6540 ;
  assign n22200 = n22199 ^ n22195 ;
  assign n22201 = n20725 & ~n22200 ;
  assign n22202 = n22196 & n22201 ;
  assign n22203 = n22202 ^ n22196 ;
  assign n22204 = n22203 ^ n20802 ;
  assign n22205 = ~n7838 & ~n22204 ;
  assign n22207 = n22206 ^ n22205 ;
  assign n22188 = n20716 ^ n20713 ;
  assign n22189 = n22188 ^ n20713 ;
  assign n22190 = n20713 ^ n6540 ;
  assign n22191 = n22190 ^ n20713 ;
  assign n22192 = n22189 & n22191 ;
  assign n22193 = n22192 ^ n20713 ;
  assign n22194 = ~n6391 & n22193 ;
  assign n22208 = n22207 ^ n22194 ;
  assign n22210 = n22209 ^ n22208 ;
  assign n22723 = n22477 ^ n22210 ;
  assign n22724 = n22723 ^ x11 ;
  assign n22722 = n7151 & ~n20702 ;
  assign n22725 = n22724 ^ n22722 ;
  assign n22721 = n7148 & ~n20706 ;
  assign n22726 = n22725 ^ n22721 ;
  assign n22078 = n21151 ^ n20808 ;
  assign n22079 = n22078 ^ n20702 ;
  assign n22720 = n20240 & n22079 ;
  assign n22727 = n22726 ^ n22720 ;
  assign n22729 = n22728 ^ n22727 ;
  assign n23011 = n22931 ^ n22729 ;
  assign n23012 = n23011 ^ x8 ;
  assign n23010 = n8484 & ~n20690 ;
  assign n23013 = n23012 ^ n23010 ;
  assign n23009 = n8144 & ~n20694 ;
  assign n23014 = n23013 ^ n23009 ;
  assign n21244 = n21154 ^ n20811 ;
  assign n21246 = n21244 ^ n20690 ;
  assign n23008 = n8150 & n21246 ;
  assign n23015 = n23014 ^ n23008 ;
  assign n23017 = n23016 ^ n23015 ;
  assign n23026 = n8139 & ~n20694 ;
  assign n23021 = n22928 ^ n22739 ;
  assign n23022 = n23021 ^ x8 ;
  assign n23020 = n8484 & ~n20693 ;
  assign n23023 = n23022 ^ n23020 ;
  assign n23019 = n8144 & ~n20702 ;
  assign n23024 = n23023 ^ n23019 ;
  assign n22090 = n21153 ^ n20810 ;
  assign n22091 = n22090 ^ n20693 ;
  assign n23018 = n8150 & n22091 ;
  assign n23025 = n23024 ^ n23018 ;
  assign n23027 = n23026 ^ n23025 ;
  assign n23039 = n8144 & ~n20705 ;
  assign n23037 = n8139 & ~n20702 ;
  assign n23034 = n22925 ^ n22749 ;
  assign n23035 = n23034 ^ x8 ;
  assign n22112 = n21152 ^ n20809 ;
  assign n23029 = n20694 ^ n9896 ;
  assign n23030 = n23029 ^ n20694 ;
  assign n23031 = ~n22112 & n23030 ;
  assign n23032 = n23031 ^ n20694 ;
  assign n23033 = n8137 & ~n23032 ;
  assign n23036 = n23035 ^ n23033 ;
  assign n23038 = n23037 ^ n23036 ;
  assign n23040 = n23039 ^ n23038 ;
  assign n23049 = n8139 & ~n20705 ;
  assign n23046 = n8144 & ~n20706 ;
  assign n23044 = n8484 & ~n20702 ;
  assign n23042 = n22922 ^ n22759 ;
  assign n23043 = n23042 ^ x8 ;
  assign n23045 = n23044 ^ n23043 ;
  assign n23047 = n23046 ^ n23045 ;
  assign n23041 = n8150 & n22079 ;
  assign n23048 = n23047 ^ n23041 ;
  assign n23050 = n23049 ^ n23048 ;
  assign n23056 = n8484 & ~n20706 ;
  assign n23055 = n8144 & n20716 ;
  assign n23057 = n23056 ^ n23055 ;
  assign n23058 = n23057 ^ x8 ;
  assign n23054 = n8150 & n21782 ;
  assign n23059 = n23058 ^ n23054 ;
  assign n23053 = n8139 & n20713 ;
  assign n23060 = n23059 ^ n23053 ;
  assign n23052 = n22916 ^ n22905 ;
  assign n23061 = n23060 ^ n23052 ;
  assign n23066 = n8484 & n20713 ;
  assign n23065 = n8144 & n20725 ;
  assign n23067 = n23066 ^ n23065 ;
  assign n23068 = n23067 ^ x8 ;
  assign n23064 = n8150 & n21793 ;
  assign n23069 = n23068 ^ n23064 ;
  assign n23063 = n8139 & n20716 ;
  assign n23070 = n23069 ^ n23063 ;
  assign n23062 = n22901 ^ n22900 ;
  assign n23071 = n23070 ^ n23062 ;
  assign n23076 = n8484 & n20716 ;
  assign n23075 = n8144 & n20729 ;
  assign n23077 = n23076 ^ n23075 ;
  assign n23078 = n23077 ^ x8 ;
  assign n23074 = n8150 & n21754 ;
  assign n23079 = n23078 ^ n23074 ;
  assign n23073 = n8139 & n20725 ;
  assign n23080 = n23079 ^ n23073 ;
  assign n23072 = n22889 ^ n22879 ;
  assign n23081 = n23080 ^ n23072 ;
  assign n23222 = n22875 ^ n22780 ;
  assign n23209 = n22872 ^ n22790 ;
  assign n23091 = n8139 & n20745 ;
  assign n23088 = n8144 & ~n20739 ;
  assign n23086 = n8484 & ~n20743 ;
  assign n23084 = n22866 ^ n22811 ;
  assign n23085 = n23084 ^ x8 ;
  assign n23087 = n23086 ^ n23085 ;
  assign n23089 = n23088 ^ n23087 ;
  assign n23083 = n8150 & n21440 ;
  assign n23090 = n23089 ^ n23083 ;
  assign n23092 = n23091 ^ n23090 ;
  assign n23181 = n22863 ^ n22855 ;
  assign n23100 = n8139 & ~n20738 ;
  assign n23098 = n8150 & n21316 ;
  assign n23095 = n8484 & ~n20739 ;
  assign n23094 = n8144 & n20100 ;
  assign n23096 = n23095 ^ n23094 ;
  assign n23097 = n23096 ^ x8 ;
  assign n23099 = n23098 ^ n23097 ;
  assign n23101 = n23100 ^ n23099 ;
  assign n23093 = n22851 ^ n22847 ;
  assign n23102 = n23101 ^ n23093 ;
  assign n23164 = n22837 ^ n22812 ;
  assign n23165 = n23164 ^ n22828 ;
  assign n23115 = n7140 & n20757 ;
  assign n23116 = n8137 & n20748 ;
  assign n23117 = n8143 & ~n20757 ;
  assign n23118 = ~n23116 & n23117 ;
  assign n23119 = n23118 ^ n8143 ;
  assign n23120 = n23119 ^ x8 ;
  assign n23125 = n8150 & n21286 ;
  assign n23124 = n8144 & n20757 ;
  assign n23126 = n23125 ^ n23124 ;
  assign n23122 = n8484 & ~n20747 ;
  assign n23121 = n8139 & n20748 ;
  assign n23123 = n23122 ^ n23121 ;
  assign n23127 = n23126 ^ n23123 ;
  assign n23128 = n23120 & ~n23127 ;
  assign n23129 = ~n23115 & ~n23128 ;
  assign n23136 = n8139 & ~n20747 ;
  assign n23134 = n8150 & ~n21276 ;
  assign n23131 = n8484 & n20750 ;
  assign n23130 = n8144 & n20748 ;
  assign n23132 = n23131 ^ n23130 ;
  assign n23133 = n23132 ^ x8 ;
  assign n23135 = n23134 ^ n23133 ;
  assign n23137 = n23136 ^ n23135 ;
  assign n23138 = n23129 & n23137 ;
  assign n23139 = n23138 ^ n23137 ;
  assign n23113 = n7140 & n20748 ;
  assign n23112 = n7139 & n20757 ;
  assign n23114 = n23113 ^ n23112 ;
  assign n23140 = n23139 ^ n23114 ;
  assign n23147 = n8139 & n20750 ;
  assign n23145 = n8150 & n21308 ;
  assign n23142 = n8484 & n20746 ;
  assign n23141 = n8144 & ~n20747 ;
  assign n23143 = n23142 ^ n23141 ;
  assign n23144 = n23143 ^ x8 ;
  assign n23146 = n23145 ^ n23144 ;
  assign n23148 = n23147 ^ n23146 ;
  assign n23149 = n23148 ^ n23139 ;
  assign n23150 = n23140 & n23149 ;
  assign n23151 = n23150 ^ n23139 ;
  assign n23107 = ~n21285 & n22827 ;
  assign n23108 = n23107 ^ n20748 ;
  assign n23109 = n7142 & n23108 ;
  assign n23110 = n23109 ^ n22826 ;
  assign n23103 = x11 & n22813 ;
  assign n23111 = n23110 ^ n23103 ;
  assign n23152 = n23151 ^ n23111 ;
  assign n23159 = n8139 & n20746 ;
  assign n23157 = n8150 & ~n21381 ;
  assign n23154 = n8484 & n20100 ;
  assign n23153 = n8144 & n20750 ;
  assign n23155 = n23154 ^ n23153 ;
  assign n23156 = n23155 ^ x8 ;
  assign n23158 = n23157 ^ n23156 ;
  assign n23160 = n23159 ^ n23158 ;
  assign n23161 = n23160 ^ n23111 ;
  assign n23162 = n23152 & ~n23161 ;
  assign n23163 = n23162 ^ n23151 ;
  assign n23166 = n23165 ^ n23163 ;
  assign n23173 = n8150 & n21329 ;
  assign n23170 = n23163 ^ x8 ;
  assign n23169 = n8144 & n20746 ;
  assign n23171 = n23170 ^ n23169 ;
  assign n23168 = n8484 & ~n20738 ;
  assign n23172 = n23171 ^ n23168 ;
  assign n23174 = n23173 ^ n23172 ;
  assign n23167 = n8139 & n20100 ;
  assign n23175 = n23174 ^ n23167 ;
  assign n23176 = n23166 & ~n23175 ;
  assign n23177 = n23176 ^ n23165 ;
  assign n23178 = n23177 ^ n23093 ;
  assign n23179 = n23102 & ~n23178 ;
  assign n23180 = n23179 ^ n23101 ;
  assign n23182 = n23181 ^ n23180 ;
  assign n23190 = n8139 & ~n20739 ;
  assign n23186 = n23181 ^ x8 ;
  assign n23185 = n8484 & n20745 ;
  assign n23187 = n23186 ^ n23185 ;
  assign n23184 = n8144 & ~n20738 ;
  assign n23188 = n23187 ^ n23184 ;
  assign n23183 = n8150 & ~n21429 ;
  assign n23189 = n23188 ^ n23183 ;
  assign n23191 = n23190 ^ n23189 ;
  assign n23192 = ~n23182 & ~n23191 ;
  assign n23193 = n23192 ^ n23181 ;
  assign n23194 = n23193 ^ n23084 ;
  assign n23195 = ~n23092 & n23194 ;
  assign n23196 = n23195 ^ n23084 ;
  assign n23082 = n22869 ^ n22800 ;
  assign n23197 = n23196 ^ n23082 ;
  assign n23204 = n8139 & ~n20743 ;
  assign n23202 = n8150 & n21575 ;
  assign n23199 = n8484 & n20737 ;
  assign n23198 = n8144 & n20745 ;
  assign n23200 = n23199 ^ n23198 ;
  assign n23201 = n23200 ^ x8 ;
  assign n23203 = n23202 ^ n23201 ;
  assign n23205 = n23204 ^ n23203 ;
  assign n23206 = n23205 ^ n23082 ;
  assign n23207 = ~n23197 & ~n23206 ;
  assign n23208 = n23207 ^ n23196 ;
  assign n23210 = n23209 ^ n23208 ;
  assign n23214 = n8484 & n20729 ;
  assign n23213 = n8144 & ~n20743 ;
  assign n23215 = n23214 ^ n23213 ;
  assign n23216 = n23215 ^ x8 ;
  assign n23212 = n8150 & ~n21593 ;
  assign n23217 = n23216 ^ n23212 ;
  assign n23211 = n8139 & n20737 ;
  assign n23218 = n23217 ^ n23211 ;
  assign n23219 = n23218 ^ n23208 ;
  assign n23220 = n23210 & ~n23219 ;
  assign n23221 = n23220 ^ n23218 ;
  assign n23223 = n23222 ^ n23221 ;
  assign n23230 = n8150 & n21736 ;
  assign n23228 = n8484 & n20725 ;
  assign n23226 = n8144 & n20737 ;
  assign n23225 = n23221 ^ x8 ;
  assign n23227 = n23226 ^ n23225 ;
  assign n23229 = n23228 ^ n23227 ;
  assign n23231 = n23230 ^ n23229 ;
  assign n23224 = n8139 & n20729 ;
  assign n23232 = n23231 ^ n23224 ;
  assign n23233 = ~n23223 & ~n23232 ;
  assign n23234 = n23233 ^ n23222 ;
  assign n23235 = n23234 ^ n23080 ;
  assign n23236 = ~n23081 & ~n23235 ;
  assign n23237 = n23236 ^ n23080 ;
  assign n23238 = n23237 ^ n23070 ;
  assign n23239 = ~n23071 & n23238 ;
  assign n23240 = n23239 ^ n23070 ;
  assign n23241 = n23240 ^ n23060 ;
  assign n23242 = n23061 & n23241 ;
  assign n23243 = n23242 ^ n23060 ;
  assign n23051 = n22919 ^ n22769 ;
  assign n23244 = n23243 ^ n23051 ;
  assign n23252 = n8139 & ~n20706 ;
  assign n23248 = n23051 ^ x8 ;
  assign n23247 = n8484 & ~n20705 ;
  assign n23249 = n23248 ^ n23247 ;
  assign n23246 = n8144 & n20713 ;
  assign n23250 = n23249 ^ n23246 ;
  assign n23245 = n8150 & n21770 ;
  assign n23251 = n23250 ^ n23245 ;
  assign n23253 = n23252 ^ n23251 ;
  assign n23254 = ~n23244 & n23253 ;
  assign n23255 = n23254 ^ n23243 ;
  assign n23256 = n23255 ^ n23042 ;
  assign n23257 = n23050 & n23256 ;
  assign n23258 = n23257 ^ n23042 ;
  assign n23259 = n23258 ^ n23034 ;
  assign n23260 = ~n23040 & ~n23259 ;
  assign n23261 = n23260 ^ n23034 ;
  assign n23262 = n23261 ^ n23021 ;
  assign n23263 = ~n23027 & n23262 ;
  assign n23264 = n23263 ^ n23021 ;
  assign n23265 = n23264 ^ n23011 ;
  assign n23266 = n23017 & ~n23265 ;
  assign n23267 = n23266 ^ n23011 ;
  assign n22932 = n22931 ^ n22723 ;
  assign n22933 = n22729 & n22932 ;
  assign n22934 = n22933 ^ n22723 ;
  assign n22718 = n7142 & ~n20702 ;
  assign n22478 = n22477 ^ n22208 ;
  assign n22479 = n22210 & n22478 ;
  assign n22480 = n22479 ^ n22477 ;
  assign n22172 = ~n6529 & n20713 ;
  assign n22171 = ~n6547 & n20716 ;
  assign n22173 = n22172 ^ n22171 ;
  assign n22174 = n22173 ^ n6537 ;
  assign n22175 = n22174 ^ x14 ;
  assign n22176 = n22173 ^ x14 ;
  assign n22177 = n22176 ^ n6539 ;
  assign n22184 = n20706 & n22177 ;
  assign n22178 = n22177 ^ n17173 ;
  assign n22179 = n22178 ^ n17173 ;
  assign n22180 = ~x13 & ~n22179 ;
  assign n22181 = n22180 ^ n17173 ;
  assign n22182 = ~n21781 & ~n22181 ;
  assign n22183 = n22182 ^ n6539 ;
  assign n22185 = n22184 ^ n22183 ;
  assign n22186 = ~n22175 & ~n22185 ;
  assign n21970 = n20437 & n20737 ;
  assign n21968 = n6143 & n20729 ;
  assign n21961 = n21736 ^ x17 ;
  assign n21962 = n21961 ^ x16 ;
  assign n21963 = n21962 ^ n21736 ;
  assign n21964 = n20800 & ~n21963 ;
  assign n21965 = n21964 ^ n21736 ;
  assign n21966 = n6141 & n21965 ;
  assign n21967 = n21966 ^ x17 ;
  assign n21969 = n21968 ^ n21967 ;
  assign n21971 = n21970 ^ n21969 ;
  assign n21565 = n21564 ^ n21466 ;
  assign n21566 = n21467 & n21565 ;
  assign n21567 = n21566 ^ n21466 ;
  assign n21451 = n13433 & ~n20739 ;
  assign n21449 = n5426 & n20745 ;
  assign n21442 = n20743 ^ x20 ;
  assign n21443 = n21442 ^ x19 ;
  assign n21444 = n21443 ^ n20743 ;
  assign n21445 = ~n21439 & n21444 ;
  assign n21446 = n21445 ^ n20743 ;
  assign n21447 = n5215 & ~n21446 ;
  assign n21448 = n21447 ^ x20 ;
  assign n21450 = n21449 ^ n21448 ;
  assign n21452 = n21451 ^ n21450 ;
  assign n21387 = n21386 ^ n21374 ;
  assign n21388 = ~n21384 & n21387 ;
  assign n21389 = n21388 ^ n21386 ;
  assign n21332 = ~n40 & n20100 ;
  assign n21330 = n4656 & n21329 ;
  assign n21325 = n4655 & ~n20738 ;
  assign n21324 = n4651 & n20746 ;
  assign n21326 = n21325 ^ n21324 ;
  assign n21327 = n21326 ^ x23 ;
  assign n21331 = n21330 ^ n21327 ;
  assign n21333 = n21332 ^ n21331 ;
  assign n21295 = n3833 & n20757 ;
  assign n21294 = n21283 & ~n21293 ;
  assign n21322 = n21295 ^ n21294 ;
  assign n21277 = ~n4435 & ~n21276 ;
  assign n21273 = ~n4434 & n20750 ;
  assign n21270 = n4600 & ~n20747 ;
  assign n21269 = n20603 & n20748 ;
  assign n21271 = n21270 ^ n21269 ;
  assign n21272 = n21271 ^ x26 ;
  assign n21274 = n21273 ^ n21272 ;
  assign n21278 = n21277 ^ n21274 ;
  assign n21323 = n21322 ^ n21278 ;
  assign n21334 = n21333 ^ n21323 ;
  assign n21436 = n21389 ^ n21334 ;
  assign n21453 = n21452 ^ n21436 ;
  assign n21959 = n21567 ^ n21453 ;
  assign n21956 = n21955 ^ n21946 ;
  assign n21957 = ~n21947 & n21956 ;
  assign n21958 = n21957 ^ n21955 ;
  assign n21960 = n21959 ^ n21958 ;
  assign n22170 = n21971 ^ n21960 ;
  assign n22187 = n22186 ^ n22170 ;
  assign n22713 = n22480 ^ n22187 ;
  assign n22714 = n22713 ^ x11 ;
  assign n22712 = n7151 & ~n20694 ;
  assign n22715 = n22714 ^ n22712 ;
  assign n22711 = n7148 & ~n20705 ;
  assign n22716 = n22715 ^ n22711 ;
  assign n22601 = n22112 ^ n20694 ;
  assign n22710 = n20240 & n22601 ;
  assign n22717 = n22716 ^ n22710 ;
  assign n22719 = n22718 ^ n22717 ;
  assign n23007 = n22934 ^ n22719 ;
  assign n23269 = n23267 ^ n23007 ;
  assign n23268 = n23007 & n23267 ;
  assign n23270 = n23269 ^ n23268 ;
  assign n22617 = n21155 ^ n20812 ;
  assign n22618 = n22617 ^ n20683 ;
  assign n23275 = n8150 & n22618 ;
  assign n23274 = n8139 & ~n20690 ;
  assign n23276 = n23275 ^ n23274 ;
  assign n23272 = n8484 & ~n20683 ;
  assign n23271 = n8144 & ~n20693 ;
  assign n23273 = n23272 ^ n23271 ;
  assign n23277 = n23276 ^ n23273 ;
  assign n23278 = n23277 ^ x8 ;
  assign n22661 = n21156 ^ n20813 ;
  assign n22662 = n22661 ^ n20680 ;
  assign n23285 = n8150 & ~n22662 ;
  assign n23284 = n8139 & ~n20683 ;
  assign n23286 = n23285 ^ n23284 ;
  assign n23282 = n8484 & n20680 ;
  assign n23281 = n8144 & ~n20690 ;
  assign n23283 = n23282 ^ n23281 ;
  assign n23287 = n23286 ^ n23283 ;
  assign n22935 = n22934 ^ n22713 ;
  assign n22936 = ~n22719 & n22935 ;
  assign n22937 = n22936 ^ n22934 ;
  assign n22706 = n7150 & ~n20693 ;
  assign n22704 = n7148 & ~n20702 ;
  assign n22481 = n22480 ^ n22186 ;
  assign n22482 = n22187 & n22481 ;
  assign n22483 = n22482 ^ n22480 ;
  assign n22153 = ~n6547 & n20713 ;
  assign n22152 = ~n6529 & ~n20706 ;
  assign n22154 = n22153 ^ n22152 ;
  assign n22155 = n22154 ^ n6537 ;
  assign n22156 = n22155 ^ x14 ;
  assign n22158 = n22154 ^ x14 ;
  assign n22159 = n22158 ^ n6539 ;
  assign n22166 = n20705 & n22159 ;
  assign n22160 = n22159 ^ n17173 ;
  assign n22161 = n22160 ^ n17173 ;
  assign n22162 = ~x13 & ~n22161 ;
  assign n22163 = n22162 ^ n17173 ;
  assign n22164 = ~n21769 & ~n22163 ;
  assign n22165 = n22164 ^ n6539 ;
  assign n22167 = n22166 ^ n22165 ;
  assign n22168 = ~n22156 & ~n22167 ;
  assign n21972 = n21971 ^ n21958 ;
  assign n21973 = ~n21960 & n21972 ;
  assign n21974 = n21973 ^ n21971 ;
  assign n21812 = n20437 & n20729 ;
  assign n21810 = n6143 & n20725 ;
  assign n21803 = n20716 ^ x17 ;
  assign n21804 = n21803 ^ x16 ;
  assign n21805 = n21804 ^ n20716 ;
  assign n21806 = n20801 & n21805 ;
  assign n21807 = n21806 ^ n20716 ;
  assign n21808 = n6141 & n21807 ;
  assign n21809 = n21808 ^ x17 ;
  assign n21811 = n21810 ^ n21809 ;
  assign n21813 = n21812 ^ n21811 ;
  assign n21586 = n13433 & n20745 ;
  assign n21584 = n5426 & ~n20743 ;
  assign n21577 = n21575 ^ x20 ;
  assign n21578 = n21577 ^ x19 ;
  assign n21579 = n21578 ^ n21575 ;
  assign n21580 = n21574 & ~n21579 ;
  assign n21581 = n21580 ^ n21575 ;
  assign n21582 = n5215 & n21581 ;
  assign n21583 = n21582 ^ x20 ;
  assign n21585 = n21584 ^ n21583 ;
  assign n21587 = n21586 ^ n21585 ;
  assign n21390 = n21389 ^ n21333 ;
  assign n21391 = n21334 & n21390 ;
  assign n21392 = n21391 ^ n21333 ;
  assign n21319 = ~n40 & ~n20738 ;
  assign n21317 = n4656 & n21316 ;
  assign n21313 = n4655 & ~n20739 ;
  assign n21312 = n4651 & n20100 ;
  assign n21314 = n21313 ^ n21312 ;
  assign n21315 = n21314 ^ x23 ;
  assign n21318 = n21317 ^ n21315 ;
  assign n21320 = n21319 ^ n21318 ;
  assign n21309 = ~n4435 & n21308 ;
  assign n21305 = ~n4434 & n20746 ;
  assign n21302 = n4600 & n20750 ;
  assign n21301 = n20603 & ~n20747 ;
  assign n21303 = n21302 ^ n21301 ;
  assign n21304 = n21303 ^ x26 ;
  assign n21306 = n21305 ^ n21304 ;
  assign n21310 = n21309 ^ n21306 ;
  assign n21296 = ~n21294 & ~n21295 ;
  assign n21297 = n21278 & n21296 ;
  assign n21298 = n21297 ^ n21278 ;
  assign n21268 = n3833 & n20748 ;
  assign n21299 = n21298 ^ n21268 ;
  assign n21267 = n3832 & n20757 ;
  assign n21300 = n21299 ^ n21267 ;
  assign n21311 = n21310 ^ n21300 ;
  assign n21321 = n21320 ^ n21311 ;
  assign n21571 = n21392 ^ n21321 ;
  assign n21568 = n21567 ^ n21452 ;
  assign n21569 = ~n21453 & n21568 ;
  assign n21570 = n21569 ^ n21567 ;
  assign n21572 = n21571 ^ n21570 ;
  assign n21802 = n21587 ^ n21572 ;
  assign n21814 = n21813 ^ n21802 ;
  assign n22151 = n21974 ^ n21814 ;
  assign n22169 = n22168 ^ n22151 ;
  assign n22702 = n22483 ^ n22169 ;
  assign n22703 = n22702 ^ x11 ;
  assign n22705 = n22704 ^ n22703 ;
  assign n22707 = n22706 ^ n22705 ;
  assign n22700 = n7149 & n22091 ;
  assign n22699 = n7141 & ~n22090 ;
  assign n22701 = n22700 ^ n22699 ;
  assign n22708 = n22707 ^ n22701 ;
  assign n22698 = n7142 & ~n20694 ;
  assign n22709 = n22708 ^ n22698 ;
  assign n23279 = n22937 ^ n22709 ;
  assign n23280 = n23279 ^ n23277 ;
  assign n23288 = n23287 ^ n23280 ;
  assign n23289 = n23278 & ~n23288 ;
  assign n23290 = n23270 & n23289 ;
  assign n23291 = n23279 ^ n23268 ;
  assign n23292 = n23287 ^ x8 ;
  assign n23293 = n23292 ^ n23279 ;
  assign n23294 = n23291 & n23293 ;
  assign n23295 = n23294 ^ n23279 ;
  assign n23296 = ~n23290 & ~n23295 ;
  assign n23005 = n8139 & n20680 ;
  assign n22938 = n22937 ^ n22702 ;
  assign n22939 = n22709 & n22938 ;
  assign n22940 = n22939 ^ n22702 ;
  assign n22696 = n7142 & ~n20693 ;
  assign n22484 = n22483 ^ n22168 ;
  assign n22485 = ~n22169 & n22484 ;
  assign n22486 = n22485 ^ n22168 ;
  assign n22131 = ~n6529 & ~n20705 ;
  assign n22130 = ~n6547 & ~n20706 ;
  assign n22132 = n22131 ^ n22130 ;
  assign n22133 = n22132 ^ n6537 ;
  assign n22134 = n22133 ^ x14 ;
  assign n22145 = x13 & ~n22079 ;
  assign n22144 = n8856 & ~n20702 ;
  assign n22146 = n22145 ^ n22144 ;
  assign n22147 = ~n6539 & n22146 ;
  assign n22142 = n22078 ^ n8856 ;
  assign n22135 = n22132 ^ x14 ;
  assign n22137 = n20702 ^ x13 ;
  assign n22138 = n22137 ^ n20702 ;
  assign n22139 = ~n22078 & ~n22138 ;
  assign n22140 = n22139 ^ n20702 ;
  assign n22141 = ~n22135 & n22140 ;
  assign n22143 = n22142 ^ n22141 ;
  assign n22148 = n22147 ^ n22143 ;
  assign n22149 = ~n22134 & n22148 ;
  assign n21975 = n21974 ^ n21813 ;
  assign n21976 = n21814 & n21975 ;
  assign n21977 = n21976 ^ n21813 ;
  assign n21796 = n6148 & n20713 ;
  assign n21795 = n6143 & n20716 ;
  assign n21797 = n21796 ^ n21795 ;
  assign n21798 = n21797 ^ x17 ;
  assign n21794 = n6163 & n21793 ;
  assign n21799 = n21798 ^ n21794 ;
  assign n21792 = n20437 & n20725 ;
  assign n21800 = n21799 ^ n21792 ;
  assign n21604 = n13433 & ~n20743 ;
  assign n21602 = n5426 & n20737 ;
  assign n21595 = n20729 ^ x20 ;
  assign n21596 = n21595 ^ x19 ;
  assign n21597 = n21596 ^ n20729 ;
  assign n21598 = ~n21594 & n21597 ;
  assign n21599 = n21598 ^ n20729 ;
  assign n21600 = n5215 & n21599 ;
  assign n21601 = n21600 ^ x20 ;
  assign n21603 = n21602 ^ n21601 ;
  assign n21605 = n21604 ^ n21603 ;
  assign n21588 = n21587 ^ n21570 ;
  assign n21589 = ~n21572 & n21588 ;
  assign n21590 = n21589 ^ n21587 ;
  assign n21432 = ~n40 & ~n20739 ;
  assign n21430 = n4656 & ~n21429 ;
  assign n21423 = n4655 & n20745 ;
  assign n21422 = n4651 & ~n20738 ;
  assign n21424 = n21423 ^ n21422 ;
  assign n21425 = n21424 ^ x23 ;
  assign n21431 = n21430 ^ n21425 ;
  assign n21433 = n21432 ^ n21431 ;
  assign n21419 = ~n4435 & ~n21381 ;
  assign n21411 = n3983 & n21286 ;
  assign n21410 = n4369 & ~n20747 ;
  assign n21412 = n21411 ^ n21410 ;
  assign n21408 = n3985 & n20748 ;
  assign n21407 = n3837 & n20757 ;
  assign n21409 = n21408 ^ n21407 ;
  assign n21413 = n21412 ^ n21409 ;
  assign n21402 = x29 & ~n21268 ;
  assign n21403 = n3835 & n20757 ;
  assign n21404 = n21402 & n21403 ;
  assign n21405 = n21404 ^ n21402 ;
  assign n21406 = n21405 ^ x29 ;
  assign n21414 = n21413 ^ n21406 ;
  assign n21415 = n21414 ^ x26 ;
  assign n21401 = n4600 & n20746 ;
  assign n21416 = n21415 ^ n21401 ;
  assign n21400 = n20603 & n20750 ;
  assign n21417 = n21416 ^ n21400 ;
  assign n21399 = ~n4434 & n20100 ;
  assign n21418 = n21417 ^ n21399 ;
  assign n21420 = n21419 ^ n21418 ;
  assign n21396 = n21310 ^ n21298 ;
  assign n21397 = ~n21300 & n21396 ;
  assign n21398 = n21397 ^ n21310 ;
  assign n21421 = n21420 ^ n21398 ;
  assign n21434 = n21433 ^ n21421 ;
  assign n21393 = n21392 ^ n21320 ;
  assign n21394 = ~n21321 & n21393 ;
  assign n21395 = n21394 ^ n21392 ;
  assign n21435 = n21434 ^ n21395 ;
  assign n21591 = n21590 ^ n21435 ;
  assign n21791 = n21605 ^ n21591 ;
  assign n21801 = n21800 ^ n21791 ;
  assign n22129 = n21977 ^ n21801 ;
  assign n22150 = n22149 ^ n22129 ;
  assign n22691 = n22486 ^ n22150 ;
  assign n22692 = n22691 ^ x11 ;
  assign n22690 = n7151 & ~n20690 ;
  assign n22693 = n22692 ^ n22690 ;
  assign n22689 = n7148 & ~n20694 ;
  assign n22694 = n22693 ^ n22689 ;
  assign n22688 = n20240 & n21246 ;
  assign n22695 = n22694 ^ n22688 ;
  assign n22697 = n22696 ^ n22695 ;
  assign n23000 = n22940 ^ n22697 ;
  assign n23001 = n23000 ^ x8 ;
  assign n22999 = n8484 & n20631 ;
  assign n23002 = n23001 ^ n22999 ;
  assign n22998 = n8144 & ~n20683 ;
  assign n23003 = n23002 ^ n22998 ;
  assign n22649 = n21157 ^ n20814 ;
  assign n22653 = n22649 ^ n20631 ;
  assign n22997 = n8150 & ~n22653 ;
  assign n23004 = n23003 ^ n22997 ;
  assign n23006 = n23005 ^ n23004 ;
  assign n23860 = n23296 ^ n23006 ;
  assign n23542 = ~n10334 & n20680 ;
  assign n21236 = n21158 ^ n20815 ;
  assign n21237 = n21236 ^ n20819 ;
  assign n23540 = n10342 & ~n21237 ;
  assign n23537 = n10425 & n20819 ;
  assign n23536 = n10327 & n20631 ;
  assign n23538 = n23537 ^ n23536 ;
  assign n23539 = n23538 ^ x5 ;
  assign n23541 = n23540 ^ n23539 ;
  assign n23543 = n23542 ^ n23541 ;
  assign n23535 = n23278 ^ n23269 ;
  assign n23544 = n23543 ^ n23535 ;
  assign n23553 = ~n10334 & ~n20683 ;
  assign n23548 = n23264 ^ n23017 ;
  assign n23549 = n23548 ^ x5 ;
  assign n23547 = n10425 & n20631 ;
  assign n23550 = n23549 ^ n23547 ;
  assign n23546 = n10327 & n20680 ;
  assign n23551 = n23550 ^ n23546 ;
  assign n23545 = n10342 & ~n22653 ;
  assign n23552 = n23551 ^ n23545 ;
  assign n23554 = n23553 ^ n23552 ;
  assign n23563 = ~n10334 & ~n20690 ;
  assign n23560 = n10327 & ~n20683 ;
  assign n23558 = n10425 & n20680 ;
  assign n23556 = n23261 ^ n23027 ;
  assign n23557 = n23556 ^ x5 ;
  assign n23559 = n23558 ^ n23557 ;
  assign n23561 = n23560 ^ n23559 ;
  assign n23555 = n10342 & ~n22662 ;
  assign n23562 = n23561 ^ n23555 ;
  assign n23564 = n23563 ^ n23562 ;
  assign n23573 = ~n10334 & ~n20693 ;
  assign n23570 = n10327 & ~n20690 ;
  assign n23568 = n10425 & ~n20683 ;
  assign n23566 = n23258 ^ n23040 ;
  assign n23567 = n23566 ^ x5 ;
  assign n23569 = n23568 ^ n23567 ;
  assign n23571 = n23570 ^ n23569 ;
  assign n23565 = n10342 & n22618 ;
  assign n23572 = n23571 ^ n23565 ;
  assign n23574 = n23573 ^ n23572 ;
  assign n23583 = ~n10334 & ~n20694 ;
  assign n23580 = n10327 & ~n20693 ;
  assign n23578 = n10425 & ~n20690 ;
  assign n23576 = n23255 ^ n23050 ;
  assign n23577 = n23576 ^ x5 ;
  assign n23579 = n23578 ^ n23577 ;
  assign n23581 = n23580 ^ n23579 ;
  assign n23575 = n10342 & n21246 ;
  assign n23582 = n23581 ^ n23575 ;
  assign n23584 = n23583 ^ n23582 ;
  assign n23590 = n10425 & ~n20694 ;
  assign n23589 = n10327 & ~n20702 ;
  assign n23591 = n23590 ^ n23589 ;
  assign n23592 = n23591 ^ x5 ;
  assign n23588 = n10342 & n22601 ;
  assign n23593 = n23592 ^ n23588 ;
  assign n23587 = ~n10334 & ~n20705 ;
  assign n23594 = n23593 ^ n23587 ;
  assign n23586 = n23240 ^ n23061 ;
  assign n23595 = n23594 ^ n23586 ;
  assign n23600 = n10425 & ~n20702 ;
  assign n23599 = n10327 & ~n20705 ;
  assign n23601 = n23600 ^ n23599 ;
  assign n23602 = n23601 ^ x5 ;
  assign n23598 = n10342 & n22079 ;
  assign n23603 = n23602 ^ n23598 ;
  assign n23597 = ~n10334 & ~n20706 ;
  assign n23604 = n23603 ^ n23597 ;
  assign n23596 = n23237 ^ n23071 ;
  assign n23605 = n23604 ^ n23596 ;
  assign n23610 = n10425 & ~n20705 ;
  assign n23609 = n10327 & ~n20706 ;
  assign n23611 = n23610 ^ n23609 ;
  assign n23612 = n23611 ^ x5 ;
  assign n23608 = n10342 & n21770 ;
  assign n23613 = n23612 ^ n23608 ;
  assign n23607 = ~n10334 & n20713 ;
  assign n23614 = n23613 ^ n23607 ;
  assign n23606 = n23234 ^ n23081 ;
  assign n23615 = n23614 ^ n23606 ;
  assign n23799 = n23232 ^ n23222 ;
  assign n23621 = n10327 & n20725 ;
  assign n23620 = n10425 & n20716 ;
  assign n23622 = n23621 ^ n23620 ;
  assign n23623 = n23622 ^ x5 ;
  assign n23619 = n10342 & n21754 ;
  assign n23624 = n23623 ^ n23619 ;
  assign n23618 = ~n10334 & n20729 ;
  assign n23625 = n23624 ^ n23618 ;
  assign n23617 = n23205 ^ n23197 ;
  assign n23626 = n23625 ^ n23617 ;
  assign n23635 = n23193 ^ n23092 ;
  assign n23630 = n10425 & n20725 ;
  assign n23629 = n10327 & n20729 ;
  assign n23631 = n23630 ^ n23629 ;
  assign n23632 = n23631 ^ x5 ;
  assign n23628 = n10342 & n21736 ;
  assign n23633 = n23632 ^ n23628 ;
  assign n23627 = ~n10334 & n20737 ;
  assign n23634 = n23633 ^ n23627 ;
  assign n23636 = n23635 ^ n23634 ;
  assign n23646 = ~n10334 & n20745 ;
  assign n23643 = n10327 & ~n20743 ;
  assign n23641 = n10425 & n20737 ;
  assign n23639 = n23177 ^ n23102 ;
  assign n23640 = n23639 ^ x5 ;
  assign n23642 = n23641 ^ n23640 ;
  assign n23644 = n23643 ^ n23642 ;
  assign n23638 = n10342 & n21575 ;
  assign n23645 = n23644 ^ n23638 ;
  assign n23647 = n23646 ^ n23645 ;
  assign n23656 = ~n10334 & ~n20739 ;
  assign n23653 = n10327 & n20745 ;
  assign n23651 = n10425 & ~n20743 ;
  assign n23649 = n23175 ^ n23165 ;
  assign n23650 = n23649 ^ x5 ;
  assign n23652 = n23651 ^ n23650 ;
  assign n23654 = n23653 ^ n23652 ;
  assign n23648 = n10342 & n21440 ;
  assign n23655 = n23654 ^ n23648 ;
  assign n23657 = n23656 ^ n23655 ;
  assign n23665 = ~n10334 & ~n20738 ;
  assign n23663 = n10342 & ~n21429 ;
  assign n23660 = n10425 & n20745 ;
  assign n23659 = n10327 & ~n20739 ;
  assign n23661 = n23660 ^ n23659 ;
  assign n23662 = n23661 ^ x5 ;
  assign n23664 = n23663 ^ n23662 ;
  assign n23666 = n23665 ^ n23664 ;
  assign n23658 = n23160 ^ n23152 ;
  assign n23667 = n23666 ^ n23658 ;
  assign n23675 = ~n10334 & n20100 ;
  assign n23673 = n10342 & n21316 ;
  assign n23670 = n10425 & ~n20739 ;
  assign n23669 = n10327 & ~n20738 ;
  assign n23671 = n23670 ^ n23669 ;
  assign n23672 = n23671 ^ x5 ;
  assign n23674 = n23673 ^ n23672 ;
  assign n23676 = n23675 ^ n23674 ;
  assign n23668 = n23148 ^ n23140 ;
  assign n23677 = n23676 ^ n23668 ;
  assign n23686 = ~n10334 & n20746 ;
  assign n23684 = n10342 & n21329 ;
  assign n23681 = n10425 & ~n20738 ;
  assign n23680 = n10327 & n20100 ;
  assign n23682 = n23681 ^ n23680 ;
  assign n23683 = n23682 ^ x5 ;
  assign n23685 = n23684 ^ n23683 ;
  assign n23687 = n23686 ^ n23685 ;
  assign n23678 = n23128 ^ n23115 ;
  assign n23679 = n23678 ^ n23137 ;
  assign n23688 = n23687 ^ n23679 ;
  assign n23691 = n8137 & n20757 ;
  assign n23692 = n10322 & n20748 ;
  assign n23693 = x5 & ~n23692 ;
  assign n23694 = n20757 & n23693 ;
  assign n23695 = n10333 & n23694 ;
  assign n23696 = n23695 ^ n23693 ;
  assign n23697 = n23696 ^ x5 ;
  assign n23698 = n23697 ^ x5 ;
  assign n23709 = n10327 & n20748 ;
  assign n23707 = n10322 & ~n20747 ;
  assign n23703 = n10329 & n23692 ;
  assign n23704 = n23703 ^ n10334 ;
  assign n23705 = ~n20757 & ~n23704 ;
  assign n23706 = n23705 ^ n10334 ;
  assign n23708 = n23707 ^ n23706 ;
  assign n23710 = n23709 ^ n23708 ;
  assign n23711 = n23698 & n23710 ;
  assign n23712 = ~n23691 & ~n23711 ;
  assign n23716 = n10342 & ~n21276 ;
  assign n23715 = ~n10334 & n20748 ;
  assign n23717 = n23716 ^ n23715 ;
  assign n23718 = n23717 ^ x5 ;
  assign n23714 = n10327 & ~n20747 ;
  assign n23719 = n23718 ^ n23714 ;
  assign n23713 = n10425 & n20750 ;
  assign n23720 = n23719 ^ n23713 ;
  assign n23721 = n23712 & n23720 ;
  assign n23722 = n23721 ^ n23720 ;
  assign n23689 = n8136 & n20757 ;
  assign n23690 = n23689 ^ n23116 ;
  assign n23724 = n23722 ^ n23690 ;
  assign n23723 = n23690 & n23722 ;
  assign n23725 = n23724 ^ n23723 ;
  assign n23730 = n10342 & n21308 ;
  assign n23729 = ~n10334 & ~n20747 ;
  assign n23731 = n23730 ^ n23729 ;
  assign n23727 = n10425 & n20746 ;
  assign n23726 = n10327 & n20750 ;
  assign n23728 = n23727 ^ n23726 ;
  assign n23732 = n23731 ^ n23728 ;
  assign n23733 = n23732 ^ x5 ;
  assign n23741 = n23127 ^ n23119 ;
  assign n23742 = n23741 ^ n23732 ;
  assign n23738 = n10342 & ~n21381 ;
  assign n23737 = ~n10334 & n20750 ;
  assign n23739 = n23738 ^ n23737 ;
  assign n23735 = n10425 & n20100 ;
  assign n23734 = n10327 & n20746 ;
  assign n23736 = n23735 ^ n23734 ;
  assign n23740 = n23739 ^ n23736 ;
  assign n23743 = n23742 ^ n23740 ;
  assign n23744 = n23733 & ~n23743 ;
  assign n23745 = n23725 & n23744 ;
  assign n23746 = n23741 ^ n23723 ;
  assign n23747 = n23740 ^ x5 ;
  assign n23748 = n23747 ^ n23723 ;
  assign n23749 = n23746 & n23748 ;
  assign n23750 = n23749 ^ n23723 ;
  assign n23751 = ~n23745 & ~n23750 ;
  assign n23752 = n23751 ^ n23687 ;
  assign n23753 = n23688 & ~n23752 ;
  assign n23754 = n23753 ^ n23687 ;
  assign n23755 = n23754 ^ n23676 ;
  assign n23756 = n23677 & n23755 ;
  assign n23757 = n23756 ^ n23676 ;
  assign n23758 = n23757 ^ n23666 ;
  assign n23759 = n23667 & n23758 ;
  assign n23760 = n23759 ^ n23666 ;
  assign n23761 = n23760 ^ n23649 ;
  assign n23762 = n23657 & n23761 ;
  assign n23763 = n23762 ^ n23649 ;
  assign n23764 = n23763 ^ n23639 ;
  assign n23765 = n23647 & n23764 ;
  assign n23766 = n23765 ^ n23639 ;
  assign n23637 = n23191 ^ n23180 ;
  assign n23767 = n23766 ^ n23637 ;
  assign n23771 = n10425 & n20729 ;
  assign n23770 = n10327 & n20737 ;
  assign n23772 = n23771 ^ n23770 ;
  assign n23773 = n23772 ^ x5 ;
  assign n23769 = n10342 & ~n21593 ;
  assign n23774 = n23773 ^ n23769 ;
  assign n23768 = ~n10334 & ~n20743 ;
  assign n23775 = n23774 ^ n23768 ;
  assign n23776 = n23775 ^ n23637 ;
  assign n23777 = ~n23767 & n23776 ;
  assign n23778 = n23777 ^ n23766 ;
  assign n23779 = n23778 ^ n23634 ;
  assign n23780 = n23636 & ~n23779 ;
  assign n23781 = n23780 ^ n23635 ;
  assign n23782 = n23781 ^ n23625 ;
  assign n23783 = ~n23626 & n23782 ;
  assign n23784 = n23783 ^ n23625 ;
  assign n23616 = n23218 ^ n23210 ;
  assign n23785 = n23784 ^ n23616 ;
  assign n23794 = ~n10334 & n20725 ;
  assign n23792 = n10327 & n20716 ;
  assign n23791 = n23616 ^ x5 ;
  assign n23793 = n23792 ^ n23791 ;
  assign n23795 = n23794 ^ n23793 ;
  assign n22063 = n21793 ^ n20713 ;
  assign n23786 = n20713 ^ n10329 ;
  assign n23787 = n23786 ^ n20713 ;
  assign n23788 = n22063 & n23787 ;
  assign n23789 = n23788 ^ n20713 ;
  assign n23790 = n10322 & n23789 ;
  assign n23796 = n23795 ^ n23790 ;
  assign n23797 = ~n23785 & n23796 ;
  assign n23798 = n23797 ^ n23784 ;
  assign n23800 = n23799 ^ n23798 ;
  assign n23810 = n10327 & n20713 ;
  assign n23808 = ~n10334 & n20716 ;
  assign n23807 = n23799 ^ x5 ;
  assign n23809 = n23808 ^ n23807 ;
  assign n23811 = n23810 ^ n23809 ;
  assign n23801 = n21782 ^ n20706 ;
  assign n23802 = n20706 ^ n10329 ;
  assign n23803 = n23802 ^ n20706 ;
  assign n23804 = ~n23801 & n23803 ;
  assign n23805 = n23804 ^ n20706 ;
  assign n23806 = n10322 & ~n23805 ;
  assign n23812 = n23811 ^ n23806 ;
  assign n23813 = ~n23800 & ~n23812 ;
  assign n23814 = n23813 ^ n23799 ;
  assign n23815 = n23814 ^ n23614 ;
  assign n23816 = n23615 & ~n23815 ;
  assign n23817 = n23816 ^ n23614 ;
  assign n23818 = n23817 ^ n23604 ;
  assign n23819 = ~n23605 & n23818 ;
  assign n23820 = n23819 ^ n23604 ;
  assign n23821 = n23820 ^ n23594 ;
  assign n23822 = n23595 & n23821 ;
  assign n23823 = n23822 ^ n23594 ;
  assign n23585 = n23253 ^ n23243 ;
  assign n23824 = n23823 ^ n23585 ;
  assign n23832 = ~n10334 & ~n20702 ;
  assign n23828 = n23585 ^ x5 ;
  assign n23827 = n10425 & ~n20693 ;
  assign n23829 = n23828 ^ n23827 ;
  assign n23826 = n10327 & ~n20694 ;
  assign n23830 = n23829 ^ n23826 ;
  assign n23825 = n10342 & n22091 ;
  assign n23831 = n23830 ^ n23825 ;
  assign n23833 = n23832 ^ n23831 ;
  assign n23834 = ~n23824 & n23833 ;
  assign n23835 = n23834 ^ n23823 ;
  assign n23836 = n23835 ^ n23576 ;
  assign n23837 = n23584 & n23836 ;
  assign n23838 = n23837 ^ n23576 ;
  assign n23839 = n23838 ^ n23566 ;
  assign n23840 = ~n23574 & ~n23839 ;
  assign n23841 = n23840 ^ n23566 ;
  assign n23842 = n23841 ^ n23556 ;
  assign n23843 = n23564 & ~n23842 ;
  assign n23844 = n23843 ^ n23556 ;
  assign n23845 = n23844 ^ n23548 ;
  assign n23846 = ~n23554 & ~n23845 ;
  assign n23847 = n23846 ^ n23548 ;
  assign n23848 = n23847 ^ n23543 ;
  assign n23849 = n23544 & ~n23848 ;
  assign n23850 = n23849 ^ n23543 ;
  assign n23530 = n10327 & n20819 ;
  assign n23529 = n10425 & ~n20628 ;
  assign n23531 = n23530 ^ n23529 ;
  assign n23532 = n23531 ^ x5 ;
  assign n23306 = n21159 ^ n20820 ;
  assign n23307 = n23306 ^ n20628 ;
  assign n23528 = n10342 & n23307 ;
  assign n23533 = n23532 ^ n23528 ;
  assign n23527 = ~n10334 & n20631 ;
  assign n23534 = n23533 ^ n23527 ;
  assign n23851 = n23850 ^ n23534 ;
  assign n23854 = n23287 ^ n23279 ;
  assign n23855 = n23854 ^ n23277 ;
  assign n23856 = n23855 ^ n23534 ;
  assign n23852 = n23278 ^ n23007 ;
  assign n23853 = ~n23269 & n23852 ;
  assign n23857 = n23856 ^ n23853 ;
  assign n23858 = n23851 & ~n23857 ;
  assign n23859 = n23858 ^ n23850 ;
  assign n23861 = n23860 ^ n23859 ;
  assign n23869 = ~n10334 & n20819 ;
  assign n23865 = n23860 ^ x5 ;
  assign n23864 = n10425 & n20829 ;
  assign n23866 = n23865 ^ n23864 ;
  assign n23863 = n10327 & ~n20628 ;
  assign n23867 = n23866 ^ n23863 ;
  assign n22978 = n21160 ^ n20821 ;
  assign n22979 = n22978 ^ n20829 ;
  assign n23862 = n10342 & ~n22979 ;
  assign n23868 = n23867 ^ n23862 ;
  assign n23870 = n23869 ^ n23868 ;
  assign n23871 = ~n23861 & ~n23870 ;
  assign n23872 = n23871 ^ n23860 ;
  assign n23525 = ~n10334 & ~n20628 ;
  assign n23297 = n23296 ^ n23000 ;
  assign n23298 = n23006 & ~n23297 ;
  assign n23299 = n23298 ^ n23000 ;
  assign n22994 = n8139 & n20631 ;
  assign n22991 = n8144 & n20680 ;
  assign n22989 = n8484 & n20819 ;
  assign n22941 = n22940 ^ n22691 ;
  assign n22942 = ~n22697 & n22941 ;
  assign n22943 = n22942 ^ n22940 ;
  assign n22684 = n7142 & ~n20690 ;
  assign n22681 = n7148 & ~n20693 ;
  assign n22679 = n7151 & ~n20683 ;
  assign n22487 = n22486 ^ n22149 ;
  assign n22488 = n22150 & n22487 ;
  assign n22489 = n22488 ^ n22486 ;
  assign n21978 = n21977 ^ n21800 ;
  assign n21979 = ~n21801 & n21978 ;
  assign n21980 = n21979 ^ n21977 ;
  assign n21785 = n6143 & n20713 ;
  assign n21784 = n6148 & ~n20706 ;
  assign n21786 = n21785 ^ n21784 ;
  assign n21787 = n21786 ^ x17 ;
  assign n21783 = n6163 & n21782 ;
  assign n21788 = n21787 ^ n21783 ;
  assign n21780 = n20437 & n20716 ;
  assign n21789 = n21788 ^ n21780 ;
  assign n21747 = n13433 & n20737 ;
  assign n21745 = n5426 & n20729 ;
  assign n21738 = n21736 ^ x20 ;
  assign n21739 = n21738 ^ x19 ;
  assign n21740 = n21739 ^ n21736 ;
  assign n21741 = n20800 & ~n21740 ;
  assign n21742 = n21741 ^ n21736 ;
  assign n21743 = n5215 & n21742 ;
  assign n21744 = n21743 ^ x20 ;
  assign n21746 = n21745 ^ n21744 ;
  assign n21748 = n21747 ^ n21746 ;
  assign n21647 = ~n40 & n20745 ;
  assign n21645 = n4656 & n21440 ;
  assign n21642 = n4655 & ~n20743 ;
  assign n21641 = n4651 & ~n20739 ;
  assign n21643 = n21642 ^ n21641 ;
  assign n21644 = n21643 ^ x23 ;
  assign n21646 = n21645 ^ n21644 ;
  assign n21648 = n21647 ^ n21646 ;
  assign n21637 = n21414 ^ n21398 ;
  assign n21638 = n21420 & n21637 ;
  assign n21639 = n21638 ^ n21414 ;
  assign n21634 = ~n4435 & n21329 ;
  assign n21632 = ~n4434 & ~n20738 ;
  assign n21629 = n4600 & n20100 ;
  assign n21628 = n20603 & n20746 ;
  assign n21630 = n21629 ^ n21628 ;
  assign n21631 = n21630 ^ x26 ;
  assign n21633 = n21632 ^ n21631 ;
  assign n21635 = n21634 ^ n21633 ;
  assign n21624 = n3837 & n20748 ;
  assign n21622 = n3985 & ~n20747 ;
  assign n21615 = n20750 ^ x29 ;
  assign n21616 = n21615 ^ x28 ;
  assign n21617 = n21616 ^ n20750 ;
  assign n21618 = ~n21275 & n21617 ;
  assign n21619 = n21618 ^ n20750 ;
  assign n21620 = n3833 & n21619 ;
  assign n21621 = n21620 ^ x29 ;
  assign n21623 = n21622 ^ n21621 ;
  assign n21625 = n21624 ^ n21623 ;
  assign n21613 = n21405 & ~n21413 ;
  assign n21626 = n21625 ^ n21613 ;
  assign n21612 = n3518 & n20757 ;
  assign n21627 = n21626 ^ n21612 ;
  assign n21636 = n21635 ^ n21627 ;
  assign n21640 = n21639 ^ n21636 ;
  assign n21649 = n21648 ^ n21640 ;
  assign n21609 = n21433 ^ n21395 ;
  assign n21610 = n21434 & n21609 ;
  assign n21611 = n21610 ^ n21433 ;
  assign n21650 = n21649 ^ n21611 ;
  assign n21606 = n21605 ^ n21590 ;
  assign n21607 = ~n21591 & n21606 ;
  assign n21608 = n21607 ^ n21605 ;
  assign n21651 = n21650 ^ n21608 ;
  assign n21779 = n21748 ^ n21651 ;
  assign n21790 = n21789 ^ n21779 ;
  assign n22127 = n21980 ^ n21790 ;
  assign n22106 = ~n6529 & ~n20702 ;
  assign n22105 = ~n6547 & ~n20705 ;
  assign n22107 = n22106 ^ n22105 ;
  assign n22108 = n22107 ^ n6537 ;
  assign n22109 = n22108 ^ x14 ;
  assign n22110 = n22107 ^ x14 ;
  assign n22116 = n22110 ^ n6539 ;
  assign n22115 = n22110 & ~n22112 ;
  assign n22117 = n22116 ^ n22115 ;
  assign n22111 = n20694 ^ n17173 ;
  assign n22118 = n22111 ^ n20694 ;
  assign n22119 = ~n22112 & ~n22118 ;
  assign n22120 = n22119 ^ n20694 ;
  assign n22121 = ~n22116 & n22120 ;
  assign n22122 = ~n22117 & n22121 ;
  assign n22123 = n22122 ^ n22119 ;
  assign n22124 = n22123 ^ n6539 ;
  assign n22125 = n22124 ^ n20694 ;
  assign n22126 = ~n22109 & ~n22125 ;
  assign n22128 = n22127 ^ n22126 ;
  assign n22677 = n22489 ^ n22128 ;
  assign n22678 = n22677 ^ x11 ;
  assign n22680 = n22679 ^ n22678 ;
  assign n22682 = n22681 ^ n22680 ;
  assign n22676 = n20240 & n22618 ;
  assign n22683 = n22682 ^ n22676 ;
  assign n22685 = n22684 ^ n22683 ;
  assign n22987 = n22943 ^ n22685 ;
  assign n22988 = n22987 ^ x8 ;
  assign n22990 = n22989 ^ n22988 ;
  assign n22992 = n22991 ^ n22990 ;
  assign n22986 = n8150 & ~n21237 ;
  assign n22993 = n22992 ^ n22986 ;
  assign n22995 = n22994 ^ n22993 ;
  assign n23520 = n23299 ^ n22995 ;
  assign n23521 = n23520 ^ x5 ;
  assign n23519 = n10425 & n20624 ;
  assign n23522 = n23521 ^ n23519 ;
  assign n23518 = n10327 & n20829 ;
  assign n23523 = n23522 ^ n23518 ;
  assign n21231 = n21161 ^ n20830 ;
  assign n21232 = n21231 ^ n20624 ;
  assign n23517 = n10342 & ~n21232 ;
  assign n23524 = n23523 ^ n23517 ;
  assign n23526 = n23525 ^ n23524 ;
  assign n24148 = n23872 ^ n23526 ;
  assign n24743 = n24742 ^ n24148 ;
  assign n23479 = n21164 ^ n20833 ;
  assign n24134 = n20614 ^ x1 ;
  assign n24136 = n24135 ^ n24134 ;
  assign n24137 = n23479 & n24136 ;
  assign n24138 = n24137 ^ n24134 ;
  assign n24149 = n24148 ^ n24138 ;
  assign n24139 = n20617 ^ x2 ;
  assign n24142 = n24139 ^ n20617 ;
  assign n24143 = ~n20620 & n24142 ;
  assign n24144 = n24143 ^ n20617 ;
  assign n24145 = ~x1 & ~n24144 ;
  assign n24140 = n24139 ^ n24138 ;
  assign n24146 = n24145 ^ n24140 ;
  assign n24147 = ~x0 & n24146 ;
  assign n24150 = n24149 ^ n24147 ;
  assign n23490 = n21163 ^ n20832 ;
  assign n24706 = n20617 ^ x1 ;
  assign n24707 = n24706 ^ n24139 ;
  assign n24708 = n23490 & n24707 ;
  assign n24709 = n24708 ^ n24706 ;
  assign n24152 = n20620 ^ x2 ;
  assign n24712 = n24709 ^ n24152 ;
  assign n24713 = n24712 ^ n24709 ;
  assign n24714 = n24713 ^ n20620 ;
  assign n24715 = n20624 & n24714 ;
  assign n24716 = n24715 ^ n20620 ;
  assign n24717 = ~x1 & ~n24716 ;
  assign n24718 = n24717 ^ n24712 ;
  assign n24719 = ~x0 & n24718 ;
  assign n24720 = n24719 ^ n24709 ;
  assign n24725 = n24720 ^ n24148 ;
  assign n24183 = n23847 ^ n23544 ;
  assign n24170 = n20624 ^ x1 ;
  assign n24158 = n20624 ^ x2 ;
  assign n24171 = n24170 ^ n24158 ;
  assign n24172 = n21231 & n24171 ;
  assign n24173 = n24172 ^ n24170 ;
  assign n24184 = n24183 ^ n24173 ;
  assign n24168 = n20829 ^ n20628 ;
  assign n24169 = n24168 ^ n20829 ;
  assign n24174 = n20829 ^ x2 ;
  assign n24177 = n24174 ^ n20829 ;
  assign n24178 = ~n24169 & n24177 ;
  assign n24179 = n24178 ^ n20829 ;
  assign n24180 = ~x1 & n24179 ;
  assign n24175 = n24174 ^ n24173 ;
  assign n24181 = n24180 ^ n24175 ;
  assign n24182 = ~x0 & n24181 ;
  assign n24185 = n24184 ^ n24182 ;
  assign n24682 = n20819 ^ n20628 ;
  assign n24683 = n24682 ^ n20628 ;
  assign n24677 = n20829 ^ x1 ;
  assign n24678 = n24677 ^ x2 ;
  assign n24679 = n24678 ^ n20829 ;
  assign n24680 = n22978 & n24679 ;
  assign n24681 = n24680 ^ n24677 ;
  assign n24189 = n20628 ^ x2 ;
  assign n24684 = n24681 ^ n24189 ;
  assign n24685 = n24684 ^ n24681 ;
  assign n24686 = n24685 ^ n20628 ;
  assign n24687 = n24683 & n24686 ;
  assign n24688 = n24687 ^ n20628 ;
  assign n24689 = ~x1 & ~n24688 ;
  assign n24690 = n24689 ^ n24684 ;
  assign n24691 = ~x0 & ~n24690 ;
  assign n24692 = n24691 ^ n24681 ;
  assign n24697 = n24692 ^ n24183 ;
  assign n24202 = n23841 ^ n23564 ;
  assign n24188 = n20628 ^ x1 ;
  assign n24190 = n24189 ^ n24188 ;
  assign n24191 = n23306 & n24190 ;
  assign n24192 = n24191 ^ n24188 ;
  assign n24203 = n24202 ^ n24192 ;
  assign n24186 = n20819 ^ n20631 ;
  assign n24187 = n24186 ^ n20819 ;
  assign n24193 = n20819 ^ x2 ;
  assign n24196 = n24193 ^ n20819 ;
  assign n24197 = n24187 & n24196 ;
  assign n24198 = n24197 ^ n20819 ;
  assign n24199 = ~x1 & n24198 ;
  assign n24194 = n24193 ^ n24192 ;
  assign n24200 = n24199 ^ n24194 ;
  assign n24201 = ~x0 & ~n24200 ;
  assign n24204 = n24203 ^ n24201 ;
  assign n24658 = n20680 ^ n20631 ;
  assign n24659 = n24658 ^ n20631 ;
  assign n24653 = n20819 ^ x1 ;
  assign n24654 = n24653 ^ x2 ;
  assign n24655 = n24654 ^ n20819 ;
  assign n24656 = n21236 & n24655 ;
  assign n24657 = n24656 ^ n24653 ;
  assign n24208 = n20631 ^ x2 ;
  assign n24660 = n24657 ^ n24208 ;
  assign n24661 = n24660 ^ n24657 ;
  assign n24662 = n24661 ^ n20631 ;
  assign n24663 = n24659 & n24662 ;
  assign n24664 = n24663 ^ n20631 ;
  assign n24665 = ~x1 & n24664 ;
  assign n24666 = n24665 ^ n24660 ;
  assign n24667 = ~x0 & n24666 ;
  assign n24668 = n24667 ^ n24657 ;
  assign n24673 = n24668 ^ n24202 ;
  assign n24221 = n23835 ^ n23584 ;
  assign n24207 = n20631 ^ x1 ;
  assign n24209 = n24208 ^ n24207 ;
  assign n24210 = n22649 & n24209 ;
  assign n24211 = n24210 ^ n24207 ;
  assign n24222 = n24221 ^ n24211 ;
  assign n24212 = n20680 ^ x2 ;
  assign n24215 = n24212 ^ n20680 ;
  assign n24216 = ~n20683 & n24215 ;
  assign n24217 = n24216 ^ n20680 ;
  assign n24218 = ~x1 & n24217 ;
  assign n24213 = n24212 ^ n24211 ;
  assign n24219 = n24218 ^ n24213 ;
  assign n24220 = ~x0 & n24219 ;
  assign n24223 = n24222 ^ n24220 ;
  assign n24228 = n20680 ^ x1 ;
  assign n24229 = n24228 ^ n24212 ;
  assign n24230 = n22661 & n24229 ;
  assign n24231 = n24230 ^ n24228 ;
  assign n24224 = n23833 ^ n23823 ;
  assign n24241 = n24231 ^ n24224 ;
  assign n24232 = n20683 ^ x2 ;
  assign n24235 = n24232 ^ n20683 ;
  assign n24236 = ~n20690 & n24235 ;
  assign n24237 = n24236 ^ n20683 ;
  assign n24238 = ~x1 & ~n24237 ;
  assign n24233 = n24232 ^ n24231 ;
  assign n24239 = n24238 ^ n24233 ;
  assign n24240 = ~x0 & ~n24239 ;
  assign n24242 = n24241 ^ n24240 ;
  assign n24247 = n20683 ^ x1 ;
  assign n24248 = n24247 ^ n24232 ;
  assign n24249 = n22617 & n24248 ;
  assign n24250 = n24249 ^ n24247 ;
  assign n24243 = n23820 ^ n23595 ;
  assign n24260 = n24250 ^ n24243 ;
  assign n24251 = n20690 ^ x2 ;
  assign n24254 = n24251 ^ n20690 ;
  assign n24255 = ~n20693 & n24254 ;
  assign n24256 = n24255 ^ n20690 ;
  assign n24257 = ~x1 & ~n24256 ;
  assign n24252 = n24251 ^ n24250 ;
  assign n24258 = n24257 ^ n24252 ;
  assign n24259 = ~x0 & n24258 ;
  assign n24261 = n24260 ^ n24259 ;
  assign n24294 = n23814 ^ n23615 ;
  assign n24268 = n20693 ^ x2 ;
  assign n24271 = n24268 ^ n20693 ;
  assign n24272 = ~n20694 & n24271 ;
  assign n24273 = n24272 ^ n20693 ;
  assign n24274 = ~x1 & ~n24273 ;
  assign n24262 = n20690 ^ x1 ;
  assign n24263 = n24262 ^ n24251 ;
  assign n24264 = n21244 & n24263 ;
  assign n24265 = n24264 ^ n24262 ;
  assign n24269 = n24268 ^ n24265 ;
  assign n24275 = n24274 ^ n24269 ;
  assign n24276 = ~x0 & n24275 ;
  assign n24277 = n24276 ^ n24265 ;
  assign n24641 = n24294 ^ n24277 ;
  assign n24281 = n20693 ^ x1 ;
  assign n24282 = n24281 ^ n24268 ;
  assign n24283 = n22090 & n24282 ;
  assign n24284 = n24283 ^ n24281 ;
  assign n24295 = n24294 ^ n24284 ;
  assign n24285 = n20694 ^ x2 ;
  assign n24288 = n24285 ^ n20694 ;
  assign n24289 = ~n20702 & n24288 ;
  assign n24290 = n24289 ^ n20694 ;
  assign n24291 = ~x1 & ~n24290 ;
  assign n24286 = n24285 ^ n24284 ;
  assign n24292 = n24291 ^ n24286 ;
  assign n24293 = ~x0 & n24292 ;
  assign n24296 = n24295 ^ n24293 ;
  assign n24305 = n20694 ^ x1 ;
  assign n24299 = n20702 ^ x2 ;
  assign n24300 = n24299 ^ n20702 ;
  assign n24301 = ~n20705 & n24300 ;
  assign n24302 = n24301 ^ n20702 ;
  assign n24303 = ~x1 & ~n24302 ;
  assign n24304 = n24303 ^ n24299 ;
  assign n24306 = n24305 ^ n24304 ;
  assign n24307 = n24306 ^ x2 ;
  assign n24308 = n24307 ^ x1 ;
  assign n24309 = n24308 ^ n24306 ;
  assign n24310 = n24306 ^ n22112 ;
  assign n24311 = n24310 ^ n24306 ;
  assign n24312 = n24309 & n24311 ;
  assign n24313 = n24312 ^ n24306 ;
  assign n24314 = x0 & n24313 ;
  assign n24315 = n24314 ^ n24304 ;
  assign n24638 = n24315 ^ n24294 ;
  assign n24326 = n23778 ^ n23636 ;
  assign n24316 = n23781 ^ n23626 ;
  assign n24595 = n24326 ^ n24316 ;
  assign n24328 = n20713 ^ x2 ;
  assign n24322 = n20706 ^ x2 ;
  assign n24321 = n20706 ^ x1 ;
  assign n24323 = n24322 ^ n24321 ;
  assign n24324 = n21781 & n24323 ;
  assign n24325 = n24324 ^ n24321 ;
  assign n24329 = n24328 ^ n24325 ;
  assign n24330 = n24329 ^ n24325 ;
  assign n24331 = n24330 ^ n20713 ;
  assign n24332 = n22189 & n24331 ;
  assign n24333 = n24332 ^ n20713 ;
  assign n24334 = ~x1 & n24333 ;
  assign n24335 = n24334 ^ n24329 ;
  assign n24336 = ~x0 & ~n24335 ;
  assign n24327 = n24326 ^ n24325 ;
  assign n24337 = n24336 ^ n24327 ;
  assign n24354 = n23775 ^ n23767 ;
  assign n24343 = n20726 ^ n20716 ;
  assign n24344 = n20716 ^ x2 ;
  assign n24347 = n24344 ^ n20716 ;
  assign n24348 = n24343 & n24347 ;
  assign n24349 = n24348 ^ n20716 ;
  assign n24350 = ~x1 & n24349 ;
  assign n24338 = n20713 ^ x1 ;
  assign n24339 = n24338 ^ x2 ;
  assign n24340 = n24339 ^ n20713 ;
  assign n24341 = ~n20802 & n24340 ;
  assign n24342 = n24341 ^ n24338 ;
  assign n24345 = n24344 ^ n24342 ;
  assign n24351 = n24350 ^ n24345 ;
  assign n24352 = ~x0 & n24351 ;
  assign n24353 = n24352 ^ n24342 ;
  assign n24355 = n24354 ^ n24353 ;
  assign n24364 = n23760 ^ n23657 ;
  assign n24357 = n23763 ^ n23647 ;
  assign n24568 = n24364 ^ n24357 ;
  assign n24367 = n20729 ^ x2 ;
  assign n24370 = n24367 ^ n20729 ;
  assign n24371 = n20737 & n24370 ;
  assign n24372 = n24371 ^ n20729 ;
  assign n24373 = ~x1 & n24372 ;
  assign n24359 = n20725 ^ x1 ;
  assign n24360 = n24359 ^ x2 ;
  assign n24361 = n24360 ^ n20725 ;
  assign n24362 = ~n20800 & n24361 ;
  assign n24363 = n24362 ^ n24359 ;
  assign n24368 = n24367 ^ n24363 ;
  assign n24374 = n24373 ^ n24368 ;
  assign n24375 = ~x0 & n24374 ;
  assign n24365 = n24364 ^ n24363 ;
  assign n24376 = n24375 ^ n24365 ;
  assign n24393 = n23757 ^ n23667 ;
  assign n24379 = n20729 ^ x1 ;
  assign n24378 = n21593 ^ x2 ;
  assign n24380 = n24379 ^ n24378 ;
  assign n24381 = n20798 & ~n24380 ;
  assign n24382 = n24381 ^ n24379 ;
  assign n24383 = n24382 ^ x2 ;
  assign n24384 = n24383 ^ n20737 ;
  assign n24385 = n24384 ^ n24382 ;
  assign n24386 = n24385 ^ n20780 ;
  assign n24387 = ~n20743 & ~n24386 ;
  assign n24388 = n24387 ^ n20780 ;
  assign n24389 = ~x1 & ~n24388 ;
  assign n24390 = n24389 ^ n24384 ;
  assign n24391 = ~x0 & n24390 ;
  assign n24392 = n24391 ^ n24382 ;
  assign n24394 = n24393 ^ n24392 ;
  assign n24522 = n23751 ^ n23688 ;
  assign n24396 = n23754 ^ n23677 ;
  assign n24544 = n24522 ^ n24396 ;
  assign n24425 = n20745 ^ x1 ;
  assign n24417 = n20739 ^ x2 ;
  assign n24418 = n24417 ^ n20739 ;
  assign n24419 = n20739 ^ n20738 ;
  assign n24420 = n24419 ^ n20739 ;
  assign n24421 = n24418 & ~n24420 ;
  assign n24422 = n24421 ^ n20739 ;
  assign n24423 = ~x1 & ~n24422 ;
  assign n24424 = n24423 ^ n24417 ;
  assign n24426 = n24425 ^ n24424 ;
  assign n24427 = n24426 ^ x2 ;
  assign n24428 = n24427 ^ x1 ;
  assign n24429 = n24428 ^ n24426 ;
  assign n24430 = n24426 ^ n21428 ;
  assign n24431 = n24430 ^ n24426 ;
  assign n24432 = n24429 & n24431 ;
  assign n24433 = n24432 ^ n24426 ;
  assign n24434 = x0 & ~n24433 ;
  assign n24435 = n24434 ^ n24424 ;
  assign n24523 = n24522 ^ n24435 ;
  assign n24415 = n23733 ^ n23724 ;
  assign n24403 = n20738 ^ n20100 ;
  assign n24404 = n24403 ^ n20738 ;
  assign n24405 = n20738 ^ x2 ;
  assign n24408 = n24405 ^ n20738 ;
  assign n24409 = n24404 & n24408 ;
  assign n24410 = n24409 ^ n20738 ;
  assign n24411 = ~x1 & ~n24410 ;
  assign n24398 = n20739 ^ x1 ;
  assign n24399 = n24398 ^ x2 ;
  assign n24400 = n24399 ^ n20739 ;
  assign n24401 = n20774 & n24400 ;
  assign n24402 = n24401 ^ n24398 ;
  assign n24406 = n24405 ^ n24402 ;
  assign n24412 = n24411 ^ n24406 ;
  assign n24413 = ~x0 & n24412 ;
  assign n24414 = n24413 ^ n24402 ;
  assign n24416 = n24415 ^ n24414 ;
  assign n24451 = x2 & n20746 ;
  assign n24452 = n24451 ^ n20100 ;
  assign n24453 = ~x1 & n24452 ;
  assign n24447 = n20100 ^ x2 ;
  assign n24440 = n20738 ^ x1 ;
  assign n24441 = n24440 ^ n24405 ;
  assign n24442 = n21328 & n24441 ;
  assign n24443 = n24442 ^ n24440 ;
  assign n24448 = n24447 ^ n24443 ;
  assign n24454 = n24453 ^ n24448 ;
  assign n24455 = ~x0 & ~n24454 ;
  assign n24437 = n23720 ^ n23711 ;
  assign n24438 = n24437 ^ n23691 ;
  assign n24444 = n24443 ^ n24438 ;
  assign n24456 = n24455 ^ n24444 ;
  assign n24498 = n11141 & n20746 ;
  assign n24497 = n11139 & n20750 ;
  assign n24499 = n24498 ^ n24497 ;
  assign n24492 = n20100 ^ n11012 ;
  assign n24493 = n24492 ^ n20100 ;
  assign n24494 = ~n21380 & n24493 ;
  assign n24495 = n24494 ^ n20100 ;
  assign n24496 = x0 & n24495 ;
  assign n24500 = n24499 ^ n24496 ;
  assign n24489 = n23710 ^ n23697 ;
  assign n24501 = n24500 ^ n24489 ;
  assign n24502 = n24501 ^ n24500 ;
  assign n24510 = n24502 ^ n24438 ;
  assign n24484 = n11395 & n20757 ;
  assign n24485 = n24484 ^ n23692 ;
  assign n24504 = n24502 ^ n24500 ;
  assign n24481 = n11141 & n20750 ;
  assign n24480 = n11139 & ~n20747 ;
  assign n24482 = n24481 ^ n24480 ;
  assign n24477 = n11012 & n21307 ;
  assign n24478 = n24477 ^ n20746 ;
  assign n24479 = x0 & n24478 ;
  assign n24483 = n24482 ^ n24479 ;
  assign n24505 = n24504 ^ n24483 ;
  assign n24506 = n24485 & n24505 ;
  assign n24458 = n20750 ^ n11012 ;
  assign n24459 = n24458 ^ n20750 ;
  assign n24460 = ~n21275 & n24459 ;
  assign n24461 = n24460 ^ n20750 ;
  assign n24462 = x0 & n24461 ;
  assign n24467 = n24462 ^ x3 ;
  assign n24466 = n11141 & ~n20747 ;
  assign n24468 = n24467 ^ n24466 ;
  assign n24465 = n11139 & n20748 ;
  assign n24469 = n24468 ^ n24465 ;
  assign n24470 = n10322 & ~n24469 ;
  assign n24471 = n20757 & n24470 ;
  assign n24457 = x2 & n20747 ;
  assign n24463 = n21284 & ~n24462 ;
  assign n24464 = n24457 & n24463 ;
  assign n24472 = n24471 ^ n24464 ;
  assign n24486 = n24485 ^ n24483 ;
  assign n24487 = n24486 ^ x2 ;
  assign n24488 = n24472 & n24487 ;
  assign n24503 = n24502 ^ n24488 ;
  assign n24507 = n24506 ^ n24503 ;
  assign n24508 = n24504 ^ x2 ;
  assign n24509 = ~n24507 & ~n24508 ;
  assign n24511 = n24510 ^ n24509 ;
  assign n24512 = ~n24456 & ~n24511 ;
  assign n24439 = n24438 ^ n24435 ;
  assign n24513 = n24512 ^ n24439 ;
  assign n24436 = n24435 ^ n24414 ;
  assign n24514 = n24513 ^ n24436 ;
  assign n24515 = n24416 & ~n24514 ;
  assign n24516 = n24515 ^ n24513 ;
  assign n24519 = n24435 ^ n23743 ;
  assign n24517 = n23733 ^ n23722 ;
  assign n24518 = ~n23724 & n24517 ;
  assign n24520 = n24519 ^ n24518 ;
  assign n24521 = ~n24516 & ~n24520 ;
  assign n24524 = n24523 ^ n24521 ;
  assign n24531 = n20745 ^ n20739 ;
  assign n24532 = n24531 ^ n20745 ;
  assign n24533 = n20745 ^ x2 ;
  assign n24526 = n20743 ^ x2 ;
  assign n24525 = n20743 ^ x1 ;
  assign n24527 = n24526 ^ n24525 ;
  assign n24528 = n21439 & n24527 ;
  assign n24529 = n24528 ^ n24525 ;
  assign n24534 = n24533 ^ n24529 ;
  assign n24535 = n24534 ^ n24529 ;
  assign n24536 = n24535 ^ n20745 ;
  assign n24537 = ~n24532 & n24536 ;
  assign n24538 = n24537 ^ n20745 ;
  assign n24539 = ~x1 & n24538 ;
  assign n24540 = n24539 ^ n24534 ;
  assign n24541 = ~x0 & ~n24540 ;
  assign n24530 = n24529 ^ n24522 ;
  assign n24542 = n24541 ^ n24530 ;
  assign n24543 = n24524 & n24542 ;
  assign n24545 = n24544 ^ n24543 ;
  assign n24546 = n20737 ^ x1 ;
  assign n24547 = n24546 ^ x2 ;
  assign n24548 = n24547 ^ n20737 ;
  assign n24549 = ~n21574 & n24548 ;
  assign n24550 = n24549 ^ n24546 ;
  assign n24553 = n24550 ^ n24526 ;
  assign n24554 = n24553 ^ n24550 ;
  assign n24555 = n24554 ^ n20743 ;
  assign n24556 = n20745 & n24555 ;
  assign n24557 = n24556 ^ n20743 ;
  assign n24558 = ~x1 & ~n24557 ;
  assign n24559 = n24558 ^ n24553 ;
  assign n24560 = ~x0 & ~n24559 ;
  assign n24551 = n24550 ^ n24396 ;
  assign n24561 = n24560 ^ n24551 ;
  assign n24562 = ~n24545 & n24561 ;
  assign n24397 = n24396 ^ n24364 ;
  assign n24563 = n24562 ^ n24397 ;
  assign n24395 = n24392 ^ n24364 ;
  assign n24564 = n24563 ^ n24395 ;
  assign n24565 = ~n24394 & n24564 ;
  assign n24566 = n24565 ^ n24563 ;
  assign n24567 = n24376 & n24566 ;
  assign n24569 = n24568 ^ n24567 ;
  assign n24570 = n20725 ^ x2 ;
  assign n24571 = n24570 ^ n20725 ;
  assign n24572 = n24570 ^ n20730 ;
  assign n24573 = n24571 & n24572 ;
  assign n24574 = n24573 ^ n24570 ;
  assign n24575 = ~x1 & n24574 ;
  assign n24576 = n24575 ^ n24570 ;
  assign n24587 = n24576 ^ n24357 ;
  assign n24577 = n20716 ^ x1 ;
  assign n24578 = n24577 ^ n24576 ;
  assign n24579 = n24578 ^ x2 ;
  assign n24580 = n24579 ^ x1 ;
  assign n24581 = n24580 ^ n24578 ;
  assign n24582 = n24578 ^ n20801 ;
  assign n24583 = n24582 ^ n24578 ;
  assign n24584 = n24581 & ~n24583 ;
  assign n24585 = n24584 ^ n24578 ;
  assign n24586 = x0 & n24585 ;
  assign n24588 = n24587 ^ n24586 ;
  assign n24589 = n24569 & n24588 ;
  assign n24358 = n24357 ^ n24326 ;
  assign n24590 = n24589 ^ n24358 ;
  assign n24356 = n24353 ^ n24326 ;
  assign n24591 = n24590 ^ n24356 ;
  assign n24592 = n24355 & n24591 ;
  assign n24593 = n24592 ^ n24590 ;
  assign n24594 = ~n24337 & n24593 ;
  assign n24596 = n24595 ^ n24594 ;
  assign n24603 = n20713 ^ n20706 ;
  assign n24604 = n24603 ^ n20706 ;
  assign n24598 = n20705 ^ x1 ;
  assign n24597 = n20705 ^ x2 ;
  assign n24599 = n24598 ^ n24597 ;
  assign n24600 = n21769 & n24599 ;
  assign n24601 = n24600 ^ n24598 ;
  assign n24605 = n24601 ^ n24322 ;
  assign n24606 = n24605 ^ n24601 ;
  assign n24607 = n24606 ^ n20706 ;
  assign n24608 = n24604 & n24607 ;
  assign n24609 = n24608 ^ n20706 ;
  assign n24610 = ~x1 & ~n24609 ;
  assign n24611 = n24610 ^ n24605 ;
  assign n24612 = ~x0 & n24611 ;
  assign n24602 = n24601 ^ n24316 ;
  assign n24613 = n24612 ^ n24602 ;
  assign n24614 = ~n24596 & n24613 ;
  assign n24318 = n23796 ^ n23784 ;
  assign n24319 = n24318 ^ n24315 ;
  assign n24317 = n24316 ^ n24315 ;
  assign n24320 = n24319 ^ n24317 ;
  assign n24615 = n24614 ^ n24320 ;
  assign n24616 = n20702 ^ x1 ;
  assign n24617 = n24616 ^ n24299 ;
  assign n24618 = n22078 & n24617 ;
  assign n24619 = n24618 ^ n24616 ;
  assign n24624 = n24619 ^ n24597 ;
  assign n24625 = n24624 ^ n24619 ;
  assign n24626 = n24625 ^ n20705 ;
  assign n24627 = ~n20706 & n24626 ;
  assign n24628 = n24627 ^ n20705 ;
  assign n24629 = ~x1 & ~n24628 ;
  assign n24630 = n24629 ^ n24624 ;
  assign n24631 = ~x0 & n24630 ;
  assign n24620 = n24319 ^ n24315 ;
  assign n24621 = n24620 ^ n24619 ;
  assign n24632 = n24631 ^ n24621 ;
  assign n24633 = n24615 & n24632 ;
  assign n24634 = n24633 ^ n24319 ;
  assign n24635 = n24315 ^ n23812 ;
  assign n24636 = n24635 ^ n23798 ;
  assign n24637 = n24634 & n24636 ;
  assign n24639 = n24638 ^ n24637 ;
  assign n24640 = n24296 & n24639 ;
  assign n24642 = n24641 ^ n24640 ;
  assign n24643 = n24277 ^ n23817 ;
  assign n24644 = n24643 ^ n23605 ;
  assign n24645 = n24642 & n24644 ;
  assign n24278 = n24277 ^ n24243 ;
  assign n24646 = n24645 ^ n24278 ;
  assign n24647 = ~n24261 & ~n24646 ;
  assign n24244 = n24243 ^ n24224 ;
  assign n24648 = n24647 ^ n24244 ;
  assign n24649 = ~n24242 & ~n24648 ;
  assign n24225 = n24224 ^ n24221 ;
  assign n24650 = n24649 ^ n24225 ;
  assign n24651 = n24223 & ~n24650 ;
  assign n24652 = n24651 ^ n24221 ;
  assign n24669 = n24668 ^ n24652 ;
  assign n24670 = n23838 ^ n23574 ;
  assign n24671 = n24670 ^ n24652 ;
  assign n24672 = n24669 & n24671 ;
  assign n24674 = n24673 ^ n24672 ;
  assign n24675 = n24204 & ~n24674 ;
  assign n24676 = n24675 ^ n24202 ;
  assign n24693 = n24692 ^ n24676 ;
  assign n24694 = n23844 ^ n23554 ;
  assign n24695 = n24694 ^ n24676 ;
  assign n24696 = ~n24693 & ~n24695 ;
  assign n24698 = n24697 ^ n24696 ;
  assign n24699 = ~n24185 & ~n24698 ;
  assign n24700 = n24699 ^ n24183 ;
  assign n24161 = n24158 ^ n20624 ;
  assign n24162 = n20829 & n24161 ;
  assign n24163 = n24162 ^ n20624 ;
  assign n24164 = ~x1 & n24163 ;
  assign n22963 = n21162 ^ n20831 ;
  assign n24151 = n20620 ^ x1 ;
  assign n24153 = n24152 ^ n24151 ;
  assign n24154 = n22963 & n24153 ;
  assign n24155 = n24154 ^ n24151 ;
  assign n24159 = n24158 ^ n24155 ;
  assign n24165 = n24164 ^ n24159 ;
  assign n24166 = ~x0 & ~n24165 ;
  assign n24167 = n24166 ^ n24155 ;
  assign n24701 = n24700 ^ n24167 ;
  assign n24702 = n23857 ^ n23850 ;
  assign n24703 = n24702 ^ n24167 ;
  assign n24704 = n24701 & n24703 ;
  assign n24705 = n24704 ^ n24700 ;
  assign n24721 = n24720 ^ n24705 ;
  assign n24722 = n23870 ^ n23859 ;
  assign n24723 = n24722 ^ n24705 ;
  assign n24724 = n24721 & ~n24723 ;
  assign n24726 = n24725 ^ n24724 ;
  assign n24727 = n24150 & n24726 ;
  assign n24744 = n24743 ^ n24727 ;
  assign n23513 = ~n10334 & n20829 ;
  assign n23310 = n8484 & ~n20628 ;
  assign n23309 = n8144 & n20631 ;
  assign n23311 = n23310 ^ n23309 ;
  assign n23312 = n23311 ^ x8 ;
  assign n23308 = n8150 & n23307 ;
  assign n23313 = n23312 ^ n23308 ;
  assign n23305 = n8139 & n20819 ;
  assign n23314 = n23313 ^ n23305 ;
  assign n22673 = n7148 & ~n20690 ;
  assign n22671 = n7142 & ~n20683 ;
  assign n22664 = n20680 ^ x11 ;
  assign n22665 = n22664 ^ x10 ;
  assign n22666 = n22665 ^ n20680 ;
  assign n22667 = ~n22661 & n22666 ;
  assign n22668 = n22667 ^ n20680 ;
  assign n22669 = n7140 & n22668 ;
  assign n22670 = n22669 ^ x11 ;
  assign n22672 = n22671 ^ n22670 ;
  assign n22674 = n22673 ^ n22672 ;
  assign n22686 = n22677 ^ n22674 ;
  assign n22687 = n22686 ^ n22674 ;
  assign n22944 = n22943 ^ n22687 ;
  assign n22945 = n22685 & n22944 ;
  assign n22946 = n22945 ^ n22686 ;
  assign n22099 = ~n6529 & ~n20694 ;
  assign n22098 = ~n6547 & ~n20702 ;
  assign n22100 = n22099 ^ n22098 ;
  assign n22101 = n22100 ^ x14 ;
  assign n22092 = n22091 ^ n20693 ;
  assign n22093 = n20693 ^ n7310 ;
  assign n22094 = n22093 ^ n20693 ;
  assign n22095 = ~n22092 & n22094 ;
  assign n22096 = n22095 ^ n20693 ;
  assign n22097 = n6391 & ~n22096 ;
  assign n22102 = n22101 ^ n22097 ;
  assign n22490 = n22127 ^ n22102 ;
  assign n22491 = n22490 ^ n22489 ;
  assign n22492 = n22491 ^ n22102 ;
  assign n22493 = ~n22128 & ~n22492 ;
  assign n22494 = n22493 ^ n22490 ;
  assign n21981 = n21980 ^ n21789 ;
  assign n21982 = n21790 & n21981 ;
  assign n21983 = n21982 ^ n21789 ;
  assign n21773 = n6148 & ~n20705 ;
  assign n21772 = n6143 & ~n20706 ;
  assign n21774 = n21773 ^ n21772 ;
  assign n21775 = n21774 ^ x17 ;
  assign n21771 = n6163 & n21770 ;
  assign n21776 = n21775 ^ n21771 ;
  assign n21768 = n20437 & n20713 ;
  assign n21777 = n21776 ^ n21768 ;
  assign n21765 = n13433 & n20729 ;
  assign n21763 = n5426 & n20725 ;
  assign n21756 = n20716 ^ x20 ;
  assign n21757 = n21756 ^ x19 ;
  assign n21758 = n21757 ^ n20716 ;
  assign n21759 = n20801 & n21758 ;
  assign n21760 = n21759 ^ n20716 ;
  assign n21761 = n5215 & n21760 ;
  assign n21762 = n21761 ^ x20 ;
  assign n21764 = n21763 ^ n21762 ;
  assign n21766 = n21765 ^ n21764 ;
  assign n21751 = n21748 ^ n21608 ;
  assign n21752 = ~n21651 & n21751 ;
  assign n21731 = ~n4435 & n21316 ;
  assign n21729 = ~n4434 & ~n20739 ;
  assign n21726 = n4600 & ~n20738 ;
  assign n21725 = n20100 & n20603 ;
  assign n21727 = n21726 ^ n21725 ;
  assign n21728 = n21727 ^ x26 ;
  assign n21730 = n21729 ^ n21728 ;
  assign n21732 = n21731 ^ n21730 ;
  assign n21720 = n3985 & n20750 ;
  assign n21719 = n3837 & ~n20747 ;
  assign n21721 = n21720 ^ n21719 ;
  assign n21722 = n21721 ^ n3978 ;
  assign n21712 = n20746 ^ x29 ;
  assign n21711 = n20746 ^ x28 ;
  assign n21713 = n21712 ^ n21711 ;
  assign n21714 = n21712 ^ n21307 ;
  assign n21715 = n21714 ^ n21712 ;
  assign n21716 = n21713 & n21715 ;
  assign n21717 = n21716 ^ n21712 ;
  assign n21718 = n3833 & n21717 ;
  assign n21723 = n21722 ^ n21718 ;
  assign n21707 = ~n21613 & n21625 ;
  assign n21708 = ~n21612 & n21707 ;
  assign n21709 = n21708 ^ n21625 ;
  assign n21703 = n20748 ^ n3518 ;
  assign n21702 = ~n3518 & ~n20748 ;
  assign n21704 = n21703 ^ n21702 ;
  assign n21701 = ~n3801 & n20757 ;
  assign n21705 = n21704 ^ n21701 ;
  assign n21694 = n13480 ^ n1630 ;
  assign n21695 = n21694 ^ n3401 ;
  assign n21692 = n675 ^ n272 ;
  assign n21691 = n1689 ^ n560 ;
  assign n21693 = n21692 ^ n21691 ;
  assign n21696 = n21695 ^ n21693 ;
  assign n21690 = n13366 ^ n4870 ;
  assign n21697 = n21696 ^ n21690 ;
  assign n21688 = n4026 ^ n4003 ;
  assign n21687 = n2604 ^ n2040 ;
  assign n21689 = n21688 ^ n21687 ;
  assign n21698 = n21697 ^ n21689 ;
  assign n21681 = n1925 ^ n256 ;
  assign n21682 = n21681 ^ n150 ;
  assign n21683 = n21682 ^ n1497 ;
  assign n21684 = n21683 ^ n14721 ;
  assign n21678 = n1844 ^ n1822 ;
  assign n21677 = n2316 ^ n711 ;
  assign n21679 = n21678 ^ n21677 ;
  assign n21675 = n13569 ^ n3719 ;
  assign n21676 = n21675 ^ n4230 ;
  assign n21680 = n21679 ^ n21676 ;
  assign n21685 = n21684 ^ n21680 ;
  assign n21671 = n14487 ^ n192 ;
  assign n21672 = n21671 ^ n1360 ;
  assign n21670 = n3746 ^ n354 ;
  assign n21673 = n21672 ^ n21670 ;
  assign n21668 = n4288 ^ n1180 ;
  assign n21667 = n2378 ^ n343 ;
  assign n21669 = n21668 ^ n21667 ;
  assign n21674 = n21673 ^ n21669 ;
  assign n21686 = n21685 ^ n21674 ;
  assign n21699 = n21698 ^ n21686 ;
  assign n21700 = ~n14648 & ~n21699 ;
  assign n21706 = n21705 ^ n21700 ;
  assign n21710 = n21709 ^ n21706 ;
  assign n21724 = n21723 ^ n21710 ;
  assign n21733 = n21732 ^ n21724 ;
  assign n21664 = n21639 ^ n21635 ;
  assign n21665 = ~n21636 & n21664 ;
  assign n21666 = n21665 ^ n21639 ;
  assign n21734 = n21733 ^ n21666 ;
  assign n21661 = n4656 & n21575 ;
  assign n21655 = n21648 ^ n21611 ;
  assign n21656 = n21649 & n21655 ;
  assign n21657 = n21656 ^ n21648 ;
  assign n21658 = n21657 ^ x23 ;
  assign n21654 = n4651 & n20745 ;
  assign n21659 = n21658 ^ n21654 ;
  assign n21653 = n4655 & n20737 ;
  assign n21660 = n21659 ^ n21653 ;
  assign n21662 = n21661 ^ n21660 ;
  assign n21652 = ~n40 & ~n20743 ;
  assign n21663 = n21662 ^ n21652 ;
  assign n21735 = n21734 ^ n21663 ;
  assign n21749 = n21748 ^ n21735 ;
  assign n21753 = n21752 ^ n21749 ;
  assign n21767 = n21766 ^ n21753 ;
  assign n21778 = n21777 ^ n21767 ;
  assign n22103 = n21983 ^ n21778 ;
  assign n22660 = n22494 ^ n22103 ;
  assign n22996 = n22946 ^ n22660 ;
  assign n23300 = n23299 ^ n22996 ;
  assign n23301 = n23300 ^ n22987 ;
  assign n23302 = n23301 ^ n22996 ;
  assign n23303 = ~n22995 & n23302 ;
  assign n23304 = n23303 ^ n23300 ;
  assign n23509 = n23314 ^ n23304 ;
  assign n23510 = n23509 ^ x5 ;
  assign n23504 = n20620 ^ n10329 ;
  assign n23505 = n23504 ^ n20620 ;
  assign n23506 = ~n22963 & n23505 ;
  assign n23507 = n23506 ^ n20620 ;
  assign n23508 = n10322 & ~n23507 ;
  assign n23511 = n23510 ^ n23508 ;
  assign n23500 = n10327 & n20624 ;
  assign n23512 = n23511 ^ n23500 ;
  assign n23514 = n23513 ^ n23512 ;
  assign n24745 = n24742 ^ n23514 ;
  assign n23873 = n23872 ^ n23520 ;
  assign n23874 = ~n23526 & ~n23873 ;
  assign n23875 = n23874 ^ n23872 ;
  assign n24746 = n24745 ^ n23875 ;
  assign n24747 = n24744 & n24746 ;
  assign n24748 = n24747 ^ n24742 ;
  assign n24115 = n24114 ^ n20613 ;
  assign n24118 = ~n20614 & n24115 ;
  assign n24119 = n24118 ^ n20613 ;
  assign n24120 = ~x1 & ~n24119 ;
  assign n24121 = n24120 ^ n24114 ;
  assign n24749 = n24748 ^ n24121 ;
  assign n24122 = n24121 ^ x1 ;
  assign n24123 = n24122 ^ n20612 ;
  assign n24124 = n24123 ^ x2 ;
  assign n24125 = n24124 ^ x1 ;
  assign n24126 = n24125 ^ n24123 ;
  assign n23892 = n21166 ^ n20835 ;
  assign n24127 = n24123 ^ n23892 ;
  assign n24128 = n24127 ^ n24123 ;
  assign n24129 = n24126 & n24128 ;
  assign n24130 = n24129 ^ n24123 ;
  assign n24131 = x0 & n24130 ;
  assign n24750 = n24749 ^ n24131 ;
  assign n22675 = n22674 ^ n22660 ;
  assign n22947 = n22675 & n22946 ;
  assign n22948 = n22947 ^ n22674 ;
  assign n22104 = n22103 ^ n22102 ;
  assign n22495 = n22104 & ~n22494 ;
  assign n22496 = n22495 ^ n22103 ;
  assign n22082 = n6148 & ~n20702 ;
  assign n22081 = n6143 & ~n20705 ;
  assign n22083 = n22082 ^ n22081 ;
  assign n22084 = n22083 ^ x17 ;
  assign n22080 = n6163 & n22079 ;
  assign n22085 = n22084 ^ n22080 ;
  assign n22077 = n20437 & ~n20706 ;
  assign n22086 = n22085 ^ n22077 ;
  assign n22073 = n5426 & n20716 ;
  assign n22071 = n13433 & n20725 ;
  assign n22064 = n20713 ^ x20 ;
  assign n22065 = n22064 ^ x19 ;
  assign n22066 = n22065 ^ n20713 ;
  assign n22067 = n22063 & n22066 ;
  assign n22068 = n22067 ^ n20713 ;
  assign n22069 = n5215 & n22068 ;
  assign n22070 = n22069 ^ x20 ;
  assign n22072 = n22071 ^ n22070 ;
  assign n22074 = n22073 ^ n22072 ;
  assign n22057 = n4655 & n20729 ;
  assign n22056 = n4651 & ~n20743 ;
  assign n22058 = n22057 ^ n22056 ;
  assign n22059 = n22058 ^ x23 ;
  assign n22055 = n4656 & ~n21593 ;
  assign n22060 = n22059 ^ n22055 ;
  assign n22054 = ~n40 & n20737 ;
  assign n22061 = n22060 ^ n22054 ;
  assign n22049 = ~n4435 & ~n21429 ;
  assign n22047 = ~n4434 & n20745 ;
  assign n22044 = n4600 & ~n20739 ;
  assign n22043 = n20603 & ~n20738 ;
  assign n22045 = n22044 ^ n22043 ;
  assign n22046 = n22045 ^ x26 ;
  assign n22048 = n22047 ^ n22046 ;
  assign n22050 = n22049 ^ n22048 ;
  assign n22040 = n3837 & n20750 ;
  assign n22038 = n3985 & n20746 ;
  assign n22033 = ~n21700 & ~n21705 ;
  assign n22026 = n12899 ^ n2281 ;
  assign n22027 = n22026 ^ n4547 ;
  assign n22028 = n22027 ^ n5596 ;
  assign n22029 = n22028 ^ n1484 ;
  assign n22021 = n1160 ^ n464 ;
  assign n22020 = n1066 ^ n157 ;
  assign n22022 = n22021 ^ n22020 ;
  assign n22019 = n1329 ^ n1086 ;
  assign n22023 = n22022 ^ n22019 ;
  assign n22017 = n890 ^ n472 ;
  assign n22016 = n12837 ^ n2828 ;
  assign n22018 = n22017 ^ n22016 ;
  assign n22024 = n22023 ^ n22018 ;
  assign n22025 = n22024 ^ n4510 ;
  assign n22030 = n22029 ^ n22025 ;
  assign n22031 = n22030 ^ n6782 ;
  assign n22032 = ~n14649 & ~n22031 ;
  assign n22034 = n22033 ^ n22032 ;
  assign n22012 = n22543 ^ n20747 ;
  assign n22011 = ~n3518 & n20747 ;
  assign n22013 = n22012 ^ n22011 ;
  assign n22006 = n20748 ^ n5280 ;
  assign n22007 = n22006 ^ n5280 ;
  assign n22008 = n22005 & ~n22007 ;
  assign n22009 = n22008 ^ n5280 ;
  assign n22010 = ~n20757 & n22009 ;
  assign n22014 = n22013 ^ n22010 ;
  assign n22004 = ~n3802 & ~n21702 ;
  assign n22015 = n22014 ^ n22004 ;
  assign n22035 = n22034 ^ n22015 ;
  assign n22036 = n22035 ^ x29 ;
  assign n22001 = n5065 & ~n21380 ;
  assign n22002 = n22001 ^ n20100 ;
  assign n22003 = n3833 & n22002 ;
  assign n22037 = n22036 ^ n22003 ;
  assign n22039 = n22038 ^ n22037 ;
  assign n22041 = n22040 ^ n22039 ;
  assign n21996 = n21723 ^ n21709 ;
  assign n21997 = ~n21710 & n21996 ;
  assign n21998 = n21997 ^ n21723 ;
  assign n22042 = n22041 ^ n21998 ;
  assign n22051 = n22050 ^ n22042 ;
  assign n21993 = n21732 ^ n21666 ;
  assign n21994 = n21733 & n21993 ;
  assign n21995 = n21994 ^ n21732 ;
  assign n22052 = n22051 ^ n21995 ;
  assign n21990 = n21734 ^ n21657 ;
  assign n21991 = ~n21663 & n21990 ;
  assign n21992 = n21991 ^ n21734 ;
  assign n22053 = n22052 ^ n21992 ;
  assign n22062 = n22061 ^ n22053 ;
  assign n22075 = n22074 ^ n22062 ;
  assign n21987 = n21766 ^ n21735 ;
  assign n21988 = ~n21753 & n21987 ;
  assign n21989 = n21988 ^ n21766 ;
  assign n22076 = n22075 ^ n21989 ;
  assign n22087 = n22086 ^ n22076 ;
  assign n21984 = n21983 ^ n21777 ;
  assign n21985 = ~n21778 & n21984 ;
  assign n21986 = n21985 ^ n21983 ;
  assign n22088 = n22087 ^ n21986 ;
  assign n21240 = ~n6529 & ~n20693 ;
  assign n21239 = ~n6547 & ~n20694 ;
  assign n21241 = n21240 ^ n21239 ;
  assign n21242 = n21241 ^ n6537 ;
  assign n21243 = n21242 ^ x14 ;
  assign n21264 = ~n17173 & ~n21244 ;
  assign n21257 = n20690 ^ n6539 ;
  assign n21245 = n21241 ^ n6538 ;
  assign n21247 = n21246 ^ n20690 ;
  assign n21248 = n21247 ^ n20690 ;
  assign n21249 = n21248 ^ n20690 ;
  assign n21250 = n20690 ^ n17173 ;
  assign n21251 = n21250 ^ n20690 ;
  assign n21252 = ~n21249 & ~n21251 ;
  assign n21253 = n21252 ^ n20690 ;
  assign n21254 = ~n21245 & n21253 ;
  assign n21258 = n21257 ^ n21254 ;
  assign n21265 = n21264 ^ n21258 ;
  assign n21266 = ~n21243 & ~n21265 ;
  assign n22089 = n22088 ^ n21266 ;
  assign n22658 = n22496 ^ n22089 ;
  assign n22644 = n7142 & n20680 ;
  assign n22643 = n7148 & ~n20683 ;
  assign n22645 = n22644 ^ n22643 ;
  assign n22646 = n22645 ^ n7149 ;
  assign n22647 = n22646 ^ x11 ;
  assign n22650 = ~x10 & ~n22649 ;
  assign n22654 = n22653 ^ n22650 ;
  assign n22655 = n7150 & ~n22654 ;
  assign n22648 = n22645 ^ x11 ;
  assign n22651 = n22650 ^ n20631 ;
  assign n22652 = n22648 & ~n22651 ;
  assign n22656 = n22655 ^ n22652 ;
  assign n22657 = ~n22647 & ~n22656 ;
  assign n22659 = n22658 ^ n22657 ;
  assign n22984 = n22948 ^ n22659 ;
  assign n23316 = n22996 ^ n22984 ;
  assign n23315 = n23314 ^ n22984 ;
  assign n23317 = n23316 ^ n23315 ;
  assign n23318 = n23304 & n23317 ;
  assign n23319 = n23318 ^ n23316 ;
  assign n22982 = n8139 & ~n20628 ;
  assign n22980 = n8150 & ~n22979 ;
  assign n22975 = n8484 & n20829 ;
  assign n22974 = n8144 & n20819 ;
  assign n22976 = n22975 ^ n22974 ;
  assign n22977 = n22976 ^ x8 ;
  assign n22981 = n22980 ^ n22977 ;
  assign n22983 = n22982 ^ n22981 ;
  assign n23488 = n23319 ^ n22983 ;
  assign n24751 = n24748 ^ n23488 ;
  assign n23494 = n10327 & ~n20620 ;
  assign n23493 = n10425 & ~n20617 ;
  assign n23495 = n23494 ^ n23493 ;
  assign n23496 = n23495 ^ x5 ;
  assign n23491 = n23490 ^ n20617 ;
  assign n23492 = n10342 & n23491 ;
  assign n23497 = n23496 ^ n23492 ;
  assign n23489 = ~n10334 & n20624 ;
  assign n23498 = n23497 ^ n23489 ;
  assign n23515 = n23509 ^ n23498 ;
  assign n23516 = n23515 ^ n23498 ;
  assign n23876 = n23875 ^ n23516 ;
  assign n23877 = n23514 & ~n23876 ;
  assign n23878 = n23877 ^ n23515 ;
  assign n24752 = n24751 ^ n23878 ;
  assign n24753 = n24750 & n24752 ;
  assign n24754 = n24753 ^ n24748 ;
  assign n24756 = n24113 & ~n24754 ;
  assign n24755 = n24754 ^ n24113 ;
  assign n24757 = n24756 ^ n24755 ;
  assign n22985 = n22984 ^ n22983 ;
  assign n23320 = ~n22985 & ~n23319 ;
  assign n23321 = n23320 ^ n22984 ;
  assign n22957 = n8139 & n20829 ;
  assign n22949 = n22948 ^ n22658 ;
  assign n22950 = ~n22659 & n22949 ;
  assign n22951 = n22950 ^ n22658 ;
  assign n22641 = n7142 & n20631 ;
  assign n22638 = n7148 & n20680 ;
  assign n22636 = n7151 & n20819 ;
  assign n22612 = ~n6529 & ~n20690 ;
  assign n22611 = ~n6547 & ~n20693 ;
  assign n22613 = n22612 ^ n22611 ;
  assign n22614 = n22613 ^ n6537 ;
  assign n22615 = n22614 ^ x14 ;
  assign n22628 = x13 & ~n22618 ;
  assign n22627 = n8856 & ~n20683 ;
  assign n22629 = n22628 ^ n22627 ;
  assign n22630 = ~n6539 & n22629 ;
  assign n22625 = n22617 ^ n8856 ;
  assign n22616 = n22613 ^ x14 ;
  assign n22620 = n20683 ^ x13 ;
  assign n22621 = n22620 ^ n20683 ;
  assign n22622 = ~n22617 & ~n22621 ;
  assign n22623 = n22622 ^ n20683 ;
  assign n22624 = ~n22616 & n22623 ;
  assign n22626 = n22625 ^ n22624 ;
  assign n22631 = n22630 ^ n22626 ;
  assign n22632 = ~n22615 & n22631 ;
  assign n22604 = n6148 & ~n20694 ;
  assign n22603 = n6143 & ~n20702 ;
  assign n22605 = n22604 ^ n22603 ;
  assign n22606 = n22605 ^ x17 ;
  assign n22602 = n6163 & n22601 ;
  assign n22607 = n22606 ^ n22602 ;
  assign n22600 = n20437 & ~n20705 ;
  assign n22608 = n22607 ^ n22600 ;
  assign n22596 = n22074 ^ n21989 ;
  assign n22597 = ~n22075 & n22596 ;
  assign n22598 = n22597 ^ n22074 ;
  assign n22593 = n5426 & n20713 ;
  assign n22591 = n5220 & ~n20706 ;
  assign n22588 = n5221 & n21782 ;
  assign n22587 = n13433 & n20716 ;
  assign n22589 = n22588 ^ n22587 ;
  assign n22590 = n22589 ^ x20 ;
  assign n22592 = n22591 ^ n22590 ;
  assign n22594 = n22593 ^ n22592 ;
  assign n22584 = n4651 & n20737 ;
  assign n22582 = ~n40 & n20729 ;
  assign n22575 = n21736 ^ x23 ;
  assign n22576 = n22575 ^ x22 ;
  assign n22577 = n22576 ^ n21736 ;
  assign n22578 = n20800 & ~n22577 ;
  assign n22579 = n22578 ^ n21736 ;
  assign n22580 = n35 & n22579 ;
  assign n22581 = n22580 ^ x23 ;
  assign n22583 = n22582 ^ n22581 ;
  assign n22585 = n22584 ^ n22583 ;
  assign n22570 = ~n4435 & n21440 ;
  assign n22568 = ~n4434 & ~n20743 ;
  assign n22565 = n4600 & n20745 ;
  assign n22564 = n20603 & ~n20739 ;
  assign n22566 = n22565 ^ n22564 ;
  assign n22567 = n22566 ^ x26 ;
  assign n22569 = n22568 ^ n22567 ;
  assign n22571 = n22570 ^ n22569 ;
  assign n22560 = n22035 ^ n21998 ;
  assign n22561 = ~n22041 & ~n22560 ;
  assign n22562 = n22561 ^ n22035 ;
  assign n22557 = n3837 & n20746 ;
  assign n22555 = n3985 & n20100 ;
  assign n22548 = n20738 ^ x29 ;
  assign n22549 = n22548 ^ x28 ;
  assign n22550 = n22549 ^ n20738 ;
  assign n22551 = ~n21328 & n22550 ;
  assign n22552 = n22551 ^ n20738 ;
  assign n22553 = n3833 & ~n22552 ;
  assign n22554 = n22553 ^ x29 ;
  assign n22556 = n22555 ^ n22554 ;
  assign n22558 = n22557 ^ n22556 ;
  assign n22544 = ~n20748 & n22543 ;
  assign n22540 = n20747 ^ x31 ;
  assign n22541 = ~n22011 & ~n22540 ;
  assign n22536 = n20747 ^ n3803 ;
  assign n22535 = ~n61 & ~n20747 ;
  assign n22537 = n22536 ^ n22535 ;
  assign n22538 = n22537 ^ x31 ;
  assign n22530 = n20750 ^ x31 ;
  assign n22531 = n22530 ^ n20750 ;
  assign n22532 = n21275 & n22531 ;
  assign n22533 = n22532 ^ n20750 ;
  assign n22534 = n3518 & n22533 ;
  assign n22539 = n22538 ^ n22534 ;
  assign n22542 = n22541 ^ n22539 ;
  assign n22545 = n22544 ^ n22542 ;
  assign n22520 = n348 ^ n270 ;
  assign n22521 = n22520 ^ n138 ;
  assign n22522 = n22521 ^ n398 ;
  assign n22519 = n842 ^ n124 ;
  assign n22523 = n22522 ^ n22519 ;
  assign n22517 = n1367 ^ n571 ;
  assign n22516 = n4288 ^ n427 ;
  assign n22518 = n22517 ^ n22516 ;
  assign n22524 = n22523 ^ n22518 ;
  assign n22513 = n1084 ^ n684 ;
  assign n22514 = n22513 ^ n2338 ;
  assign n22512 = n5496 ^ n3571 ;
  assign n22515 = n22514 ^ n22512 ;
  assign n22525 = n22524 ^ n22515 ;
  assign n22526 = n22525 ^ n4539 ;
  assign n22527 = n22526 ^ n5649 ;
  assign n22528 = ~n1818 & ~n22527 ;
  assign n22529 = ~n1251 & n22528 ;
  assign n22546 = n22545 ^ n22529 ;
  assign n22509 = n22033 ^ n22015 ;
  assign n22510 = ~n22034 & n22509 ;
  assign n22511 = n22510 ^ n22033 ;
  assign n22547 = n22546 ^ n22511 ;
  assign n22559 = n22558 ^ n22547 ;
  assign n22563 = n22562 ^ n22559 ;
  assign n22572 = n22571 ^ n22563 ;
  assign n22506 = n22050 ^ n21995 ;
  assign n22507 = ~n22051 & n22506 ;
  assign n22508 = n22507 ^ n22050 ;
  assign n22573 = n22572 ^ n22508 ;
  assign n22503 = n22061 ^ n21992 ;
  assign n22504 = n22053 & n22503 ;
  assign n22505 = n22504 ^ n22061 ;
  assign n22574 = n22573 ^ n22505 ;
  assign n22586 = n22585 ^ n22574 ;
  assign n22595 = n22594 ^ n22586 ;
  assign n22599 = n22598 ^ n22595 ;
  assign n22609 = n22608 ^ n22599 ;
  assign n22500 = n22086 ^ n21986 ;
  assign n22501 = ~n22087 & n22500 ;
  assign n22502 = n22501 ^ n22086 ;
  assign n22610 = n22609 ^ n22502 ;
  assign n22633 = n22632 ^ n22610 ;
  assign n22497 = n22496 ^ n22088 ;
  assign n22498 = ~n22089 & ~n22497 ;
  assign n22499 = n22498 ^ n22496 ;
  assign n22634 = n22633 ^ n22499 ;
  assign n22635 = n22634 ^ x11 ;
  assign n22637 = n22636 ^ n22635 ;
  assign n22639 = n22638 ^ n22637 ;
  assign n21238 = n20240 & ~n21237 ;
  assign n22640 = n22639 ^ n21238 ;
  assign n22642 = n22641 ^ n22640 ;
  assign n22952 = n22951 ^ n22642 ;
  assign n22953 = n22952 ^ x8 ;
  assign n21235 = n8484 & n20624 ;
  assign n22954 = n22953 ^ n21235 ;
  assign n21234 = n8144 & ~n20628 ;
  assign n22955 = n22954 ^ n21234 ;
  assign n21233 = n8150 & ~n21232 ;
  assign n22956 = n22955 ^ n21233 ;
  assign n22958 = n22957 ^ n22956 ;
  assign n23486 = n23321 ^ n22958 ;
  assign n23483 = ~n10334 & ~n20620 ;
  assign n23480 = n23479 ^ n20614 ;
  assign n23481 = n10342 & n23480 ;
  assign n23476 = n10425 & ~n20614 ;
  assign n23475 = n10327 & ~n20617 ;
  assign n23477 = n23476 ^ n23475 ;
  assign n23478 = n23477 ^ x5 ;
  assign n23482 = n23481 ^ n23478 ;
  assign n23484 = n23483 ^ n23482 ;
  assign n24767 = n23486 ^ n23484 ;
  assign n23499 = n23498 ^ n23488 ;
  assign n23879 = ~n23499 & n23878 ;
  assign n23880 = n23879 ^ n23498 ;
  assign n24768 = n24767 ^ n23880 ;
  assign n24778 = ~n24757 & ~n24768 ;
  assign n24779 = n23484 & n23880 ;
  assign n23473 = ~n10334 & ~n20617 ;
  assign n23463 = n22610 ^ n22499 ;
  assign n23464 = n22633 & ~n23463 ;
  assign n23465 = n23464 ^ n22610 ;
  assign n23338 = ~x13 & ~n22661 ;
  assign n23339 = n23338 ^ n20680 ;
  assign n23460 = n23339 ^ n22661 ;
  assign n23461 = n6539 & ~n23460 ;
  assign n23453 = n6143 & ~n20694 ;
  assign n23450 = n20437 & ~n20702 ;
  assign n23448 = n16849 & n22091 ;
  assign n23446 = ~n22090 & n23445 ;
  assign n23440 = n5426 & ~n20706 ;
  assign n23438 = n13433 & n20713 ;
  assign n23431 = n20705 ^ x20 ;
  assign n23432 = n23431 ^ x19 ;
  assign n23433 = n23432 ^ n20705 ;
  assign n23434 = ~n21769 & n23433 ;
  assign n23435 = n23434 ^ n20705 ;
  assign n23436 = n5215 & ~n23435 ;
  assign n23437 = n23436 ^ x20 ;
  assign n23439 = n23438 ^ n23437 ;
  assign n23441 = n23440 ^ n23439 ;
  assign n23426 = n4651 & n20729 ;
  assign n23424 = ~n40 & n20725 ;
  assign n23417 = n20716 ^ x23 ;
  assign n23418 = n23417 ^ x22 ;
  assign n23419 = n23418 ^ n20716 ;
  assign n23420 = n20801 & n23419 ;
  assign n23421 = n23420 ^ n20716 ;
  assign n23422 = n35 & n23421 ;
  assign n23423 = n23422 ^ x23 ;
  assign n23425 = n23424 ^ n23423 ;
  assign n23427 = n23426 ^ n23425 ;
  assign n23413 = ~n4435 & n21575 ;
  assign n23411 = ~n4434 & n20737 ;
  assign n23408 = n4600 & ~n20743 ;
  assign n23407 = n20603 & n20745 ;
  assign n23409 = n23408 ^ n23407 ;
  assign n23410 = n23409 ^ x26 ;
  assign n23412 = n23411 ^ n23410 ;
  assign n23414 = n23413 ^ n23412 ;
  assign n23404 = n22571 ^ n22508 ;
  assign n23405 = ~n22572 & n23404 ;
  assign n23406 = n23405 ^ n22571 ;
  assign n23415 = n23414 ^ n23406 ;
  assign n23400 = n3837 & n20100 ;
  assign n23398 = n3985 & ~n20738 ;
  assign n23391 = n20739 ^ x28 ;
  assign n23392 = n23391 ^ x29 ;
  assign n23393 = n23392 ^ n20739 ;
  assign n23394 = ~n20774 & n23393 ;
  assign n23395 = n23394 ^ n20739 ;
  assign n23396 = n3833 & ~n23395 ;
  assign n23397 = n23396 ^ x29 ;
  assign n23399 = n23398 ^ n23397 ;
  assign n23401 = n23400 ^ n23399 ;
  assign n23387 = n22545 ^ n22511 ;
  assign n23388 = n22546 & ~n23387 ;
  assign n23389 = n23388 ^ n22545 ;
  assign n23384 = x31 & n22535 ;
  assign n23381 = n21308 ^ n20750 ;
  assign n23382 = ~n3967 & n23381 ;
  assign n23378 = n20750 ^ n3807 ;
  assign n23377 = ~n61 & n20750 ;
  assign n23379 = n23378 ^ n23377 ;
  assign n23371 = n21307 ^ n3807 ;
  assign n23372 = n23371 ^ n21307 ;
  assign n23373 = n21308 ^ n21307 ;
  assign n23374 = ~n23372 & ~n23373 ;
  assign n23375 = n23374 ^ n21307 ;
  assign n23376 = ~x31 & ~n23375 ;
  assign n23380 = n23379 ^ n23376 ;
  assign n23383 = n23382 ^ n23380 ;
  assign n23385 = n23384 ^ n23383 ;
  assign n23363 = n13622 ^ n778 ;
  assign n23364 = n23363 ^ n479 ;
  assign n23362 = n2331 ^ n721 ;
  assign n23365 = n23364 ^ n23362 ;
  assign n23359 = n3317 ^ n737 ;
  assign n23360 = n23359 ^ n637 ;
  assign n23357 = n905 ^ n845 ;
  assign n23358 = n23357 ^ n610 ;
  assign n23361 = n23360 ^ n23358 ;
  assign n23366 = n23365 ^ n23361 ;
  assign n23356 = n14576 ^ n12496 ;
  assign n23367 = n23366 ^ n23356 ;
  assign n23368 = n23367 ^ n12465 ;
  assign n23369 = n23368 ^ n12700 ;
  assign n23370 = ~n14682 & ~n23369 ;
  assign n23386 = n23385 ^ n23370 ;
  assign n23390 = n23389 ^ n23386 ;
  assign n23402 = n23401 ^ n23390 ;
  assign n23353 = n22562 ^ n22558 ;
  assign n23354 = ~n22559 & ~n23353 ;
  assign n23355 = n23354 ^ n22562 ;
  assign n23403 = n23402 ^ n23355 ;
  assign n23416 = n23415 ^ n23403 ;
  assign n23428 = n23427 ^ n23416 ;
  assign n23350 = n22585 ^ n22505 ;
  assign n23351 = n22574 & n23350 ;
  assign n23352 = n23351 ^ n22585 ;
  assign n23429 = n23428 ^ n23352 ;
  assign n23442 = n23441 ^ n23429 ;
  assign n23347 = n22598 ^ n22594 ;
  assign n23348 = n22595 & n23347 ;
  assign n23349 = n23348 ^ n22598 ;
  assign n23443 = n23442 ^ n23349 ;
  assign n23444 = n23443 ^ x17 ;
  assign n23447 = n23446 ^ n23444 ;
  assign n23449 = n23448 ^ n23447 ;
  assign n23451 = n23450 ^ n23449 ;
  assign n23346 = n6147 & ~n20693 ;
  assign n23452 = n23451 ^ n23346 ;
  assign n23454 = n23453 ^ n23452 ;
  assign n23343 = n22608 ^ n22502 ;
  assign n23344 = ~n22609 & n23343 ;
  assign n23345 = n23344 ^ n22608 ;
  assign n23455 = n23454 ^ n23345 ;
  assign n23456 = n23455 ^ x14 ;
  assign n23342 = ~n6529 & ~n20683 ;
  assign n23457 = n23456 ^ n23342 ;
  assign n23341 = ~n6547 & ~n20690 ;
  assign n23458 = n23457 ^ n23341 ;
  assign n23340 = n6537 & n23339 ;
  assign n23459 = n23458 ^ n23340 ;
  assign n23462 = n23461 ^ n23459 ;
  assign n23466 = n23465 ^ n23462 ;
  assign n23328 = n7151 & ~n20628 ;
  assign n23327 = n7148 & n20631 ;
  assign n23329 = n23328 ^ n23327 ;
  assign n23330 = n23329 ^ x11 ;
  assign n23326 = n20240 & n23307 ;
  assign n23331 = n23330 ^ n23326 ;
  assign n23325 = n7142 & n20819 ;
  assign n23332 = n23331 ^ n23325 ;
  assign n23333 = n23332 ^ n22951 ;
  assign n23334 = n23333 ^ n22634 ;
  assign n23335 = n23334 ^ n23332 ;
  assign n23336 = ~n22642 & n23335 ;
  assign n23337 = n23336 ^ n23333 ;
  assign n23467 = n23466 ^ n23337 ;
  assign n22968 = n22963 ^ n20620 ;
  assign n22964 = ~x7 & ~n22963 ;
  assign n22969 = n22968 ^ n22964 ;
  assign n22970 = n8146 & n22969 ;
  assign n22965 = n22964 ^ n20620 ;
  assign n22966 = n8145 & ~n22965 ;
  assign n22960 = n8139 & n20624 ;
  assign n22959 = n8144 & n20829 ;
  assign n22961 = n22960 ^ n22959 ;
  assign n22962 = n22961 ^ x8 ;
  assign n22967 = n22966 ^ n22962 ;
  assign n22971 = n22970 ^ n22967 ;
  assign n22972 = n22971 ^ n22952 ;
  assign n22973 = n22972 ^ n22971 ;
  assign n23322 = n23321 ^ n22973 ;
  assign n23323 = n22958 & ~n23322 ;
  assign n23324 = n23323 ^ n22972 ;
  assign n23468 = n23467 ^ n23324 ;
  assign n23469 = n23468 ^ x5 ;
  assign n21230 = n10425 & ~n20613 ;
  assign n23470 = n23469 ^ n21230 ;
  assign n21229 = n10327 & ~n20614 ;
  assign n23471 = n23470 ^ n21229 ;
  assign n21227 = n21226 ^ n20613 ;
  assign n21228 = n10342 & n21227 ;
  assign n23472 = n23471 ^ n21228 ;
  assign n23474 = n23473 ^ n23472 ;
  assign n24780 = n24779 ^ n23474 ;
  assign n24781 = n24778 & n24780 ;
  assign n24759 = n23486 ^ n23474 ;
  assign n24761 = n24759 ^ n23484 ;
  assign n24782 = n24761 ^ n23880 ;
  assign n24783 = n24782 ^ n24759 ;
  assign n24784 = n24767 ^ n24759 ;
  assign n24785 = n24784 ^ n24759 ;
  assign n24786 = ~n24783 & ~n24785 ;
  assign n24787 = n24786 ^ n24759 ;
  assign n24788 = n24756 & ~n24787 ;
  assign n24789 = ~n24781 & ~n24788 ;
  assign n24084 = n20908 ^ n20612 ;
  assign n24085 = n24084 ^ n20908 ;
  assign n24086 = n20908 ^ x2 ;
  assign n24089 = n24086 ^ n20908 ;
  assign n24090 = ~n24085 & n24089 ;
  assign n24091 = n24090 ^ n20908 ;
  assign n24092 = ~x1 & n24091 ;
  assign n21168 = ~n20908 & ~n21167 ;
  assign n20909 = ~n20836 & n20908 ;
  assign n24078 = n21168 ^ n20909 ;
  assign n21141 = ~n56 & n3833 ;
  assign n21142 = ~n14140 & n21141 ;
  assign n21136 = n3833 & ~n14140 ;
  assign n21133 = n3835 ^ n3830 ;
  assign n21135 = n12204 & ~n21133 ;
  assign n21137 = n21136 ^ n21135 ;
  assign n21138 = n21137 ^ n3835 ;
  assign n21139 = x29 & n21138 ;
  assign n21134 = n21133 ^ n300 ;
  assign n21140 = n21139 ^ n21134 ;
  assign n21143 = n21142 ^ n21140 ;
  assign n21128 = n3518 & n13052 ;
  assign n21127 = n3807 & ~n13051 ;
  assign n21129 = n21128 ^ n21127 ;
  assign n21125 = n5465 ^ n61 ;
  assign n21126 = n12419 & ~n21125 ;
  assign n21130 = n21129 ^ n21126 ;
  assign n21118 = n3502 ^ n330 ;
  assign n21119 = n21118 ^ n230 ;
  assign n21120 = n21119 ^ n362 ;
  assign n21121 = n21120 ^ n426 ;
  assign n21122 = n21121 ^ n161 ;
  assign n21123 = n21122 ^ n404 ;
  assign n21124 = n21123 ^ n20600 ;
  assign n21131 = n21130 ^ n21124 ;
  assign n21116 = n20877 ^ n20594 ;
  assign n21117 = ~n20878 & ~n21116 ;
  assign n21132 = n21131 ^ n21117 ;
  assign n21144 = n21143 ^ n21132 ;
  assign n21066 = n20580 ^ n20563 ;
  assign n21090 = n21066 ^ n20566 ;
  assign n21058 = n20878 ^ n20566 ;
  assign n21081 = n21058 ^ n20563 ;
  assign n21087 = n21081 ^ n20580 ;
  assign n21088 = n21087 ^ n20552 ;
  assign n21075 = n20881 ^ n20566 ;
  assign n21089 = n21088 ^ n21075 ;
  assign n21091 = n21090 ^ n21089 ;
  assign n21038 = n20881 ^ n20878 ;
  assign n21039 = n21038 ^ n20566 ;
  assign n21040 = n21039 ^ n20580 ;
  assign n21076 = n21075 ^ n21040 ;
  assign n21079 = n21076 ^ n20563 ;
  assign n21080 = n21079 ^ n21040 ;
  assign n21082 = n21081 ^ n21080 ;
  assign n21049 = n21038 ^ n20880 ;
  assign n21050 = n21049 ^ n21038 ;
  assign n21051 = n21050 ^ n20566 ;
  assign n21052 = n21051 ^ n20563 ;
  assign n21053 = n21052 ^ n20566 ;
  assign n21055 = n21053 ^ n21049 ;
  assign n21061 = n21055 ^ n20878 ;
  assign n21062 = n21061 ^ n21058 ;
  assign n21064 = n20878 & n21055 ;
  assign n21067 = n21064 ^ n20878 ;
  assign n21068 = ~n21062 & ~n21067 ;
  assign n21060 = n21081 ^ n21049 ;
  assign n21071 = n21068 ^ n21060 ;
  assign n21065 = n21081 ^ n21064 ;
  assign n21069 = ~n21066 & ~n21068 ;
  assign n21070 = n21065 & n21069 ;
  assign n21072 = n21071 ^ n21070 ;
  assign n21073 = n21072 ^ n21058 ;
  assign n21063 = n21062 ^ n21060 ;
  assign n21074 = n21073 ^ n21063 ;
  assign n21083 = n21082 ^ n21074 ;
  assign n21037 = n20878 ^ n20567 ;
  assign n21084 = n21083 ^ n21037 ;
  assign n21041 = n21040 ^ n21037 ;
  assign n21044 = n21041 ^ n20563 ;
  assign n21045 = n21044 ^ n21040 ;
  assign n21036 = n20879 ^ n20563 ;
  assign n21046 = n21045 ^ n21036 ;
  assign n21085 = n21084 ^ n21046 ;
  assign n21086 = n21085 ^ n20878 ;
  assign n21092 = n21091 ^ n21086 ;
  assign n21093 = n20594 & n21092 ;
  assign n21094 = ~n20594 & n20878 ;
  assign n21095 = n21094 ^ n20563 ;
  assign n21096 = n21095 ^ n21094 ;
  assign n21097 = n21094 ^ n20552 ;
  assign n21098 = n21097 ^ n21094 ;
  assign n21099 = n21096 & n21098 ;
  assign n21100 = n21099 ^ n21094 ;
  assign n21108 = n21098 ^ n21096 ;
  assign n21109 = n21108 ^ n21094 ;
  assign n21102 = n21094 ^ n20580 ;
  assign n21101 = n21094 ^ n20566 ;
  assign n21103 = n21102 ^ n21101 ;
  assign n21104 = n21102 ^ n21097 ;
  assign n21105 = n21104 ^ n21095 ;
  assign n21106 = n21105 ^ n21094 ;
  assign n21107 = n21103 & n21106 ;
  assign n21110 = n21109 ^ n21107 ;
  assign n21111 = n21100 & n21110 ;
  assign n21112 = n21111 ^ n21094 ;
  assign n21115 = ~n21093 & ~n21112 ;
  assign n21145 = n21144 ^ n21115 ;
  assign n21032 = n20886 ^ n20850 ;
  assign n21033 = n20886 ^ n20600 ;
  assign n21034 = ~n21032 & n21033 ;
  assign n21035 = n21034 ^ n20600 ;
  assign n21146 = n21145 ^ n21035 ;
  assign n20910 = ~n20899 & ~n20901 ;
  assign n20915 = n20605 & n20608 ;
  assign n20916 = n20915 ^ n20900 ;
  assign n20911 = n20904 ^ n20887 ;
  assign n20917 = n20916 ^ n20911 ;
  assign n20918 = n20917 ^ n20538 ;
  assign n21016 = n20918 ^ n20916 ;
  assign n21015 = n20916 ^ n20904 ;
  assign n21017 = n21016 ^ n21015 ;
  assign n20919 = n20918 ^ n20911 ;
  assign n21007 = n20919 ^ n20900 ;
  assign n21008 = n21007 ^ n20919 ;
  assign n21009 = n21008 ^ n20911 ;
  assign n21005 = n20919 ^ n20915 ;
  assign n21006 = n21005 ^ n20911 ;
  assign n21010 = n21009 ^ n21006 ;
  assign n20935 = n20900 ^ n20538 ;
  assign n20995 = n20935 ^ n20917 ;
  assign n20912 = n20911 ^ n20900 ;
  assign n20996 = n20995 ^ n20912 ;
  assign n20997 = n20996 ^ n20904 ;
  assign n20999 = n20997 ^ n20995 ;
  assign n20940 = n20915 ^ n20912 ;
  assign n20984 = n20940 ^ n20935 ;
  assign n20985 = n20984 ^ n20912 ;
  assign n20986 = n20985 ^ n20904 ;
  assign n20988 = n20986 ^ n20984 ;
  assign n20936 = n20935 ^ n20911 ;
  assign n20981 = n20940 ^ n20936 ;
  assign n20951 = n20940 ^ n20538 ;
  assign n20952 = n20951 ^ n20911 ;
  assign n20948 = n20940 ^ n20915 ;
  assign n20949 = n20948 ^ n20911 ;
  assign n20960 = n20952 ^ n20949 ;
  assign n20953 = n20952 ^ n20948 ;
  assign n20961 = n20960 ^ n20953 ;
  assign n20941 = n20940 ^ n20911 ;
  assign n20955 = n20953 ^ n20941 ;
  assign n20957 = n20955 ^ n20887 ;
  assign n20962 = n20957 ^ n20941 ;
  assign n20963 = n20962 ^ n20960 ;
  assign n20964 = n20961 & n20963 ;
  assign n20965 = n20964 ^ n20949 ;
  assign n20966 = n20965 ^ n20941 ;
  assign n20959 = n20957 ^ n20955 ;
  assign n20967 = n20966 ^ n20959 ;
  assign n20968 = n20960 ^ n20941 ;
  assign n20969 = n20968 ^ n20959 ;
  assign n20970 = n20967 & ~n20969 ;
  assign n20971 = n20955 ^ n20952 ;
  assign n20972 = n20971 ^ n20957 ;
  assign n20973 = n20955 ^ n20949 ;
  assign n20974 = n20973 ^ n20957 ;
  assign n20975 = ~n20972 & n20974 ;
  assign n20976 = n20970 & n20975 ;
  assign n20977 = n20976 ^ n20964 ;
  assign n20978 = n20977 ^ n20960 ;
  assign n20958 = n20957 ^ n20953 ;
  assign n20979 = n20978 ^ n20958 ;
  assign n20980 = n20979 ^ n20957 ;
  assign n20982 = n20981 ^ n20980 ;
  assign n20989 = n20988 ^ n20982 ;
  assign n20990 = n20989 ^ n20538 ;
  assign n20991 = n20990 ^ n20986 ;
  assign n20937 = n20936 ^ n20917 ;
  assign n20938 = n20937 ^ n20912 ;
  assign n20939 = n20938 ^ n20911 ;
  assign n20943 = n20940 ^ n20939 ;
  assign n20913 = n20912 ^ n20911 ;
  assign n20944 = n20943 ^ n20913 ;
  assign n20946 = n20944 ^ n20887 ;
  assign n20947 = n20946 ^ n20943 ;
  assign n20992 = n20991 ^ n20947 ;
  assign n20993 = n20992 ^ n20946 ;
  assign n20994 = n20993 ^ n20937 ;
  assign n21000 = n20999 ^ n20994 ;
  assign n21001 = n21000 ^ n20997 ;
  assign n20926 = n20917 ^ n20915 ;
  assign n20927 = n20926 ^ n20911 ;
  assign n20934 = n20927 ^ n20919 ;
  assign n21002 = n21001 ^ n20934 ;
  assign n20929 = n20927 ^ n20918 ;
  assign n20930 = n20929 ^ n20916 ;
  assign n20932 = n20930 ^ n20887 ;
  assign n20933 = n20932 ^ n20929 ;
  assign n21003 = n21002 ^ n20933 ;
  assign n21004 = n21003 ^ n20932 ;
  assign n21011 = n21010 ^ n21004 ;
  assign n21018 = n21017 ^ n21011 ;
  assign n21019 = n21018 ^ n21007 ;
  assign n21020 = n21019 ^ n21015 ;
  assign n20920 = n20919 ^ n20912 ;
  assign n20922 = n20920 ^ n20916 ;
  assign n20924 = n20922 ^ n20887 ;
  assign n20925 = n20924 ^ n20920 ;
  assign n21021 = n21020 ^ n20925 ;
  assign n21022 = n21021 ^ n20924 ;
  assign n21023 = n21022 ^ n20937 ;
  assign n21024 = n21023 ^ n20999 ;
  assign n21025 = n21024 ^ n20887 ;
  assign n21026 = n21025 ^ n20997 ;
  assign n21027 = n20915 ^ n20887 ;
  assign n21028 = n21027 ^ n20609 ;
  assign n21029 = n21026 & n21028 ;
  assign n21030 = n20910 & n21029 ;
  assign n21031 = n21030 ^ n21026 ;
  assign n21147 = n21146 ^ n21031 ;
  assign n24079 = n21147 ^ x1 ;
  assign n24080 = n24079 ^ x2 ;
  assign n24081 = n24080 ^ n21147 ;
  assign n24082 = n24078 & n24081 ;
  assign n24083 = n24082 ^ n24079 ;
  assign n24087 = n24086 ^ n24083 ;
  assign n24093 = n24092 ^ n24087 ;
  assign n24094 = ~x0 & n24093 ;
  assign n24095 = n24094 ^ n24083 ;
  assign n24791 = n24789 ^ n24095 ;
  assign n24790 = ~n24095 & n24789 ;
  assign n24792 = n24791 ^ n24790 ;
  assign n24758 = n23484 ^ n23474 ;
  assign n24760 = n24759 ^ n24758 ;
  assign n24762 = ~n23880 & ~n24761 ;
  assign n24763 = n24762 ^ n24759 ;
  assign n24764 = ~n24760 & n24763 ;
  assign n24765 = n24764 ^ n24759 ;
  assign n24766 = n24757 & n24765 ;
  assign n24769 = ~n24756 & n24768 ;
  assign n24773 = ~n23484 & ~n23880 ;
  assign n24774 = n24773 ^ n23474 ;
  assign n24775 = n24769 & n24774 ;
  assign n24776 = ~n24766 & ~n24775 ;
  assign n24777 = ~n24095 & ~n24776 ;
  assign n24793 = n24792 ^ n24777 ;
  assign n24070 = n8484 & ~n20617 ;
  assign n24069 = n8144 & n20624 ;
  assign n24071 = n24070 ^ n24069 ;
  assign n24072 = n24071 ^ x8 ;
  assign n24068 = n8150 & n23491 ;
  assign n24073 = n24072 ^ n24068 ;
  assign n24067 = n8139 & ~n20620 ;
  assign n24074 = n24073 ^ n24067 ;
  assign n24056 = n20437 & ~n20694 ;
  assign n24048 = n23441 ^ n23349 ;
  assign n24049 = ~n23442 & n24048 ;
  assign n24050 = n24049 ^ n23441 ;
  assign n24046 = n13433 & ~n20706 ;
  assign n24044 = n5426 & ~n20705 ;
  assign n23960 = ~n23352 & ~n23427 ;
  assign n23959 = n23427 ^ n23352 ;
  assign n23961 = n23960 ^ n23959 ;
  assign n24036 = n23416 & n23961 ;
  assign n24022 = n23414 ^ n23403 ;
  assign n24014 = ~n23403 & n23414 ;
  assign n24023 = n24022 ^ n24014 ;
  assign n24012 = ~n4435 & ~n21593 ;
  assign n24004 = n23401 ^ n23355 ;
  assign n24005 = n23402 & ~n24004 ;
  assign n24006 = n24005 ^ n23401 ;
  assign n24001 = n3837 & ~n20738 ;
  assign n23999 = n3985 & ~n20739 ;
  assign n23992 = n20745 ^ x29 ;
  assign n23993 = n23992 ^ x28 ;
  assign n23994 = n23993 ^ n20745 ;
  assign n23995 = ~n21428 & n23994 ;
  assign n23996 = n23995 ^ n20745 ;
  assign n23997 = n3833 & n23996 ;
  assign n23998 = n23997 ^ x29 ;
  assign n24000 = n23999 ^ n23998 ;
  assign n24002 = n24001 ^ n24000 ;
  assign n23986 = n23377 ^ n3518 ;
  assign n23985 = n3518 & n21381 ;
  assign n23987 = n23986 ^ n23985 ;
  assign n23988 = x31 & n23987 ;
  assign n23983 = n3807 & n20100 ;
  assign n23982 = ~n3850 & n20746 ;
  assign n23984 = n23983 ^ n23982 ;
  assign n23989 = n23988 ^ n23984 ;
  assign n23975 = n2583 ^ n776 ;
  assign n23976 = n23975 ^ n955 ;
  assign n23973 = n794 ^ n615 ;
  assign n23974 = n23973 ^ n5351 ;
  assign n23977 = n23976 ^ n23974 ;
  assign n23978 = n23977 ^ n4286 ;
  assign n23969 = n13627 ^ n1107 ;
  assign n23968 = n3573 ^ n2025 ;
  assign n23970 = n23969 ^ n23968 ;
  assign n23971 = n23970 ^ n12776 ;
  assign n23972 = n23971 ^ n5313 ;
  assign n23979 = n23978 ^ n23972 ;
  assign n23980 = n23979 ^ n4787 ;
  assign n23981 = ~n12855 & ~n23980 ;
  assign n23990 = n23989 ^ n23981 ;
  assign n23965 = n23389 ^ n23385 ;
  assign n23966 = n23386 & ~n23965 ;
  assign n23967 = n23966 ^ n23389 ;
  assign n23991 = n23990 ^ n23967 ;
  assign n24003 = n24002 ^ n23991 ;
  assign n24007 = n24006 ^ n24003 ;
  assign n24008 = n24007 ^ x26 ;
  assign n23964 = ~n4434 & n20729 ;
  assign n24009 = n24008 ^ n23964 ;
  assign n23963 = n20603 & ~n20743 ;
  assign n24010 = n24009 ^ n23963 ;
  assign n23962 = n4600 & n20737 ;
  assign n24011 = n24010 ^ n23962 ;
  assign n24013 = n24012 ^ n24011 ;
  assign n24025 = n24023 ^ n24013 ;
  assign n24019 = n23406 ^ n23403 ;
  assign n24020 = n23415 & n24019 ;
  assign n24021 = n24020 ^ n23414 ;
  assign n24031 = n24021 ^ n24014 ;
  assign n24015 = n24014 ^ n24013 ;
  assign n24032 = n24015 ^ n24014 ;
  assign n24033 = ~n24031 & ~n24032 ;
  assign n24034 = n24033 ^ n24014 ;
  assign n24035 = n23960 & n24034 ;
  assign n24037 = n24025 & ~n24035 ;
  assign n24038 = n24036 & n24037 ;
  assign n24039 = n24038 ^ n24035 ;
  assign n24016 = ~n23416 & ~n23960 ;
  assign n24017 = n24015 & n24016 ;
  assign n24018 = ~n23961 & ~n24017 ;
  assign n24024 = n24023 ^ n24021 ;
  assign n24026 = n24025 ^ n24023 ;
  assign n24027 = n24024 & ~n24026 ;
  assign n24028 = n24027 ^ n24023 ;
  assign n24029 = n24018 & n24028 ;
  assign n24030 = n24029 ^ n24017 ;
  assign n24040 = n24039 ^ n24030 ;
  assign n23955 = n4656 & n21793 ;
  assign n23954 = ~n40 & n20716 ;
  assign n23956 = n23955 ^ n23954 ;
  assign n23952 = n4655 & n20713 ;
  assign n23951 = n4651 & n20725 ;
  assign n23953 = n23952 ^ n23951 ;
  assign n23957 = n23956 ^ n23953 ;
  assign n23958 = n23957 ^ x23 ;
  assign n24041 = n24040 ^ n23958 ;
  assign n24042 = n24041 ^ x20 ;
  assign n23946 = n20702 ^ n5224 ;
  assign n23947 = n23946 ^ n20702 ;
  assign n23948 = ~n22078 & n23947 ;
  assign n23949 = n23948 ^ n20702 ;
  assign n23950 = n5215 & ~n23949 ;
  assign n24043 = n24042 ^ n23950 ;
  assign n24045 = n24044 ^ n24043 ;
  assign n24047 = n24046 ^ n24045 ;
  assign n24051 = n24050 ^ n24047 ;
  assign n24052 = n24051 ^ x17 ;
  assign n23945 = n6148 & ~n20690 ;
  assign n24053 = n24052 ^ n23945 ;
  assign n23944 = n6143 & ~n20693 ;
  assign n24054 = n24053 ^ n23944 ;
  assign n23943 = n6163 & n21246 ;
  assign n24055 = n24054 ^ n23943 ;
  assign n24057 = n24056 ^ n24055 ;
  assign n23940 = n23443 ^ n23345 ;
  assign n23941 = ~n23454 & ~n23940 ;
  assign n23942 = n23941 ^ n23443 ;
  assign n24058 = n24057 ^ n23942 ;
  assign n23916 = x13 & ~n22649 ;
  assign n23935 = n23916 ^ n22653 ;
  assign n23936 = n6537 & n23935 ;
  assign n23917 = n23916 ^ n20631 ;
  assign n23921 = x13 & ~x14 ;
  assign n23922 = ~n6392 & ~n20683 ;
  assign n23923 = n23921 & n23922 ;
  assign n23924 = n23923 ^ n6392 ;
  assign n23918 = n6390 & n15585 ;
  assign n23919 = ~n20683 & n23918 ;
  assign n23920 = n23919 ^ n6390 ;
  assign n23925 = n23924 ^ n23920 ;
  assign n23928 = n23920 ^ x13 ;
  assign n23929 = ~n20680 & ~n23928 ;
  assign n23930 = n23929 ^ x13 ;
  assign n23931 = ~n23925 & ~n23930 ;
  assign n23932 = n23931 ^ n23924 ;
  assign n23933 = n23932 ^ x14 ;
  assign n23934 = n23917 & n23933 ;
  assign n23937 = n23936 ^ n23934 ;
  assign n23938 = n23932 ^ n6538 ;
  assign n23939 = ~n23937 & ~n23938 ;
  assign n24059 = n24058 ^ n23939 ;
  assign n23913 = n23465 ^ n23455 ;
  assign n23914 = n23462 & n23913 ;
  assign n23915 = n23914 ^ n23465 ;
  assign n24060 = n24059 ^ n23915 ;
  assign n23906 = n7142 & ~n20628 ;
  assign n23904 = n20240 & ~n22979 ;
  assign n23901 = n7151 & n20829 ;
  assign n23900 = n7148 & n20819 ;
  assign n23902 = n23901 ^ n23900 ;
  assign n23903 = n23902 ^ x11 ;
  assign n23905 = n23904 ^ n23903 ;
  assign n23907 = n23906 ^ n23905 ;
  assign n23909 = n23907 ^ n23332 ;
  assign n23908 = n23907 ^ n23466 ;
  assign n23910 = n23909 ^ n23908 ;
  assign n23911 = n23337 & n23910 ;
  assign n23912 = n23911 ^ n23909 ;
  assign n24061 = n24060 ^ n23912 ;
  assign n24063 = n24061 ^ n22971 ;
  assign n24062 = n24061 ^ n23467 ;
  assign n24064 = n24063 ^ n24062 ;
  assign n24065 = n23324 & n24064 ;
  assign n24066 = n24065 ^ n24063 ;
  assign n24075 = n24074 ^ n24066 ;
  assign n23896 = ~n10334 & ~n20614 ;
  assign n23893 = n23892 ^ n20612 ;
  assign n23894 = n10342 & n23893 ;
  assign n23889 = n10425 & ~n20612 ;
  assign n23888 = n10327 & ~n20613 ;
  assign n23890 = n23889 ^ n23888 ;
  assign n23891 = n23890 ^ x5 ;
  assign n23895 = n23894 ^ n23891 ;
  assign n23897 = n23896 ^ n23895 ;
  assign n23898 = n23897 ^ n23468 ;
  assign n23485 = n23484 ^ n23468 ;
  assign n23487 = n23486 ^ n23485 ;
  assign n23881 = n23880 ^ n23487 ;
  assign n23882 = n23881 ^ n23485 ;
  assign n23883 = n23486 ^ n23468 ;
  assign n23884 = n23883 ^ n23485 ;
  assign n23885 = n23882 & ~n23884 ;
  assign n23886 = n23885 ^ n23485 ;
  assign n23887 = n23474 & n23886 ;
  assign n23899 = n23898 ^ n23887 ;
  assign n24076 = n24075 ^ n23899 ;
  assign n21223 = n11139 & ~n20908 ;
  assign n21221 = n21147 ^ x2 ;
  assign n21222 = n11141 & n21221 ;
  assign n21224 = n21223 ^ n21222 ;
  assign n21209 = n21035 ^ n21031 ;
  assign n21171 = ~n21132 & n21143 ;
  assign n21172 = ~n21115 & n21171 ;
  assign n21210 = n21172 ^ n21035 ;
  assign n21211 = n21209 & n21210 ;
  assign n21174 = n21143 ^ n21115 ;
  assign n21175 = n21144 & ~n21174 ;
  assign n21177 = n21175 ^ n21115 ;
  assign n21173 = n21172 ^ n21144 ;
  assign n21176 = n21175 ^ n21173 ;
  assign n21178 = n21177 ^ n21176 ;
  assign n21197 = n3807 & ~n12204 ;
  assign n21196 = ~n3850 & ~n12209 ;
  assign n21198 = n21197 ^ n21196 ;
  assign n21199 = n21198 ^ x31 ;
  assign n21194 = x31 & ~n12422 ;
  assign n21195 = ~n20872 & n21194 ;
  assign n21200 = n21199 ^ n21195 ;
  assign n21191 = n21119 ^ n361 ;
  assign n21192 = n21191 ^ n220 ;
  assign n21188 = n20600 ^ n20594 ;
  assign n21189 = n21124 & n21188 ;
  assign n21190 = n21189 ^ n20600 ;
  assign n21193 = n21192 ^ n21190 ;
  assign n21201 = n21200 ^ n21193 ;
  assign n21180 = n21124 ^ n21117 ;
  assign n21181 = n21133 ^ n3836 ;
  assign n21182 = n21181 ^ n21130 ;
  assign n21183 = n21182 ^ n20594 ;
  assign n21184 = n21183 ^ n21117 ;
  assign n21185 = n21184 ^ n21181 ;
  assign n21186 = n21180 & n21185 ;
  assign n21187 = n21186 ^ n21182 ;
  assign n21202 = n21201 ^ n21187 ;
  assign n21179 = n21177 ^ n21031 ;
  assign n21203 = n21202 ^ n21179 ;
  assign n21204 = n21203 ^ n21176 ;
  assign n21205 = n21204 ^ n21202 ;
  assign n21206 = n21205 ^ n21035 ;
  assign n21207 = ~n21178 & n21206 ;
  assign n21208 = n21207 ^ n21203 ;
  assign n21212 = n21211 ^ n21208 ;
  assign n21213 = n21212 ^ x2 ;
  assign n21169 = n21147 & ~n21168 ;
  assign n21148 = ~n20909 & ~n21147 ;
  assign n21170 = n21169 ^ n21148 ;
  assign n21214 = n21213 ^ n21170 ;
  assign n21215 = n21214 ^ n21213 ;
  assign n21216 = n21213 ^ n11012 ;
  assign n21217 = n21216 ^ n21213 ;
  assign n21218 = ~n21215 & n21217 ;
  assign n21219 = n21218 ^ n21213 ;
  assign n21220 = x0 & ~n21219 ;
  assign n21225 = n21224 ^ n21220 ;
  assign n24077 = n24076 ^ n21225 ;
  assign n24794 = n24793 ^ n24077 ;
  assign n25056 = n24096 ^ n20908 ;
  assign n25052 = ~x4 & ~n24096 ;
  assign n25057 = n25056 ^ n25052 ;
  assign n25058 = n18778 & ~n25057 ;
  assign n25053 = n25052 ^ n20908 ;
  assign n25054 = n25051 & n25053 ;
  assign n25049 = n10327 & ~n20612 ;
  assign n25047 = ~n10334 & ~n20613 ;
  assign n25043 = n8139 & ~n20617 ;
  assign n25041 = n8150 & n23480 ;
  assign n25038 = n8484 & ~n20614 ;
  assign n25037 = n8144 & ~n20620 ;
  assign n25039 = n25038 ^ n25037 ;
  assign n25040 = n25039 ^ x8 ;
  assign n25042 = n25041 ^ n25040 ;
  assign n25044 = n25043 ^ n25042 ;
  assign n25019 = n7142 & n20829 ;
  assign n25018 = n7148 & ~n20628 ;
  assign n25020 = n25019 ^ n25018 ;
  assign n25021 = n25020 ^ n7149 ;
  assign n25022 = n25021 ^ x11 ;
  assign n25024 = ~x10 & ~n21231 ;
  assign n25027 = n25024 ^ n21232 ;
  assign n25028 = n7150 & ~n25027 ;
  assign n25023 = n25020 ^ x11 ;
  assign n25025 = n25024 ^ n20624 ;
  assign n25026 = n25023 & ~n25025 ;
  assign n25029 = n25028 ^ n25026 ;
  assign n25030 = ~n25022 & ~n25029 ;
  assign n25009 = n24058 ^ n23915 ;
  assign n25010 = ~n24059 & ~n25009 ;
  assign n25011 = n25010 ^ n24058 ;
  assign n24859 = ~n6529 & n20631 ;
  assign n24858 = ~n6547 & n20680 ;
  assign n24860 = n24859 ^ n24858 ;
  assign n24999 = n20437 & ~n20693 ;
  assign n24996 = n6143 & ~n20690 ;
  assign n24994 = n6148 & ~n20683 ;
  assign n24990 = n13433 & ~n20705 ;
  assign n24988 = n5426 & ~n20702 ;
  assign n24982 = ~n23957 & ~n24030 ;
  assign n24971 = n24021 ^ n24007 ;
  assign n24972 = n24013 & n24971 ;
  assign n24973 = n24972 ^ n24007 ;
  assign n24968 = n3837 & ~n20739 ;
  assign n24966 = n3985 & n20745 ;
  assign n24959 = n20743 ^ x29 ;
  assign n24960 = n24959 ^ x28 ;
  assign n24961 = n24960 ^ n20743 ;
  assign n24962 = ~n21439 & n24961 ;
  assign n24963 = n24962 ^ n20743 ;
  assign n24964 = n3833 & ~n24963 ;
  assign n24965 = n24964 ^ x29 ;
  assign n24967 = n24966 ^ n24965 ;
  assign n24969 = n24968 ^ n24967 ;
  assign n24933 = ~n61 & n20100 ;
  assign n24932 = n3849 ^ x31 ;
  assign n24934 = n24933 ^ n24932 ;
  assign n24943 = n24934 ^ x31 ;
  assign n24944 = n24943 ^ n20738 ;
  assign n24945 = n24944 ^ n24934 ;
  assign n24946 = n24945 ^ n20738 ;
  assign n24947 = ~n20771 & n24946 ;
  assign n24948 = n24947 ^ n20738 ;
  assign n24949 = n3518 & ~n24948 ;
  assign n24950 = n24949 ^ n24943 ;
  assign n24935 = n24934 ^ n24933 ;
  assign n24936 = n24933 ^ n20746 ;
  assign n24937 = n24936 ^ n24933 ;
  assign n24938 = ~n24935 & n24937 ;
  assign n24939 = n24938 ^ n24933 ;
  assign n24940 = n12812 & ~n24939 ;
  assign n24951 = n24950 ^ n24940 ;
  assign n24928 = n23985 ^ n3801 ;
  assign n24929 = ~n12812 & ~n24928 ;
  assign n24930 = n24929 ^ n3801 ;
  assign n24931 = ~n20100 & ~n24930 ;
  assign n24952 = n24951 ^ n24931 ;
  assign n24910 = n13666 ^ n924 ;
  assign n24920 = n4159 ^ n2025 ;
  assign n24921 = n24920 ^ n1204 ;
  assign n24919 = n2304 ^ n1067 ;
  assign n24922 = n24921 ^ n24919 ;
  assign n24923 = n24922 ^ n6802 ;
  assign n24915 = n5301 ^ n277 ;
  assign n24914 = n385 ^ n188 ;
  assign n24916 = n24915 ^ n24914 ;
  assign n24912 = n2145 ^ n1616 ;
  assign n24911 = n13619 ^ n2267 ;
  assign n24913 = n24912 ^ n24911 ;
  assign n24917 = n24916 ^ n24913 ;
  assign n24918 = n24917 ^ n6933 ;
  assign n24924 = n24923 ^ n24918 ;
  assign n24925 = n24924 ^ n3246 ;
  assign n24926 = ~n24910 & ~n24925 ;
  assign n24907 = n23981 ^ n23967 ;
  assign n24908 = ~n23990 & ~n24907 ;
  assign n24909 = n24908 ^ n23989 ;
  assign n24927 = n24926 ^ n24909 ;
  assign n24953 = n24952 ^ n24927 ;
  assign n24954 = n24953 ^ n24006 ;
  assign n24955 = n24954 ^ n24002 ;
  assign n24956 = n24955 ^ n24953 ;
  assign n24957 = ~n24003 & n24956 ;
  assign n24958 = n24957 ^ n24954 ;
  assign n24970 = n24969 ^ n24958 ;
  assign n24974 = n24973 ^ n24970 ;
  assign n24892 = n4600 & n20729 ;
  assign n24891 = n20603 & n20737 ;
  assign n24893 = n24892 ^ n24891 ;
  assign n24894 = n24893 ^ x26 ;
  assign n24896 = n24894 ^ n20725 ;
  assign n24897 = n24896 ^ n13110 ;
  assign n24898 = n24897 ^ n24896 ;
  assign n24899 = n24896 ^ n20800 ;
  assign n24900 = n24899 ^ n24896 ;
  assign n24901 = ~n24898 & n24900 ;
  assign n24902 = n24901 ^ n24896 ;
  assign n24903 = ~n24893 & n24902 ;
  assign n24904 = n24903 ^ x26 ;
  assign n24905 = n96 & n24904 ;
  assign n24906 = n24905 ^ n24894 ;
  assign n24975 = n24974 ^ n24906 ;
  assign n24889 = n4656 & n21782 ;
  assign n24888 = ~n40 & n20713 ;
  assign n24890 = n24889 ^ n24888 ;
  assign n24976 = n24975 ^ n24890 ;
  assign n24887 = n4651 & n20716 ;
  assign n24977 = n24976 ^ n24887 ;
  assign n24886 = n4655 & ~n20706 ;
  assign n24978 = n24977 ^ n24886 ;
  assign n24885 = n24039 ^ x23 ;
  assign n24979 = n24978 ^ n24885 ;
  assign n24980 = n24979 ^ n24030 ;
  assign n24981 = n24980 ^ n24978 ;
  assign n24983 = n24982 ^ n24981 ;
  assign n24984 = ~n24040 & n24983 ;
  assign n24985 = n24984 ^ n24979 ;
  assign n24986 = n24985 ^ x20 ;
  assign n24880 = n20694 ^ n5224 ;
  assign n24881 = n24880 ^ n20694 ;
  assign n24882 = ~n22112 & n24881 ;
  assign n24883 = n24882 ^ n20694 ;
  assign n24884 = n5215 & ~n24883 ;
  assign n24987 = n24986 ^ n24884 ;
  assign n24989 = n24988 ^ n24987 ;
  assign n24991 = n24990 ^ n24989 ;
  assign n24877 = n24050 ^ n24041 ;
  assign n24878 = n24047 & ~n24877 ;
  assign n24879 = n24878 ^ n24050 ;
  assign n24992 = n24991 ^ n24879 ;
  assign n24993 = n24992 ^ x17 ;
  assign n24995 = n24994 ^ n24993 ;
  assign n24997 = n24996 ^ n24995 ;
  assign n24876 = n6163 & n22618 ;
  assign n24998 = n24997 ^ n24876 ;
  assign n25000 = n24999 ^ n24998 ;
  assign n24873 = n24051 ^ n23942 ;
  assign n24874 = ~n24057 & n24873 ;
  assign n24875 = n24874 ^ n24051 ;
  assign n25001 = n25000 ^ n24875 ;
  assign n25002 = n25001 ^ x14 ;
  assign n24861 = n21237 ^ x13 ;
  assign n24862 = n24861 ^ n21237 ;
  assign n24866 = ~n21236 & ~n24862 ;
  assign n24867 = n24866 ^ n21237 ;
  assign n24868 = n6539 & ~n24867 ;
  assign n25003 = n25002 ^ n24868 ;
  assign n25004 = n25003 ^ n25001 ;
  assign n24869 = ~n21236 & n24862 ;
  assign n24870 = n24869 ^ n21237 ;
  assign n24871 = n6537 & n24870 ;
  assign n24872 = n24871 ^ n15618 ;
  assign n25005 = n25004 ^ n24872 ;
  assign n25006 = n25005 ^ n24868 ;
  assign n25007 = ~n24860 & ~n25006 ;
  assign n25008 = n25007 ^ n25003 ;
  assign n25012 = n25011 ^ n25008 ;
  assign n25014 = n25012 ^ n23907 ;
  assign n25013 = n25012 ^ n24060 ;
  assign n25015 = n25014 ^ n25013 ;
  assign n25016 = n23912 & n25015 ;
  assign n25017 = n25016 ^ n25014 ;
  assign n25031 = n25030 ^ n25017 ;
  assign n25033 = n25031 ^ n24061 ;
  assign n25032 = n25031 ^ n24074 ;
  assign n25034 = n25033 ^ n25032 ;
  assign n25035 = n24066 & n25034 ;
  assign n25036 = n25035 ^ n25033 ;
  assign n25045 = n25044 ^ n25036 ;
  assign n25046 = n25045 ^ x5 ;
  assign n25048 = n25047 ^ n25046 ;
  assign n25050 = n25049 ^ n25048 ;
  assign n25055 = n25054 ^ n25050 ;
  assign n25059 = n25058 ^ n25055 ;
  assign n24855 = n24075 ^ n23897 ;
  assign n24856 = ~n23899 & n24855 ;
  assign n24857 = n24856 ^ n24075 ;
  assign n25060 = n25059 ^ n24857 ;
  assign n24809 = ~n21169 & n21212 ;
  assign n24808 = ~n21148 & ~n21212 ;
  assign n24810 = n24809 ^ n24808 ;
  assign n24833 = n12209 & n22543 ;
  assign n24834 = n24833 ^ n52 ;
  assign n24835 = x31 & ~n15160 ;
  assign n24836 = ~n24834 & n24835 ;
  assign n24837 = n24836 ^ n24834 ;
  assign n24838 = n24837 ^ n21181 ;
  assign n24830 = n21201 ^ n21181 ;
  assign n24831 = n21187 & n24830 ;
  assign n24832 = n24831 ^ n21181 ;
  assign n24839 = n24838 ^ n24832 ;
  assign n24825 = n21200 ^ n21190 ;
  assign n24823 = n21190 & ~n21200 ;
  assign n24826 = n24825 ^ n24823 ;
  assign n24827 = n21192 & n24826 ;
  assign n24824 = ~n21192 & n24823 ;
  assign n24828 = n24827 ^ n24824 ;
  assign n24822 = n364 ^ n304 ;
  assign n24829 = n24828 ^ n24822 ;
  assign n24840 = n24839 ^ n24829 ;
  assign n24811 = ~n21176 & n21202 ;
  assign n24812 = n21031 & n21035 ;
  assign n24813 = n21209 ^ n21202 ;
  assign n24814 = n24813 ^ n24812 ;
  assign n24815 = n21177 & n24814 ;
  assign n24816 = ~n24812 & ~n24815 ;
  assign n24817 = ~n21172 & n24816 ;
  assign n24820 = n24811 & n24817 ;
  assign n24818 = n24817 ^ n24815 ;
  assign n24821 = n24820 ^ n24818 ;
  assign n24841 = n24840 ^ n24821 ;
  assign n24842 = n24841 ^ x1 ;
  assign n24843 = n24842 ^ x2 ;
  assign n24844 = n24843 ^ n24841 ;
  assign n24845 = n24810 & n24844 ;
  assign n24846 = n24845 ^ n24842 ;
  assign n25061 = n25060 ^ n24846 ;
  assign n24806 = n21212 ^ n21147 ;
  assign n24807 = n24806 ^ n21212 ;
  assign n24847 = n24846 ^ n21213 ;
  assign n24848 = n24847 ^ n24846 ;
  assign n24849 = n24848 ^ n21212 ;
  assign n24850 = n24807 & n24849 ;
  assign n24851 = n24850 ^ n21212 ;
  assign n24852 = ~x1 & ~n24851 ;
  assign n24853 = n24852 ^ n24847 ;
  assign n24854 = ~x0 & ~n24853 ;
  assign n25062 = n25061 ^ n24854 ;
  assign n24795 = n24790 ^ n24776 ;
  assign n24796 = n24795 ^ n24777 ;
  assign n24803 = n24796 ^ n21225 ;
  assign n24804 = n24077 & ~n24803 ;
  assign n24805 = n24804 ^ n24076 ;
  assign n25063 = n25062 ^ n24805 ;
  assign n24797 = n24796 ^ n24792 ;
  assign n24798 = n24792 ^ n24077 ;
  assign n24799 = n24798 ^ n24792 ;
  assign n24800 = ~n24797 & n24799 ;
  assign n24801 = n24800 ^ n24792 ;
  assign n24802 = ~n24777 & n24801 ;
  assign n25064 = n25063 ^ n24802 ;
  assign n25283 = n24841 ^ n21212 ;
  assign n25284 = n25283 ^ n24841 ;
  assign n25285 = n24841 ^ x2 ;
  assign n25286 = n25285 ^ n24841 ;
  assign n25287 = ~n25284 & n25286 ;
  assign n25288 = n25287 ^ n24841 ;
  assign n25289 = ~x1 & n25288 ;
  assign n25290 = n25289 ^ n25285 ;
  assign n25291 = n25290 ^ x1 ;
  assign n25281 = n24827 & n24829 ;
  assign n25264 = n24832 ^ n24821 ;
  assign n25265 = n25264 ^ n24837 ;
  assign n25267 = ~n24832 & n24837 ;
  assign n25266 = n24839 ^ n21181 ;
  assign n25268 = n25267 ^ n25266 ;
  assign n25269 = n25265 & ~n25268 ;
  assign n25275 = n25269 ^ n25265 ;
  assign n25276 = n24829 ^ n21181 ;
  assign n25277 = n25265 ^ n24829 ;
  assign n25278 = n25276 & ~n25277 ;
  assign n25279 = ~n25275 & n25278 ;
  assign n25272 = n24821 & n25267 ;
  assign n25263 = n24829 ^ n3799 ;
  assign n25270 = n25269 ^ n25263 ;
  assign n25261 = n367 & n24823 ;
  assign n25271 = n25270 ^ n25261 ;
  assign n25273 = n25272 ^ n25271 ;
  assign n25259 = n24822 ^ n367 ;
  assign n25260 = ~n24824 & n25259 ;
  assign n25274 = n25273 ^ n25260 ;
  assign n25280 = n25279 ^ n25274 ;
  assign n25282 = n25281 ^ n25280 ;
  assign n25292 = n25291 ^ n25282 ;
  assign n25293 = n25292 ^ x1 ;
  assign n25294 = n25293 ^ x2 ;
  assign n25295 = n25294 ^ n25292 ;
  assign n25297 = ~n24808 & ~n24841 ;
  assign n25298 = n25297 ^ n24841 ;
  assign n25296 = n24809 & n24841 ;
  assign n25299 = n25298 ^ n25296 ;
  assign n25302 = n25295 & n25299 ;
  assign n25303 = n25302 ^ n25292 ;
  assign n25304 = x0 & ~n25303 ;
  assign n25305 = n25304 ^ n25290 ;
  assign n25255 = n25060 ^ n24805 ;
  assign n25256 = ~n25062 & ~n25255 ;
  assign n25257 = n25256 ^ n25060 ;
  assign n25250 = n25044 ^ n25031 ;
  assign n25251 = ~n25036 & ~n25250 ;
  assign n25252 = n25251 ^ n25031 ;
  assign n25248 = n8139 & ~n20614 ;
  assign n25225 = ~n6529 & n20819 ;
  assign n25224 = ~n6547 & n20631 ;
  assign n25226 = n25225 ^ n25224 ;
  assign n25227 = n25226 ^ n6537 ;
  assign n25228 = n25227 ^ x14 ;
  assign n25238 = n6539 & n23306 ;
  assign n25229 = n25226 ^ n6538 ;
  assign n25230 = n23307 ^ n20628 ;
  assign n25233 = n20628 ^ x13 ;
  assign n25234 = n25233 ^ n20628 ;
  assign n25235 = ~n25230 & ~n25234 ;
  assign n25236 = n25235 ^ n20628 ;
  assign n25237 = n25229 & n25236 ;
  assign n25239 = n25238 ^ n25237 ;
  assign n25240 = ~n25228 & ~n25239 ;
  assign n25220 = n24992 ^ n24875 ;
  assign n25221 = n25000 & ~n25220 ;
  assign n25222 = n25221 ^ n24992 ;
  assign n25218 = n20437 & ~n20690 ;
  assign n25215 = n6143 & ~n20683 ;
  assign n25213 = n6148 & n20680 ;
  assign n25209 = n13433 & ~n20702 ;
  assign n25207 = n5426 & ~n20694 ;
  assign n25197 = n24978 ^ n23957 ;
  assign n25198 = ~n24030 & ~n24039 ;
  assign n25199 = ~n25197 & n25198 ;
  assign n25192 = n24975 ^ n24039 ;
  assign n25200 = n25199 ^ n25192 ;
  assign n25201 = x23 & n25200 ;
  assign n25202 = n25201 ^ n24975 ;
  assign n25193 = n25192 ^ n24975 ;
  assign n25194 = ~n24982 & ~n25193 ;
  assign n25195 = n25194 ^ n24975 ;
  assign n25196 = ~n24978 & ~n25195 ;
  assign n25203 = n25202 ^ n25196 ;
  assign n25188 = ~n40 & ~n20706 ;
  assign n25167 = n4600 & n20725 ;
  assign n25166 = n20603 & n20729 ;
  assign n25168 = n25167 ^ n25166 ;
  assign n25169 = n25168 ^ n97 ;
  assign n25179 = ~n13110 & ~n20801 ;
  assign n25170 = n25168 ^ n99 ;
  assign n25171 = n25170 ^ x26 ;
  assign n25172 = n20716 ^ x25 ;
  assign n25173 = ~n99 & n25172 ;
  assign n25174 = n25173 ^ n20716 ;
  assign n25175 = n20801 & ~n25174 ;
  assign n25176 = n25175 ^ n20716 ;
  assign n25177 = ~n25171 & ~n25176 ;
  assign n25178 = n25177 ^ n25172 ;
  assign n25180 = n25179 ^ n25178 ;
  assign n25181 = ~n25169 & ~n25180 ;
  assign n25162 = n3985 & ~n20743 ;
  assign n25157 = n24969 ^ n24953 ;
  assign n25158 = ~n24958 & ~n25157 ;
  assign n25159 = n25158 ^ n24953 ;
  assign n25160 = n25159 ^ x29 ;
  assign n25152 = n21575 ^ n5065 ;
  assign n25153 = n25152 ^ n21575 ;
  assign n25154 = n21574 & ~n25153 ;
  assign n25155 = n25154 ^ n21575 ;
  assign n25156 = n3833 & n25155 ;
  assign n25161 = n25160 ^ n25156 ;
  assign n25163 = n25162 ^ n25161 ;
  assign n25151 = n3837 & n20745 ;
  assign n25164 = n25163 ^ n25151 ;
  assign n25147 = n24952 ^ n24909 ;
  assign n25148 = n24927 & n25147 ;
  assign n25149 = n25148 ^ n24952 ;
  assign n25143 = ~n3850 & ~n20738 ;
  assign n25142 = x31 & n24933 ;
  assign n25144 = n25143 ^ n25142 ;
  assign n25139 = x31 & ~n20774 ;
  assign n25140 = n25139 ^ n20739 ;
  assign n25141 = n3518 & ~n25140 ;
  assign n25145 = n25144 ^ n25141 ;
  assign n25130 = n12876 ^ n2496 ;
  assign n25127 = n14293 ^ n2569 ;
  assign n25128 = n25127 ^ n1136 ;
  assign n25125 = n1233 ^ n479 ;
  assign n25124 = n4103 ^ n839 ;
  assign n25126 = n25125 ^ n25124 ;
  assign n25129 = n25128 ^ n25126 ;
  assign n25131 = n25130 ^ n25129 ;
  assign n25120 = n1308 ^ n250 ;
  assign n25121 = n25120 ^ n753 ;
  assign n25118 = n3296 ^ n357 ;
  assign n25119 = n25118 ^ n1554 ;
  assign n25122 = n25121 ^ n25119 ;
  assign n25123 = n25122 ^ n4269 ;
  assign n25132 = n25131 ^ n25123 ;
  assign n25133 = n25132 ^ n4251 ;
  assign n25134 = ~n2659 & ~n25133 ;
  assign n25146 = n25145 ^ n25134 ;
  assign n25150 = n25149 ^ n25146 ;
  assign n25165 = n25164 ^ n25150 ;
  assign n25182 = n25181 ^ n25165 ;
  assign n25115 = n24973 ^ n24906 ;
  assign n25116 = ~n24974 & n25115 ;
  assign n25117 = n25116 ^ n24973 ;
  assign n25183 = n25182 ^ n25117 ;
  assign n25184 = n25183 ^ x23 ;
  assign n25114 = n4655 & ~n20705 ;
  assign n25185 = n25184 ^ n25114 ;
  assign n25113 = n4651 & n20713 ;
  assign n25186 = n25185 ^ n25113 ;
  assign n25112 = n4656 & n21770 ;
  assign n25187 = n25186 ^ n25112 ;
  assign n25189 = n25188 ^ n25187 ;
  assign n25204 = n25203 ^ n25189 ;
  assign n25205 = n25204 ^ x20 ;
  assign n25107 = n20693 ^ n5224 ;
  assign n25108 = n25107 ^ n20693 ;
  assign n25109 = ~n22092 & n25108 ;
  assign n25110 = n25109 ^ n20693 ;
  assign n25111 = n5215 & ~n25110 ;
  assign n25206 = n25205 ^ n25111 ;
  assign n25208 = n25207 ^ n25206 ;
  assign n25210 = n25209 ^ n25208 ;
  assign n25104 = n24985 ^ n24879 ;
  assign n25105 = ~n24991 & n25104 ;
  assign n25106 = n25105 ^ n24879 ;
  assign n25211 = n25210 ^ n25106 ;
  assign n25212 = n25211 ^ x17 ;
  assign n25214 = n25213 ^ n25212 ;
  assign n25216 = n25215 ^ n25214 ;
  assign n25103 = n6163 & ~n22662 ;
  assign n25217 = n25216 ^ n25103 ;
  assign n25219 = n25218 ^ n25217 ;
  assign n25223 = n25222 ^ n25219 ;
  assign n25241 = n25240 ^ n25223 ;
  assign n25100 = n25011 ^ n25001 ;
  assign n25101 = ~n25008 & ~n25100 ;
  assign n25102 = n25101 ^ n25011 ;
  assign n25242 = n25241 ^ n25102 ;
  assign n25093 = n7142 & n20624 ;
  assign n25091 = n20240 & n22968 ;
  assign n25088 = n7151 & ~n20620 ;
  assign n25087 = n7148 & n20829 ;
  assign n25089 = n25088 ^ n25087 ;
  assign n25090 = n25089 ^ x11 ;
  assign n25092 = n25091 ^ n25090 ;
  assign n25094 = n25093 ^ n25092 ;
  assign n25096 = n25094 ^ n25012 ;
  assign n25095 = n25094 ^ n25030 ;
  assign n25097 = n25096 ^ n25095 ;
  assign n25098 = n25017 & ~n25097 ;
  assign n25099 = n25098 ^ n25096 ;
  assign n25243 = n25242 ^ n25099 ;
  assign n25244 = n25243 ^ x8 ;
  assign n25086 = n8484 & ~n20613 ;
  assign n25245 = n25244 ^ n25086 ;
  assign n25085 = n8144 & ~n20617 ;
  assign n25246 = n25245 ^ n25085 ;
  assign n25084 = n8150 & n21227 ;
  assign n25247 = n25246 ^ n25084 ;
  assign n25249 = n25248 ^ n25247 ;
  assign n25253 = n25252 ^ n25249 ;
  assign n25073 = n24078 ^ n21147 ;
  assign n25070 = ~x4 & ~n24078 ;
  assign n25074 = n25073 ^ n25070 ;
  assign n25075 = n18778 & ~n25074 ;
  assign n25067 = n10327 & n20908 ;
  assign n25066 = ~n10334 & ~n20612 ;
  assign n25068 = n25067 ^ n25066 ;
  assign n25069 = n25068 ^ x5 ;
  assign n25071 = n25070 ^ n21147 ;
  assign n25072 = n25069 & ~n25071 ;
  assign n25076 = n25075 ^ n25072 ;
  assign n25077 = n25068 ^ n10340 ;
  assign n25078 = ~n25076 & ~n25077 ;
  assign n25079 = n25078 ^ n25045 ;
  assign n25080 = n25079 ^ n25078 ;
  assign n25081 = n25080 ^ n24857 ;
  assign n25082 = ~n25059 & ~n25081 ;
  assign n25083 = n25082 ^ n25079 ;
  assign n25254 = n25253 ^ n25083 ;
  assign n25258 = n25257 ^ n25254 ;
  assign n25306 = n25305 ^ n25258 ;
  assign n25065 = n24802 & ~n25063 ;
  assign n25307 = n25306 ^ n25065 ;
  assign n25502 = ~n10334 & n20908 ;
  assign n25491 = n7151 & ~n20617 ;
  assign n25490 = n7148 & n20624 ;
  assign n25492 = n25491 ^ n25490 ;
  assign n25493 = n25492 ^ x11 ;
  assign n25489 = n20240 & n23491 ;
  assign n25494 = n25493 ^ n25489 ;
  assign n25488 = n7142 & ~n20620 ;
  assign n25495 = n25494 ^ n25488 ;
  assign n25479 = n25223 ^ n25102 ;
  assign n25480 = ~n25241 & n25479 ;
  assign n25481 = n25480 ^ n25223 ;
  assign n25472 = n20437 & ~n20683 ;
  assign n25465 = n13433 & ~n20694 ;
  assign n25463 = n5426 & ~n20693 ;
  assign n25458 = ~n40 & ~n20705 ;
  assign n25389 = n20603 & n20725 ;
  assign n25388 = n4600 & n20716 ;
  assign n25390 = n25389 ^ n25388 ;
  assign n25450 = n25390 ^ x26 ;
  assign n25447 = n3837 & ~n20743 ;
  assign n25445 = n3985 & n20737 ;
  assign n25438 = n20729 ^ x29 ;
  assign n25439 = n25438 ^ x28 ;
  assign n25440 = n25439 ^ n20729 ;
  assign n25441 = ~n21594 & n25440 ;
  assign n25442 = n25441 ^ n20729 ;
  assign n25443 = n3833 & n25442 ;
  assign n25444 = n25443 ^ x29 ;
  assign n25446 = n25445 ^ n25444 ;
  assign n25448 = n25447 ^ n25446 ;
  assign n25430 = ~n61 & ~n20745 ;
  assign n25431 = n25430 ^ n20745 ;
  assign n25429 = ~n61 & n20739 ;
  assign n25432 = n25431 ^ n25429 ;
  assign n25433 = ~n3800 & n25432 ;
  assign n25420 = n21429 ^ n20738 ;
  assign n25419 = n21429 ^ n20739 ;
  assign n25421 = n25420 ^ n25419 ;
  assign n25424 = ~x30 & n25421 ;
  assign n25425 = n25424 ^ n25420 ;
  assign n25426 = ~n3518 & n25425 ;
  assign n25427 = n25426 ^ n21429 ;
  assign n25428 = x31 & ~n25427 ;
  assign n25434 = n25433 ^ n25428 ;
  assign n25412 = n5304 ^ n2956 ;
  assign n25413 = n25412 ^ n4758 ;
  assign n25414 = n25413 ^ n14484 ;
  assign n25409 = n1040 ^ n126 ;
  assign n25410 = n25409 ^ n919 ;
  assign n25407 = n2468 ^ n658 ;
  assign n25405 = n4280 ^ n575 ;
  assign n25406 = n25405 ^ n3920 ;
  assign n25408 = n25407 ^ n25406 ;
  assign n25411 = n25410 ^ n25408 ;
  assign n25415 = n25414 ^ n25411 ;
  assign n25416 = n25415 ^ n2760 ;
  assign n25417 = n25416 ^ n6925 ;
  assign n25418 = ~n6905 & ~n25417 ;
  assign n25435 = n25434 ^ n25418 ;
  assign n25402 = n25149 ^ n25145 ;
  assign n25403 = n25146 & n25402 ;
  assign n25404 = n25403 ^ n25149 ;
  assign n25436 = n25435 ^ n25404 ;
  assign n25399 = n25159 ^ n25150 ;
  assign n25400 = ~n25164 & n25399 ;
  assign n25401 = n25400 ^ n25159 ;
  assign n25437 = n25436 ^ n25401 ;
  assign n25449 = n25448 ^ n25437 ;
  assign n25451 = n25450 ^ n25449 ;
  assign n25392 = n20713 ^ n285 ;
  assign n25391 = n25390 ^ n20713 ;
  assign n25393 = n25392 ^ n25391 ;
  assign n25394 = n25392 ^ n20802 ;
  assign n25395 = n25394 ^ n25392 ;
  assign n25396 = n25393 & ~n25395 ;
  assign n25397 = n25396 ^ n25392 ;
  assign n25398 = n96 & n25397 ;
  assign n25452 = n25451 ^ n25398 ;
  assign n25385 = n25181 ^ n25117 ;
  assign n25386 = ~n25182 & ~n25385 ;
  assign n25387 = n25386 ^ n25181 ;
  assign n25453 = n25452 ^ n25387 ;
  assign n25454 = n25453 ^ x23 ;
  assign n25384 = n4655 & ~n20702 ;
  assign n25455 = n25454 ^ n25384 ;
  assign n25383 = n4651 & ~n20706 ;
  assign n25456 = n25455 ^ n25383 ;
  assign n25382 = n4656 & n22079 ;
  assign n25457 = n25456 ^ n25382 ;
  assign n25459 = n25458 ^ n25457 ;
  assign n25379 = n25203 ^ n25183 ;
  assign n25380 = n25189 & n25379 ;
  assign n25381 = n25380 ^ n25203 ;
  assign n25460 = n25459 ^ n25381 ;
  assign n25461 = n25460 ^ x20 ;
  assign n25374 = n20690 ^ n5224 ;
  assign n25375 = n25374 ^ n20690 ;
  assign n25376 = ~n21247 & n25375 ;
  assign n25377 = n25376 ^ n20690 ;
  assign n25378 = n5215 & ~n25377 ;
  assign n25462 = n25461 ^ n25378 ;
  assign n25464 = n25463 ^ n25462 ;
  assign n25466 = n25465 ^ n25464 ;
  assign n25371 = n25204 ^ n25106 ;
  assign n25372 = n25210 & n25371 ;
  assign n25373 = n25372 ^ n25204 ;
  assign n25467 = n25466 ^ n25373 ;
  assign n25468 = n25467 ^ x17 ;
  assign n25370 = n6148 & n20631 ;
  assign n25469 = n25468 ^ n25370 ;
  assign n25369 = n6143 & n20680 ;
  assign n25470 = n25469 ^ n25369 ;
  assign n25368 = n6163 & ~n22653 ;
  assign n25471 = n25470 ^ n25368 ;
  assign n25473 = n25472 ^ n25471 ;
  assign n25365 = n25222 ^ n25211 ;
  assign n25366 = ~n25219 & n25365 ;
  assign n25367 = n25366 ^ n25222 ;
  assign n25474 = n25473 ^ n25367 ;
  assign n25475 = n25474 ^ x14 ;
  assign n25364 = ~n6529 & ~n20628 ;
  assign n25476 = n25475 ^ n25364 ;
  assign n25363 = ~n6547 & n20819 ;
  assign n25477 = n25476 ^ n25363 ;
  assign n25358 = n22979 ^ n7310 ;
  assign n25359 = n25358 ^ n22979 ;
  assign n25360 = ~n22978 & ~n25359 ;
  assign n25361 = n25360 ^ n22979 ;
  assign n25362 = n6391 & ~n25361 ;
  assign n25478 = n25477 ^ n25362 ;
  assign n25482 = n25481 ^ n25478 ;
  assign n25484 = n25482 ^ n25094 ;
  assign n25483 = n25482 ^ n25242 ;
  assign n25485 = n25484 ^ n25483 ;
  assign n25486 = n25099 & ~n25485 ;
  assign n25487 = n25486 ^ n25484 ;
  assign n25496 = n25495 ^ n25487 ;
  assign n25354 = n25252 ^ n25243 ;
  assign n25355 = n25249 & n25354 ;
  assign n25356 = n25355 ^ n25252 ;
  assign n25497 = n25496 ^ n25356 ;
  assign n25350 = n8150 & n23893 ;
  assign n25349 = n8139 & ~n20613 ;
  assign n25351 = n25350 ^ n25349 ;
  assign n25347 = n8484 & ~n20612 ;
  assign n25346 = n8144 & ~n20614 ;
  assign n25348 = n25347 ^ n25346 ;
  assign n25352 = n25351 ^ n25348 ;
  assign n25353 = n25352 ^ x8 ;
  assign n25498 = n25497 ^ n25353 ;
  assign n25499 = n25498 ^ x5 ;
  assign n25339 = n21212 ^ n10329 ;
  assign n25340 = n25339 ^ n21212 ;
  assign n25341 = n21212 ^ n21170 ;
  assign n25342 = n25341 ^ n21212 ;
  assign n25343 = n25340 & ~n25342 ;
  assign n25344 = n25343 ^ n21212 ;
  assign n25345 = n10322 & ~n25344 ;
  assign n25500 = n25499 ^ n25345 ;
  assign n25338 = n10327 & n21147 ;
  assign n25501 = n25500 ^ n25338 ;
  assign n25503 = n25502 ^ n25501 ;
  assign n25335 = n25253 ^ n25078 ;
  assign n25336 = n25083 & ~n25335 ;
  assign n25337 = n25336 ^ n25078 ;
  assign n25504 = n25503 ^ n25337 ;
  assign n25332 = n25305 ^ n25257 ;
  assign n25333 = n25258 & ~n25332 ;
  assign n25334 = n25333 ^ n25305 ;
  assign n25505 = n25504 ^ n25334 ;
  assign n25330 = n25065 & ~n25306 ;
  assign n25318 = ~x0 & n25282 ;
  assign n25326 = n25318 ^ n11664 ;
  assign n25310 = ~n25282 & ~n25297 ;
  assign n25311 = ~n25296 & ~n25310 ;
  assign n25317 = n25311 ^ x2 ;
  assign n25319 = n25318 ^ n25317 ;
  assign n25320 = n25319 ^ n25311 ;
  assign n25321 = n25311 ^ n24841 ;
  assign n25322 = n25321 ^ n25311 ;
  assign n25323 = n25320 & n25322 ;
  assign n25324 = n25323 ^ n25311 ;
  assign n25325 = n11138 & ~n25324 ;
  assign n25327 = n25326 ^ n25325 ;
  assign n25315 = x0 & ~x2 ;
  assign n25316 = n25311 & n25315 ;
  assign n25328 = n25327 ^ n25316 ;
  assign n25308 = ~n24841 & n25282 ;
  assign n25312 = n25311 ^ n25308 ;
  assign n25313 = ~x1 & n25312 ;
  assign n25309 = n11663 & n25308 ;
  assign n25314 = n25313 ^ n25309 ;
  assign n25329 = n25328 ^ n25314 ;
  assign n25331 = n25330 ^ n25329 ;
  assign n25506 = n25505 ^ n25331 ;
  assign n25692 = ~n10334 & n21147 ;
  assign n25682 = n7142 & ~n20617 ;
  assign n25680 = n20240 & n23480 ;
  assign n25677 = n7151 & ~n20614 ;
  assign n25676 = n7148 & ~n20620 ;
  assign n25678 = n25677 ^ n25676 ;
  assign n25679 = n25678 ^ x11 ;
  assign n25681 = n25680 ^ n25679 ;
  assign n25683 = n25682 ^ n25681 ;
  assign n25672 = n25495 ^ n25482 ;
  assign n25673 = n25487 & n25672 ;
  assign n25674 = n25673 ^ n25482 ;
  assign n25668 = n25481 ^ n25474 ;
  assign n25669 = n25478 & n25668 ;
  assign n25670 = n25669 ^ n25474 ;
  assign n25660 = n25467 ^ n25367 ;
  assign n25661 = n25473 & n25660 ;
  assign n25662 = n25661 ^ n25467 ;
  assign n25658 = n20437 & n20680 ;
  assign n25655 = n6143 & n20631 ;
  assign n25653 = n6148 & n20819 ;
  assign n25649 = n13433 & ~n20693 ;
  assign n25647 = n5426 & ~n20690 ;
  assign n25640 = n20683 ^ x20 ;
  assign n25641 = n25640 ^ x19 ;
  assign n25642 = n25641 ^ n20683 ;
  assign n25643 = ~n22617 & n25642 ;
  assign n25644 = n25643 ^ n20683 ;
  assign n25645 = n5215 & ~n25644 ;
  assign n25646 = n25645 ^ x20 ;
  assign n25648 = n25647 ^ n25646 ;
  assign n25650 = n25649 ^ n25648 ;
  assign n25631 = n25453 ^ n25381 ;
  assign n25632 = ~n25459 & n25631 ;
  assign n25633 = n25632 ^ n25453 ;
  assign n25629 = ~n40 & ~n20702 ;
  assign n25621 = ~n4435 & n21782 ;
  assign n25619 = ~n4434 & ~n20706 ;
  assign n25616 = n4600 & n20713 ;
  assign n25615 = n20603 & n20716 ;
  assign n25617 = n25616 ^ n25615 ;
  assign n25618 = n25617 ^ x26 ;
  assign n25620 = n25619 ^ n25618 ;
  assign n25622 = n25621 ^ n25620 ;
  assign n25610 = n25434 ^ n25404 ;
  assign n25611 = ~n25435 & n25610 ;
  assign n25612 = n25611 ^ n25434 ;
  assign n25601 = n5732 ^ n413 ;
  assign n25602 = n25601 ^ n1503 ;
  assign n25599 = n2425 ^ n995 ;
  assign n25598 = n1837 ^ n1273 ;
  assign n25600 = n25599 ^ n25598 ;
  assign n25603 = n25602 ^ n25600 ;
  assign n25604 = n25603 ^ n2698 ;
  assign n25596 = n3884 ^ n2044 ;
  assign n25594 = n241 ^ n114 ;
  assign n25593 = n6319 ^ n649 ;
  assign n25595 = n25594 ^ n25593 ;
  assign n25597 = n25596 ^ n25595 ;
  assign n25605 = n25604 ^ n25597 ;
  assign n25590 = n14683 ^ n4257 ;
  assign n25587 = n785 ^ n250 ;
  assign n25588 = n25587 ^ n476 ;
  assign n25586 = n459 ^ n411 ;
  assign n25589 = n25588 ^ n25586 ;
  assign n25591 = n25590 ^ n25589 ;
  assign n25592 = n25591 ^ n24919 ;
  assign n25606 = n25605 ^ n25592 ;
  assign n25607 = n25606 ^ n4226 ;
  assign n25608 = ~n4812 & ~n25607 ;
  assign n25576 = x31 & ~n25429 ;
  assign n25579 = ~x30 & ~n20745 ;
  assign n25580 = n25579 ^ n21440 ;
  assign n25581 = ~n3518 & ~n25580 ;
  assign n25582 = n25581 ^ n21440 ;
  assign n25583 = n25576 & ~n25582 ;
  assign n25584 = n25583 ^ n25576 ;
  assign n25571 = n20745 ^ n61 ;
  assign n25572 = n25571 ^ n20745 ;
  assign n25573 = ~n20781 & n25572 ;
  assign n25574 = n25573 ^ n20745 ;
  assign n25575 = ~n3800 & n25574 ;
  assign n25585 = n25584 ^ n25575 ;
  assign n25609 = n25608 ^ n25585 ;
  assign n25613 = n25612 ^ n25609 ;
  assign n25569 = n3837 & n20737 ;
  assign n25567 = n3985 & n20729 ;
  assign n25562 = n25448 ^ n25401 ;
  assign n25563 = ~n25437 & ~n25562 ;
  assign n25564 = n25563 ^ n25448 ;
  assign n25565 = n25564 ^ x29 ;
  assign n25557 = n21736 ^ n5065 ;
  assign n25558 = n25557 ^ n21736 ;
  assign n25559 = n20800 & ~n25558 ;
  assign n25560 = n25559 ^ n21736 ;
  assign n25561 = n3833 & n25560 ;
  assign n25566 = n25565 ^ n25561 ;
  assign n25568 = n25567 ^ n25566 ;
  assign n25570 = n25569 ^ n25568 ;
  assign n25614 = n25613 ^ n25570 ;
  assign n25623 = n25622 ^ n25614 ;
  assign n25554 = n25449 ^ n25387 ;
  assign n25555 = n25452 & ~n25554 ;
  assign n25556 = n25555 ^ n25449 ;
  assign n25624 = n25623 ^ n25556 ;
  assign n25625 = n25624 ^ x23 ;
  assign n25553 = n4655 & ~n20694 ;
  assign n25626 = n25625 ^ n25553 ;
  assign n25552 = n4651 & ~n20705 ;
  assign n25627 = n25626 ^ n25552 ;
  assign n25551 = n4656 & n22601 ;
  assign n25628 = n25627 ^ n25551 ;
  assign n25630 = n25629 ^ n25628 ;
  assign n25634 = n25633 ^ n25630 ;
  assign n25635 = n25634 ^ n25460 ;
  assign n25636 = n25635 ^ n25373 ;
  assign n25637 = n25636 ^ n25634 ;
  assign n25638 = n25466 & n25637 ;
  assign n25639 = n25638 ^ n25635 ;
  assign n25651 = n25650 ^ n25639 ;
  assign n25652 = n25651 ^ x17 ;
  assign n25654 = n25653 ^ n25652 ;
  assign n25656 = n25655 ^ n25654 ;
  assign n25550 = n6163 & ~n21237 ;
  assign n25657 = n25656 ^ n25550 ;
  assign n25659 = n25658 ^ n25657 ;
  assign n25663 = n25662 ^ n25659 ;
  assign n25664 = n25663 ^ x14 ;
  assign n25549 = ~n6547 & ~n20628 ;
  assign n25665 = n25664 ^ n25549 ;
  assign n25548 = ~n6529 & n20829 ;
  assign n25666 = n25665 ^ n25548 ;
  assign n25542 = n20624 ^ n7310 ;
  assign n25543 = n25542 ^ n20624 ;
  assign n25545 = ~n21231 & n25543 ;
  assign n25546 = n25545 ^ n20624 ;
  assign n25547 = n6391 & n25546 ;
  assign n25667 = n25666 ^ n25547 ;
  assign n25671 = n25670 ^ n25667 ;
  assign n25675 = n25674 ^ n25671 ;
  assign n25684 = n25683 ^ n25675 ;
  assign n25685 = n25684 ^ n25352 ;
  assign n25539 = n8150 & ~n25056 ;
  assign n25538 = n8139 & ~n20612 ;
  assign n25540 = n25539 ^ n25538 ;
  assign n25536 = n8484 & n20908 ;
  assign n25535 = n8144 & ~n20613 ;
  assign n25537 = n25536 ^ n25535 ;
  assign n25541 = n25540 ^ n25537 ;
  assign n25686 = n25685 ^ n25541 ;
  assign n25532 = n25496 ^ n25353 ;
  assign n25533 = n25356 ^ n25353 ;
  assign n25534 = n25532 & ~n25533 ;
  assign n25687 = n25686 ^ n25534 ;
  assign n25688 = n25687 ^ x5 ;
  assign n25531 = n10425 & n24841 ;
  assign n25689 = n25688 ^ n25531 ;
  assign n25530 = n10327 & ~n21212 ;
  assign n25690 = n25689 ^ n25530 ;
  assign n25528 = n24841 ^ n24810 ;
  assign n25529 = n10342 & ~n25528 ;
  assign n25691 = n25690 ^ n25529 ;
  assign n25693 = n25692 ^ n25691 ;
  assign n25525 = n25498 ^ n25337 ;
  assign n25526 = ~n25503 & n25525 ;
  assign n25527 = n25526 ^ n25498 ;
  assign n25694 = n25693 ^ n25527 ;
  assign n25512 = n25318 ^ n25308 ;
  assign n25513 = x1 & ~n25512 ;
  assign n25514 = n11663 ^ n11657 ;
  assign n25515 = n25310 ^ n25308 ;
  assign n25516 = n25514 & ~n25515 ;
  assign n25517 = n25516 ^ n11657 ;
  assign n25518 = n25513 ^ n25318 ;
  assign n25519 = n25518 ^ x2 ;
  assign n25520 = ~n25517 & ~n25519 ;
  assign n25521 = ~n25513 & n25520 ;
  assign n25522 = ~x2 & n25521 ;
  assign n25523 = n25522 ^ n25520 ;
  assign n25524 = n25523 ^ n25517 ;
  assign n25695 = n25694 ^ n25524 ;
  assign n25509 = n25334 ^ n25329 ;
  assign n25510 = n25331 & n25509 ;
  assign n25507 = n25334 ^ n25331 ;
  assign n25508 = ~n25504 & ~n25507 ;
  assign n25511 = n25510 ^ n25508 ;
  assign n25696 = n25695 ^ n25511 ;
  assign n25882 = n25694 ^ n25329 ;
  assign n25881 = n25524 ^ n25334 ;
  assign n25883 = n25882 ^ n25881 ;
  assign n25884 = n25882 ^ n25505 ;
  assign n25885 = n25884 ^ n25882 ;
  assign n25886 = ~n25883 & ~n25885 ;
  assign n25887 = n25886 ^ n25882 ;
  assign n25888 = ~n25695 & n25887 ;
  assign n25889 = n25888 ^ n25694 ;
  assign n25879 = n11139 & n25308 ;
  assign n25880 = n25879 ^ x2 ;
  assign n25890 = n25889 ^ n25880 ;
  assign n25875 = n10425 & ~n25282 ;
  assign n25871 = n10327 & n24841 ;
  assign n25872 = n25871 ^ x5 ;
  assign n25870 = ~n10334 & ~n21212 ;
  assign n25873 = n25872 ^ n25870 ;
  assign n25868 = n25299 ^ n25282 ;
  assign n25869 = n10342 & n25868 ;
  assign n25874 = n25873 ^ n25869 ;
  assign n25876 = n25875 ^ n25874 ;
  assign n25865 = n8139 & n20908 ;
  assign n25856 = n25670 ^ n25663 ;
  assign n25857 = n25667 & n25856 ;
  assign n25858 = n25857 ^ n25663 ;
  assign n25851 = n20437 & n20631 ;
  assign n25842 = n25650 ^ n25634 ;
  assign n25843 = n25639 & n25842 ;
  assign n25844 = n25843 ^ n25634 ;
  assign n25839 = ~n40 & ~n20694 ;
  assign n25831 = n25622 ^ n25556 ;
  assign n25832 = ~n25623 & n25831 ;
  assign n25833 = n25832 ^ n25622 ;
  assign n25828 = ~n4435 & n21770 ;
  assign n25826 = ~n4434 & ~n20705 ;
  assign n25823 = n20603 & n20713 ;
  assign n25822 = n4600 & ~n20706 ;
  assign n25824 = n25823 ^ n25822 ;
  assign n25825 = n25824 ^ x26 ;
  assign n25827 = n25826 ^ n25825 ;
  assign n25829 = n25828 ^ n25827 ;
  assign n25818 = n3837 & n20729 ;
  assign n25816 = n3985 & n20725 ;
  assign n25809 = n20716 ^ x29 ;
  assign n25810 = n25809 ^ x28 ;
  assign n25811 = n25810 ^ n20716 ;
  assign n25812 = n20801 & n25811 ;
  assign n25813 = n25812 ^ n20716 ;
  assign n25814 = n3833 & n25813 ;
  assign n25815 = n25814 ^ x29 ;
  assign n25817 = n25816 ^ n25815 ;
  assign n25819 = n25818 ^ n25817 ;
  assign n25803 = n4124 ^ n4055 ;
  assign n25799 = n6062 ^ n1471 ;
  assign n25800 = n25799 ^ n2358 ;
  assign n25801 = n25800 ^ n1097 ;
  assign n25796 = n1011 ^ n716 ;
  assign n25797 = n25796 ^ n341 ;
  assign n25794 = n1027 ^ n188 ;
  assign n25793 = n1568 ^ n436 ;
  assign n25795 = n25794 ^ n25793 ;
  assign n25798 = n25797 ^ n25795 ;
  assign n25802 = n25801 ^ n25798 ;
  assign n25804 = n25803 ^ n25802 ;
  assign n25805 = n25804 ^ n14735 ;
  assign n25806 = ~n5689 & ~n25805 ;
  assign n25783 = x31 & ~n25430 ;
  assign n25786 = ~x30 & n20743 ;
  assign n25787 = n25786 ^ n21575 ;
  assign n25788 = ~n3518 & ~n25787 ;
  assign n25789 = n25788 ^ n21575 ;
  assign n25790 = n25783 & ~n25789 ;
  assign n25791 = n25790 ^ n25783 ;
  assign n25780 = n61 & ~n20780 ;
  assign n25781 = n25780 ^ n20743 ;
  assign n25782 = ~n3800 & ~n25781 ;
  assign n25792 = n25791 ^ n25782 ;
  assign n25807 = n25806 ^ n25792 ;
  assign n25775 = n25612 ^ n25585 ;
  assign n25776 = n25609 & n25775 ;
  assign n25777 = n25776 ^ n25612 ;
  assign n25808 = n25807 ^ n25777 ;
  assign n25820 = n25819 ^ n25808 ;
  assign n25772 = n25613 ^ n25564 ;
  assign n25773 = ~n25570 & ~n25772 ;
  assign n25774 = n25773 ^ n25613 ;
  assign n25821 = n25820 ^ n25774 ;
  assign n25830 = n25829 ^ n25821 ;
  assign n25834 = n25833 ^ n25830 ;
  assign n25835 = n25834 ^ x23 ;
  assign n25771 = n4655 & ~n20693 ;
  assign n25836 = n25835 ^ n25771 ;
  assign n25770 = n4651 & ~n20702 ;
  assign n25837 = n25836 ^ n25770 ;
  assign n25769 = n4656 & n22091 ;
  assign n25838 = n25837 ^ n25769 ;
  assign n25840 = n25839 ^ n25838 ;
  assign n25766 = n25633 ^ n25624 ;
  assign n25767 = n25630 & n25766 ;
  assign n25768 = n25767 ^ n25633 ;
  assign n25841 = n25840 ^ n25768 ;
  assign n25845 = n25844 ^ n25841 ;
  assign n25762 = n5220 & ~n22661 ;
  assign n25761 = n5215 & ~n22662 ;
  assign n25763 = n25762 ^ n25761 ;
  assign n25759 = n5426 & ~n20683 ;
  assign n25758 = n13433 & ~n20690 ;
  assign n25760 = n25759 ^ n25758 ;
  assign n25764 = n25763 ^ n25760 ;
  assign n25765 = n25764 ^ x20 ;
  assign n25846 = n25845 ^ n25765 ;
  assign n25847 = n25846 ^ x17 ;
  assign n25757 = n6143 & n20819 ;
  assign n25848 = n25847 ^ n25757 ;
  assign n25756 = n6148 & ~n20628 ;
  assign n25849 = n25848 ^ n25756 ;
  assign n25755 = n6163 & n23307 ;
  assign n25850 = n25849 ^ n25755 ;
  assign n25852 = n25851 ^ n25850 ;
  assign n25752 = n25662 ^ n25651 ;
  assign n25753 = ~n25659 & n25752 ;
  assign n25754 = n25753 ^ n25662 ;
  assign n25853 = n25852 ^ n25754 ;
  assign n25744 = n20620 ^ x14 ;
  assign n25743 = n20620 ^ x13 ;
  assign n25745 = n25744 ^ n25743 ;
  assign n25746 = n22963 & n25745 ;
  assign n25747 = n25746 ^ n25743 ;
  assign n25854 = n25853 ^ n25747 ;
  assign n25748 = n20624 ^ x14 ;
  assign n25749 = n25748 ^ n25747 ;
  assign n25740 = n20829 & n25543 ;
  assign n25741 = n25740 ^ n20624 ;
  assign n25742 = ~n6540 & n25741 ;
  assign n25750 = n25749 ^ n25742 ;
  assign n25751 = ~n6391 & ~n25750 ;
  assign n25855 = n25854 ^ n25751 ;
  assign n25859 = n25858 ^ n25855 ;
  assign n25733 = n7148 & ~n20617 ;
  assign n25731 = n7142 & ~n20614 ;
  assign n25724 = n20613 ^ x11 ;
  assign n25725 = n25724 ^ x10 ;
  assign n25726 = n25725 ^ n20613 ;
  assign n25727 = ~n21226 & n25726 ;
  assign n25728 = n25727 ^ n20613 ;
  assign n25729 = n7140 & ~n25728 ;
  assign n25730 = n25729 ^ x11 ;
  assign n25732 = n25731 ^ n25730 ;
  assign n25734 = n25733 ^ n25732 ;
  assign n25735 = n25734 ^ n25683 ;
  assign n25736 = n25735 ^ n25674 ;
  assign n25737 = n25736 ^ n25734 ;
  assign n25738 = ~n25675 & n25737 ;
  assign n25739 = n25738 ^ n25735 ;
  assign n25860 = n25859 ^ n25739 ;
  assign n25861 = n25860 ^ x8 ;
  assign n25722 = n8484 & n21147 ;
  assign n25862 = n25861 ^ n25722 ;
  assign n25721 = n8144 & ~n20612 ;
  assign n25863 = n25862 ^ n25721 ;
  assign n25720 = n8150 & ~n25073 ;
  assign n25864 = n25863 ^ n25720 ;
  assign n25866 = n25865 ^ n25864 ;
  assign n25710 = ~n25356 & n25496 ;
  assign n25711 = n25710 ^ n25497 ;
  assign n25712 = n25353 & ~n25686 ;
  assign n25713 = ~n25711 & n25712 ;
  assign n25714 = n25710 ^ n25684 ;
  assign n25715 = n25541 ^ x8 ;
  assign n25716 = n25715 ^ n25684 ;
  assign n25717 = n25714 & n25716 ;
  assign n25718 = n25717 ^ n25684 ;
  assign n25719 = ~n25713 & ~n25718 ;
  assign n25867 = n25866 ^ n25719 ;
  assign n25877 = n25876 ^ n25867 ;
  assign n25707 = n25687 ^ n25527 ;
  assign n25708 = ~n25693 & ~n25707 ;
  assign n25709 = n25708 ^ n25527 ;
  assign n25878 = n25877 ^ n25709 ;
  assign n25891 = n25890 ^ n25878 ;
  assign n25697 = n25504 ^ n25329 ;
  assign n25698 = n25697 ^ n25334 ;
  assign n25699 = n25330 & ~n25698 ;
  assign n25700 = n25695 ^ n25334 ;
  assign n25701 = n25700 ^ n25695 ;
  assign n25702 = n25695 ^ n25329 ;
  assign n25703 = n25702 ^ n25695 ;
  assign n25704 = n25701 & ~n25703 ;
  assign n25705 = n25704 ^ n25695 ;
  assign n25706 = n25699 & ~n25705 ;
  assign n25892 = n25891 ^ n25706 ;
  assign n25893 = n25878 ^ n25706 ;
  assign n25894 = n25893 ^ n25706 ;
  assign n25895 = n25880 & ~n25889 ;
  assign n25896 = n25895 ^ n25706 ;
  assign n25897 = n25896 ^ n25706 ;
  assign n25898 = ~n25894 & ~n25897 ;
  assign n25899 = n25898 ^ n25706 ;
  assign n26077 = n25895 ^ n25890 ;
  assign n26069 = n10342 & n25311 ;
  assign n26068 = ~n10334 & n24841 ;
  assign n26070 = n26069 ^ n26068 ;
  assign n26071 = n26070 ^ n10327 ;
  assign n26065 = n10425 & ~n24841 ;
  assign n26066 = n26065 ^ n10327 ;
  assign n26067 = n25282 & n26066 ;
  assign n26072 = n26071 ^ n26067 ;
  assign n26073 = n26072 ^ n6053 ;
  assign n26055 = n8484 & ~n21212 ;
  assign n26054 = n8144 & n20908 ;
  assign n26056 = n26055 ^ n26054 ;
  assign n26057 = n26056 ^ x8 ;
  assign n26053 = n8150 & n25341 ;
  assign n26058 = n26057 ^ n26053 ;
  assign n26052 = n8139 & n21147 ;
  assign n26059 = n26058 ^ n26052 ;
  assign n26048 = n25860 ^ n25719 ;
  assign n26049 = n25866 & ~n26048 ;
  assign n26050 = n26049 ^ n25860 ;
  assign n26045 = n7142 & ~n20613 ;
  assign n26042 = n7148 & ~n20614 ;
  assign n26040 = n7151 & ~n20612 ;
  assign n26032 = n25846 ^ n25754 ;
  assign n26033 = ~n25852 & ~n26032 ;
  assign n26034 = n26033 ^ n25846 ;
  assign n26030 = n20437 & n20819 ;
  assign n26023 = n25841 ^ n25765 ;
  assign n26024 = n25845 & ~n26023 ;
  assign n26017 = n5221 & ~n22653 ;
  assign n26016 = n13433 & ~n20683 ;
  assign n26018 = n26017 ^ n26016 ;
  assign n26015 = n5220 & n20631 ;
  assign n26019 = n26018 ^ n26015 ;
  assign n26014 = n5426 & n20680 ;
  assign n26020 = n26019 ^ n26014 ;
  assign n26021 = n26020 ^ n25764 ;
  assign n26010 = n25834 ^ n25768 ;
  assign n26011 = n25840 & ~n26010 ;
  assign n26012 = n26011 ^ n25834 ;
  assign n26008 = ~n40 & ~n20693 ;
  assign n26005 = n13745 & ~n20690 ;
  assign n26003 = n4651 & ~n20694 ;
  assign n25998 = ~n4435 & n22079 ;
  assign n25996 = ~n4434 & ~n20702 ;
  assign n25993 = n4600 & ~n20705 ;
  assign n25992 = n20603 & ~n20706 ;
  assign n25994 = n25993 ^ n25992 ;
  assign n25995 = n25994 ^ x26 ;
  assign n25997 = n25996 ^ n25995 ;
  assign n25999 = n25998 ^ n25997 ;
  assign n25988 = n25819 ^ n25774 ;
  assign n25989 = ~n25820 & ~n25988 ;
  assign n25990 = n25989 ^ n25819 ;
  assign n25985 = n3985 & n20716 ;
  assign n25983 = n3837 & n20725 ;
  assign n25976 = n20713 ^ x29 ;
  assign n25977 = n25976 ^ x28 ;
  assign n25978 = n25977 ^ n20713 ;
  assign n25979 = n22063 & n25978 ;
  assign n25980 = n25979 ^ n20713 ;
  assign n25981 = n3833 & n25980 ;
  assign n25982 = n25981 ^ x29 ;
  assign n25984 = n25983 ^ n25982 ;
  assign n25986 = n25985 ^ n25984 ;
  assign n25972 = n25792 ^ n25777 ;
  assign n25973 = n25807 & n25972 ;
  assign n25974 = n25973 ^ n25777 ;
  assign n25962 = n14271 ^ n2679 ;
  assign n25961 = n2176 ^ n1180 ;
  assign n25963 = n25962 ^ n25961 ;
  assign n25964 = n25963 ^ n13625 ;
  assign n25965 = n25964 ^ n25410 ;
  assign n25957 = n3370 ^ n1680 ;
  assign n25958 = n25957 ^ n2277 ;
  assign n25955 = n5551 ^ n149 ;
  assign n25956 = n25955 ^ n575 ;
  assign n25959 = n25958 ^ n25956 ;
  assign n25952 = n1461 ^ n322 ;
  assign n25951 = n1735 ^ n495 ;
  assign n25953 = n25952 ^ n25951 ;
  assign n25950 = n23973 ^ n4867 ;
  assign n25954 = n25953 ^ n25950 ;
  assign n25960 = n25959 ^ n25954 ;
  assign n25966 = n25965 ^ n25960 ;
  assign n25967 = n14052 ^ n5503 ;
  assign n25968 = n25967 ^ n3246 ;
  assign n25969 = ~n25966 & ~n25968 ;
  assign n25944 = n20729 ^ n3518 ;
  assign n25943 = ~n3518 & ~n20729 ;
  assign n25945 = n25944 ^ n25943 ;
  assign n25942 = ~n61 & n20737 ;
  assign n25946 = n25945 ^ n25942 ;
  assign n25970 = n25969 ^ n25946 ;
  assign n25947 = n25946 ^ n21593 ;
  assign n25935 = n21593 ^ n20743 ;
  assign n25934 = n21593 ^ n20737 ;
  assign n25936 = n25935 ^ n25934 ;
  assign n25939 = ~x30 & ~n25936 ;
  assign n25940 = n25939 ^ n25935 ;
  assign n25941 = ~n3518 & n25940 ;
  assign n25948 = n25947 ^ n25941 ;
  assign n25949 = x31 & n25948 ;
  assign n25971 = n25970 ^ n25949 ;
  assign n25975 = n25974 ^ n25971 ;
  assign n25987 = n25986 ^ n25975 ;
  assign n25991 = n25990 ^ n25987 ;
  assign n26000 = n25999 ^ n25991 ;
  assign n25931 = n25833 ^ n25829 ;
  assign n25932 = ~n25830 & n25931 ;
  assign n25933 = n25932 ^ n25833 ;
  assign n26001 = n26000 ^ n25933 ;
  assign n26002 = n26001 ^ x23 ;
  assign n26004 = n26003 ^ n26002 ;
  assign n26006 = n26005 ^ n26004 ;
  assign n25929 = n13744 & n21246 ;
  assign n25928 = n38 & ~n21244 ;
  assign n25930 = n25929 ^ n25928 ;
  assign n26007 = n26006 ^ n25930 ;
  assign n26009 = n26008 ^ n26007 ;
  assign n26013 = n26012 ^ n26009 ;
  assign n26022 = n26021 ^ n26013 ;
  assign n26025 = n26024 ^ n26022 ;
  assign n26026 = n26025 ^ x17 ;
  assign n25927 = n6148 & n20829 ;
  assign n26027 = n26026 ^ n25927 ;
  assign n25926 = n6143 & ~n20628 ;
  assign n26028 = n26027 ^ n25926 ;
  assign n25925 = n6163 & ~n22979 ;
  assign n26029 = n26028 ^ n25925 ;
  assign n26031 = n26030 ^ n26029 ;
  assign n26035 = n26034 ^ n26031 ;
  assign n25909 = n25744 ^ x13 ;
  assign n25910 = n25909 ^ n20620 ;
  assign n25911 = n20624 & n25910 ;
  assign n25912 = n25911 ^ n20620 ;
  assign n25913 = ~n6540 & ~n25912 ;
  assign n25914 = n25913 ^ n25744 ;
  assign n26036 = n26035 ^ n25914 ;
  assign n25915 = n20617 ^ x13 ;
  assign n25916 = n25915 ^ n25914 ;
  assign n25917 = n25916 ^ x13 ;
  assign n25918 = n25917 ^ x14 ;
  assign n25919 = n25918 ^ n25916 ;
  assign n25920 = n25916 ^ n23490 ;
  assign n25921 = n25920 ^ n25916 ;
  assign n25922 = n25919 & n25921 ;
  assign n25923 = n25922 ^ n25916 ;
  assign n25924 = n6391 & n25923 ;
  assign n26037 = n26036 ^ n25924 ;
  assign n25906 = n25858 ^ n25853 ;
  assign n25907 = ~n25855 & ~n25906 ;
  assign n25908 = n25907 ^ n25858 ;
  assign n26038 = n26037 ^ n25908 ;
  assign n26039 = n26038 ^ x11 ;
  assign n26041 = n26040 ^ n26039 ;
  assign n26043 = n26042 ^ n26041 ;
  assign n25905 = n20240 & n23893 ;
  assign n26044 = n26043 ^ n25905 ;
  assign n26046 = n26045 ^ n26044 ;
  assign n25902 = n25859 ^ n25734 ;
  assign n25903 = n25739 & n25902 ;
  assign n25904 = n25903 ^ n25734 ;
  assign n26047 = n26046 ^ n25904 ;
  assign n26051 = n26050 ^ n26047 ;
  assign n26060 = n26059 ^ n26051 ;
  assign n26074 = n26073 ^ n26060 ;
  assign n26075 = n26074 ^ n25867 ;
  assign n25900 = n25867 ^ n25709 ;
  assign n25901 = ~n25877 & n25900 ;
  assign n26076 = n26075 ^ n25901 ;
  assign n26078 = n26077 ^ n26076 ;
  assign n26079 = n26078 ^ n25706 ;
  assign n26080 = n26079 ^ n26076 ;
  assign n26081 = n25899 & ~n26080 ;
  assign n26082 = n26081 ^ n26078 ;
  assign n26274 = n8484 & n24841 ;
  assign n26273 = n8144 & n21147 ;
  assign n26275 = n26274 ^ n26273 ;
  assign n26276 = n26275 ^ x8 ;
  assign n26272 = n8150 & ~n25528 ;
  assign n26277 = n26276 ^ n26272 ;
  assign n26271 = n8139 & ~n21212 ;
  assign n26278 = n26277 ^ n26271 ;
  assign n26266 = n26035 ^ n25908 ;
  assign n26267 = n26037 & ~n26266 ;
  assign n26268 = n26267 ^ n26035 ;
  assign n26263 = n7142 & ~n20612 ;
  assign n26261 = n20240 & ~n25056 ;
  assign n26258 = n7151 & n20908 ;
  assign n26257 = n7148 & ~n20613 ;
  assign n26259 = n26258 ^ n26257 ;
  assign n26260 = n26259 ^ x11 ;
  assign n26262 = n26261 ^ n26260 ;
  assign n26264 = n26263 ^ n26262 ;
  assign n26235 = ~n6547 & ~n20620 ;
  assign n26234 = ~n6529 & ~n20617 ;
  assign n26236 = n26235 ^ n26234 ;
  assign n26237 = n26236 ^ n6537 ;
  assign n26238 = n26237 ^ x14 ;
  assign n26239 = n26236 ^ x14 ;
  assign n26244 = n26239 ^ n6539 ;
  assign n26240 = n20614 ^ n17173 ;
  assign n26241 = n26240 ^ n23479 ;
  assign n26242 = n26241 ^ n26240 ;
  assign n26243 = n26239 & ~n26242 ;
  assign n26245 = n26244 ^ n26243 ;
  assign n26246 = n26240 ^ n20614 ;
  assign n26247 = ~n26242 & ~n26246 ;
  assign n26248 = n26247 ^ n20614 ;
  assign n26249 = ~n26244 & n26248 ;
  assign n26250 = ~n26245 & n26249 ;
  assign n26251 = n26250 ^ n26247 ;
  assign n26252 = n26251 ^ n6539 ;
  assign n26253 = n26252 ^ n20614 ;
  assign n26254 = ~n26238 & ~n26253 ;
  assign n26228 = n6148 & n20624 ;
  assign n26227 = n6143 & n20829 ;
  assign n26229 = n26228 ^ n26227 ;
  assign n26230 = n26229 ^ x17 ;
  assign n26226 = n6163 & ~n21232 ;
  assign n26231 = n26230 ^ n26226 ;
  assign n26225 = n20437 & ~n20628 ;
  assign n26232 = n26231 ^ n26225 ;
  assign n26221 = n13433 & n20680 ;
  assign n26219 = n5426 & n20631 ;
  assign n26213 = ~n4435 & n22601 ;
  assign n26211 = ~n4434 & ~n20694 ;
  assign n26208 = n4600 & ~n20702 ;
  assign n26207 = n20603 & ~n20705 ;
  assign n26209 = n26208 ^ n26207 ;
  assign n26210 = n26209 ^ x26 ;
  assign n26212 = n26211 ^ n26210 ;
  assign n26214 = n26213 ^ n26212 ;
  assign n26203 = n3837 & n20716 ;
  assign n26201 = n3985 & n20713 ;
  assign n26194 = n20706 ^ x29 ;
  assign n26195 = n26194 ^ x28 ;
  assign n26196 = n26195 ^ n20706 ;
  assign n26197 = ~n23801 & n26196 ;
  assign n26198 = n26197 ^ n20706 ;
  assign n26199 = n3833 & ~n26198 ;
  assign n26200 = n26199 ^ x29 ;
  assign n26202 = n26201 ^ n26200 ;
  assign n26204 = n26203 ^ n26202 ;
  assign n26186 = x31 & n25942 ;
  assign n26184 = n12664 & ~n25943 ;
  assign n26182 = ~n61 & n20729 ;
  assign n26179 = ~x31 & n20800 ;
  assign n26180 = n26179 ^ n21736 ;
  assign n26181 = n3518 & ~n26180 ;
  assign n26183 = n26182 ^ n26181 ;
  assign n26185 = n26184 ^ n26183 ;
  assign n26187 = n26186 ^ n26185 ;
  assign n26169 = n5678 ^ n3603 ;
  assign n26170 = n26169 ^ n13502 ;
  assign n26171 = n26170 ^ n12481 ;
  assign n26172 = n26171 ^ n2579 ;
  assign n26163 = n12575 ^ n1065 ;
  assign n26164 = n26163 ^ n3880 ;
  assign n26160 = n389 ^ n379 ;
  assign n26161 = n26160 ^ n362 ;
  assign n26159 = n813 ^ n735 ;
  assign n26162 = n26161 ^ n26159 ;
  assign n26165 = n26164 ^ n26162 ;
  assign n26166 = n12756 ^ n2949 ;
  assign n26167 = n26166 ^ n169 ;
  assign n26168 = ~n26165 & n26167 ;
  assign n26173 = n26172 ^ n26168 ;
  assign n26174 = ~n2980 & n26173 ;
  assign n26175 = ~n696 & n26174 ;
  assign n26176 = n26175 ^ x2 ;
  assign n26188 = n26187 ^ n26176 ;
  assign n26189 = n26188 ^ n25974 ;
  assign n26190 = n26189 ^ n25969 ;
  assign n26191 = n26190 ^ n26188 ;
  assign n26192 = ~n25971 & ~n26191 ;
  assign n26193 = n26192 ^ n26189 ;
  assign n26205 = n26204 ^ n26193 ;
  assign n26156 = n25990 ^ n25986 ;
  assign n26157 = ~n25987 & n26156 ;
  assign n26158 = n26157 ^ n25990 ;
  assign n26206 = n26205 ^ n26158 ;
  assign n26215 = n26214 ^ n26206 ;
  assign n26149 = n13743 & ~n22617 ;
  assign n26147 = ~n40 & ~n20690 ;
  assign n26143 = n38 ^ n35 ;
  assign n26144 = ~n20683 & n26143 ;
  assign n26142 = n4651 & ~n20693 ;
  assign n26145 = n26144 ^ n26142 ;
  assign n26140 = n38 & n22618 ;
  assign n26139 = x23 & n22617 ;
  assign n26141 = n26140 ^ n26139 ;
  assign n26146 = n26145 ^ n26141 ;
  assign n26148 = n26147 ^ n26146 ;
  assign n26150 = n26149 ^ n26148 ;
  assign n26151 = n26150 ^ n25999 ;
  assign n26152 = n26151 ^ n26150 ;
  assign n26153 = n26152 ^ n25933 ;
  assign n26154 = n26000 & n26153 ;
  assign n26155 = n26154 ^ n26151 ;
  assign n26216 = n26215 ^ n26155 ;
  assign n26217 = n26216 ^ x20 ;
  assign n26134 = n21237 ^ n5224 ;
  assign n26135 = n26134 ^ n21237 ;
  assign n26136 = ~n21236 & ~n26135 ;
  assign n26137 = n26136 ^ n21237 ;
  assign n26138 = n5215 & ~n26137 ;
  assign n26218 = n26217 ^ n26138 ;
  assign n26220 = n26219 ^ n26218 ;
  assign n26222 = n26221 ^ n26220 ;
  assign n26131 = n26012 ^ n26001 ;
  assign n26132 = ~n26009 & n26131 ;
  assign n26133 = n26132 ^ n26012 ;
  assign n26223 = n26222 ^ n26133 ;
  assign n26121 = ~n25841 & n25844 ;
  assign n26122 = n26121 ^ n25845 ;
  assign n26123 = n25765 & ~n26022 ;
  assign n26124 = ~n26122 & n26123 ;
  assign n26125 = n26121 ^ n26013 ;
  assign n26126 = n26020 ^ x20 ;
  assign n26127 = n26126 ^ n26013 ;
  assign n26128 = n26125 & n26127 ;
  assign n26129 = n26128 ^ n26013 ;
  assign n26130 = ~n26124 & ~n26129 ;
  assign n26224 = n26223 ^ n26130 ;
  assign n26233 = n26232 ^ n26224 ;
  assign n26255 = n26254 ^ n26233 ;
  assign n26118 = n26034 ^ n26025 ;
  assign n26119 = ~n26031 & ~n26118 ;
  assign n26120 = n26119 ^ n26034 ;
  assign n26256 = n26255 ^ n26120 ;
  assign n26265 = n26264 ^ n26256 ;
  assign n26269 = n26268 ^ n26265 ;
  assign n26115 = n26038 ^ n25904 ;
  assign n26116 = n26046 & n26115 ;
  assign n26117 = n26116 ^ n26038 ;
  assign n26270 = n26269 ^ n26117 ;
  assign n26279 = n26278 ^ n26270 ;
  assign n26110 = n26060 ^ x2 ;
  assign n26111 = n26072 ^ x5 ;
  assign n26112 = n26111 ^ n26060 ;
  assign n26113 = n26110 & ~n26112 ;
  assign n26114 = n26113 ^ x2 ;
  assign n26284 = n26279 ^ n26114 ;
  assign n26280 = ~n26114 & n26279 ;
  assign n26285 = n26284 ^ n26280 ;
  assign n26106 = n26059 ^ n26050 ;
  assign n26107 = ~n26051 & n26106 ;
  assign n26108 = n26107 ^ n26059 ;
  assign n26104 = n10342 & n25515 ;
  assign n26100 = n10332 ^ n10322 ;
  assign n26101 = n26100 ^ n25871 ;
  assign n26102 = n25282 & ~n26101 ;
  assign n26099 = n10334 ^ x5 ;
  assign n26103 = n26102 ^ n26099 ;
  assign n26105 = n26104 ^ n26103 ;
  assign n26282 = n26108 ^ n26105 ;
  assign n26109 = ~n26105 & n26108 ;
  assign n26283 = n26282 ^ n26109 ;
  assign n26286 = n26285 ^ n26283 ;
  assign n26281 = n26280 ^ n26109 ;
  assign n26287 = n26286 ^ n26281 ;
  assign n26086 = n26074 ^ n25876 ;
  assign n26087 = n26074 ^ n25709 ;
  assign n26088 = n26086 & ~n26087 ;
  assign n26089 = ~n26075 & n26088 ;
  assign n26090 = n26089 ^ n26075 ;
  assign n26091 = n26090 ^ n25867 ;
  assign n26092 = ~n26077 & n26091 ;
  assign n26093 = n26074 ^ n25895 ;
  assign n26096 = ~n26076 & n26093 ;
  assign n26097 = n26096 ^ n26074 ;
  assign n26098 = ~n26092 & ~n26097 ;
  assign n26288 = n26287 ^ n26098 ;
  assign n26083 = n26076 ^ n25895 ;
  assign n26084 = n25706 & ~n25891 ;
  assign n26085 = ~n26083 & n26084 ;
  assign n26289 = n26288 ^ n26085 ;
  assign n26477 = n7151 & n21147 ;
  assign n26476 = n7148 & ~n20612 ;
  assign n26478 = n26477 ^ n26476 ;
  assign n26479 = n26478 ^ x11 ;
  assign n26475 = n20240 & ~n25073 ;
  assign n26480 = n26479 ^ n26475 ;
  assign n26474 = n7142 & n20908 ;
  assign n26481 = n26480 ^ n26474 ;
  assign n26449 = n6538 & ~n20613 ;
  assign n26451 = ~n6529 & ~n20614 ;
  assign n26450 = ~n6547 & ~n20617 ;
  assign n26452 = n26451 ^ n26450 ;
  assign n26453 = x14 & n26452 ;
  assign n26454 = n26449 & ~n26453 ;
  assign n26456 = ~x14 & n21226 ;
  assign n26455 = ~x13 & ~n21226 ;
  assign n26457 = n26456 ^ n26455 ;
  assign n26458 = n26452 ^ n6537 ;
  assign n26459 = n26458 ^ x14 ;
  assign n26460 = n26449 ^ n6538 ;
  assign n26461 = n26456 ^ n26453 ;
  assign n26462 = ~n26455 & ~n26461 ;
  assign n26463 = n26460 & n26462 ;
  assign n26464 = ~n26459 & ~n26463 ;
  assign n26465 = n26457 & n26464 ;
  assign n26466 = n26454 & n26465 ;
  assign n26467 = n26466 ^ n26464 ;
  assign n26445 = n20437 & n20829 ;
  assign n26443 = n6163 & n22968 ;
  assign n26440 = n6148 & ~n20620 ;
  assign n26439 = n6143 & n20624 ;
  assign n26441 = n26440 ^ n26439 ;
  assign n26442 = n26441 ^ x17 ;
  assign n26444 = n26443 ^ n26442 ;
  assign n26446 = n26445 ^ n26444 ;
  assign n26435 = n26216 ^ n26133 ;
  assign n26436 = ~n26222 & ~n26435 ;
  assign n26437 = n26436 ^ n26216 ;
  assign n26432 = n5426 & n20819 ;
  assign n26430 = n5220 & ~n20628 ;
  assign n26427 = n5221 & n23307 ;
  assign n26426 = n13433 & n20631 ;
  assign n26428 = n26427 ^ n26426 ;
  assign n26429 = n26428 ^ x20 ;
  assign n26431 = n26430 ^ n26429 ;
  assign n26433 = n26432 ^ n26431 ;
  assign n26418 = ~n40 & ~n20683 ;
  assign n26416 = n4656 & ~n22662 ;
  assign n26413 = n4655 & n20680 ;
  assign n26412 = n4651 & ~n20690 ;
  assign n26414 = n26413 ^ n26412 ;
  assign n26415 = n26414 ^ x23 ;
  assign n26417 = n26416 ^ n26415 ;
  assign n26419 = n26418 ^ n26417 ;
  assign n26408 = n3985 & ~n20706 ;
  assign n26399 = n26187 ^ n26175 ;
  assign n26400 = ~n26176 & n26399 ;
  assign n26401 = n26400 ^ x2 ;
  assign n26380 = n5302 ^ n637 ;
  assign n26378 = n13017 ^ n818 ;
  assign n26379 = n26378 ^ n438 ;
  assign n26381 = n26380 ^ n26379 ;
  assign n26382 = n26381 ^ n1980 ;
  assign n26392 = n4025 ^ n2956 ;
  assign n26391 = n3997 ^ n1465 ;
  assign n26393 = n26392 ^ n26391 ;
  assign n26389 = n1834 ^ n1291 ;
  assign n26388 = n1702 ^ n1260 ;
  assign n26390 = n26389 ^ n26388 ;
  assign n26394 = n26393 ^ n26390 ;
  assign n26385 = n1298 ^ n1008 ;
  assign n26383 = n3647 ^ n430 ;
  assign n26384 = n26383 ^ n435 ;
  assign n26386 = n26385 ^ n26384 ;
  assign n26387 = n26386 ^ n2544 ;
  assign n26395 = n26394 ^ n26387 ;
  assign n26396 = n26395 ^ n3269 ;
  assign n26397 = ~n14837 & ~n26396 ;
  assign n26398 = ~n26382 & n26397 ;
  assign n26402 = n26401 ^ n26398 ;
  assign n26403 = n26402 ^ x2 ;
  assign n26368 = n21754 ^ n3807 ;
  assign n26369 = n26368 ^ n26182 ;
  assign n26367 = ~n61 & n20725 ;
  assign n26370 = n26369 ^ n26367 ;
  assign n26365 = n21754 ^ n20725 ;
  assign n26366 = ~n22005 & n26365 ;
  assign n26371 = n26370 ^ n26366 ;
  assign n26357 = n26182 ^ n20725 ;
  assign n26358 = n26357 ^ n3807 ;
  assign n26359 = n26358 ^ n26357 ;
  assign n26360 = n26357 ^ n20716 ;
  assign n26361 = n26360 ^ n26357 ;
  assign n26362 = n26359 & ~n26361 ;
  assign n26363 = n26362 ^ n26357 ;
  assign n26364 = ~x31 & n26363 ;
  assign n26372 = n26371 ^ n26364 ;
  assign n26374 = n26372 ^ n26188 ;
  assign n26373 = n26372 ^ n26204 ;
  assign n26375 = n26374 ^ n26373 ;
  assign n26376 = ~n26193 & ~n26375 ;
  assign n26377 = n26376 ^ n26374 ;
  assign n26404 = n26403 ^ n26377 ;
  assign n26405 = n26404 ^ x29 ;
  assign n26351 = n21770 ^ n20705 ;
  assign n26352 = n20705 ^ n5065 ;
  assign n26353 = n26352 ^ n20705 ;
  assign n26354 = ~n26351 & n26353 ;
  assign n26355 = n26354 ^ n20705 ;
  assign n26356 = n3833 & ~n26355 ;
  assign n26406 = n26405 ^ n26356 ;
  assign n26349 = n3837 & n20713 ;
  assign n26407 = n26406 ^ n26349 ;
  assign n26409 = n26408 ^ n26407 ;
  assign n26328 = n4600 & ~n20694 ;
  assign n26327 = n20603 & ~n20702 ;
  assign n26329 = n26328 ^ n26327 ;
  assign n26330 = n26329 ^ n97 ;
  assign n26331 = n26329 ^ x26 ;
  assign n26332 = n26331 ^ n99 ;
  assign n26333 = n26332 ^ x25 ;
  assign n26334 = n26333 ^ n20693 ;
  assign n26335 = n26334 ^ n26331 ;
  assign n26336 = n26335 ^ n22090 ;
  assign n26337 = n26336 ^ n26335 ;
  assign n26338 = n26331 & ~n26337 ;
  assign n26339 = n26338 ^ n26332 ;
  assign n26340 = n26335 ^ n20693 ;
  assign n26341 = ~n26337 & ~n26340 ;
  assign n26342 = n26341 ^ n20693 ;
  assign n26343 = ~n26332 & n26342 ;
  assign n26344 = ~n26339 & n26343 ;
  assign n26345 = n26344 ^ n26341 ;
  assign n26346 = n26345 ^ n99 ;
  assign n26347 = n26346 ^ n20693 ;
  assign n26348 = ~n26330 & ~n26347 ;
  assign n26410 = n26409 ^ n26348 ;
  assign n26324 = n26214 ^ n26158 ;
  assign n26325 = n26206 & n26324 ;
  assign n26326 = n26325 ^ n26214 ;
  assign n26411 = n26410 ^ n26326 ;
  assign n26420 = n26419 ^ n26411 ;
  assign n26422 = n26420 ^ n26150 ;
  assign n26421 = n26420 ^ n26215 ;
  assign n26423 = n26422 ^ n26421 ;
  assign n26424 = n26155 & ~n26423 ;
  assign n26425 = n26424 ^ n26422 ;
  assign n26434 = n26433 ^ n26425 ;
  assign n26438 = n26437 ^ n26434 ;
  assign n26447 = n26446 ^ n26438 ;
  assign n26321 = n26232 ^ n26223 ;
  assign n26322 = ~n26224 & ~n26321 ;
  assign n26323 = n26322 ^ n26232 ;
  assign n26448 = n26447 ^ n26323 ;
  assign n26468 = n26467 ^ n26448 ;
  assign n26469 = n26468 ^ n26254 ;
  assign n26470 = n26469 ^ n26468 ;
  assign n26471 = n26470 ^ n26120 ;
  assign n26472 = ~n26255 & n26471 ;
  assign n26473 = n26472 ^ n26469 ;
  assign n26482 = n26481 ^ n26473 ;
  assign n26301 = n8139 & n24841 ;
  assign n26300 = n8144 & ~n21212 ;
  assign n26302 = n26301 ^ n26300 ;
  assign n26303 = n26302 ^ n8145 ;
  assign n26304 = n26303 ^ x8 ;
  assign n26305 = n26302 ^ x8 ;
  assign n26306 = n26305 ^ n8146 ;
  assign n26313 = n25282 & n26306 ;
  assign n26309 = ~x7 & ~n26306 ;
  assign n26310 = n26309 ^ n8147 ;
  assign n26311 = ~n25299 & ~n26310 ;
  assign n26312 = n26311 ^ n8146 ;
  assign n26314 = n26313 ^ n26312 ;
  assign n26315 = ~n26304 & ~n26314 ;
  assign n26316 = n26315 ^ n26268 ;
  assign n26317 = n26316 ^ n26264 ;
  assign n26318 = n26317 ^ n26315 ;
  assign n26319 = ~n26265 & ~n26318 ;
  assign n26320 = n26319 ^ n26316 ;
  assign n26483 = n26482 ^ n26320 ;
  assign n26293 = ~n10334 & n25308 ;
  assign n26294 = n26293 ^ x5 ;
  assign n26295 = n26294 ^ n26278 ;
  assign n26296 = n26295 ^ n26294 ;
  assign n26297 = n26296 ^ n26117 ;
  assign n26298 = n26270 & n26297 ;
  assign n26299 = n26298 ^ n26295 ;
  assign n26484 = n26483 ^ n26299 ;
  assign n26485 = n26484 ^ n26281 ;
  assign n26291 = n26282 ^ n26098 ;
  assign n26292 = n26287 & ~n26291 ;
  assign n26486 = n26485 ^ n26292 ;
  assign n26290 = n26085 & ~n26288 ;
  assign n26487 = n26486 ^ n26290 ;
  assign n26674 = n26484 ^ n26285 ;
  assign n26675 = n26484 ^ n26105 ;
  assign n26676 = n26675 ^ n26098 ;
  assign n26677 = n26676 ^ n26108 ;
  assign n26678 = n26677 ^ n26675 ;
  assign n26679 = n26484 ^ n26098 ;
  assign n26680 = n26679 ^ n26675 ;
  assign n26681 = n26678 & n26680 ;
  assign n26682 = n26681 ^ n26675 ;
  assign n26683 = n26674 & n26682 ;
  assign n26684 = n26683 ^ n26285 ;
  assign n26685 = n26484 ^ n26108 ;
  assign n26686 = ~n26679 & n26685 ;
  assign n26687 = ~n26675 & n26686 ;
  assign n26688 = n26687 ^ n26675 ;
  assign n26689 = n26688 ^ n26105 ;
  assign n26690 = ~n26280 & n26689 ;
  assign n26691 = ~n26684 & ~n26690 ;
  assign n26670 = n26483 ^ n26294 ;
  assign n26671 = n26299 & n26670 ;
  assign n26672 = n26671 ^ n26294 ;
  assign n26664 = n8144 ^ x8 ;
  assign n26657 = n25282 ^ n8144 ;
  assign n26658 = n26657 ^ n8144 ;
  assign n26659 = n8484 ^ n8144 ;
  assign n26660 = n26659 ^ n8144 ;
  assign n26661 = n26658 & n26660 ;
  assign n26662 = n26661 ^ n8144 ;
  assign n26663 = ~n24841 & n26662 ;
  assign n26665 = n26664 ^ n26663 ;
  assign n26655 = n8150 & n25311 ;
  assign n26654 = n8139 & ~n25282 ;
  assign n26656 = n26655 ^ n26654 ;
  assign n26666 = n26665 ^ n26656 ;
  assign n26643 = n7151 & ~n21212 ;
  assign n26642 = n7148 & n20908 ;
  assign n26644 = n26643 ^ n26642 ;
  assign n26645 = n26644 ^ x11 ;
  assign n26641 = n20240 & n25341 ;
  assign n26646 = n26645 ^ n26641 ;
  assign n26640 = n7142 & n21147 ;
  assign n26647 = n26646 ^ n26640 ;
  assign n26618 = ~n6529 & ~n20613 ;
  assign n26617 = ~n6547 & ~n20614 ;
  assign n26619 = n26618 ^ n26617 ;
  assign n26620 = n26619 ^ n6537 ;
  assign n26621 = n26620 ^ x14 ;
  assign n26622 = n26619 ^ x14 ;
  assign n26627 = n26622 ^ n6539 ;
  assign n26623 = n20612 ^ n17173 ;
  assign n26624 = n26623 ^ n23892 ;
  assign n26625 = n26624 ^ n26623 ;
  assign n26626 = n26622 & ~n26625 ;
  assign n26628 = n26627 ^ n26626 ;
  assign n26629 = n26623 ^ n20612 ;
  assign n26630 = ~n26625 & ~n26629 ;
  assign n26631 = n26630 ^ n20612 ;
  assign n26632 = ~n26627 & n26631 ;
  assign n26633 = ~n26628 & n26632 ;
  assign n26634 = n26633 ^ n26630 ;
  assign n26635 = n26634 ^ n6539 ;
  assign n26636 = n26635 ^ n20612 ;
  assign n26637 = ~n26621 & ~n26636 ;
  assign n26607 = n26433 ^ n26420 ;
  assign n26608 = ~n26425 & ~n26607 ;
  assign n26609 = n26608 ^ n26420 ;
  assign n26599 = ~x16 & ~n23490 ;
  assign n26602 = n26599 ^ n23491 ;
  assign n26603 = n6147 & n26602 ;
  assign n26596 = n6143 & ~n20620 ;
  assign n26595 = n20437 & n20624 ;
  assign n26597 = n26596 ^ n26595 ;
  assign n26598 = n26597 ^ x17 ;
  assign n26600 = n26599 ^ n20617 ;
  assign n26601 = n26598 & n26600 ;
  assign n26604 = n26603 ^ n26601 ;
  assign n26605 = n26597 ^ n6145 ;
  assign n26606 = ~n26604 & ~n26605 ;
  assign n26610 = n26609 ^ n26606 ;
  assign n26592 = n5426 & ~n20628 ;
  assign n26590 = n13433 & n20819 ;
  assign n26583 = n22979 ^ x20 ;
  assign n26584 = n26583 ^ x19 ;
  assign n26585 = n26584 ^ n22979 ;
  assign n26586 = ~n22978 & ~n26585 ;
  assign n26587 = n26586 ^ n22979 ;
  assign n26588 = n5215 & ~n26587 ;
  assign n26589 = n26588 ^ x20 ;
  assign n26591 = n26590 ^ n26589 ;
  assign n26593 = n26592 ^ n26591 ;
  assign n26572 = n4655 & n20631 ;
  assign n26571 = n4651 & ~n20683 ;
  assign n26573 = n26572 ^ n26571 ;
  assign n26574 = n26573 ^ x23 ;
  assign n26570 = n4656 & ~n22653 ;
  assign n26575 = n26574 ^ n26570 ;
  assign n26569 = ~n40 & n20680 ;
  assign n26576 = n26575 ^ n26569 ;
  assign n26561 = n3837 & ~n20706 ;
  assign n26559 = n3985 & ~n20705 ;
  assign n26555 = n5065 & ~n22078 ;
  assign n26556 = n26555 ^ n20702 ;
  assign n26557 = n3833 & ~n26556 ;
  assign n26558 = n26557 ^ x29 ;
  assign n26560 = n26559 ^ n26558 ;
  assign n26562 = n26561 ^ n26560 ;
  assign n26549 = ~n4435 & n21246 ;
  assign n26547 = ~n4434 & ~n20690 ;
  assign n26544 = n4600 & ~n20693 ;
  assign n26543 = n20603 & ~n20694 ;
  assign n26545 = n26544 ^ n26543 ;
  assign n26546 = n26545 ^ x26 ;
  assign n26548 = n26547 ^ n26546 ;
  assign n26550 = n26549 ^ n26548 ;
  assign n26539 = n26398 ^ n26175 ;
  assign n26540 = n26400 & ~n26539 ;
  assign n26532 = n4082 ^ n779 ;
  assign n26531 = n1906 ^ n485 ;
  assign n26533 = n26532 ^ n26531 ;
  assign n26534 = n26533 ^ n14277 ;
  assign n26526 = n2028 ^ n918 ;
  assign n26527 = n26526 ^ n584 ;
  assign n26525 = n667 ^ n637 ;
  assign n26528 = n26527 ^ n26525 ;
  assign n26524 = n3203 ^ n3098 ;
  assign n26529 = n26528 ^ n26524 ;
  assign n26530 = n26529 ^ n5584 ;
  assign n26535 = n26534 ^ n26530 ;
  assign n26536 = n26535 ^ n1431 ;
  assign n26537 = n26536 ^ n2746 ;
  assign n26538 = ~n1599 & ~n26537 ;
  assign n26541 = n26540 ^ n26538 ;
  assign n26495 = n20803 ^ n20713 ;
  assign n26496 = ~n52 & n26495 ;
  assign n26514 = n3803 & n20716 ;
  assign n26517 = n26496 & n26514 ;
  assign n26502 = n26367 ^ n20716 ;
  assign n26503 = n26502 ^ n26367 ;
  assign n26508 = n3518 & n26495 ;
  assign n26509 = ~n26503 & n26508 ;
  assign n26510 = n26509 ^ n26503 ;
  assign n26511 = n26510 ^ n26502 ;
  assign n26512 = x31 & n26511 ;
  assign n26497 = n20716 ^ n61 ;
  assign n26498 = n26497 ^ n20716 ;
  assign n26499 = n22188 & n26498 ;
  assign n26500 = n26499 ^ n20716 ;
  assign n26501 = ~n3800 & n26500 ;
  assign n26513 = n26512 ^ n26501 ;
  assign n26515 = n26514 ^ n26513 ;
  assign n26518 = n26517 ^ n26515 ;
  assign n26520 = n26518 ^ n26372 ;
  assign n26519 = n26518 ^ n26403 ;
  assign n26521 = n26520 ^ n26519 ;
  assign n26522 = ~n26377 & ~n26521 ;
  assign n26523 = n26522 ^ n26520 ;
  assign n26542 = n26541 ^ n26523 ;
  assign n26551 = n26550 ^ n26542 ;
  assign n26563 = n26562 ^ n26551 ;
  assign n26564 = n26563 ^ n26404 ;
  assign n26565 = n26564 ^ n26348 ;
  assign n26566 = n26565 ^ n26563 ;
  assign n26567 = n26409 & ~n26566 ;
  assign n26568 = n26567 ^ n26564 ;
  assign n26577 = n26576 ^ n26568 ;
  assign n26578 = n26577 ^ n26419 ;
  assign n26579 = n26578 ^ n26326 ;
  assign n26580 = n26579 ^ n26577 ;
  assign n26581 = n26411 & n26580 ;
  assign n26582 = n26581 ^ n26578 ;
  assign n26594 = n26593 ^ n26582 ;
  assign n26611 = n26610 ^ n26594 ;
  assign n26612 = n26611 ^ n26446 ;
  assign n26613 = n26612 ^ n26437 ;
  assign n26614 = n26613 ^ n26611 ;
  assign n26615 = ~n26438 & ~n26614 ;
  assign n26616 = n26615 ^ n26612 ;
  assign n26638 = n26637 ^ n26616 ;
  assign n26492 = n26467 ^ n26323 ;
  assign n26493 = ~n26448 & ~n26492 ;
  assign n26494 = n26493 ^ n26467 ;
  assign n26639 = n26638 ^ n26494 ;
  assign n26648 = n26647 ^ n26639 ;
  assign n26650 = n26648 ^ n26468 ;
  assign n26649 = n26648 ^ n26481 ;
  assign n26651 = n26650 ^ n26649 ;
  assign n26652 = n26473 & ~n26651 ;
  assign n26653 = n26652 ^ n26650 ;
  assign n26667 = n26666 ^ n26653 ;
  assign n26668 = n26667 ^ x5 ;
  assign n26489 = n26482 ^ n26315 ;
  assign n26490 = n26320 & ~n26489 ;
  assign n26491 = n26490 ^ n26315 ;
  assign n26669 = n26668 ^ n26491 ;
  assign n26673 = n26672 ^ n26669 ;
  assign n26692 = n26691 ^ n26673 ;
  assign n26488 = n26290 & ~n26486 ;
  assign n26693 = n26692 ^ n26488 ;
  assign n26871 = n26672 ^ n26488 ;
  assign n26872 = n26673 & ~n26871 ;
  assign n26869 = n26673 ^ n26488 ;
  assign n26870 = n26691 & ~n26869 ;
  assign n26873 = n26872 ^ n26870 ;
  assign n26694 = n26667 ^ n26491 ;
  assign n26860 = n26666 ^ n26648 ;
  assign n26861 = n26653 & ~n26860 ;
  assign n26862 = n26861 ^ n26648 ;
  assign n26857 = n8150 & n25515 ;
  assign n26853 = n8144 ^ n8139 ;
  assign n26854 = n26853 ^ n26301 ;
  assign n26855 = n25282 & n26854 ;
  assign n26856 = n26855 ^ n26664 ;
  assign n26858 = n26857 ^ n26856 ;
  assign n26846 = n7151 & n24841 ;
  assign n26845 = n7148 & n21147 ;
  assign n26847 = n26846 ^ n26845 ;
  assign n26848 = n26847 ^ x11 ;
  assign n26844 = n20240 & ~n25528 ;
  assign n26849 = n26848 ^ n26844 ;
  assign n26843 = n7142 & ~n21212 ;
  assign n26850 = n26849 ^ n26843 ;
  assign n26838 = n20437 & ~n20620 ;
  assign n26836 = n6163 & n23480 ;
  assign n26833 = n6148 & ~n20614 ;
  assign n26832 = n6143 & ~n20617 ;
  assign n26834 = n26833 ^ n26832 ;
  assign n26835 = n26834 ^ x17 ;
  assign n26837 = n26836 ^ n26835 ;
  assign n26839 = n26838 ^ n26837 ;
  assign n26827 = n26593 ^ n26577 ;
  assign n26828 = ~n26582 & ~n26827 ;
  assign n26829 = n26828 ^ n26577 ;
  assign n26823 = n4656 & ~n21237 ;
  assign n26821 = n4655 & n20819 ;
  assign n26819 = n4651 & n20680 ;
  assign n26815 = n26576 ^ n26563 ;
  assign n26816 = ~n26568 & ~n26815 ;
  assign n26817 = n26816 ^ n26563 ;
  assign n26818 = n26817 ^ x23 ;
  assign n26820 = n26819 ^ n26818 ;
  assign n26822 = n26821 ^ n26820 ;
  assign n26824 = n26823 ^ n26822 ;
  assign n26814 = ~n40 & n20631 ;
  assign n26825 = n26824 ^ n26814 ;
  assign n26799 = n611 ^ n511 ;
  assign n26800 = n26799 ^ n563 ;
  assign n26797 = n657 ^ n211 ;
  assign n26798 = n26797 ^ n459 ;
  assign n26801 = n26800 ^ n26798 ;
  assign n26796 = n5495 ^ n5343 ;
  assign n26802 = n26801 ^ n26796 ;
  assign n26793 = n3880 ^ n995 ;
  assign n26794 = n26793 ^ n2965 ;
  assign n26795 = n26794 ^ n12882 ;
  assign n26803 = n26802 ^ n26795 ;
  assign n26804 = n26803 ^ n21674 ;
  assign n26805 = n26804 ^ n4149 ;
  assign n26806 = ~n2499 & ~n26805 ;
  assign n26807 = n26806 ^ x5 ;
  assign n26785 = x30 & n24604 ;
  assign n26786 = n26785 ^ n20706 ;
  assign n26787 = ~n3518 & ~n26786 ;
  assign n26788 = n26787 ^ n20706 ;
  assign n26789 = n26788 ^ n21782 ;
  assign n26776 = n21782 ^ n20716 ;
  assign n26775 = n21782 ^ n20713 ;
  assign n26777 = n26776 ^ n26775 ;
  assign n26780 = ~x30 & n26777 ;
  assign n26781 = n26780 ^ n26776 ;
  assign n26782 = ~n3518 & n26781 ;
  assign n26790 = n26789 ^ n26782 ;
  assign n26791 = x31 & ~n26790 ;
  assign n26792 = n26791 ^ n26788 ;
  assign n26808 = n26807 ^ n26792 ;
  assign n26760 = n26398 & ~n26401 ;
  assign n26761 = n26538 & n26760 ;
  assign n26809 = n26808 ^ n26761 ;
  assign n26773 = n3837 & ~n20705 ;
  assign n26771 = n3985 & ~n20702 ;
  assign n26764 = n20694 ^ x29 ;
  assign n26765 = n26764 ^ x28 ;
  assign n26766 = n26765 ^ n20694 ;
  assign n26767 = ~n22112 & n26766 ;
  assign n26768 = n26767 ^ n20694 ;
  assign n26769 = n3833 & ~n26768 ;
  assign n26770 = n26769 ^ x29 ;
  assign n26772 = n26771 ^ n26770 ;
  assign n26774 = n26773 ^ n26772 ;
  assign n26810 = n26809 ^ n26774 ;
  assign n26758 = ~n26398 & n26401 ;
  assign n26759 = ~n26538 & n26758 ;
  assign n26762 = n26761 ^ n26759 ;
  assign n26763 = ~x2 & n26762 ;
  assign n26811 = n26810 ^ n26763 ;
  assign n26755 = n26541 ^ n26518 ;
  assign n26756 = n26523 & ~n26755 ;
  assign n26757 = n26756 ^ n26518 ;
  assign n26812 = n26811 ^ n26757 ;
  assign n26729 = n4600 & ~n20690 ;
  assign n26728 = n20603 & ~n20693 ;
  assign n26730 = n26729 ^ n26728 ;
  assign n26731 = n26730 ^ n97 ;
  assign n26732 = n26730 ^ x26 ;
  assign n26733 = n26732 ^ n99 ;
  assign n26734 = n26733 ^ x25 ;
  assign n26735 = n26734 ^ n20683 ;
  assign n26736 = n26735 ^ n26732 ;
  assign n26737 = n26736 ^ n22617 ;
  assign n26738 = n26737 ^ n26736 ;
  assign n26739 = n26732 & ~n26738 ;
  assign n26740 = n26739 ^ n26733 ;
  assign n26741 = n26736 ^ n20683 ;
  assign n26742 = ~n26738 & ~n26741 ;
  assign n26743 = n26742 ^ n20683 ;
  assign n26744 = ~n26733 & n26743 ;
  assign n26745 = ~n26740 & n26744 ;
  assign n26746 = n26745 ^ n26742 ;
  assign n26747 = n26746 ^ n99 ;
  assign n26748 = n26747 ^ n20683 ;
  assign n26749 = ~n26731 & ~n26748 ;
  assign n26750 = n26749 ^ n26562 ;
  assign n26751 = n26750 ^ n26550 ;
  assign n26752 = n26751 ^ n26749 ;
  assign n26753 = n26551 & n26752 ;
  assign n26754 = n26753 ^ n26750 ;
  assign n26813 = n26812 ^ n26754 ;
  assign n26826 = n26825 ^ n26813 ;
  assign n26830 = n26829 ^ n26826 ;
  assign n26724 = ~x20 & n21231 ;
  assign n26723 = n13433 & ~n20628 ;
  assign n26725 = n26724 ^ n26723 ;
  assign n26721 = ~n5218 & ~n21231 ;
  assign n26720 = n5217 & n20624 ;
  assign n26722 = n26721 ^ n26720 ;
  assign n26726 = n26725 ^ n26722 ;
  assign n26718 = n5216 & ~n21232 ;
  assign n26717 = n5426 & n20829 ;
  assign n26719 = n26718 ^ n26717 ;
  assign n26727 = n26726 ^ n26719 ;
  assign n26831 = n26830 ^ n26727 ;
  assign n26840 = n26839 ^ n26831 ;
  assign n26714 = n26609 ^ n26594 ;
  assign n26715 = n26610 & n26714 ;
  assign n26716 = n26715 ^ n26609 ;
  assign n26841 = n26840 ^ n26716 ;
  assign n26704 = ~n6529 & ~n20612 ;
  assign n26703 = ~n6547 & ~n20613 ;
  assign n26705 = n26704 ^ n26703 ;
  assign n26706 = n26705 ^ x14 ;
  assign n26698 = ~x13 & ~n24096 ;
  assign n26699 = n26698 ^ n20908 ;
  assign n26702 = n6537 & n26699 ;
  assign n26707 = n26706 ^ n26702 ;
  assign n26700 = n26699 ^ n24096 ;
  assign n26701 = n6539 & ~n26700 ;
  assign n26708 = n26707 ^ n26701 ;
  assign n26710 = n26708 ^ n26611 ;
  assign n26709 = n26708 ^ n26637 ;
  assign n26711 = n26710 ^ n26709 ;
  assign n26712 = ~n26616 & n26711 ;
  assign n26713 = n26712 ^ n26710 ;
  assign n26842 = n26841 ^ n26713 ;
  assign n26851 = n26850 ^ n26842 ;
  assign n26695 = n26647 ^ n26494 ;
  assign n26696 = n26639 & ~n26695 ;
  assign n26697 = n26696 ^ n26647 ;
  assign n26852 = n26851 ^ n26697 ;
  assign n26859 = n26858 ^ n26852 ;
  assign n26863 = n26862 ^ n26859 ;
  assign n26864 = n26863 ^ x5 ;
  assign n26865 = n26864 ^ n26491 ;
  assign n26866 = n26865 ^ n26863 ;
  assign n26867 = n26694 & ~n26866 ;
  assign n26868 = n26867 ^ n26864 ;
  assign n26874 = n26873 ^ n26868 ;
  assign n27056 = ~n26491 & n26667 ;
  assign n27065 = n27056 ^ n26863 ;
  assign n27057 = n26863 & ~n27056 ;
  assign n27066 = n27065 ^ n27057 ;
  assign n27058 = n26691 ^ x5 ;
  assign n27059 = n26691 ^ n26672 ;
  assign n27062 = ~n27058 & ~n27059 ;
  assign n27063 = n27062 ^ n26691 ;
  assign n27064 = ~n27057 & ~n27063 ;
  assign n27067 = n27066 ^ n27064 ;
  assign n27068 = n27056 ^ n26694 ;
  assign n27069 = n26863 ^ n26672 ;
  assign n27070 = n27058 & n27059 ;
  assign n27071 = ~n27069 & n27070 ;
  assign n27072 = n27071 ^ n26863 ;
  assign n27073 = ~n27068 & ~n27072 ;
  assign n27074 = ~n27067 & ~n27073 ;
  assign n27052 = n20240 & n25868 ;
  assign n27050 = n7148 & ~n21212 ;
  assign n27046 = n7151 & n25282 ;
  assign n27047 = n27046 ^ n7151 ;
  assign n27045 = n7142 & n24841 ;
  assign n27048 = n27047 ^ n27045 ;
  assign n27049 = n27048 ^ x11 ;
  assign n27051 = n27050 ^ n27049 ;
  assign n27053 = n27052 ^ n27051 ;
  assign n27038 = n20908 ^ x14 ;
  assign n27028 = n21147 ^ x13 ;
  assign n27029 = n27028 ^ x14 ;
  assign n27030 = n27029 ^ n21147 ;
  assign n27031 = n24078 & n27030 ;
  assign n27032 = n27031 ^ n27028 ;
  assign n27039 = n27038 ^ n27032 ;
  assign n27033 = n20908 ^ n7310 ;
  assign n27034 = n27033 ^ n20908 ;
  assign n27035 = ~n24085 & n27034 ;
  assign n27036 = n27035 ^ n20908 ;
  assign n27037 = ~n6540 & n27036 ;
  assign n27040 = n27039 ^ n27037 ;
  assign n27041 = ~n6391 & n27040 ;
  assign n27042 = n27041 ^ n27032 ;
  assign n27024 = n26839 ^ n26716 ;
  assign n27025 = n26840 & ~n27024 ;
  assign n27026 = n27025 ^ n26839 ;
  assign n27018 = n6148 & ~n20613 ;
  assign n27017 = n6143 & ~n20614 ;
  assign n27019 = n27018 ^ n27017 ;
  assign n27020 = n27019 ^ x17 ;
  assign n27016 = n6163 & n21227 ;
  assign n27021 = n27020 ^ n27016 ;
  assign n27015 = n20437 & ~n20617 ;
  assign n27022 = n27021 ^ n27015 ;
  assign n27011 = n13433 & n20829 ;
  assign n27009 = n5426 & n20624 ;
  assign n27002 = n20620 ^ x20 ;
  assign n27003 = n27002 ^ x19 ;
  assign n27004 = n27003 ^ n20620 ;
  assign n27005 = ~n22963 & n27004 ;
  assign n27006 = n27005 ^ n20620 ;
  assign n27007 = n5215 & ~n27006 ;
  assign n27008 = n27007 ^ x20 ;
  assign n27010 = n27009 ^ n27008 ;
  assign n27012 = n27011 ^ n27010 ;
  assign n26995 = n4655 & ~n20628 ;
  assign n26994 = n4651 & n20631 ;
  assign n26996 = n26995 ^ n26994 ;
  assign n26997 = n26996 ^ x23 ;
  assign n26993 = n4656 & n23307 ;
  assign n26998 = n26997 ^ n26993 ;
  assign n26992 = ~n40 & n20819 ;
  assign n26999 = n26998 ^ n26992 ;
  assign n26988 = ~n4435 & ~n22662 ;
  assign n26986 = ~n4434 & n20680 ;
  assign n26983 = n4600 & ~n20683 ;
  assign n26982 = n20603 & ~n20690 ;
  assign n26984 = n26983 ^ n26982 ;
  assign n26985 = n26984 ^ x26 ;
  assign n26987 = n26986 ^ n26985 ;
  assign n26989 = n26988 ^ n26987 ;
  assign n26969 = x30 & ~n20706 ;
  assign n26955 = n21770 ^ n20706 ;
  assign n26954 = n21770 ^ n20713 ;
  assign n26956 = n26955 ^ n26954 ;
  assign n26957 = n26955 ^ x30 ;
  assign n26958 = n26957 ^ n26955 ;
  assign n26959 = ~n26956 & n26958 ;
  assign n26960 = n26959 ^ n26955 ;
  assign n26961 = ~n3518 & ~n26960 ;
  assign n26962 = n26961 ^ n21770 ;
  assign n26963 = n26962 ^ n20705 ;
  assign n26964 = n26963 ^ n26962 ;
  assign n26970 = n26969 ^ n26964 ;
  assign n26971 = ~n3518 & ~n26970 ;
  assign n26972 = n26971 ^ n26963 ;
  assign n26973 = ~x31 & ~n26972 ;
  assign n26974 = n26973 ^ n26962 ;
  assign n26951 = n6053 & ~n26807 ;
  assign n26952 = n26951 ^ x2 ;
  assign n26945 = n6246 ^ n1653 ;
  assign n26946 = n26945 ^ n2035 ;
  assign n26943 = n2593 ^ n1992 ;
  assign n26944 = n26943 ^ n6909 ;
  assign n26947 = n26946 ^ n26944 ;
  assign n26939 = n12522 ^ n520 ;
  assign n26938 = n710 ^ n237 ;
  assign n26940 = n26939 ^ n26938 ;
  assign n26941 = n26940 ^ n12534 ;
  assign n26942 = n26941 ^ n1174 ;
  assign n26948 = n26947 ^ n26942 ;
  assign n26933 = n3080 ^ n637 ;
  assign n26932 = n884 ^ n668 ;
  assign n26934 = n26933 ^ n26932 ;
  assign n26931 = n6042 ^ n4085 ;
  assign n26935 = n26934 ^ n26931 ;
  assign n26936 = n26935 ^ n2180 ;
  assign n26926 = n247 ^ n189 ;
  assign n26927 = n26926 ^ n6936 ;
  assign n26928 = n26927 ^ n12626 ;
  assign n26929 = n26928 ^ n1686 ;
  assign n26925 = n4159 ^ n888 ;
  assign n26930 = n26929 ^ n26925 ;
  assign n26937 = n26936 ^ n26930 ;
  assign n26949 = n26948 ^ n26937 ;
  assign n26950 = ~n1383 & ~n26949 ;
  assign n26953 = n26952 ^ n26950 ;
  assign n26975 = n26974 ^ n26953 ;
  assign n26917 = n3837 & ~n20702 ;
  assign n26915 = n3985 & ~n20694 ;
  assign n26908 = n20693 ^ x29 ;
  assign n26909 = n26908 ^ x28 ;
  assign n26910 = n26909 ^ n20693 ;
  assign n26911 = ~n22092 & n26910 ;
  assign n26912 = n26911 ^ n20693 ;
  assign n26913 = n3833 & ~n26912 ;
  assign n26914 = n26913 ^ x29 ;
  assign n26916 = n26915 ^ n26914 ;
  assign n26918 = n26917 ^ n26916 ;
  assign n26919 = n26918 ^ n26792 ;
  assign n26901 = n26807 ^ n26759 ;
  assign n26900 = n26792 ^ n26761 ;
  assign n26902 = n26901 ^ n26900 ;
  assign n26903 = ~n26762 & n26902 ;
  assign n26904 = n26903 ^ n26900 ;
  assign n26905 = n26807 ^ x2 ;
  assign n26906 = n26905 ^ n26792 ;
  assign n26907 = n26904 & n26906 ;
  assign n26920 = n26919 ^ n26907 ;
  assign n26976 = n26975 ^ n26920 ;
  assign n26977 = n26976 ^ n26774 ;
  assign n26978 = n26977 ^ n26757 ;
  assign n26979 = n26978 ^ n26976 ;
  assign n26980 = n26811 & n26979 ;
  assign n26981 = n26980 ^ n26977 ;
  assign n26990 = n26989 ^ n26981 ;
  assign n26897 = n26812 ^ n26749 ;
  assign n26898 = ~n26754 & ~n26897 ;
  assign n26899 = n26898 ^ n26749 ;
  assign n26991 = n26990 ^ n26899 ;
  assign n27000 = n26999 ^ n26991 ;
  assign n26894 = n26817 ^ n26813 ;
  assign n26895 = ~n26825 & n26894 ;
  assign n26896 = n26895 ^ n26817 ;
  assign n27001 = n27000 ^ n26896 ;
  assign n27013 = n27012 ^ n27001 ;
  assign n26891 = n26829 ^ n26727 ;
  assign n26892 = ~n26830 & n26891 ;
  assign n26893 = n26892 ^ n26829 ;
  assign n27014 = n27013 ^ n26893 ;
  assign n27023 = n27022 ^ n27014 ;
  assign n27027 = n27026 ^ n27023 ;
  assign n27043 = n27042 ^ n27027 ;
  assign n26888 = n26841 ^ n26708 ;
  assign n26889 = ~n26713 & ~n26888 ;
  assign n26890 = n26889 ^ n26708 ;
  assign n27044 = n27043 ^ n26890 ;
  assign n27054 = n27053 ^ n27044 ;
  assign n26885 = n8144 & n25308 ;
  assign n26886 = n26885 ^ x8 ;
  assign n26882 = n26842 ^ n26697 ;
  assign n26883 = n26851 & ~n26882 ;
  assign n26884 = n26883 ^ n26850 ;
  assign n26887 = n26886 ^ n26884 ;
  assign n27055 = n27054 ^ n26887 ;
  assign n27075 = n27074 ^ n27055 ;
  assign n26878 = n26488 & n26692 ;
  assign n26879 = n26868 ^ n26691 ;
  assign n26880 = n26878 & n26879 ;
  assign n26875 = n26862 ^ n26858 ;
  assign n26876 = ~n26859 & ~n26875 ;
  assign n26877 = n26876 ^ n26862 ;
  assign n26881 = n26880 ^ n26877 ;
  assign n27076 = n27075 ^ n26881 ;
  assign n27077 = n27055 ^ n26877 ;
  assign n27078 = n27077 ^ n27074 ;
  assign n27225 = ~n6547 & n20908 ;
  assign n27224 = ~n6529 & n21147 ;
  assign n27226 = n27225 ^ n27224 ;
  assign n27227 = n27226 ^ n6537 ;
  assign n27228 = n27227 ^ x14 ;
  assign n27244 = ~n17173 & ~n21170 ;
  assign n27230 = n27226 ^ n6538 ;
  assign n27231 = n21212 ^ n17173 ;
  assign n27232 = n27231 ^ n21212 ;
  assign n27233 = ~n25342 & ~n27232 ;
  assign n27234 = n27233 ^ n21212 ;
  assign n27235 = ~n27230 & n27234 ;
  assign n27229 = n21212 ^ n6539 ;
  assign n27236 = n27235 ^ n27229 ;
  assign n27245 = n27244 ^ n27236 ;
  assign n27246 = ~n27228 & ~n27245 ;
  assign n27216 = n20437 & ~n20614 ;
  assign n27214 = n6163 & n23893 ;
  assign n27211 = n6148 & ~n20612 ;
  assign n27210 = n6143 & ~n20613 ;
  assign n27212 = n27211 ^ n27210 ;
  assign n27213 = n27212 ^ x17 ;
  assign n27215 = n27214 ^ n27213 ;
  assign n27217 = n27216 ^ n27215 ;
  assign n27198 = n5426 & ~n20620 ;
  assign n27197 = n5217 & ~n20617 ;
  assign n27199 = n27198 ^ n27197 ;
  assign n27200 = n27199 ^ x20 ;
  assign n27196 = n5216 & n23491 ;
  assign n27201 = n27200 ^ n27196 ;
  assign n27195 = n13433 & n20624 ;
  assign n27202 = n27201 ^ n27195 ;
  assign n27194 = ~n23490 & n27193 ;
  assign n27203 = n27202 ^ n27194 ;
  assign n27185 = ~n40 & ~n20628 ;
  assign n27183 = n4656 & ~n22979 ;
  assign n27180 = n4655 & n20829 ;
  assign n27179 = n4651 & n20819 ;
  assign n27181 = n27180 ^ n27179 ;
  assign n27182 = n27181 ^ x23 ;
  assign n27184 = n27183 ^ n27182 ;
  assign n27186 = n27185 ^ n27184 ;
  assign n27165 = ~x25 & ~n22649 ;
  assign n27168 = n27165 ^ n22653 ;
  assign n27169 = n99 & ~n27168 ;
  assign n27162 = n4600 & n20680 ;
  assign n27161 = n20603 & ~n20683 ;
  assign n27163 = n27162 ^ n27161 ;
  assign n27164 = n27163 ^ x26 ;
  assign n27166 = n27165 ^ n20631 ;
  assign n27167 = n27164 & ~n27166 ;
  assign n27170 = n27169 ^ n27167 ;
  assign n27171 = n27163 ^ n97 ;
  assign n27172 = ~n27170 & ~n27171 ;
  assign n27159 = n3837 & ~n20694 ;
  assign n27157 = n3985 & ~n20693 ;
  assign n27144 = n22079 ^ n20705 ;
  assign n27143 = n22079 ^ n20706 ;
  assign n27145 = n27144 ^ n27143 ;
  assign n27148 = x30 & n27145 ;
  assign n27149 = n27148 ^ n27144 ;
  assign n27150 = ~n3518 & ~n27149 ;
  assign n27151 = n27150 ^ n22079 ;
  assign n27152 = x31 & n27151 ;
  assign n27139 = n26974 ^ n26952 ;
  assign n27140 = ~n26953 & n27139 ;
  assign n27130 = n2732 ^ n468 ;
  assign n27131 = n27130 ^ n905 ;
  assign n27132 = n27131 ^ n547 ;
  assign n27129 = n735 ^ n464 ;
  assign n27133 = n27132 ^ n27129 ;
  assign n27127 = n1424 ^ n1330 ;
  assign n27126 = n1628 ^ n1308 ;
  assign n27128 = n27127 ^ n27126 ;
  assign n27134 = n27133 ^ n27128 ;
  assign n27122 = n788 ^ n524 ;
  assign n27120 = n1754 ^ n117 ;
  assign n27121 = n27120 ^ n1008 ;
  assign n27123 = n27122 ^ n27121 ;
  assign n27124 = n27123 ^ n916 ;
  assign n27125 = n27124 ^ n4153 ;
  assign n27135 = n27134 ^ n27125 ;
  assign n27136 = n27135 ^ n4006 ;
  assign n27115 = n1957 ^ n1162 ;
  assign n27116 = n27115 ^ n1776 ;
  assign n27117 = n27116 ^ n3746 ;
  assign n27118 = n27117 ^ n2959 ;
  assign n27112 = n2428 ^ n750 ;
  assign n27110 = n3677 ^ n575 ;
  assign n27111 = n27110 ^ n3226 ;
  assign n27113 = n27112 ^ n27111 ;
  assign n27109 = n13385 ^ n4770 ;
  assign n27114 = n27113 ^ n27109 ;
  assign n27119 = n27118 ^ n27114 ;
  assign n27137 = n27136 ^ n27119 ;
  assign n27138 = ~n12910 & ~n27137 ;
  assign n27141 = n27140 ^ n27138 ;
  assign n24297 = n20705 ^ n20702 ;
  assign n27106 = ~n61 & n24297 ;
  assign n27107 = n27106 ^ n20702 ;
  assign n27108 = ~n3800 & ~n27107 ;
  assign n27142 = n27141 ^ n27108 ;
  assign n27153 = n27152 ^ n27142 ;
  assign n27100 = n26975 ^ n26918 ;
  assign n27101 = ~n26920 & ~n27100 ;
  assign n27102 = n27101 ^ n26918 ;
  assign n27154 = n27153 ^ n27102 ;
  assign n27155 = n27154 ^ x29 ;
  assign n27095 = n20690 ^ n5065 ;
  assign n27096 = n27095 ^ n20690 ;
  assign n27097 = ~n21247 & n27096 ;
  assign n27098 = n27097 ^ n20690 ;
  assign n27099 = n3833 & ~n27098 ;
  assign n27156 = n27155 ^ n27099 ;
  assign n27158 = n27157 ^ n27156 ;
  assign n27160 = n27159 ^ n27158 ;
  assign n27173 = n27172 ^ n27160 ;
  assign n27175 = n27173 ^ n26976 ;
  assign n27174 = n27173 ^ n26989 ;
  assign n27176 = n27175 ^ n27174 ;
  assign n27177 = n26981 & n27176 ;
  assign n27178 = n27177 ^ n27175 ;
  assign n27187 = n27186 ^ n27178 ;
  assign n27188 = n27187 ^ n26999 ;
  assign n27189 = n27188 ^ n26899 ;
  assign n27190 = n27189 ^ n27187 ;
  assign n27191 = n26991 & ~n27190 ;
  assign n27192 = n27191 ^ n27188 ;
  assign n27204 = n27203 ^ n27192 ;
  assign n27205 = n27204 ^ n27012 ;
  assign n27206 = n27205 ^ n27204 ;
  assign n27207 = n27206 ^ n26896 ;
  assign n27208 = ~n27001 & ~n27207 ;
  assign n27209 = n27208 ^ n27205 ;
  assign n27218 = n27217 ^ n27209 ;
  assign n27219 = n27218 ^ n27022 ;
  assign n27220 = n27219 ^ n27218 ;
  assign n27221 = n27220 ^ n26893 ;
  assign n27222 = n27014 & ~n27221 ;
  assign n27223 = n27222 ^ n27219 ;
  assign n27247 = n27246 ^ n27223 ;
  assign n27092 = n27042 ^ n27026 ;
  assign n27093 = n27027 & n27092 ;
  assign n27094 = n27093 ^ n27042 ;
  assign n27248 = n27247 ^ n27094 ;
  assign n27089 = n27046 ^ n7148 ;
  assign n27090 = ~n24841 & n27089 ;
  assign n27087 = n7148 ^ x11 ;
  assign n27085 = n20240 & n25311 ;
  assign n27084 = n7142 & ~n25282 ;
  assign n27086 = n27085 ^ n27084 ;
  assign n27088 = n27087 ^ n27086 ;
  assign n27091 = n27090 ^ n27088 ;
  assign n27249 = n27248 ^ n27091 ;
  assign n27250 = n27249 ^ x8 ;
  assign n27081 = n27053 ^ n26890 ;
  assign n27082 = n27044 & n27081 ;
  assign n27083 = n27082 ^ n27053 ;
  assign n27251 = n27250 ^ n27083 ;
  assign n27252 = n27251 ^ n27054 ;
  assign n27253 = n27252 ^ n27251 ;
  assign n27254 = n27253 ^ n26884 ;
  assign n27255 = ~n26887 & ~n27254 ;
  assign n27256 = n27255 ^ n27252 ;
  assign n27079 = ~n27055 & ~n27074 ;
  assign n27080 = n27079 ^ n27075 ;
  assign n27257 = n27256 ^ n27080 ;
  assign n27258 = n27257 ^ n26880 ;
  assign n27259 = n27258 ^ n27079 ;
  assign n27260 = n27259 ^ n27256 ;
  assign n27261 = ~n27078 & n27260 ;
  assign n27262 = n27261 ^ n27257 ;
  assign n27439 = n20240 & n25515 ;
  assign n27435 = n7148 ^ n7142 ;
  assign n27436 = n27435 ^ n27045 ;
  assign n27437 = n25282 & n27436 ;
  assign n27438 = n27437 ^ n27087 ;
  assign n27440 = n27439 ^ n27438 ;
  assign n27412 = n26884 ^ n26877 ;
  assign n27411 = ~n26877 & n26884 ;
  assign n27413 = n27412 ^ n27411 ;
  assign n27414 = n27413 ^ n27251 ;
  assign n27415 = n26886 & ~n27054 ;
  assign n27416 = n27415 ^ n26884 ;
  assign n27417 = n27416 ^ n26877 ;
  assign n27418 = n27417 ^ n27415 ;
  assign n27419 = n27054 ^ n26886 ;
  assign n27420 = n27419 ^ n27415 ;
  assign n27421 = n27420 ^ n26884 ;
  assign n27422 = n27421 ^ n27415 ;
  assign n27423 = n27418 & n27422 ;
  assign n27424 = n27423 ^ n27415 ;
  assign n27425 = n27414 & n27424 ;
  assign n27426 = n27425 ^ n27251 ;
  assign n27429 = n27414 & ~n27415 ;
  assign n27427 = n27420 ^ n27251 ;
  assign n27428 = ~n27411 & n27427 ;
  assign n27430 = n27429 ^ n27428 ;
  assign n27431 = ~n27066 & n27430 ;
  assign n27432 = ~n27064 & n27431 ;
  assign n27433 = n27074 & n27432 ;
  assign n27434 = ~n27426 & ~n27433 ;
  assign n27441 = n27440 ^ n27434 ;
  assign n27406 = n27094 ^ n27091 ;
  assign n27407 = n27248 & n27406 ;
  assign n27408 = n27407 ^ n27091 ;
  assign n27403 = n27249 ^ n27083 ;
  assign n27404 = ~n27250 & n27403 ;
  assign n27405 = n27404 ^ x8 ;
  assign n27409 = n27408 ^ n27405 ;
  assign n27399 = n20437 & ~n20613 ;
  assign n27391 = n27203 ^ n27187 ;
  assign n27392 = n27192 & n27391 ;
  assign n27393 = n27392 ^ n27187 ;
  assign n27388 = n5426 & ~n20617 ;
  assign n27386 = n13433 & ~n20620 ;
  assign n27379 = n20614 ^ x20 ;
  assign n27380 = n27379 ^ x19 ;
  assign n27381 = n27380 ^ n20614 ;
  assign n27382 = ~n23479 & n27381 ;
  assign n27383 = n27382 ^ n20614 ;
  assign n27384 = n5215 & ~n27383 ;
  assign n27385 = n27384 ^ x20 ;
  assign n27387 = n27386 ^ n27385 ;
  assign n27389 = n27388 ^ n27387 ;
  assign n27372 = n4655 & n20624 ;
  assign n27371 = n4651 & ~n20628 ;
  assign n27373 = n27372 ^ n27371 ;
  assign n27374 = n27373 ^ x23 ;
  assign n27370 = n4656 & ~n21232 ;
  assign n27375 = n27374 ^ n27370 ;
  assign n27369 = ~n40 & n20829 ;
  assign n27376 = n27375 ^ n27369 ;
  assign n27365 = n27186 ^ n27173 ;
  assign n27366 = n27178 & n27365 ;
  assign n27367 = n27366 ^ n27173 ;
  assign n27361 = ~n4435 & ~n21237 ;
  assign n27359 = ~n4434 & n20819 ;
  assign n27356 = n4600 & n20631 ;
  assign n27355 = n20603 & n20680 ;
  assign n27357 = n27356 ^ n27355 ;
  assign n27358 = n27357 ^ x26 ;
  assign n27360 = n27359 ^ n27358 ;
  assign n27362 = n27361 ^ n27360 ;
  assign n27350 = n3985 & ~n20690 ;
  assign n27343 = n20683 ^ x29 ;
  assign n27344 = n27343 ^ x28 ;
  assign n27345 = n27344 ^ n20683 ;
  assign n27346 = ~n22617 & n27345 ;
  assign n27347 = n27346 ^ n20683 ;
  assign n27348 = n3833 & ~n27347 ;
  assign n27349 = n27348 ^ x29 ;
  assign n27351 = n27350 ^ n27349 ;
  assign n27342 = n3837 & ~n20693 ;
  assign n27352 = n27351 ^ n27342 ;
  assign n27332 = n12850 ^ n12828 ;
  assign n27330 = n799 ^ n355 ;
  assign n27331 = n27330 ^ n2184 ;
  assign n27333 = n27332 ^ n27331 ;
  assign n27328 = n14289 ^ n2951 ;
  assign n27327 = n1313 ^ n1178 ;
  assign n27329 = n27328 ^ n27327 ;
  assign n27334 = n27333 ^ n27329 ;
  assign n27335 = n27334 ^ n3076 ;
  assign n27336 = n6054 ^ n2688 ;
  assign n27337 = n27336 ^ n882 ;
  assign n27338 = ~n27335 & ~n27337 ;
  assign n27339 = n27338 ^ n26950 ;
  assign n27340 = n27339 ^ x8 ;
  assign n27303 = n22601 ^ n20702 ;
  assign n27302 = n22601 ^ n20705 ;
  assign n27304 = n27303 ^ n27302 ;
  assign n27305 = n27303 ^ x30 ;
  assign n27306 = n27305 ^ n27303 ;
  assign n27307 = n27304 & n27306 ;
  assign n27308 = n27307 ^ n27303 ;
  assign n27309 = ~n3518 & ~n27308 ;
  assign n27310 = n27309 ^ n22601 ;
  assign n27300 = ~n61 & n20702 ;
  assign n27301 = n27300 ^ x29 ;
  assign n27311 = n27310 ^ n27301 ;
  assign n27312 = n27311 ^ n20694 ;
  assign n27313 = n27312 ^ x30 ;
  assign n27314 = n27313 ^ n27311 ;
  assign n27315 = n27311 ^ x29 ;
  assign n27316 = n27315 ^ n20694 ;
  assign n27317 = n27316 ^ n27311 ;
  assign n27318 = n27314 & ~n27317 ;
  assign n27319 = n27318 ^ n27311 ;
  assign n27320 = ~x31 & n27319 ;
  assign n27321 = n27320 ^ n27310 ;
  assign n27322 = n27321 ^ n26950 ;
  assign n27323 = n27322 ^ n27138 ;
  assign n27324 = n27323 ^ n27321 ;
  assign n27325 = n27140 & ~n27324 ;
  assign n27326 = n27325 ^ n27322 ;
  assign n27341 = n27340 ^ n27326 ;
  assign n27353 = n27352 ^ n27341 ;
  assign n27297 = n27141 ^ n27102 ;
  assign n27298 = ~n27153 & ~n27297 ;
  assign n27299 = n27298 ^ n27141 ;
  assign n27354 = n27353 ^ n27299 ;
  assign n27363 = n27362 ^ n27354 ;
  assign n27294 = n27172 ^ n27154 ;
  assign n27295 = n27160 & n27294 ;
  assign n27296 = n27295 ^ n27172 ;
  assign n27364 = n27363 ^ n27296 ;
  assign n27368 = n27367 ^ n27364 ;
  assign n27377 = n27376 ^ n27368 ;
  assign n27390 = n27389 ^ n27377 ;
  assign n27394 = n27393 ^ n27390 ;
  assign n27395 = n27394 ^ x17 ;
  assign n27293 = n6148 & n20908 ;
  assign n27396 = n27395 ^ n27293 ;
  assign n27292 = n6143 & ~n20612 ;
  assign n27397 = n27396 ^ n27292 ;
  assign n27291 = n6163 & ~n25056 ;
  assign n27398 = n27397 ^ n27291 ;
  assign n27400 = n27399 ^ n27398 ;
  assign n27288 = n27217 ^ n27204 ;
  assign n27289 = n27209 & n27288 ;
  assign n27290 = n27289 ^ n27204 ;
  assign n27401 = n27400 ^ n27290 ;
  assign n27267 = ~n6529 & ~n21212 ;
  assign n27266 = ~n6547 & n21147 ;
  assign n27268 = n27267 ^ n27266 ;
  assign n27269 = n27268 ^ n6537 ;
  assign n27270 = n27269 ^ x14 ;
  assign n27280 = n6539 & n24810 ;
  assign n27271 = n27268 ^ n6538 ;
  assign n27272 = n25528 ^ n24841 ;
  assign n27275 = n24841 ^ x13 ;
  assign n27276 = n27275 ^ n24841 ;
  assign n27277 = ~n27272 & ~n27276 ;
  assign n27278 = n27277 ^ n24841 ;
  assign n27279 = n27271 & ~n27278 ;
  assign n27281 = n27280 ^ n27279 ;
  assign n27282 = ~n27270 & ~n27281 ;
  assign n27284 = n27282 ^ n27218 ;
  assign n27283 = n27282 ^ n27246 ;
  assign n27285 = n27284 ^ n27283 ;
  assign n27286 = n27223 & ~n27285 ;
  assign n27287 = n27286 ^ n27284 ;
  assign n27402 = n27401 ^ n27287 ;
  assign n27410 = n27409 ^ n27402 ;
  assign n27442 = n27441 ^ n27410 ;
  assign n27263 = n26880 & ~n27078 ;
  assign n27264 = n27256 ^ n27079 ;
  assign n27265 = n27263 & n27264 ;
  assign n27443 = n27442 ^ n27265 ;
  assign n27594 = n27265 & n27442 ;
  assign n27591 = n27405 ^ n27402 ;
  assign n27592 = ~n27409 & ~n27591 ;
  assign n27584 = n27401 ^ n27282 ;
  assign n27585 = ~n27287 & n27584 ;
  assign n27586 = n27585 ^ n27282 ;
  assign n27587 = n27586 ^ x11 ;
  assign n27583 = n7148 & n25308 ;
  assign n27588 = n27587 ^ n27583 ;
  assign n27561 = ~n6529 & n24841 ;
  assign n27560 = ~n6547 & ~n21212 ;
  assign n27562 = n27561 ^ n27560 ;
  assign n27563 = n27562 ^ n6537 ;
  assign n27564 = n27563 ^ x14 ;
  assign n27568 = n27562 ^ x14 ;
  assign n27569 = n27568 ^ n6539 ;
  assign n27565 = n25282 ^ n6539 ;
  assign n27566 = n27565 ^ x13 ;
  assign n27567 = n27566 ^ n25282 ;
  assign n27570 = n27569 ^ n27567 ;
  assign n27571 = n27570 ^ n27569 ;
  assign n27574 = ~n25299 & ~n27571 ;
  assign n27575 = ~x13 & n27574 ;
  assign n27578 = n27575 ^ n27574 ;
  assign n27576 = n27575 ^ n25282 ;
  assign n27577 = n27569 & n27576 ;
  assign n27579 = n27578 ^ n27577 ;
  assign n27580 = n27579 ^ n6539 ;
  assign n27581 = ~n27564 & ~n27580 ;
  assign n27553 = n6143 & n20908 ;
  assign n27552 = n6148 & n21147 ;
  assign n27554 = n27553 ^ n27552 ;
  assign n27555 = n27554 ^ x17 ;
  assign n27551 = n6163 & ~n25073 ;
  assign n27556 = n27555 ^ n27551 ;
  assign n27550 = n20437 & ~n20612 ;
  assign n27557 = n27556 ^ n27550 ;
  assign n27546 = n13433 & ~n20617 ;
  assign n27544 = n5426 & ~n20614 ;
  assign n27537 = n20613 ^ x20 ;
  assign n27538 = n27537 ^ x19 ;
  assign n27539 = n27538 ^ n20613 ;
  assign n27540 = ~n21226 & n27539 ;
  assign n27541 = n27540 ^ n20613 ;
  assign n27542 = n5215 & ~n27541 ;
  assign n27543 = n27542 ^ x20 ;
  assign n27545 = n27544 ^ n27543 ;
  assign n27547 = n27546 ^ n27545 ;
  assign n27529 = ~n40 & n20624 ;
  assign n27527 = n4656 & n22968 ;
  assign n27524 = n4655 & ~n20620 ;
  assign n27523 = n4651 & n20829 ;
  assign n27525 = n27524 ^ n27523 ;
  assign n27526 = n27525 ^ x23 ;
  assign n27528 = n27527 ^ n27526 ;
  assign n27530 = n27529 ^ n27528 ;
  assign n27513 = ~x25 & ~n23306 ;
  assign n27516 = n27513 ^ n23307 ;
  assign n27517 = n99 & n27516 ;
  assign n27510 = n4600 & n20819 ;
  assign n27509 = n20603 & n20631 ;
  assign n27511 = n27510 ^ n27509 ;
  assign n27512 = n27511 ^ x26 ;
  assign n27514 = n27513 ^ n20628 ;
  assign n27515 = n27512 & n27514 ;
  assign n27518 = n27517 ^ n27515 ;
  assign n27519 = n27511 ^ n97 ;
  assign n27520 = ~n27518 & ~n27519 ;
  assign n27505 = n27352 ^ n27299 ;
  assign n27506 = ~n27353 & ~n27505 ;
  assign n27507 = n27506 ^ n27352 ;
  assign n27502 = n3837 & ~n20690 ;
  assign n27500 = n3985 & ~n20683 ;
  assign n27493 = n20680 ^ x29 ;
  assign n27494 = n27493 ^ x28 ;
  assign n27495 = n27494 ^ n20680 ;
  assign n27496 = ~n22661 & n27495 ;
  assign n27497 = n27496 ^ n20680 ;
  assign n27498 = n3833 & n27497 ;
  assign n27499 = n27498 ^ x29 ;
  assign n27501 = n27500 ^ n27499 ;
  assign n27503 = n27502 ^ n27501 ;
  assign n27487 = n26950 ^ x8 ;
  assign n27488 = ~n27339 & n27487 ;
  assign n27489 = n27488 ^ x8 ;
  assign n27479 = n5354 ^ n444 ;
  assign n27480 = n27479 ^ n915 ;
  assign n27478 = n838 ^ n354 ;
  assign n27481 = n27480 ^ n27478 ;
  assign n27476 = n26926 ^ n1699 ;
  assign n27475 = n13617 ^ n1554 ;
  assign n27477 = n27476 ^ n27475 ;
  assign n27482 = n27481 ^ n27477 ;
  assign n27474 = n13466 ^ n5299 ;
  assign n27483 = n27482 ^ n27474 ;
  assign n27484 = n27483 ^ n4929 ;
  assign n27485 = n27484 ^ n1072 ;
  assign n27486 = ~n2466 & ~n27485 ;
  assign n27490 = n27489 ^ n27486 ;
  assign n27464 = x31 & ~n27300 ;
  assign n27465 = n22091 ^ n3518 ;
  assign n27466 = n27465 ^ n22091 ;
  assign n27467 = ~x30 & n20694 ;
  assign n27468 = n27467 ^ n22091 ;
  assign n27469 = ~n27466 & ~n27468 ;
  assign n27470 = n27469 ^ n22091 ;
  assign n27471 = n27464 & ~n27470 ;
  assign n27472 = n27471 ^ n27464 ;
  assign n24266 = n20694 ^ n20693 ;
  assign n27461 = ~n61 & n24266 ;
  assign n27462 = n27461 ^ n20693 ;
  assign n27463 = ~n3800 & ~n27462 ;
  assign n27473 = n27472 ^ n27463 ;
  assign n27491 = n27490 ^ n27473 ;
  assign n27455 = n27340 ^ n27321 ;
  assign n27456 = n27326 & ~n27455 ;
  assign n27457 = n27456 ^ n27321 ;
  assign n27492 = n27491 ^ n27457 ;
  assign n27504 = n27503 ^ n27492 ;
  assign n27508 = n27507 ^ n27504 ;
  assign n27521 = n27520 ^ n27508 ;
  assign n27452 = n27362 ^ n27296 ;
  assign n27453 = n27363 & ~n27452 ;
  assign n27454 = n27453 ^ n27362 ;
  assign n27522 = n27521 ^ n27454 ;
  assign n27531 = n27530 ^ n27522 ;
  assign n27532 = n27531 ^ n27376 ;
  assign n27533 = n27532 ^ n27367 ;
  assign n27534 = n27533 ^ n27531 ;
  assign n27535 = n27368 & n27534 ;
  assign n27536 = n27535 ^ n27532 ;
  assign n27548 = n27547 ^ n27536 ;
  assign n27449 = n27393 ^ n27389 ;
  assign n27450 = n27390 & n27449 ;
  assign n27451 = n27450 ^ n27393 ;
  assign n27549 = n27548 ^ n27451 ;
  assign n27558 = n27557 ^ n27549 ;
  assign n27446 = n27394 ^ n27290 ;
  assign n27447 = ~n27400 & ~n27446 ;
  assign n27448 = n27447 ^ n27394 ;
  assign n27559 = n27558 ^ n27448 ;
  assign n27582 = n27581 ^ n27559 ;
  assign n27589 = n27588 ^ n27582 ;
  assign n27444 = n27434 ^ n27410 ;
  assign n27445 = ~n27441 & n27444 ;
  assign n27590 = n27589 ^ n27445 ;
  assign n27593 = n27592 ^ n27590 ;
  assign n27595 = n27594 ^ n27593 ;
  assign n27738 = n27434 & n27589 ;
  assign n27743 = n27409 & ~n27591 ;
  assign n27744 = n27743 ^ n27408 ;
  assign n27745 = n27738 & ~n27744 ;
  assign n27746 = n27745 ^ n27434 ;
  assign n27747 = n27440 & n27746 ;
  assign n27741 = n27591 ^ n27408 ;
  assign n27748 = n27591 ^ n27440 ;
  assign n27749 = n27748 ^ n27591 ;
  assign n27750 = n27591 ^ n27434 ;
  assign n27751 = n27750 ^ n27591 ;
  assign n27752 = ~n27749 & ~n27751 ;
  assign n27753 = n27752 ^ n27591 ;
  assign n27754 = n27741 & ~n27753 ;
  assign n27755 = n27754 ^ n27591 ;
  assign n27756 = n27755 ^ n27589 ;
  assign n27757 = n27754 ^ n27589 ;
  assign n27758 = n27405 & ~n27757 ;
  assign n27759 = n27758 ^ n27589 ;
  assign n27760 = ~n27756 & ~n27759 ;
  assign n27761 = n27760 ^ n27589 ;
  assign n27762 = ~n27747 & ~n27761 ;
  assign n27763 = n27762 ^ n27747 ;
  assign n27733 = n27581 ^ n27448 ;
  assign n27734 = n27559 & n27733 ;
  assign n27735 = n27734 ^ n27581 ;
  assign n27730 = n27586 ^ n27582 ;
  assign n27731 = ~n27588 & ~n27730 ;
  assign n27732 = n27731 ^ n27586 ;
  assign n27736 = n27735 ^ n27732 ;
  assign n27724 = n25311 ^ n7047 ;
  assign n27725 = n7047 ^ x14 ;
  assign n27726 = ~n27724 & n27725 ;
  assign n27721 = ~n6547 & ~n24841 ;
  assign n27718 = n6391 & ~n7310 ;
  assign n27719 = n25308 & n27718 ;
  assign n27716 = ~n6529 & n25282 ;
  assign n27715 = n8855 ^ n6392 ;
  assign n27717 = n27716 ^ n27715 ;
  assign n27720 = n27719 ^ n27717 ;
  assign n27722 = n27721 ^ n27720 ;
  assign n27714 = n15618 & n25311 ;
  assign n27723 = n27722 ^ n27714 ;
  assign n27727 = n27726 ^ n27723 ;
  assign n27706 = n20437 & n20908 ;
  assign n27704 = n6143 & n21147 ;
  assign n27697 = n21212 ^ x16 ;
  assign n27698 = n27697 ^ x17 ;
  assign n27699 = n27698 ^ n21212 ;
  assign n27700 = ~n25342 & n27699 ;
  assign n27701 = n27700 ^ n21212 ;
  assign n27702 = n6141 & ~n27701 ;
  assign n27703 = n27702 ^ x17 ;
  assign n27705 = n27704 ^ n27703 ;
  assign n27707 = n27706 ^ n27705 ;
  assign n27689 = n13433 & ~n20614 ;
  assign n27687 = n5426 & ~n20613 ;
  assign n27680 = n20612 ^ x20 ;
  assign n27681 = n27680 ^ x19 ;
  assign n27682 = n27681 ^ n20612 ;
  assign n27683 = ~n23892 & n27682 ;
  assign n27684 = n27683 ^ n20612 ;
  assign n27685 = n5215 & ~n27684 ;
  assign n27686 = n27685 ^ x20 ;
  assign n27688 = n27687 ^ n27686 ;
  assign n27690 = n27689 ^ n27688 ;
  assign n27668 = n4655 & ~n20617 ;
  assign n27667 = n4651 & n20624 ;
  assign n27669 = n27668 ^ n27667 ;
  assign n27670 = n27669 ^ x23 ;
  assign n27666 = n4656 & n23491 ;
  assign n27671 = n27670 ^ n27666 ;
  assign n27665 = ~n40 & ~n20620 ;
  assign n27672 = n27671 ^ n27665 ;
  assign n27657 = ~n4435 & ~n22979 ;
  assign n27655 = ~n4434 & n20829 ;
  assign n27652 = n20603 & n20819 ;
  assign n27651 = n4600 & ~n20628 ;
  assign n27653 = n27652 ^ n27651 ;
  assign n27654 = n27653 ^ x26 ;
  assign n27656 = n27655 ^ n27654 ;
  assign n27658 = n27657 ^ n27656 ;
  assign n27643 = n3837 & ~n20683 ;
  assign n27641 = n3985 & n20680 ;
  assign n27634 = n20631 ^ x29 ;
  assign n27635 = n27634 ^ x28 ;
  assign n27636 = n27635 ^ n20631 ;
  assign n27637 = ~n22649 & n27636 ;
  assign n27638 = n27637 ^ n20631 ;
  assign n27639 = n3833 & n27638 ;
  assign n27640 = n27639 ^ x29 ;
  assign n27642 = n27641 ^ n27640 ;
  assign n27644 = n27643 ^ n27642 ;
  assign n27628 = n27489 ^ n27473 ;
  assign n27629 = ~n27490 & n27628 ;
  assign n27620 = n1581 ^ n527 ;
  assign n27621 = n27620 ^ n524 ;
  assign n27618 = n2032 ^ n969 ;
  assign n27619 = n27618 ^ n1778 ;
  assign n27622 = n27621 ^ n27619 ;
  assign n27617 = n13570 ^ n843 ;
  assign n27623 = n27622 ^ n27617 ;
  assign n27615 = n5327 ^ n2073 ;
  assign n27614 = n4859 ^ n2735 ;
  assign n27616 = n27615 ^ n27614 ;
  assign n27624 = n27623 ^ n27616 ;
  assign n27613 = n14320 ^ n12824 ;
  assign n27625 = n27624 ^ n27613 ;
  assign n27626 = ~n26948 & ~n27625 ;
  assign n27627 = ~n5689 & n27626 ;
  assign n27630 = n27629 ^ n27627 ;
  assign n27607 = n20690 ^ n3518 ;
  assign n27606 = ~n3518 & n20690 ;
  assign n27608 = n27607 ^ n27606 ;
  assign n27605 = ~n61 & ~n20693 ;
  assign n27609 = n27608 ^ n27605 ;
  assign n27631 = n27630 ^ n27609 ;
  assign n27610 = n27609 ^ n21246 ;
  assign n27598 = n21246 ^ n20693 ;
  assign n27597 = n21246 ^ n20694 ;
  assign n27599 = n27598 ^ n27597 ;
  assign n27600 = n27598 ^ x30 ;
  assign n27601 = n27600 ^ n27598 ;
  assign n27602 = n27599 & n27601 ;
  assign n27603 = n27602 ^ n27598 ;
  assign n27604 = ~n3518 & ~n27603 ;
  assign n27611 = n27610 ^ n27604 ;
  assign n27612 = x31 & n27611 ;
  assign n27632 = n27631 ^ n27612 ;
  assign n27645 = n27644 ^ n27632 ;
  assign n27646 = n27645 ^ n27503 ;
  assign n27647 = n27646 ^ n27457 ;
  assign n27648 = n27647 ^ n27645 ;
  assign n27649 = n27492 & n27648 ;
  assign n27650 = n27649 ^ n27646 ;
  assign n27659 = n27658 ^ n27650 ;
  assign n27660 = n27659 ^ n27520 ;
  assign n27661 = n27660 ^ n27507 ;
  assign n27662 = n27661 ^ n27659 ;
  assign n27663 = n27508 & ~n27662 ;
  assign n27664 = n27663 ^ n27660 ;
  assign n27673 = n27672 ^ n27664 ;
  assign n27674 = n27673 ^ n27530 ;
  assign n27675 = n27674 ^ n27454 ;
  assign n27676 = n27675 ^ n27673 ;
  assign n27677 = ~n27522 & n27676 ;
  assign n27678 = n27677 ^ n27674 ;
  assign n27691 = n27690 ^ n27678 ;
  assign n27693 = n27691 ^ n27531 ;
  assign n27692 = n27691 ^ n27547 ;
  assign n27694 = n27693 ^ n27692 ;
  assign n27695 = n27536 & n27694 ;
  assign n27696 = n27695 ^ n27693 ;
  assign n27708 = n27707 ^ n27696 ;
  assign n27709 = n27708 ^ n27557 ;
  assign n27710 = n27709 ^ n27708 ;
  assign n27711 = n27710 ^ n27451 ;
  assign n27712 = ~n27549 & n27711 ;
  assign n27713 = n27712 ^ n27709 ;
  assign n27728 = n27727 ^ n27713 ;
  assign n27729 = n27728 ^ x11 ;
  assign n27737 = n27736 ^ n27729 ;
  assign n27764 = n27763 ^ n27737 ;
  assign n27596 = n27593 & n27594 ;
  assign n27765 = n27764 ^ n27596 ;
  assign n27912 = n27596 & ~n27764 ;
  assign n27906 = n27727 ^ n27708 ;
  assign n27907 = n27713 & ~n27906 ;
  assign n27908 = n27907 ^ n27708 ;
  assign n27883 = n25282 ^ x13 ;
  assign n27893 = n6390 & ~n27883 ;
  assign n27885 = n24841 ^ x14 ;
  assign n27896 = ~n25282 & ~n27885 ;
  assign n27897 = n27896 ^ n24841 ;
  assign n27898 = n27893 & ~n27897 ;
  assign n27899 = n27898 ^ x14 ;
  assign n27884 = ~n6392 & n27883 ;
  assign n27890 = n25282 & n27885 ;
  assign n27891 = n27890 ^ x14 ;
  assign n27892 = n27884 & ~n27891 ;
  assign n27900 = n27899 ^ n27892 ;
  assign n27901 = n27900 ^ x13 ;
  assign n27902 = n6391 & n25515 ;
  assign n27903 = n27901 & n27902 ;
  assign n27904 = n27903 ^ n27900 ;
  assign n27879 = n27707 ^ n27691 ;
  assign n27880 = n27696 & n27879 ;
  assign n27881 = n27880 ^ n27691 ;
  assign n27873 = n6148 & n24841 ;
  assign n27872 = n6143 & ~n21212 ;
  assign n27874 = n27873 ^ n27872 ;
  assign n27875 = n27874 ^ x17 ;
  assign n27871 = n6163 & ~n25528 ;
  assign n27876 = n27875 ^ n27871 ;
  assign n27870 = n20437 & n21147 ;
  assign n27877 = n27876 ^ n27870 ;
  assign n27865 = n27672 ^ n27659 ;
  assign n27866 = n27664 & ~n27865 ;
  assign n27867 = n27866 ^ n27659 ;
  assign n27862 = ~n40 & ~n20617 ;
  assign n27860 = n4656 & n23480 ;
  assign n27857 = n4655 & ~n20614 ;
  assign n27856 = n4651 & ~n20620 ;
  assign n27858 = n27857 ^ n27856 ;
  assign n27859 = n27858 ^ x23 ;
  assign n27861 = n27860 ^ n27859 ;
  assign n27863 = n27862 ^ n27861 ;
  assign n27853 = ~n4435 & ~n21232 ;
  assign n27846 = n3985 & n20631 ;
  assign n27842 = n4368 & ~n21236 ;
  assign n27841 = n3837 & n20680 ;
  assign n27843 = n27842 ^ n27841 ;
  assign n27844 = n27843 ^ x29 ;
  assign n27838 = x28 & ~n21236 ;
  assign n27839 = n27838 ^ n21237 ;
  assign n27840 = n3833 & ~n27839 ;
  assign n27845 = n27844 ^ n27840 ;
  assign n27847 = n27846 ^ n27845 ;
  assign n27829 = n12664 & ~n27606 ;
  assign n27823 = n22618 ^ n20683 ;
  assign n27824 = n20683 ^ x31 ;
  assign n27825 = n27824 ^ n20683 ;
  assign n27826 = ~n27823 & n27825 ;
  assign n27827 = n27826 ^ n20683 ;
  assign n27828 = n3518 & n27827 ;
  assign n27830 = n27829 ^ n27828 ;
  assign n27821 = ~n61 & ~n20690 ;
  assign n27831 = n27830 ^ n27821 ;
  assign n27820 = x31 & n27605 ;
  assign n27832 = n27831 ^ n27820 ;
  assign n27807 = n27130 ^ n602 ;
  assign n27806 = n3582 ^ n567 ;
  assign n27808 = n27807 ^ n27806 ;
  assign n27805 = n2510 ^ n1315 ;
  assign n27809 = n27808 ^ n27805 ;
  assign n27804 = n5555 ^ n2714 ;
  assign n27810 = n27809 ^ n27804 ;
  assign n27811 = n27810 ^ n2113 ;
  assign n27812 = n27811 ^ n2160 ;
  assign n27814 = n5543 ^ n1175 ;
  assign n27813 = n3769 ^ n528 ;
  assign n27815 = n27814 ^ n27813 ;
  assign n27816 = n27815 ^ n1246 ;
  assign n27817 = ~n27812 & ~n27816 ;
  assign n27818 = n27817 ^ x11 ;
  assign n27795 = ~n27473 & n27489 ;
  assign n27798 = n27627 & n27795 ;
  assign n27819 = n27818 ^ n27798 ;
  assign n27833 = n27832 ^ n27819 ;
  assign n27801 = n27644 ^ n27630 ;
  assign n27802 = n27632 & ~n27801 ;
  assign n27803 = n27802 ^ n27644 ;
  assign n27834 = n27833 ^ n27803 ;
  assign n27796 = n27795 ^ n27628 ;
  assign n27797 = ~n27627 & n27796 ;
  assign n27799 = n27798 ^ n27797 ;
  assign n27800 = ~n27486 & n27799 ;
  assign n27835 = n27834 ^ n27800 ;
  assign n27848 = n27847 ^ n27835 ;
  assign n27849 = n27848 ^ x26 ;
  assign n27794 = n4600 & n20829 ;
  assign n27850 = n27849 ^ n27794 ;
  assign n27793 = n20603 & ~n20628 ;
  assign n27851 = n27850 ^ n27793 ;
  assign n27792 = ~n4434 & n20624 ;
  assign n27852 = n27851 ^ n27792 ;
  assign n27854 = n27853 ^ n27852 ;
  assign n27789 = n27658 ^ n27645 ;
  assign n27790 = ~n27650 & ~n27789 ;
  assign n27791 = n27790 ^ n27645 ;
  assign n27855 = n27854 ^ n27791 ;
  assign n27864 = n27863 ^ n27855 ;
  assign n27868 = n27867 ^ n27864 ;
  assign n27786 = n5426 & ~n20612 ;
  assign n27781 = n27690 ^ n27673 ;
  assign n27782 = n27678 & n27781 ;
  assign n27783 = n27782 ^ n27673 ;
  assign n27784 = n27783 ^ x20 ;
  assign n27776 = n20908 ^ n5224 ;
  assign n27777 = n27776 ^ n20908 ;
  assign n27778 = ~n24096 & n27777 ;
  assign n27779 = n27778 ^ n20908 ;
  assign n27780 = n5215 & n27779 ;
  assign n27785 = n27784 ^ n27780 ;
  assign n27787 = n27786 ^ n27785 ;
  assign n27774 = n13433 & ~n20613 ;
  assign n27788 = n27787 ^ n27774 ;
  assign n27869 = n27868 ^ n27788 ;
  assign n27878 = n27877 ^ n27869 ;
  assign n27882 = n27881 ^ n27878 ;
  assign n27905 = n27904 ^ n27882 ;
  assign n27909 = n27908 ^ n27905 ;
  assign n27769 = n27735 ^ x11 ;
  assign n27770 = n27735 ^ n27728 ;
  assign n27771 = n27770 ^ n27763 ;
  assign n27772 = n27771 ^ n27732 ;
  assign n27773 = n27769 & ~n27772 ;
  assign n27910 = n27909 ^ n27773 ;
  assign n27766 = n27763 ^ n27728 ;
  assign n27767 = n27732 ^ n27728 ;
  assign n27768 = n27766 & ~n27767 ;
  assign n27911 = n27910 ^ n27768 ;
  assign n27913 = n27912 ^ n27911 ;
  assign n28060 = n27911 & n27912 ;
  assign n28039 = n27728 & ~n27763 ;
  assign n28040 = n28039 ^ n27766 ;
  assign n28041 = n27909 ^ n27735 ;
  assign n28042 = n27769 & n28041 ;
  assign n28043 = n27909 ^ n27732 ;
  assign n28044 = n28042 & n28043 ;
  assign n28045 = n28044 ^ n27909 ;
  assign n28046 = ~n28040 & n28045 ;
  assign n28047 = n28039 ^ n27909 ;
  assign n28049 = n28039 ^ n27735 ;
  assign n28048 = n28039 ^ n27732 ;
  assign n28050 = n28049 ^ n28048 ;
  assign n28051 = n28049 ^ n27732 ;
  assign n28052 = n28051 ^ x11 ;
  assign n28053 = n28052 ^ n28049 ;
  assign n28054 = n28050 & n28053 ;
  assign n28055 = n28054 ^ n28049 ;
  assign n28056 = n28047 & ~n28055 ;
  assign n28057 = n28056 ^ n27909 ;
  assign n28058 = ~n28046 & ~n28057 ;
  assign n28032 = n6148 & ~n25282 ;
  assign n28028 = n6143 & n24841 ;
  assign n28029 = n28028 ^ x17 ;
  assign n28027 = n20437 & ~n21212 ;
  assign n28030 = n28029 ^ n28027 ;
  assign n28026 = n6163 & n25868 ;
  assign n28031 = n28030 ^ n28026 ;
  assign n28033 = n28032 ^ n28031 ;
  assign n28022 = n13433 & ~n20612 ;
  assign n28020 = n5426 & n20908 ;
  assign n28013 = n21147 ^ x20 ;
  assign n28014 = n28013 ^ x19 ;
  assign n28015 = n28014 ^ n21147 ;
  assign n28016 = ~n24078 & n28015 ;
  assign n28017 = n28016 ^ n21147 ;
  assign n28018 = n5215 & n28017 ;
  assign n28019 = n28018 ^ x20 ;
  assign n28021 = n28020 ^ n28019 ;
  assign n28023 = n28022 ^ n28021 ;
  assign n28005 = n4655 & ~n20613 ;
  assign n28004 = n4651 & ~n20617 ;
  assign n28006 = n28005 ^ n28004 ;
  assign n28007 = n28006 ^ x23 ;
  assign n28003 = n4656 & n21227 ;
  assign n28008 = n28007 ^ n28003 ;
  assign n28002 = ~n40 & ~n20614 ;
  assign n28009 = n28008 ^ n28002 ;
  assign n27994 = ~n4435 & n22968 ;
  assign n27992 = ~n4434 & ~n20620 ;
  assign n27989 = n4600 & n20624 ;
  assign n27988 = n20603 & n20829 ;
  assign n27990 = n27989 ^ n27988 ;
  assign n27991 = n27990 ^ x26 ;
  assign n27993 = n27992 ^ n27991 ;
  assign n27995 = n27994 ^ n27993 ;
  assign n27984 = n3837 & n20631 ;
  assign n27982 = n3985 & n20819 ;
  assign n27975 = n20628 ^ x29 ;
  assign n27976 = n27975 ^ x28 ;
  assign n27977 = n27976 ^ n20628 ;
  assign n27978 = ~n25230 & n27977 ;
  assign n27979 = n27978 ^ n20628 ;
  assign n27980 = n3833 & ~n27979 ;
  assign n27981 = n27980 ^ x29 ;
  assign n27983 = n27982 ^ n27981 ;
  assign n27985 = n27984 ^ n27983 ;
  assign n27963 = n22662 ^ n20683 ;
  assign n27962 = n22662 ^ n20690 ;
  assign n27964 = n27963 ^ n27962 ;
  assign n27967 = x30 & n27964 ;
  assign n27968 = n27967 ^ n27963 ;
  assign n27969 = ~n3518 & n27968 ;
  assign n27970 = n27969 ^ n22662 ;
  assign n27971 = x31 & ~n27970 ;
  assign n27960 = n3807 & n20680 ;
  assign n27959 = ~n3805 & ~n20683 ;
  assign n27961 = n27960 ^ n27959 ;
  assign n27972 = n27971 ^ n27961 ;
  assign n27946 = n4710 ^ n744 ;
  assign n27945 = n3214 ^ n900 ;
  assign n27947 = n27946 ^ n27945 ;
  assign n27948 = n27947 ^ n12583 ;
  assign n27949 = n27948 ^ n14322 ;
  assign n27952 = n2243 ^ n218 ;
  assign n27950 = n2153 ^ n716 ;
  assign n27951 = n27950 ^ n1103 ;
  assign n27953 = n27952 ^ n27951 ;
  assign n27954 = n27953 ^ n25959 ;
  assign n27955 = n27954 ^ n25592 ;
  assign n27956 = n27955 ^ n12527 ;
  assign n27957 = ~n27949 & ~n27956 ;
  assign n27941 = n27817 ^ n27486 ;
  assign n27942 = n27486 ^ x11 ;
  assign n27943 = ~n27941 & n27942 ;
  assign n27944 = n27943 ^ x11 ;
  assign n27958 = n27957 ^ n27944 ;
  assign n27973 = n27972 ^ n27958 ;
  assign n27931 = n27832 ^ n27818 ;
  assign n27932 = ~n27799 & n27931 ;
  assign n27930 = n27832 ^ n27797 ;
  assign n27933 = n27932 ^ n27930 ;
  assign n27934 = n27832 ^ n27486 ;
  assign n27935 = n27934 ^ n27818 ;
  assign n27936 = n27933 & ~n27935 ;
  assign n27937 = n27936 ^ n27832 ;
  assign n27974 = n27973 ^ n27937 ;
  assign n27986 = n27985 ^ n27974 ;
  assign n27927 = n27847 ^ n27803 ;
  assign n27928 = n27835 & n27927 ;
  assign n27929 = n27928 ^ n27847 ;
  assign n27987 = n27986 ^ n27929 ;
  assign n27996 = n27995 ^ n27987 ;
  assign n27997 = n27996 ^ n27848 ;
  assign n27998 = n27997 ^ n27791 ;
  assign n27999 = n27998 ^ n27996 ;
  assign n28000 = ~n27854 & n27999 ;
  assign n28001 = n28000 ^ n27997 ;
  assign n28010 = n28009 ^ n28001 ;
  assign n27924 = n27867 ^ n27863 ;
  assign n27925 = ~n27864 & ~n27924 ;
  assign n27926 = n27925 ^ n27867 ;
  assign n28011 = n28010 ^ n27926 ;
  assign n28024 = n28023 ^ n28011 ;
  assign n27921 = n27868 ^ n27783 ;
  assign n27922 = ~n27788 & ~n27921 ;
  assign n27923 = n27922 ^ n27868 ;
  assign n28025 = n28024 ^ n27923 ;
  assign n28034 = n28033 ^ n28025 ;
  assign n28035 = n28034 ^ x14 ;
  assign n27920 = ~n6547 & n25308 ;
  assign n28036 = n28035 ^ n27920 ;
  assign n27917 = n27881 ^ n27877 ;
  assign n27918 = n27878 & n27917 ;
  assign n27919 = n27918 ^ n27881 ;
  assign n28037 = n28036 ^ n27919 ;
  assign n27914 = n27908 ^ n27904 ;
  assign n27915 = n27905 & n27914 ;
  assign n27916 = n27915 ^ n27908 ;
  assign n28038 = n28037 ^ n27916 ;
  assign n28059 = n28058 ^ n28038 ;
  assign n28061 = n28060 ^ n28059 ;
  assign n28187 = n28059 & n28060 ;
  assign n28184 = n28034 ^ n27919 ;
  assign n28185 = n28036 & n28184 ;
  assign n28186 = n28185 ^ n28034 ;
  assign n28188 = n28187 ^ n28186 ;
  assign n28177 = n20437 & n24841 ;
  assign n28175 = n6143 ^ x17 ;
  assign n28174 = n6163 & n25311 ;
  assign n28176 = n28175 ^ n28174 ;
  assign n28178 = n28177 ^ n28176 ;
  assign n28171 = n6148 & ~n24841 ;
  assign n28172 = n28171 ^ n6143 ;
  assign n28173 = n25282 & n28172 ;
  assign n28179 = n28178 ^ n28173 ;
  assign n28159 = n13433 & n20908 ;
  assign n28157 = n5426 & n21147 ;
  assign n28150 = n21212 ^ x19 ;
  assign n28151 = n28150 ^ x20 ;
  assign n28152 = n28151 ^ n21212 ;
  assign n28153 = ~n25342 & n28152 ;
  assign n28154 = n28153 ^ n21212 ;
  assign n28155 = n5215 & ~n28154 ;
  assign n28156 = n28155 ^ x20 ;
  assign n28158 = n28157 ^ n28156 ;
  assign n28160 = n28159 ^ n28158 ;
  assign n28142 = n4651 & ~n20614 ;
  assign n28140 = ~n40 & ~n20613 ;
  assign n28133 = n20612 ^ x23 ;
  assign n28134 = n28133 ^ x22 ;
  assign n28135 = n28134 ^ n20612 ;
  assign n28136 = ~n23892 & n28135 ;
  assign n28137 = n28136 ^ n20612 ;
  assign n28138 = n35 & ~n28137 ;
  assign n28139 = n28138 ^ x23 ;
  assign n28141 = n28140 ^ n28139 ;
  assign n28143 = n28142 ^ n28141 ;
  assign n28125 = ~n4435 & n23491 ;
  assign n28123 = n4600 & ~n20620 ;
  assign n28120 = ~n4434 & ~n20617 ;
  assign n28119 = n20603 & n20624 ;
  assign n28121 = n28120 ^ n28119 ;
  assign n28122 = n28121 ^ x26 ;
  assign n28124 = n28123 ^ n28122 ;
  assign n28126 = n28125 ^ n28124 ;
  assign n28117 = n3985 & ~n20628 ;
  assign n28115 = n3837 & n20819 ;
  assign n28109 = n27937 & n27985 ;
  assign n28107 = ~n27944 & n27957 ;
  assign n28108 = n28107 ^ n27958 ;
  assign n28110 = n28109 ^ n28108 ;
  assign n28089 = n3518 & n22653 ;
  assign n28090 = n20631 ^ n3518 ;
  assign n28091 = n28090 ^ n20631 ;
  assign n28092 = x30 & n24659 ;
  assign n28093 = n28092 ^ n20631 ;
  assign n28094 = ~n28091 & n28093 ;
  assign n28095 = n28094 ^ n20631 ;
  assign n28096 = ~x31 & n28095 ;
  assign n28101 = n28096 ^ x31 ;
  assign n24205 = n20683 ^ n20680 ;
  assign n28097 = n27493 ^ n20680 ;
  assign n28098 = ~n24205 & n28097 ;
  assign n28099 = n28098 ^ n20680 ;
  assign n28100 = n3967 & ~n28099 ;
  assign n28102 = n28101 ^ n28100 ;
  assign n28103 = n28102 ^ n28096 ;
  assign n28104 = n28089 & n28103 ;
  assign n28105 = n28104 ^ n28102 ;
  assign n28084 = n3581 ^ n824 ;
  assign n28085 = n28084 ^ n5596 ;
  assign n28079 = n3188 ^ n2018 ;
  assign n28078 = n1148 ^ n611 ;
  assign n28080 = n28079 ^ n28078 ;
  assign n28077 = n3620 ^ n711 ;
  assign n28081 = n28080 ^ n28077 ;
  assign n28076 = n3675 ^ n2716 ;
  assign n28082 = n28081 ^ n28076 ;
  assign n28083 = n28082 ^ n2997 ;
  assign n28086 = n28085 ^ n28083 ;
  assign n28087 = ~n12769 & ~n28086 ;
  assign n28088 = n28087 ^ n27957 ;
  assign n28106 = n28105 ^ n28088 ;
  assign n28111 = n28110 ^ n28106 ;
  assign n28073 = n27985 ^ n27937 ;
  assign n28074 = n28073 ^ n27958 ;
  assign n28075 = ~n27973 & ~n28074 ;
  assign n28112 = n28111 ^ n28075 ;
  assign n28113 = n28112 ^ x29 ;
  assign n28068 = n22979 ^ n5065 ;
  assign n28069 = n28068 ^ n22979 ;
  assign n28070 = ~n22978 & ~n28069 ;
  assign n28071 = n28070 ^ n22979 ;
  assign n28072 = n3833 & ~n28071 ;
  assign n28114 = n28113 ^ n28072 ;
  assign n28116 = n28115 ^ n28114 ;
  assign n28118 = n28117 ^ n28116 ;
  assign n28127 = n28126 ^ n28118 ;
  assign n28128 = n28127 ^ n27995 ;
  assign n28129 = n28128 ^ n27929 ;
  assign n28130 = n28129 ^ n28127 ;
  assign n28131 = n27987 & n28130 ;
  assign n28132 = n28131 ^ n28128 ;
  assign n28144 = n28143 ^ n28132 ;
  assign n28146 = n28144 ^ n27996 ;
  assign n28145 = n28144 ^ n28009 ;
  assign n28147 = n28146 ^ n28145 ;
  assign n28148 = n28001 & ~n28147 ;
  assign n28149 = n28148 ^ n28146 ;
  assign n28161 = n28160 ^ n28149 ;
  assign n28162 = n28161 ^ n28023 ;
  assign n28163 = n28162 ^ n28161 ;
  assign n28164 = n28163 ^ n27926 ;
  assign n28165 = n28011 & ~n28164 ;
  assign n28166 = n28165 ^ n28162 ;
  assign n28180 = n28179 ^ n28166 ;
  assign n28065 = n28033 ^ n27923 ;
  assign n28066 = ~n28025 & ~n28065 ;
  assign n28067 = n28066 ^ n28033 ;
  assign n28181 = n28180 ^ n28067 ;
  assign n28182 = n28181 ^ x14 ;
  assign n28062 = n28058 ^ n27916 ;
  assign n28063 = ~n28038 & n28062 ;
  assign n28064 = n28063 ^ n28058 ;
  assign n28183 = n28182 ^ n28064 ;
  assign n28189 = n28188 ^ n28183 ;
  assign n28323 = n28186 ^ n28182 ;
  assign n28326 = n28183 & n28323 ;
  assign n28324 = n28323 ^ n28064 ;
  assign n28325 = ~n28187 & ~n28324 ;
  assign n28327 = n28326 ^ n28325 ;
  assign n28314 = n28179 ^ n28161 ;
  assign n28315 = ~n28166 & ~n28314 ;
  assign n28316 = n28315 ^ n28161 ;
  assign n28311 = n6163 & n25515 ;
  assign n28307 = n20437 ^ n6143 ;
  assign n28308 = n28307 ^ n28028 ;
  assign n28309 = n25282 & n28308 ;
  assign n28306 = n20437 ^ x17 ;
  assign n28310 = n28309 ^ n28306 ;
  assign n28312 = n28311 ^ n28310 ;
  assign n28302 = n28160 ^ n28144 ;
  assign n28303 = ~n28149 & n28302 ;
  assign n28304 = n28303 ^ n28144 ;
  assign n28299 = n13433 & n21147 ;
  assign n28297 = n5426 & ~n21212 ;
  assign n28290 = n24841 ^ x20 ;
  assign n28291 = n28290 ^ x19 ;
  assign n28292 = n28291 ^ n24841 ;
  assign n28293 = ~n27272 & n28292 ;
  assign n28294 = n28293 ^ n24841 ;
  assign n28295 = n5215 & n28294 ;
  assign n28296 = n28295 ^ x20 ;
  assign n28298 = n28297 ^ n28296 ;
  assign n28300 = n28299 ^ n28298 ;
  assign n28287 = ~n40 & ~n20612 ;
  assign n28285 = n4656 & ~n25056 ;
  assign n28282 = n4655 & n20908 ;
  assign n28281 = n4651 & ~n20613 ;
  assign n28283 = n28282 ^ n28281 ;
  assign n28284 = n28283 ^ x23 ;
  assign n28286 = n28285 ^ n28284 ;
  assign n28288 = n28287 ^ n28286 ;
  assign n28277 = n28143 ^ n28127 ;
  assign n28278 = n28132 & n28277 ;
  assign n28279 = n28278 ^ n28127 ;
  assign n28274 = ~n4435 & n23480 ;
  assign n28272 = ~n4434 & ~n20614 ;
  assign n28269 = n20603 & ~n20620 ;
  assign n28268 = n4600 & ~n20617 ;
  assign n28270 = n28269 ^ n28268 ;
  assign n28271 = n28270 ^ x26 ;
  assign n28273 = n28272 ^ n28271 ;
  assign n28275 = n28274 ^ n28273 ;
  assign n28259 = n28105 ^ n28087 ;
  assign n28260 = ~n28088 & n28259 ;
  assign n28247 = n21237 ^ n20631 ;
  assign n28246 = n21237 ^ n20680 ;
  assign n28248 = n28247 ^ n28246 ;
  assign n28251 = x30 & n28248 ;
  assign n28252 = n28251 ^ n28247 ;
  assign n28253 = ~n3518 & ~n28252 ;
  assign n28254 = n28253 ^ n21237 ;
  assign n28255 = x31 & ~n28254 ;
  assign n28244 = n3807 & n20819 ;
  assign n28243 = ~n3805 & n20631 ;
  assign n28245 = n28244 ^ n28243 ;
  assign n28256 = n28255 ^ n28245 ;
  assign n28237 = n5347 ^ n1492 ;
  assign n28233 = n2352 ^ n247 ;
  assign n28234 = n28233 ^ n429 ;
  assign n28231 = n4138 ^ n240 ;
  assign n28232 = n28231 ^ n1837 ;
  assign n28235 = n28234 ^ n28232 ;
  assign n28230 = n13579 ^ n3025 ;
  assign n28236 = n28235 ^ n28230 ;
  assign n28238 = n28237 ^ n28236 ;
  assign n28239 = n28238 ^ n6890 ;
  assign n28240 = n28239 ^ n13373 ;
  assign n28241 = ~n2094 & ~n28240 ;
  assign n28242 = n28241 ^ x14 ;
  assign n28257 = n28256 ^ n28242 ;
  assign n28209 = n27972 & n28107 ;
  assign n28202 = n28106 ^ n27972 ;
  assign n28201 = n28106 ^ n27944 ;
  assign n28203 = n28202 ^ n28201 ;
  assign n28204 = n28201 ^ n27958 ;
  assign n28205 = n28204 ^ n28201 ;
  assign n28206 = ~n28203 & ~n28205 ;
  assign n28207 = n28206 ^ n28201 ;
  assign n28208 = n28109 & n28207 ;
  assign n28210 = n28109 ^ n28073 ;
  assign n28211 = ~n28208 & n28210 ;
  assign n28212 = n28209 & n28211 ;
  assign n28213 = n28212 ^ n28208 ;
  assign n28214 = n28210 ^ n27958 ;
  assign n28215 = ~n27973 & ~n28214 ;
  assign n28216 = n28215 ^ n27958 ;
  assign n28217 = ~n28106 & n28216 ;
  assign n28218 = n28217 ^ n28106 ;
  assign n28219 = n28218 ^ n27957 ;
  assign n28220 = n28219 ^ n28218 ;
  assign n28223 = n28218 ^ n28215 ;
  assign n28224 = n28223 ^ n28218 ;
  assign n28225 = n28217 & ~n28224 ;
  assign n28226 = n28220 & n28225 ;
  assign n28227 = n28226 ^ n28220 ;
  assign n28228 = n28227 ^ n28219 ;
  assign n28229 = ~n28213 & n28228 ;
  assign n28258 = n28257 ^ n28229 ;
  assign n28261 = n28260 ^ n28258 ;
  assign n28199 = n3837 & ~n20628 ;
  assign n28197 = n3985 & n20829 ;
  assign n28190 = n20624 ^ x29 ;
  assign n28191 = n28190 ^ x28 ;
  assign n28192 = n28191 ^ n20624 ;
  assign n28193 = ~n21231 & n28192 ;
  assign n28194 = n28193 ^ n20624 ;
  assign n28195 = n3833 & n28194 ;
  assign n28196 = n28195 ^ x29 ;
  assign n28198 = n28197 ^ n28196 ;
  assign n28200 = n28199 ^ n28198 ;
  assign n28262 = n28261 ^ n28200 ;
  assign n28263 = n28262 ^ n28126 ;
  assign n28264 = n28263 ^ n28262 ;
  assign n28265 = n28264 ^ n28112 ;
  assign n28266 = ~n28118 & n28265 ;
  assign n28267 = n28266 ^ n28263 ;
  assign n28276 = n28275 ^ n28267 ;
  assign n28280 = n28279 ^ n28276 ;
  assign n28289 = n28288 ^ n28280 ;
  assign n28301 = n28300 ^ n28289 ;
  assign n28305 = n28304 ^ n28301 ;
  assign n28313 = n28312 ^ n28305 ;
  assign n28317 = n28316 ^ n28313 ;
  assign n28318 = n28317 ^ x14 ;
  assign n28319 = n28318 ^ n28067 ;
  assign n28320 = n28319 ^ n28317 ;
  assign n28321 = n28181 & n28320 ;
  assign n28322 = n28321 ^ n28318 ;
  assign n28328 = n28327 ^ n28322 ;
  assign n28448 = n28187 & ~n28324 ;
  assign n28449 = n28323 ^ n28322 ;
  assign n28450 = n28448 & ~n28449 ;
  assign n28429 = n28186 ^ n28180 ;
  assign n28430 = n28186 ^ x14 ;
  assign n28431 = n28429 & n28430 ;
  assign n28432 = n28431 ^ x14 ;
  assign n28433 = n28317 & ~n28432 ;
  assign n28434 = n28432 ^ n28317 ;
  assign n28435 = n28434 ^ n28433 ;
  assign n28436 = ~n28067 & ~n28435 ;
  assign n28437 = n28436 ^ n28064 ;
  assign n28441 = n28317 ^ n28064 ;
  assign n28438 = n28317 ^ n28180 ;
  assign n28439 = n28429 & ~n28430 ;
  assign n28440 = n28438 & n28439 ;
  assign n28442 = n28441 ^ n28440 ;
  assign n28443 = ~n28437 & ~n28442 ;
  assign n28444 = n28443 ^ n28064 ;
  assign n28445 = ~n28433 & n28444 ;
  assign n28421 = n5426 & n24841 ;
  assign n28419 = n5215 & n25868 ;
  assign n28418 = n5220 & ~n25299 ;
  assign n28420 = n28419 ^ n28418 ;
  assign n28422 = n28421 ^ n28420 ;
  assign n28423 = n28422 ^ x20 ;
  assign n28417 = n13433 & ~n21212 ;
  assign n28424 = n28423 ^ n28417 ;
  assign n28410 = n4655 & n21147 ;
  assign n28409 = n4651 & ~n20612 ;
  assign n28411 = n28410 ^ n28409 ;
  assign n28412 = n28411 ^ x23 ;
  assign n28408 = n4656 & ~n25073 ;
  assign n28413 = n28412 ^ n28408 ;
  assign n28407 = ~n40 & n20908 ;
  assign n28414 = n28413 ^ n28407 ;
  assign n28403 = n28275 ^ n28262 ;
  assign n28404 = n28267 & n28403 ;
  assign n28405 = n28404 ^ n28262 ;
  assign n28400 = ~n4435 & n21227 ;
  assign n28398 = ~n4434 & ~n20613 ;
  assign n28395 = n4600 & ~n20614 ;
  assign n28394 = n20603 & ~n20617 ;
  assign n28396 = n28395 ^ n28394 ;
  assign n28397 = n28396 ^ x26 ;
  assign n28399 = n28398 ^ n28397 ;
  assign n28401 = n28400 ^ n28399 ;
  assign n28380 = ~x28 & ~n22963 ;
  assign n28385 = n28380 ^ n22968 ;
  assign n28386 = n4368 & n28385 ;
  assign n28381 = n28380 ^ n20620 ;
  assign n28383 = n28381 & n28382 ;
  assign n28377 = n3985 & n20624 ;
  assign n28376 = n3837 & n20829 ;
  assign n28378 = n28377 ^ n28376 ;
  assign n28379 = n28378 ^ n3978 ;
  assign n28384 = n28383 ^ n28379 ;
  assign n28387 = n28386 ^ n28384 ;
  assign n28365 = n28256 ^ n27957 ;
  assign n28366 = n28365 ^ n28242 ;
  assign n28367 = n28256 ^ n28087 ;
  assign n28368 = n28367 ^ n28242 ;
  assign n28371 = n28259 & ~n28368 ;
  assign n28372 = n28371 ^ n28242 ;
  assign n28373 = ~n28366 & n28372 ;
  assign n28374 = n28373 ^ n28256 ;
  assign n28361 = n3518 & n23307 ;
  assign n28360 = n3807 & ~n23306 ;
  assign n28362 = n28361 ^ n28360 ;
  assign n28358 = ~n3850 & n20819 ;
  assign n28357 = n20631 & n22543 ;
  assign n28359 = n28358 ^ n28357 ;
  assign n28363 = n28362 ^ n28359 ;
  assign n28339 = n28241 ^ n27957 ;
  assign n28344 = n2173 ^ n1236 ;
  assign n28343 = n1506 ^ n511 ;
  assign n28345 = n28344 ^ n28343 ;
  assign n28346 = n28345 ^ n22520 ;
  assign n28340 = n14827 ^ n747 ;
  assign n28341 = n28340 ^ n14059 ;
  assign n28342 = n28341 ^ n828 ;
  assign n28347 = n28346 ^ n28342 ;
  assign n28348 = n28347 ^ n6059 ;
  assign n28349 = n28348 ^ n13651 ;
  assign n28350 = n28349 ^ n5567 ;
  assign n28351 = ~n3077 & ~n28350 ;
  assign n28352 = n28351 ^ x14 ;
  assign n28353 = n28352 ^ n28241 ;
  assign n28354 = n28353 ^ n28351 ;
  assign n28355 = ~n28339 & n28354 ;
  assign n28356 = n28355 ^ n28352 ;
  assign n28364 = n28363 ^ n28356 ;
  assign n28375 = n28374 ^ n28364 ;
  assign n28388 = n28387 ^ n28375 ;
  assign n28389 = n28388 ^ n28200 ;
  assign n28390 = n28389 ^ n28388 ;
  assign n28391 = n28390 ^ n28229 ;
  assign n28392 = ~n28261 & ~n28391 ;
  assign n28393 = n28392 ^ n28389 ;
  assign n28402 = n28401 ^ n28393 ;
  assign n28406 = n28405 ^ n28402 ;
  assign n28415 = n28414 ^ n28406 ;
  assign n28336 = n28288 ^ n28279 ;
  assign n28337 = ~n28280 & n28336 ;
  assign n28338 = n28337 ^ n28288 ;
  assign n28416 = n28415 ^ n28338 ;
  assign n28425 = n28424 ^ n28416 ;
  assign n28426 = n28425 ^ x17 ;
  assign n28335 = n20437 & n25308 ;
  assign n28427 = n28426 ^ n28335 ;
  assign n28332 = n28304 ^ n28300 ;
  assign n28333 = ~n28301 & n28332 ;
  assign n28334 = n28333 ^ n28304 ;
  assign n28428 = n28427 ^ n28334 ;
  assign n28446 = n28445 ^ n28428 ;
  assign n28329 = n28316 ^ n28312 ;
  assign n28330 = ~n28313 & ~n28329 ;
  assign n28331 = n28330 ^ n28316 ;
  assign n28447 = n28446 ^ n28331 ;
  assign n28451 = n28450 ^ n28447 ;
  assign n28555 = n28445 ^ n28331 ;
  assign n28556 = ~n28446 & ~n28555 ;
  assign n28557 = n28556 ^ n28445 ;
  assign n28554 = n28447 & n28450 ;
  assign n28558 = n28557 ^ n28554 ;
  assign n28548 = n13433 & n24841 ;
  assign n28546 = n5426 & ~n25282 ;
  assign n28539 = n25311 ^ x20 ;
  assign n28540 = n28539 ^ x19 ;
  assign n28541 = n28540 ^ n25311 ;
  assign n28542 = n25312 & ~n28541 ;
  assign n28543 = n28542 ^ n25311 ;
  assign n28544 = n5215 & n28543 ;
  assign n28545 = n28544 ^ x20 ;
  assign n28547 = n28546 ^ n28545 ;
  assign n28549 = n28548 ^ n28547 ;
  assign n28531 = n4651 & n20908 ;
  assign n28529 = ~n40 & n21147 ;
  assign n28522 = n21212 ^ x22 ;
  assign n28523 = n28522 ^ x23 ;
  assign n28524 = n28523 ^ n21212 ;
  assign n28525 = ~n25342 & n28524 ;
  assign n28526 = n28525 ^ n21212 ;
  assign n28527 = n35 & ~n28526 ;
  assign n28528 = n28527 ^ x23 ;
  assign n28530 = n28529 ^ n28528 ;
  assign n28532 = n28531 ^ n28530 ;
  assign n28514 = ~n4435 & n23893 ;
  assign n28512 = n20603 & ~n20614 ;
  assign n28509 = ~n4434 & ~n20612 ;
  assign n28508 = n4600 & ~n20613 ;
  assign n28510 = n28509 ^ n28508 ;
  assign n28511 = n28510 ^ x26 ;
  assign n28513 = n28512 ^ n28511 ;
  assign n28515 = n28514 ^ n28513 ;
  assign n28504 = n3837 & n20624 ;
  assign n28502 = n3985 & ~n20620 ;
  assign n28495 = n20617 ^ x29 ;
  assign n28496 = n28495 ^ x28 ;
  assign n28497 = n28496 ^ n20617 ;
  assign n28498 = ~n23490 & n28497 ;
  assign n28499 = n28498 ^ n20617 ;
  assign n28500 = n3833 & ~n28499 ;
  assign n28501 = n28500 ^ x29 ;
  assign n28503 = n28502 ^ n28501 ;
  assign n28505 = n28504 ^ n28503 ;
  assign n28486 = n22979 ^ n20819 ;
  assign n28489 = ~n61 & ~n28486 ;
  assign n28490 = n28489 ^ n22979 ;
  assign n28491 = n5280 & n28490 ;
  assign n28476 = n20829 ^ n12812 ;
  assign n28477 = n28476 ^ n20829 ;
  assign n28478 = n28477 ^ x31 ;
  assign n28481 = ~x31 & n20829 ;
  assign n28479 = n20628 ^ x31 ;
  assign n28480 = n6015 & ~n28479 ;
  assign n28482 = n28481 ^ n28480 ;
  assign n28483 = ~n28478 & n28482 ;
  assign n28484 = n28483 ^ n28481 ;
  assign n28485 = n28484 ^ x31 ;
  assign n28492 = n28491 ^ n28485 ;
  assign n28472 = n28363 ^ n28351 ;
  assign n28473 = ~n28356 & n28472 ;
  assign n28468 = n3666 ^ n3004 ;
  assign n28464 = n14736 ^ n3567 ;
  assign n28465 = n28464 ^ n6062 ;
  assign n28462 = n4838 ^ n2153 ;
  assign n28463 = n28462 ^ n2830 ;
  assign n28466 = n28465 ^ n28463 ;
  assign n28461 = n13495 ^ n673 ;
  assign n28467 = n28466 ^ n28461 ;
  assign n28469 = n28468 ^ n28467 ;
  assign n28470 = n5633 ^ n1967 ;
  assign n28471 = ~n28469 & ~n28470 ;
  assign n28474 = n28473 ^ n28471 ;
  assign n28493 = n28492 ^ n28474 ;
  assign n28506 = n28505 ^ n28493 ;
  assign n28458 = n28387 ^ n28374 ;
  assign n28459 = n28375 & n28458 ;
  assign n28460 = n28459 ^ n28387 ;
  assign n28507 = n28506 ^ n28460 ;
  assign n28516 = n28515 ^ n28507 ;
  assign n28518 = n28516 ^ n28388 ;
  assign n28517 = n28516 ^ n28401 ;
  assign n28519 = n28518 ^ n28517 ;
  assign n28520 = ~n28393 & ~n28519 ;
  assign n28521 = n28520 ^ n28518 ;
  assign n28533 = n28532 ^ n28521 ;
  assign n28534 = n28533 ^ n28414 ;
  assign n28535 = n28534 ^ n28405 ;
  assign n28536 = n28535 ^ n28533 ;
  assign n28537 = n28406 & n28536 ;
  assign n28538 = n28537 ^ n28534 ;
  assign n28550 = n28549 ^ n28538 ;
  assign n28551 = n28550 ^ x17 ;
  assign n28455 = n28424 ^ n28338 ;
  assign n28456 = n28416 & n28455 ;
  assign n28457 = n28456 ^ n28424 ;
  assign n28552 = n28551 ^ n28457 ;
  assign n28452 = n28425 ^ n28334 ;
  assign n28453 = ~n28427 & ~n28452 ;
  assign n28454 = n28453 ^ n28425 ;
  assign n28553 = n28552 ^ n28454 ;
  assign n28559 = n28558 ^ n28553 ;
  assign n28648 = n28549 ^ n28533 ;
  assign n28649 = n28538 & n28648 ;
  assign n28650 = n28649 ^ n28533 ;
  assign n28645 = n5221 & n25515 ;
  assign n28641 = n13433 ^ n5426 ;
  assign n28642 = n28641 ^ n28421 ;
  assign n28643 = n25282 & n28642 ;
  assign n28644 = n28643 ^ n13432 ;
  assign n28646 = n28645 ^ n28644 ;
  assign n28636 = n28532 ^ n28516 ;
  assign n28637 = n28521 & ~n28636 ;
  assign n28638 = n28637 ^ n28516 ;
  assign n28630 = n4655 & n24841 ;
  assign n28629 = n4651 & n21147 ;
  assign n28631 = n28630 ^ n28629 ;
  assign n28632 = n28631 ^ x23 ;
  assign n28628 = n4656 & ~n25528 ;
  assign n28633 = n28632 ^ n28628 ;
  assign n28627 = ~n40 & ~n21212 ;
  assign n28634 = n28633 ^ n28627 ;
  assign n28623 = n3985 & ~n20617 ;
  assign n28621 = n3837 & ~n20620 ;
  assign n28612 = x31 & ~n21231 ;
  assign n28613 = n28612 ^ n20624 ;
  assign n28614 = n28613 ^ n20829 ;
  assign n28609 = x31 & ~n24169 ;
  assign n28610 = n28609 ^ n20829 ;
  assign n28611 = ~n6015 & n28610 ;
  assign n28615 = n28614 ^ n28611 ;
  assign n28616 = ~n3518 & n28615 ;
  assign n28617 = n28616 ^ n28613 ;
  assign n28597 = n22513 ^ n794 ;
  assign n28596 = n2543 ^ n420 ;
  assign n28598 = n28597 ^ n28596 ;
  assign n28599 = n28598 ^ n1789 ;
  assign n28600 = n28599 ^ n12469 ;
  assign n28593 = n12522 ^ n478 ;
  assign n28592 = n801 ^ n318 ;
  assign n28594 = n28593 ^ n28592 ;
  assign n28591 = n3648 ^ n120 ;
  assign n28595 = n28594 ^ n28591 ;
  assign n28601 = n28600 ^ n28595 ;
  assign n28602 = n28601 ^ n1359 ;
  assign n28603 = n28602 ^ n5320 ;
  assign n28604 = ~n4529 & ~n28603 ;
  assign n28590 = n28471 ^ x17 ;
  assign n28605 = n28604 ^ n28590 ;
  assign n28587 = n28471 ^ n28363 ;
  assign n28588 = ~n28473 & n28587 ;
  assign n28589 = n28588 ^ n28363 ;
  assign n28606 = n28605 ^ n28589 ;
  assign n28618 = n28617 ^ n28606 ;
  assign n28619 = n28618 ^ x29 ;
  assign n28582 = n20614 ^ n5065 ;
  assign n28583 = n28582 ^ n20614 ;
  assign n28584 = ~n23479 & n28583 ;
  assign n28585 = n28584 ^ n20614 ;
  assign n28586 = n3833 & ~n28585 ;
  assign n28620 = n28619 ^ n28586 ;
  assign n28622 = n28621 ^ n28620 ;
  assign n28624 = n28623 ^ n28622 ;
  assign n28579 = n28505 ^ n28492 ;
  assign n28580 = n28493 & n28579 ;
  assign n28581 = n28580 ^ n28505 ;
  assign n28625 = n28624 ^ n28581 ;
  assign n28576 = ~n4434 & n20908 ;
  assign n28570 = n28515 ^ n28460 ;
  assign n28571 = n28507 & n28570 ;
  assign n28572 = n28571 ^ n28515 ;
  assign n28573 = n28572 ^ x26 ;
  assign n28569 = n20603 & ~n20613 ;
  assign n28574 = n28573 ^ n28569 ;
  assign n28568 = n4600 & ~n20612 ;
  assign n28575 = n28574 ^ n28568 ;
  assign n28577 = n28576 ^ n28575 ;
  assign n28567 = ~n4435 & ~n25056 ;
  assign n28578 = n28577 ^ n28567 ;
  assign n28626 = n28625 ^ n28578 ;
  assign n28635 = n28634 ^ n28626 ;
  assign n28639 = n28638 ^ n28635 ;
  assign n28647 = n28646 ^ n28639 ;
  assign n28651 = n28650 ^ n28647 ;
  assign n28652 = n28651 ^ x17 ;
  assign n28565 = n28550 ^ n28457 ;
  assign n28566 = n28551 & ~n28565 ;
  assign n28653 = n28652 ^ n28566 ;
  assign n28560 = n28554 ^ n28552 ;
  assign n28563 = n28553 & ~n28560 ;
  assign n28561 = n28560 ^ n28454 ;
  assign n28562 = ~n28557 & ~n28561 ;
  assign n28564 = n28563 ^ n28562 ;
  assign n28654 = n28653 ^ n28564 ;
  assign n28759 = n4656 & n25868 ;
  assign n28757 = n4651 & ~n21212 ;
  assign n28753 = n4655 & n25282 ;
  assign n28752 = ~n40 & n24841 ;
  assign n28754 = n28753 ^ n28752 ;
  assign n28755 = n28754 ^ n4655 ;
  assign n28756 = n28755 ^ x23 ;
  assign n28758 = n28757 ^ n28756 ;
  assign n28760 = n28759 ^ n28758 ;
  assign n28748 = ~n4435 & ~n25073 ;
  assign n28746 = ~n4434 & n21147 ;
  assign n28743 = n4600 & n20908 ;
  assign n28742 = n20603 & ~n20612 ;
  assign n28744 = n28743 ^ n28742 ;
  assign n28745 = n28744 ^ x26 ;
  assign n28747 = n28746 ^ n28745 ;
  assign n28749 = n28748 ^ n28747 ;
  assign n28734 = n3837 & ~n20617 ;
  assign n28732 = n3985 & ~n20614 ;
  assign n28725 = n20613 ^ x29 ;
  assign n28726 = n28725 ^ x28 ;
  assign n28727 = n28726 ^ n20613 ;
  assign n28728 = ~n21226 & n28727 ;
  assign n28729 = n28728 ^ n20613 ;
  assign n28730 = n3833 & ~n28729 ;
  assign n28731 = n28730 ^ x29 ;
  assign n28733 = n28732 ^ n28731 ;
  assign n28735 = n28734 ^ n28733 ;
  assign n28712 = n20620 ^ x30 ;
  assign n28713 = n28712 ^ n20620 ;
  assign n28714 = n20624 & n28713 ;
  assign n28715 = n28714 ^ n20620 ;
  assign n28716 = ~n3518 & ~n28715 ;
  assign n28717 = n28716 ^ n20620 ;
  assign n28718 = n28717 ^ n22968 ;
  assign n28705 = n22968 ^ n20624 ;
  assign n28704 = n22968 ^ n20829 ;
  assign n28706 = n28705 ^ n28704 ;
  assign n28707 = n28705 ^ x30 ;
  assign n28708 = n28707 ^ n28705 ;
  assign n28709 = n28706 & n28708 ;
  assign n28710 = n28709 ^ n28705 ;
  assign n28711 = ~n3518 & n28710 ;
  assign n28719 = n28718 ^ n28711 ;
  assign n28720 = x31 & ~n28719 ;
  assign n28721 = n28720 ^ n28717 ;
  assign n28695 = n14719 ^ n251 ;
  assign n28696 = n28695 ^ n585 ;
  assign n28694 = n1687 ^ n657 ;
  assign n28697 = n28696 ^ n28694 ;
  assign n28693 = n2924 ^ n1363 ;
  assign n28698 = n28697 ^ n28693 ;
  assign n28691 = n12628 ^ n4857 ;
  assign n28692 = n28691 ^ n6926 ;
  assign n28699 = n28698 ^ n28692 ;
  assign n28700 = n28699 ^ n1232 ;
  assign n28701 = n28700 ^ n3030 ;
  assign n28702 = n27119 ^ n6692 ;
  assign n28703 = ~n28701 & ~n28702 ;
  assign n28722 = n28721 ^ n28703 ;
  assign n28688 = n28617 ^ n28589 ;
  assign n28689 = n28606 & n28688 ;
  assign n28690 = n28689 ^ n28617 ;
  assign n28723 = n28722 ^ n28690 ;
  assign n28685 = n28604 ^ n28471 ;
  assign n28686 = n28590 & ~n28685 ;
  assign n28687 = n28686 ^ x17 ;
  assign n28724 = n28723 ^ n28687 ;
  assign n28736 = n28735 ^ n28724 ;
  assign n28737 = n28736 ^ n28618 ;
  assign n28738 = n28737 ^ n28736 ;
  assign n28739 = n28738 ^ n28581 ;
  assign n28740 = ~n28624 & ~n28739 ;
  assign n28741 = n28740 ^ n28737 ;
  assign n28750 = n28749 ^ n28741 ;
  assign n28682 = n28625 ^ n28572 ;
  assign n28683 = ~n28578 & ~n28682 ;
  assign n28684 = n28683 ^ n28625 ;
  assign n28751 = n28750 ^ n28684 ;
  assign n28761 = n28760 ^ n28751 ;
  assign n28762 = n28761 ^ x20 ;
  assign n28681 = n13433 & n25308 ;
  assign n28763 = n28762 ^ n28681 ;
  assign n28678 = n28638 ^ n28634 ;
  assign n28679 = n28635 & ~n28678 ;
  assign n28680 = n28679 ^ n28638 ;
  assign n28764 = n28763 ^ n28680 ;
  assign n28675 = n28650 ^ n28646 ;
  assign n28676 = ~n28647 & n28675 ;
  assign n28677 = n28676 ^ n28650 ;
  assign n28765 = n28764 ^ n28677 ;
  assign n28660 = n28557 ^ n28454 ;
  assign n28659 = n28454 & ~n28557 ;
  assign n28661 = n28660 ^ n28659 ;
  assign n28662 = n28651 ^ n28457 ;
  assign n28663 = n28651 ^ n28550 ;
  assign n28664 = n28652 & n28663 ;
  assign n28665 = n28662 & n28664 ;
  assign n28666 = n28665 ^ n28662 ;
  assign n28667 = n28666 ^ n28457 ;
  assign n28668 = ~n28661 & ~n28667 ;
  assign n28669 = n28659 ^ n28651 ;
  assign n28670 = n28659 ^ n28653 ;
  assign n28671 = n28670 ^ n28659 ;
  assign n28672 = ~n28669 & ~n28671 ;
  assign n28673 = n28672 ^ n28659 ;
  assign n28674 = ~n28668 & ~n28673 ;
  assign n28766 = n28765 ^ n28674 ;
  assign n28655 = n28557 ^ n28553 ;
  assign n28656 = n28554 & ~n28655 ;
  assign n28657 = n28653 ^ n28553 ;
  assign n28658 = n28656 & n28657 ;
  assign n28767 = n28766 ^ n28658 ;
  assign n28861 = n28753 ^ n4651 ;
  assign n28862 = ~n24841 & n28861 ;
  assign n28859 = n4651 ^ x23 ;
  assign n28857 = n4656 & n25311 ;
  assign n28856 = ~n40 & ~n25282 ;
  assign n28858 = n28857 ^ n28856 ;
  assign n28860 = n28859 ^ n28858 ;
  assign n28863 = n28862 ^ n28860 ;
  assign n28829 = n20603 & n20908 ;
  assign n28828 = n4600 & n21147 ;
  assign n28830 = n28829 ^ n28828 ;
  assign n28831 = n28830 ^ n97 ;
  assign n28832 = n28830 ^ x26 ;
  assign n28833 = n28832 ^ n99 ;
  assign n28834 = n28833 ^ x25 ;
  assign n28835 = n28834 ^ n28832 ;
  assign n28836 = n28835 ^ n21212 ;
  assign n28837 = n28836 ^ n21170 ;
  assign n28838 = n28837 ^ n28836 ;
  assign n28839 = n28832 & ~n28838 ;
  assign n28840 = n28839 ^ n28833 ;
  assign n28842 = ~n28835 & ~n28838 ;
  assign n28843 = n28842 ^ n21212 ;
  assign n28844 = ~n28833 & n28843 ;
  assign n28845 = ~n28840 & n28844 ;
  assign n28846 = n28845 ^ n28842 ;
  assign n28847 = n28846 ^ n99 ;
  assign n28848 = n28847 ^ n21212 ;
  assign n28849 = ~n28831 & ~n28848 ;
  assign n28826 = n3837 & ~n20614 ;
  assign n28824 = n3985 & ~n20613 ;
  assign n28787 = n28721 ^ n28690 ;
  assign n28819 = n28735 ^ n28690 ;
  assign n28820 = n28787 & ~n28819 ;
  assign n28814 = ~n3850 & n20620 ;
  assign n28806 = n20617 ^ n3518 ;
  assign n28807 = n28806 ^ n20617 ;
  assign n28808 = x30 & ~n20624 ;
  assign n28809 = n28808 ^ n20617 ;
  assign n28810 = ~n28807 & ~n28809 ;
  assign n28811 = n28810 ^ n20617 ;
  assign n28812 = n12812 & n28811 ;
  assign n28813 = n28812 ^ n3800 ;
  assign n28815 = n28814 ^ n28813 ;
  assign n28805 = n22005 & n23491 ;
  assign n28816 = n28815 ^ n28805 ;
  assign n28796 = n12902 ^ n182 ;
  assign n28797 = n28796 ^ n3061 ;
  assign n28795 = n2125 ^ n876 ;
  assign n28798 = n28797 ^ n28795 ;
  assign n28799 = n28798 ^ n26381 ;
  assign n28792 = n14736 ^ n975 ;
  assign n28793 = n28792 ^ n214 ;
  assign n28791 = n14040 ^ n1106 ;
  assign n28794 = n28793 ^ n28791 ;
  assign n28800 = n28799 ^ n28794 ;
  assign n28801 = n28800 ^ n4522 ;
  assign n28790 = n6713 ^ n4834 ;
  assign n28802 = n28801 ^ n28790 ;
  assign n28803 = ~n1383 & ~n28802 ;
  assign n28804 = n28803 ^ n28703 ;
  assign n28817 = n28816 ^ n28804 ;
  assign n28785 = n28703 ^ n28687 ;
  assign n28786 = n28735 ^ n28687 ;
  assign n28788 = n28787 ^ n28786 ;
  assign n28789 = n28785 & n28788 ;
  assign n28818 = n28817 ^ n28789 ;
  assign n28821 = n28820 ^ n28818 ;
  assign n28822 = n28821 ^ x29 ;
  assign n28780 = n20612 ^ n5065 ;
  assign n28781 = n28780 ^ n20612 ;
  assign n28782 = ~n23892 & n28781 ;
  assign n28783 = n28782 ^ n20612 ;
  assign n28784 = n3833 & ~n28783 ;
  assign n28823 = n28822 ^ n28784 ;
  assign n28825 = n28824 ^ n28823 ;
  assign n28827 = n28826 ^ n28825 ;
  assign n28850 = n28849 ^ n28827 ;
  assign n28852 = n28850 ^ n28736 ;
  assign n28851 = n28850 ^ n28749 ;
  assign n28853 = n28852 ^ n28851 ;
  assign n28854 = ~n28741 & n28853 ;
  assign n28855 = n28854 ^ n28852 ;
  assign n28864 = n28863 ^ n28855 ;
  assign n28865 = n28864 ^ x20 ;
  assign n28777 = n28760 ^ n28684 ;
  assign n28778 = ~n28751 & ~n28777 ;
  assign n28779 = n28778 ^ n28760 ;
  assign n28866 = n28865 ^ n28779 ;
  assign n28774 = n28761 ^ n28680 ;
  assign n28775 = n28763 & ~n28774 ;
  assign n28776 = n28775 ^ n28761 ;
  assign n28867 = n28866 ^ n28776 ;
  assign n28768 = n28674 ^ n28658 ;
  assign n28771 = n28677 ^ n28674 ;
  assign n28772 = ~n28768 & ~n28771 ;
  assign n28769 = n28768 ^ n28677 ;
  assign n28770 = n28764 & n28769 ;
  assign n28773 = n28772 ^ n28770 ;
  assign n28868 = n28867 ^ n28773 ;
  assign n28987 = n28864 ^ n28779 ;
  assign n28988 = n28865 & ~n28987 ;
  assign n28989 = n28988 ^ x20 ;
  assign n28984 = n4656 & n25515 ;
  assign n28980 = n4651 ^ n40 ;
  assign n28981 = n28980 ^ n28752 ;
  assign n28982 = n25282 & ~n28981 ;
  assign n28966 = ~x28 & ~n24096 ;
  assign n28974 = n28966 ^ n25056 ;
  assign n28975 = n4368 & ~n28974 ;
  assign n28970 = n3985 & ~n20612 ;
  assign n28969 = n3837 & ~n20613 ;
  assign n28971 = n28970 ^ n28969 ;
  assign n28972 = n28971 ^ n3978 ;
  assign n28967 = n28966 ^ n20908 ;
  assign n28968 = n28382 & ~n28967 ;
  assign n28973 = n28972 ^ n28968 ;
  assign n28976 = n28975 ^ n28973 ;
  assign n28947 = ~n28690 & ~n28735 ;
  assign n28948 = n28947 ^ n28819 ;
  assign n28949 = n28722 & n28785 ;
  assign n28950 = n28817 ^ n28687 ;
  assign n28951 = n28949 & ~n28950 ;
  assign n28952 = n28951 ^ n28817 ;
  assign n28953 = n28948 & ~n28952 ;
  assign n28954 = n28947 ^ n28817 ;
  assign n28956 = n28947 ^ n28721 ;
  assign n28955 = n28947 ^ n28687 ;
  assign n28957 = n28956 ^ n28955 ;
  assign n28958 = n28955 ^ n28785 ;
  assign n28959 = n28958 ^ n28955 ;
  assign n28960 = n28957 & ~n28959 ;
  assign n28961 = n28960 ^ n28955 ;
  assign n28962 = ~n28954 & ~n28961 ;
  assign n28963 = n28962 ^ n28817 ;
  assign n28964 = ~n28953 & n28963 ;
  assign n28942 = n52 & n20617 ;
  assign n28936 = x30 & ~n20617 ;
  assign n28937 = n28936 ^ n20614 ;
  assign n28938 = ~n3518 & ~n28937 ;
  assign n28939 = n28938 ^ n20614 ;
  assign n28940 = ~x31 & ~n28939 ;
  assign n28927 = n23480 ^ n3518 ;
  assign n28928 = n28927 ^ n23480 ;
  assign n28929 = x30 & n20620 ;
  assign n28930 = n28929 ^ n23480 ;
  assign n28931 = ~n28928 & ~n28930 ;
  assign n28932 = n28931 ^ n23480 ;
  assign n28933 = x31 & n28932 ;
  assign n28941 = n28940 ^ n28933 ;
  assign n28943 = n28941 ^ n28940 ;
  assign n28944 = n28942 & n28943 ;
  assign n28945 = n28944 ^ n28941 ;
  assign n28924 = n28816 ^ n28703 ;
  assign n28925 = ~n28804 & ~n28924 ;
  assign n28917 = n5637 ^ n1390 ;
  assign n28918 = n28917 ^ n1614 ;
  assign n28919 = n28918 ^ n14042 ;
  assign n28912 = n12780 ^ n717 ;
  assign n28911 = n1065 ^ n680 ;
  assign n28913 = n28912 ^ n28911 ;
  assign n28909 = n1915 ^ n429 ;
  assign n28908 = n427 ^ n157 ;
  assign n28910 = n28909 ^ n28908 ;
  assign n28914 = n28913 ^ n28910 ;
  assign n28915 = n28914 ^ n3003 ;
  assign n28916 = n28915 ^ n14726 ;
  assign n28920 = n28919 ^ n28916 ;
  assign n28921 = n28920 ^ n1477 ;
  assign n28922 = ~n4748 & ~n28921 ;
  assign n28923 = n28922 ^ x20 ;
  assign n28926 = n28925 ^ n28923 ;
  assign n28946 = n28945 ^ n28926 ;
  assign n28965 = n28964 ^ n28946 ;
  assign n28977 = n28976 ^ n28965 ;
  assign n28895 = ~x25 & ~n24810 ;
  assign n28898 = n28895 ^ n25528 ;
  assign n28899 = n99 & ~n28898 ;
  assign n28892 = n4600 & ~n21212 ;
  assign n28891 = n20603 & n21147 ;
  assign n28893 = n28892 ^ n28891 ;
  assign n28894 = n28893 ^ x26 ;
  assign n28896 = n28895 ^ n24841 ;
  assign n28897 = n28894 & ~n28896 ;
  assign n28900 = n28899 ^ n28897 ;
  assign n28901 = n28893 ^ n97 ;
  assign n28902 = ~n28900 & ~n28901 ;
  assign n28903 = n28902 ^ n28849 ;
  assign n28904 = n28903 ^ n28821 ;
  assign n28905 = n28904 ^ n28902 ;
  assign n28906 = n28827 & n28905 ;
  assign n28907 = n28906 ^ n28903 ;
  assign n28978 = n28977 ^ n28907 ;
  assign n28979 = n28978 ^ n28859 ;
  assign n28983 = n28982 ^ n28979 ;
  assign n28985 = n28984 ^ n28983 ;
  assign n28888 = n28863 ^ n28850 ;
  assign n28889 = n28855 & n28888 ;
  assign n28890 = n28889 ^ n28850 ;
  assign n28986 = n28985 ^ n28890 ;
  assign n28990 = n28989 ^ n28986 ;
  assign n28879 = n28776 ^ n28764 ;
  assign n28880 = n28879 ^ n28771 ;
  assign n28881 = n28880 ^ n28879 ;
  assign n28882 = n28776 ^ n28677 ;
  assign n28883 = n28882 ^ n28879 ;
  assign n28884 = ~n28881 & ~n28883 ;
  assign n28885 = n28884 ^ n28879 ;
  assign n28886 = n28867 & ~n28885 ;
  assign n28887 = n28886 ^ n28776 ;
  assign n28991 = n28990 ^ n28887 ;
  assign n28869 = n28764 ^ n28674 ;
  assign n28870 = n28869 ^ n28677 ;
  assign n28871 = n28658 & ~n28870 ;
  assign n28872 = n28867 ^ n28677 ;
  assign n28873 = n28872 ^ n28867 ;
  assign n28874 = n28867 ^ n28674 ;
  assign n28875 = n28874 ^ n28867 ;
  assign n28876 = n28873 & n28875 ;
  assign n28877 = n28876 ^ n28867 ;
  assign n28878 = n28871 & n28877 ;
  assign n28992 = n28991 ^ n28878 ;
  assign n29072 = ~n4435 & n25868 ;
  assign n29070 = ~n4434 & ~n25282 ;
  assign n29067 = n4600 & n24841 ;
  assign n29066 = n20603 & ~n21212 ;
  assign n29068 = n29067 ^ n29066 ;
  assign n29069 = n29068 ^ x26 ;
  assign n29071 = n29070 ^ n29069 ;
  assign n29073 = n29072 ^ n29071 ;
  assign n29056 = n20613 ^ n3518 ;
  assign n29055 = ~n3518 & n20613 ;
  assign n29057 = n29056 ^ n29055 ;
  assign n29054 = ~n61 & ~n20614 ;
  assign n29058 = n29057 ^ n29054 ;
  assign n29059 = n29058 ^ n21227 ;
  assign n29047 = n21227 ^ n20614 ;
  assign n29046 = n21227 ^ n20617 ;
  assign n29048 = n29047 ^ n29046 ;
  assign n29051 = x30 & n29048 ;
  assign n29052 = n29051 ^ n29047 ;
  assign n29053 = ~n3518 & ~n29052 ;
  assign n29060 = n29059 ^ n29053 ;
  assign n29061 = x31 & n29060 ;
  assign n29062 = n29061 ^ n29058 ;
  assign n29026 = n28922 ^ n28703 ;
  assign n29032 = n4046 ^ n1418 ;
  assign n29031 = n2349 ^ n2058 ;
  assign n29033 = n29032 ^ n29031 ;
  assign n29029 = n722 ^ n592 ;
  assign n29027 = n1128 ^ n234 ;
  assign n29028 = n29027 ^ n563 ;
  assign n29030 = n29029 ^ n29028 ;
  assign n29034 = n29033 ^ n29030 ;
  assign n29035 = n29034 ^ n2313 ;
  assign n29036 = n29035 ^ n4136 ;
  assign n29037 = n29036 ^ n13640 ;
  assign n29038 = n14830 ^ n4529 ;
  assign n29039 = n29038 ^ n2443 ;
  assign n29040 = ~n29037 & ~n29039 ;
  assign n29041 = n29040 ^ x20 ;
  assign n29042 = n29041 ^ n28922 ;
  assign n29043 = n29042 ^ n29040 ;
  assign n29044 = ~n29026 & n29043 ;
  assign n29045 = n29044 ^ n29041 ;
  assign n29063 = n29062 ^ n29045 ;
  assign n29023 = n3985 & n20908 ;
  assign n29017 = n28945 ^ n28923 ;
  assign n29018 = n29017 ^ n28703 ;
  assign n29019 = n28926 & ~n29018 ;
  assign n29020 = n29019 ^ n28945 ;
  assign n29021 = n29020 ^ x29 ;
  assign n29012 = n21147 ^ n5065 ;
  assign n29013 = n29012 ^ n21147 ;
  assign n29014 = ~n24078 & n29013 ;
  assign n29015 = n29014 ^ n21147 ;
  assign n29016 = n3833 & n29015 ;
  assign n29022 = n29021 ^ n29016 ;
  assign n29024 = n29023 ^ n29022 ;
  assign n29009 = n3837 & ~n20612 ;
  assign n29025 = n29024 ^ n29009 ;
  assign n29064 = n29063 ^ n29025 ;
  assign n29006 = n28976 ^ n28964 ;
  assign n29007 = n28965 & n29006 ;
  assign n29008 = n29007 ^ n28976 ;
  assign n29065 = n29064 ^ n29008 ;
  assign n29074 = n29073 ^ n29065 ;
  assign n29004 = n4651 & n25308 ;
  assign n29005 = n29004 ^ x23 ;
  assign n29075 = n29074 ^ n29005 ;
  assign n29001 = n28977 ^ n28902 ;
  assign n29002 = n28907 & n29001 ;
  assign n29003 = n29002 ^ n28902 ;
  assign n29076 = n29075 ^ n29003 ;
  assign n28998 = n28989 ^ n28887 ;
  assign n28999 = ~n28990 & n28998 ;
  assign n29000 = n28999 ^ n28989 ;
  assign n29077 = n29076 ^ n29000 ;
  assign n28996 = n28878 & ~n28991 ;
  assign n28993 = n28978 ^ n28890 ;
  assign n28994 = ~n28985 & ~n28993 ;
  assign n28995 = n28994 ^ n28978 ;
  assign n28997 = n28996 ^ n28995 ;
  assign n29078 = n29077 ^ n28997 ;
  assign n29151 = n29077 ^ n28996 ;
  assign n29152 = n28997 & n29151 ;
  assign n29144 = n3837 & n20908 ;
  assign n29142 = n3985 & n21147 ;
  assign n29138 = x31 & n29054 ;
  assign n29132 = n29062 ^ n29040 ;
  assign n29133 = ~n29045 & n29132 ;
  assign n29124 = n1322 ^ n236 ;
  assign n29123 = n438 ^ n108 ;
  assign n29125 = n29124 ^ n29123 ;
  assign n29122 = n14608 ^ n2962 ;
  assign n29126 = n29125 ^ n29122 ;
  assign n29120 = n2058 ^ n1631 ;
  assign n29119 = n1129 ^ n1050 ;
  assign n29121 = n29120 ^ n29119 ;
  assign n29127 = n29126 ^ n29121 ;
  assign n29128 = n29127 ^ n27124 ;
  assign n29129 = n29128 ^ n20586 ;
  assign n29130 = n29129 ^ n21698 ;
  assign n29131 = ~n4905 & ~n29130 ;
  assign n29134 = n29133 ^ n29131 ;
  assign n29118 = ~n61 & ~n20613 ;
  assign n29135 = n29134 ^ n29118 ;
  assign n29115 = x31 & ~n23892 ;
  assign n29116 = n29115 ^ n20612 ;
  assign n29117 = n3518 & n29116 ;
  assign n29136 = n29135 ^ n29117 ;
  assign n29110 = n12664 & ~n29055 ;
  assign n29137 = n29136 ^ n29110 ;
  assign n29139 = n29138 ^ n29137 ;
  assign n29107 = n29063 ^ n29020 ;
  assign n29108 = ~n29025 & ~n29107 ;
  assign n29109 = n29108 ^ n29063 ;
  assign n29140 = n29139 ^ n29109 ;
  assign n29141 = n29140 ^ x29 ;
  assign n29143 = n29142 ^ n29141 ;
  assign n29145 = n29144 ^ n29143 ;
  assign n29104 = n5065 & ~n25342 ;
  assign n29105 = n29104 ^ n21212 ;
  assign n29106 = n3833 & ~n29105 ;
  assign n29146 = n29145 ^ n29106 ;
  assign n29099 = n20603 & n24841 ;
  assign n29097 = n4600 ^ x26 ;
  assign n29096 = ~n4435 & n25311 ;
  assign n29098 = n29097 ^ n29096 ;
  assign n29100 = n29099 ^ n29098 ;
  assign n29093 = ~n4434 & ~n24841 ;
  assign n29094 = n29093 ^ n4600 ;
  assign n29095 = n25282 & n29094 ;
  assign n29101 = n29100 ^ n29095 ;
  assign n29147 = n29146 ^ n29101 ;
  assign n29086 = n29073 ^ n29008 ;
  assign n29087 = n29065 & n29086 ;
  assign n29088 = n29087 ^ n29073 ;
  assign n29148 = n29147 ^ n29088 ;
  assign n29149 = n29148 ^ x23 ;
  assign n29079 = n29005 ^ n29003 ;
  assign n29081 = n29003 ^ n29000 ;
  assign n29084 = n29079 & n29081 ;
  assign n29082 = n29081 ^ n29005 ;
  assign n29083 = ~n29074 & n29082 ;
  assign n29085 = n29084 ^ n29083 ;
  assign n29150 = n29149 ^ n29085 ;
  assign n29153 = n29152 ^ n29150 ;
  assign n29218 = n29003 ^ n28995 ;
  assign n29217 = n29074 ^ n29003 ;
  assign n29221 = n29149 ^ n29003 ;
  assign n29222 = ~n29217 & ~n29221 ;
  assign n29223 = ~n29218 & n29222 ;
  assign n29224 = n29223 ^ n29149 ;
  assign n29255 = n29224 ^ n29005 ;
  assign n29256 = n29255 ^ n29149 ;
  assign n29257 = n29256 ^ n29224 ;
  assign n29219 = n29217 & ~n29218 ;
  assign n29220 = n29219 ^ n29074 ;
  assign n29258 = n29257 ^ n29220 ;
  assign n29259 = n29258 ^ n29000 ;
  assign n29248 = n29149 ^ n29005 ;
  assign n29249 = n29248 ^ n29000 ;
  assign n29250 = n29249 ^ n29220 ;
  assign n29226 = n29005 ^ n29000 ;
  assign n29230 = n29226 ^ n29000 ;
  assign n29231 = n29230 ^ n29224 ;
  assign n29234 = n29231 ^ n29149 ;
  assign n29235 = n29234 ^ n29224 ;
  assign n29232 = n29231 ^ n29220 ;
  assign n29233 = n29232 ^ n29224 ;
  assign n29236 = n29235 ^ n29233 ;
  assign n29237 = n29224 & n29236 ;
  assign n29238 = n29237 ^ n29231 ;
  assign n29239 = n29224 ^ n29000 ;
  assign n29240 = n29239 ^ n29235 ;
  assign n29241 = n29236 & ~n29240 ;
  assign n29242 = n29241 ^ n29239 ;
  assign n29243 = ~n29231 & ~n29242 ;
  assign n29244 = ~n29238 & n29243 ;
  assign n29245 = n29244 ^ n29241 ;
  assign n29246 = n29245 ^ n29226 ;
  assign n29247 = n29246 ^ n29239 ;
  assign n29251 = n29250 ^ n29247 ;
  assign n29252 = n29251 ^ n29239 ;
  assign n29227 = n29226 ^ n29149 ;
  assign n29253 = n29252 ^ n29227 ;
  assign n29225 = n29224 ^ n29220 ;
  assign n29228 = n29227 ^ n29225 ;
  assign n29229 = n29228 ^ n29220 ;
  assign n29254 = n29253 ^ n29229 ;
  assign n29260 = n29259 ^ n29254 ;
  assign n29212 = n29088 ^ x23 ;
  assign n29213 = ~n29148 & n29212 ;
  assign n29214 = n29213 ^ x23 ;
  assign n29209 = n29140 ^ n29101 ;
  assign n29210 = n29146 & n29209 ;
  assign n29211 = n29210 ^ n29140 ;
  assign n29215 = n29214 ^ n29211 ;
  assign n29204 = ~n4435 & n25515 ;
  assign n29203 = n20603 & ~n25282 ;
  assign n29205 = n29204 ^ n29203 ;
  assign n29206 = n29205 ^ x26 ;
  assign n29202 = n4600 & n25308 ;
  assign n29207 = n29206 ^ n29202 ;
  assign n29198 = n3837 & n21147 ;
  assign n29196 = n3985 & ~n21212 ;
  assign n29189 = n24841 ^ x29 ;
  assign n29190 = n29189 ^ x28 ;
  assign n29191 = n29190 ^ n24841 ;
  assign n29192 = ~n27272 & n29191 ;
  assign n29193 = n29192 ^ n24841 ;
  assign n29194 = n3833 & n29193 ;
  assign n29195 = n29194 ^ x29 ;
  assign n29197 = n29196 ^ n29195 ;
  assign n29199 = n29198 ^ n29197 ;
  assign n29185 = ~n3850 & ~n20612 ;
  assign n29184 = x31 & n29118 ;
  assign n29186 = n29185 ^ n29184 ;
  assign n29178 = n25056 ^ n20908 ;
  assign n29181 = x31 & ~n29178 ;
  assign n29182 = n29181 ^ n20908 ;
  assign n29183 = n3518 & n29182 ;
  assign n29187 = n29186 ^ n29183 ;
  assign n29173 = n29131 ^ n29062 ;
  assign n29174 = ~n29133 & n29173 ;
  assign n29175 = n29174 ^ n29062 ;
  assign n29168 = n5345 ^ n1884 ;
  assign n29165 = n1935 ^ n199 ;
  assign n29166 = n29165 ^ n896 ;
  assign n29163 = n5560 ^ n1021 ;
  assign n29162 = n2126 ^ n228 ;
  assign n29164 = n29163 ^ n29162 ;
  assign n29167 = n29166 ^ n29164 ;
  assign n29169 = n29168 ^ n29167 ;
  assign n29170 = n29169 ^ n71 ;
  assign n29171 = n29170 ^ n3606 ;
  assign n29161 = n29131 ^ x23 ;
  assign n29172 = n29171 ^ n29161 ;
  assign n29176 = n29175 ^ n29172 ;
  assign n29188 = n29187 ^ n29176 ;
  assign n29200 = n29199 ^ n29188 ;
  assign n29158 = n29134 ^ n29109 ;
  assign n29159 = ~n29139 & n29158 ;
  assign n29160 = n29159 ^ n29134 ;
  assign n29201 = n29200 ^ n29160 ;
  assign n29208 = n29207 ^ n29201 ;
  assign n29216 = n29215 ^ n29208 ;
  assign n29261 = n29260 ^ n29216 ;
  assign n29154 = n29150 ^ n28995 ;
  assign n29155 = n29077 ^ n28995 ;
  assign n29156 = n28996 & ~n29155 ;
  assign n29157 = ~n29154 & n29156 ;
  assign n29262 = n29261 ^ n29157 ;
  assign n29339 = n29211 & n29214 ;
  assign n29338 = ~n29201 & ~n29207 ;
  assign n29340 = n29339 ^ n29338 ;
  assign n29317 = n3985 & n24841 ;
  assign n29316 = n3837 & ~n21212 ;
  assign n29318 = n29317 ^ n29316 ;
  assign n29319 = n29318 ^ n3978 ;
  assign n29323 = n29318 ^ x29 ;
  assign n29324 = n29323 ^ n4368 ;
  assign n29320 = n25282 ^ n4368 ;
  assign n29321 = n29320 ^ x28 ;
  assign n29322 = n29321 ^ n25282 ;
  assign n29325 = n29324 ^ n29322 ;
  assign n29326 = n29325 ^ n29324 ;
  assign n29328 = ~n25299 & ~n29326 ;
  assign n29329 = ~x28 & n29328 ;
  assign n29332 = n29329 ^ n29328 ;
  assign n29330 = n29329 ^ n25282 ;
  assign n29331 = n29324 & n29330 ;
  assign n29333 = n29332 ^ n29331 ;
  assign n29334 = n29333 ^ n4368 ;
  assign n29335 = ~n29319 & ~n29334 ;
  assign n29308 = x30 & n20908 ;
  assign n29294 = n25073 ^ n20612 ;
  assign n29293 = n25073 ^ n20908 ;
  assign n29295 = n29294 ^ n29293 ;
  assign n29298 = ~x30 & ~n29295 ;
  assign n29299 = n29298 ^ n29294 ;
  assign n29300 = ~n3518 & n29299 ;
  assign n29301 = n29300 ^ n25073 ;
  assign n29302 = n29301 ^ n21147 ;
  assign n29303 = n29302 ^ n29301 ;
  assign n29309 = n29308 ^ n29303 ;
  assign n29310 = ~n3518 & n29309 ;
  assign n29311 = n29310 ^ n29302 ;
  assign n29312 = ~x31 & ~n29311 ;
  assign n29313 = n29312 ^ n29301 ;
  assign n29289 = n29171 ^ n29131 ;
  assign n29290 = n29161 & ~n29289 ;
  assign n29291 = n29290 ^ x23 ;
  assign n29275 = n21118 ^ n14280 ;
  assign n29280 = n514 ^ n158 ;
  assign n29278 = n5539 ^ n3756 ;
  assign n29277 = n4838 ^ n2383 ;
  assign n29279 = n29278 ^ n29277 ;
  assign n29281 = n29280 ^ n29279 ;
  assign n29276 = ~n70 & ~n2206 ;
  assign n29282 = n29281 ^ n29276 ;
  assign n29283 = ~n29275 & n29282 ;
  assign n29284 = n12841 ^ n2437 ;
  assign n29285 = n29284 ^ n14008 ;
  assign n29286 = n29285 ^ n425 ;
  assign n29287 = n29283 & ~n29286 ;
  assign n29288 = ~n14635 & n29287 ;
  assign n29292 = n29291 ^ n29288 ;
  assign n29314 = n29313 ^ n29292 ;
  assign n29272 = n29187 ^ n29175 ;
  assign n29273 = n29176 & n29272 ;
  assign n29274 = n29273 ^ n29187 ;
  assign n29315 = n29314 ^ n29274 ;
  assign n29336 = n29335 ^ n29315 ;
  assign n29270 = n20603 & n25308 ;
  assign n29266 = n29199 ^ n29160 ;
  assign n29267 = ~n29200 & ~n29266 ;
  assign n29268 = n29267 ^ n29199 ;
  assign n29269 = n29268 ^ x26 ;
  assign n29271 = n29270 ^ n29269 ;
  assign n29337 = n29336 ^ n29271 ;
  assign n29341 = n29340 ^ n29337 ;
  assign n29264 = n29260 ^ n29215 ;
  assign n29265 = n29216 & n29264 ;
  assign n29342 = n29341 ^ n29265 ;
  assign n29263 = n29157 & ~n29261 ;
  assign n29343 = n29342 ^ n29263 ;
  assign n29415 = n3837 & n24841 ;
  assign n29413 = n3985 & ~n25282 ;
  assign n29406 = n25311 ^ x29 ;
  assign n29407 = n29406 ^ x28 ;
  assign n29408 = n29407 ^ n25311 ;
  assign n29409 = n25312 & ~n29408 ;
  assign n29410 = n29409 ^ n25311 ;
  assign n29411 = n3833 & n29410 ;
  assign n29412 = n29411 ^ x29 ;
  assign n29414 = n29413 ^ n29412 ;
  assign n29416 = n29415 ^ n29414 ;
  assign n29398 = n29313 ^ n29291 ;
  assign n29399 = ~n29292 & ~n29398 ;
  assign n29392 = n171 ^ n169 ;
  assign n29391 = n367 ^ n129 ;
  assign n29393 = n29392 ^ n29391 ;
  assign n29394 = n21118 ^ n295 ;
  assign n29395 = n29394 ^ n255 ;
  assign n29396 = n29393 & ~n29395 ;
  assign n29397 = ~n3542 & n29396 ;
  assign n29400 = n29399 ^ n29397 ;
  assign n29371 = n21147 ^ x31 ;
  assign n29372 = n29371 ^ n52 ;
  assign n29373 = n29372 ^ n3805 ;
  assign n29401 = n29400 ^ n29373 ;
  assign n29376 = n29373 ^ n21212 ;
  assign n29377 = n29376 ^ n29373 ;
  assign n29380 = ~n52 & ~n29377 ;
  assign n29381 = n29380 ^ n29373 ;
  assign n29382 = ~x31 & ~n29381 ;
  assign n29402 = n29401 ^ n29382 ;
  assign n29385 = n25341 ^ n20908 ;
  assign n29388 = n61 & n29385 ;
  assign n29389 = n29388 ^ n20908 ;
  assign n29390 = n5280 & ~n29389 ;
  assign n29403 = n29402 ^ n29390 ;
  assign n29374 = n29373 ^ x31 ;
  assign n29375 = n29373 ^ n21147 ;
  assign n29383 = ~n29375 & ~n29382 ;
  assign n29384 = ~n29374 & n29383 ;
  assign n29404 = n29403 ^ n29384 ;
  assign n29405 = n29404 ^ x26 ;
  assign n29417 = n29416 ^ n29405 ;
  assign n29368 = n29335 ^ n29274 ;
  assign n29369 = ~n29315 & ~n29368 ;
  assign n29370 = n29369 ^ n29335 ;
  assign n29418 = n29417 ^ n29370 ;
  assign n29349 = n29260 & ~n29339 ;
  assign n29350 = n29338 & n29349 ;
  assign n29345 = n29337 & ~n29339 ;
  assign n29351 = n29350 ^ n29345 ;
  assign n29346 = n29339 ^ n29215 ;
  assign n29347 = n29201 & n29346 ;
  assign n29348 = n29345 & n29347 ;
  assign n29352 = n29351 ^ n29348 ;
  assign n29353 = n29260 ^ n29207 ;
  assign n29354 = n29345 ^ n29201 ;
  assign n29355 = n29354 ^ n29207 ;
  assign n29356 = ~n29353 & n29355 ;
  assign n29357 = n29356 ^ n29207 ;
  assign n29358 = ~n29352 & ~n29357 ;
  assign n29360 = ~n29337 & n29346 ;
  assign n29361 = n29358 & n29360 ;
  assign n29359 = n29358 ^ n29352 ;
  assign n29362 = n29361 ^ n29359 ;
  assign n29364 = n29362 ^ n29336 ;
  assign n29363 = n29362 ^ n29268 ;
  assign n29365 = n29364 ^ n29363 ;
  assign n29366 = ~n29271 & ~n29365 ;
  assign n29367 = n29366 ^ n29364 ;
  assign n29419 = n29418 ^ n29367 ;
  assign n29344 = n29263 & n29342 ;
  assign n29420 = n29419 ^ n29344 ;
  assign n29455 = n29400 ^ n29370 ;
  assign n29427 = n29416 ^ x26 ;
  assign n29456 = n29455 ^ n29427 ;
  assign n29457 = ~n29404 & n29456 ;
  assign n29450 = n29397 ^ n29291 ;
  assign n29451 = n29399 & ~n29450 ;
  assign n29447 = n3503 ^ n363 ;
  assign n29446 = x29 ^ x26 ;
  assign n29448 = n29447 ^ n29446 ;
  assign n29434 = ~x30 & n24806 ;
  assign n29435 = n29434 ^ n21147 ;
  assign n29436 = n12812 & ~n29435 ;
  assign n29437 = n29436 ^ x30 ;
  assign n29449 = n29448 ^ n29437 ;
  assign n29452 = n29451 ^ n29449 ;
  assign n29438 = n29437 ^ n24841 ;
  assign n29441 = n29438 ^ n24810 ;
  assign n29442 = n29441 ^ n29438 ;
  assign n29443 = x31 & ~n29442 ;
  assign n29444 = n29443 ^ n29438 ;
  assign n29445 = n3518 & n29444 ;
  assign n29453 = n29452 ^ n29445 ;
  assign n29430 = n3983 & n25515 ;
  assign n29429 = n3837 & ~n25282 ;
  assign n29431 = n29430 ^ n29429 ;
  assign n29454 = n29453 ^ n29431 ;
  assign n29458 = n29457 ^ n29454 ;
  assign n29426 = n29416 ^ n29370 ;
  assign n29428 = n29426 & ~n29427 ;
  assign n29459 = n29458 ^ n29428 ;
  assign n29422 = n29418 ^ n29344 ;
  assign n29423 = n29367 ^ n29344 ;
  assign n29424 = n29422 & n29423 ;
  assign n29421 = n29362 & ~n29367 ;
  assign n29425 = n29424 ^ n29421 ;
  assign n29460 = n29459 ^ n29425 ;
  assign y0 = ~n24794 ;
  assign y1 = ~n25064 ;
  assign y2 = ~n25307 ;
  assign y3 = ~n25506 ;
  assign y4 = n25696 ;
  assign y5 = ~n25892 ;
  assign y6 = n26082 ;
  assign y7 = ~n26289 ;
  assign y8 = ~n26487 ;
  assign y9 = n26693 ;
  assign y10 = n26874 ;
  assign y11 = ~n27076 ;
  assign y12 = n27262 ;
  assign y13 = n27443 ;
  assign y14 = n27595 ;
  assign y15 = ~n27765 ;
  assign y16 = n27913 ;
  assign y17 = n28061 ;
  assign y18 = ~n28189 ;
  assign y19 = n28328 ;
  assign y20 = n28451 ;
  assign y21 = ~n28559 ;
  assign y22 = ~n28654 ;
  assign y23 = ~n28767 ;
  assign y24 = ~n28868 ;
  assign y25 = ~n28992 ;
  assign y26 = ~n29078 ;
  assign y27 = ~n29153 ;
  assign y28 = ~n29262 ;
  assign y29 = n29343 ;
  assign y30 = ~n29420 ;
  assign y31 = n29460 ;
endmodule
